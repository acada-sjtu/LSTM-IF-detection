
module leon3mp ( resetn, clk, pllref, errorn, address, datain, dataout, 
        datadir, dsutx, dsurx, dsuen, dsubre, dsuact, txd1, rxd1, txd2, rxd2, 
        ramsn, ramoen, rwen, oen, writen, read, iosn, romsn, tck, tms, tdi, 
        tdo, ic_address, ic_data, ic_wren, ic_ce, ic_q, it_address, it_data, 
        it_wren, it_ce, it_q, dc_address, dc_data, dc_wren, dc_ce, dc_q, 
        dt_address, dt_data, dt_wren, dt_ce, dt_q, clk_out, rf_ce_a, rf_addr_a, 
        rf_do_a, rf_ce_b, rf_addr_b, rf_do_b, rf_ce_w, rf_we_w, rf_addr_w, 
        rf_di_w );
  output [27:0] address;
  input [31:0] datain;
  output [31:0] dataout;
  output [3:0] datadir;
  output [4:0] ramsn;
  output [4:0] ramoen;
  output [3:0] rwen;
  output [1:0] romsn;
  output [9:0] ic_address;
  output [31:0] ic_data;
  input [31:0] ic_q;
  output [6:0] it_address;
  output [27:0] it_data;
  input [27:0] it_q;
  output [9:0] dc_address;
  output [31:0] dc_data;
  input [31:0] dc_q;
  output [6:0] dt_address;
  output [27:0] dt_data;
  input [27:0] dt_q;
  output [7:0] rf_addr_a;
  input [31:0] rf_do_a;
  output [7:0] rf_addr_b;
  input [31:0] rf_do_b;
  output [7:0] rf_addr_w;
  output [31:0] rf_di_w;
  input resetn, clk, pllref, dsurx, dsuen, dsubre, rxd1, rxd2, tck, tms, tdi;
  output errorn, dsutx, dsuact, txd1, txd2, oen, writen, read, iosn, tdo,
         ic_wren, ic_ce, it_wren, it_ce, dc_wren, dc_ce, dt_wren, dt_ce,
         clk_out, rf_ce_a, rf_ce_b, rf_ce_w, rf_we_w;
  wire   rstn, ahbso_1__HREADY_, ahbso_1__HRDATA__31_, ahbso_1__HRDATA__30_,
         ahbso_1__HRDATA__29_, ahbso_1__HRDATA__28_, ahbso_1__HRDATA__27_,
         ahbso_1__HRDATA__26_, ahbso_1__HRDATA__25_, ahbso_1__HRDATA__24_,
         ahbso_1__HRDATA__23_, ahbso_1__HRDATA__22_, ahbso_1__HRDATA__21_,
         ahbso_1__HRDATA__20_, ahbso_1__HRDATA__19_, ahbso_1__HRDATA__18_,
         ahbso_1__HRDATA__17_, ahbso_1__HRDATA__16_, ahbso_1__HRDATA__15_,
         ahbso_1__HRDATA__14_, ahbso_1__HRDATA__13_, ahbso_1__HRDATA__12_,
         ahbso_1__HRDATA__11_, ahbso_1__HRDATA__10_, ahbso_1__HRDATA__9_,
         ahbso_1__HRDATA__8_, ahbso_1__HRDATA__7_, ahbso_1__HRDATA__6_,
         ahbso_1__HRDATA__5_, ahbso_1__HRDATA__4_, ahbso_1__HRDATA__3_,
         ahbso_1__HRDATA__2_, ahbso_1__HRDATA__1_, ahbso_1__HRDATA__0_,
         ahbso_0__HRESP__0_, ahbso_0__HRDATA__31_, ahbso_0__HRDATA__30_,
         ahbso_0__HRDATA__29_, ahbso_0__HRDATA__28_, ahbso_0__HRDATA__27_,
         ahbso_0__HRDATA__26_, ahbso_0__HRDATA__25_, ahbso_0__HRDATA__24_,
         ahbso_0__HRDATA__23_, ahbso_0__HRDATA__22_, ahbso_0__HRDATA__21_,
         ahbso_0__HRDATA__20_, ahbso_0__HRDATA__19_, ahbso_0__HRDATA__18_,
         ahbso_0__HRDATA__17_, ahbso_0__HRDATA__16_, ahbso_0__HRDATA__15_,
         ahbso_0__HRDATA__14_, ahbso_0__HRDATA__13_, ahbso_0__HRDATA__12_,
         ahbso_0__HRDATA__11_, ahbso_0__HRDATA__10_, ahbso_0__HRDATA__9_,
         ahbso_0__HRDATA__8_, ahbso_0__HRDATA__7_, ahbso_0__HRDATA__6_,
         ahbso_0__HRDATA__5_, ahbso_0__HRDATA__4_, ahbso_0__HRDATA__3_,
         ahbso_0__HRDATA__2_, ahbso_0__HRDATA__1_, ahbso_0__HRDATA__0_,
         irqi_0__IRL__0_, apbo_1__PIRQ__2_, rst0_r_1_, rst0_r_3_,
         ahb0_r_HRDATAS__1_, ahb0_r_HRDATAS__4_, ahb0_r_HRDATAS__5_,
         ahb0_r_HRDATAS__6_, ahb0_r_HRDATAS__7_, ahb0_r_HRDATAS__8_,
         ahb0_r_HRDATAS__9_, ahb0_r_HRDATAS__10_, ahb0_r_HRDATAS__11_,
         ahb0_r_HRDATAS__12_, ahb0_r_HRDATAS__13_, ahb0_r_HRDATAS__14_,
         ahb0_r_HRDATAS__15_, ahb0_r_HRDATAS__16_, ahb0_r_HRDATAS__17_,
         ahb0_r_HRDATAS__24_, ahb0_r_HRDATAS__26_, ahb0_r_HRDATAS__29_,
         ahb0_r_HRDATAS__30_, ahb0_r_HRDATAS__31_, ahb0_r_HRDATAM__5_,
         ahb0_r_HRDATAM__6_, ahb0_r_HRDATAM__12_, ahb0_r_HRDATAM__13_,
         ahb0_r_HRDATAM__24_, ahb0_r_CFGA11_, ahb0_r_HADDR__2_,
         ahb0_r_HADDR__3_, ahb0_r_HADDR__5_, ahb0_r_HADDR__6_,
         ahb0_r_HADDR__7_, ahb0_r_HADDR__8_, ahb0_r_HADDR__9_,
         ahb0_r_HADDR__10_, ahb0_r_HTRANS__1_, ahb0_r_DEFSLV_,
         ahb0_r_HMASTERD_, ahb0_v_CFGSEL_, ahb0_v_HADDR__4_, ahb0_v_HREADY_,
         ahb0_v_HSLAVE__0_, u0_0_dbgo_SU_, u0_0_dbgo_OPTYPE__0_,
         u0_0_dbgo_OPTYPE__1_, u0_0_dbgo_OPTYPE__2_, u0_0_dbgo_OPTYPE__3_,
         u0_0_dbgo_OPTYPE__4_, u0_0_dbgo_OPTYPE__5_, u0_0_leon3x0_p0_dco_HIT_,
         u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__0_,
         u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__1_,
         u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DCS__1_,
         u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__IFRZ_,
         u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DFRZ_,
         u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__BURST_,
         u0_0_leon3x0_p0_dco_ICDIAG__ENABLE_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__0_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__1_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__3_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__4_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__5_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__6_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__7_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__8_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__9_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__10_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__11_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__12_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__13_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__14_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__15_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__16_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__17_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__18_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__19_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__20_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__21_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__22_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__23_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__24_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__25_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__26_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__27_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__28_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__29_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__30_,
         u0_0_leon3x0_p0_dco_ICDIAG__ADDR__31_, u0_0_leon3x0_p0_dco_WERR_,
         u0_0_leon3x0_p0_ico_DIAGRDY_, u0_0_leon3x0_p0_iu_N5495,
         u0_0_leon3x0_p0_iu_N5494, u0_0_leon3x0_p0_iu_N5493,
         u0_0_leon3x0_p0_iu_N5492, u0_0_leon3x0_p0_iu_N5491,
         u0_0_leon3x0_p0_iu_N5490, u0_0_leon3x0_p0_iu_N5489,
         u0_0_leon3x0_p0_iu_N5488, u0_0_leon3x0_p0_iu_N5487,
         u0_0_leon3x0_p0_iu_N5486, u0_0_leon3x0_p0_iu_N5485,
         u0_0_leon3x0_p0_iu_N5484, u0_0_leon3x0_p0_iu_N5483,
         u0_0_leon3x0_p0_iu_N5482, u0_0_leon3x0_p0_iu_N5481,
         u0_0_leon3x0_p0_iu_N5480, u0_0_leon3x0_p0_iu_N5479,
         u0_0_leon3x0_p0_iu_N5478, u0_0_leon3x0_p0_iu_N5477,
         u0_0_leon3x0_p0_iu_N5476, u0_0_leon3x0_p0_iu_N5475,
         u0_0_leon3x0_p0_iu_N5474, u0_0_leon3x0_p0_iu_N5473,
         u0_0_leon3x0_p0_iu_N5472, u0_0_leon3x0_p0_iu_N5471,
         u0_0_leon3x0_p0_iu_N5470, u0_0_leon3x0_p0_iu_N5469,
         u0_0_leon3x0_p0_iu_N5468, u0_0_leon3x0_p0_iu_N5467,
         u0_0_leon3x0_p0_iu_fe_npc_3_, u0_0_leon3x0_p0_iu_fe_npc_4_,
         u0_0_leon3x0_p0_iu_fe_npc_5_, u0_0_leon3x0_p0_iu_fe_npc_6_,
         u0_0_leon3x0_p0_iu_fe_npc_7_, u0_0_leon3x0_p0_iu_fe_npc_8_,
         u0_0_leon3x0_p0_iu_fe_npc_9_, u0_0_leon3x0_p0_iu_fe_npc_10_,
         u0_0_leon3x0_p0_iu_fe_npc_11_, u0_0_leon3x0_p0_iu_fe_npc_12_,
         u0_0_leon3x0_p0_iu_fe_npc_13_, u0_0_leon3x0_p0_iu_fe_npc_14_,
         u0_0_leon3x0_p0_iu_fe_npc_15_, u0_0_leon3x0_p0_iu_fe_npc_16_,
         u0_0_leon3x0_p0_iu_fe_npc_17_, u0_0_leon3x0_p0_iu_fe_npc_18_,
         u0_0_leon3x0_p0_iu_fe_npc_19_, u0_0_leon3x0_p0_iu_fe_npc_20_,
         u0_0_leon3x0_p0_iu_fe_npc_21_, u0_0_leon3x0_p0_iu_fe_npc_22_,
         u0_0_leon3x0_p0_iu_fe_npc_23_, u0_0_leon3x0_p0_iu_fe_npc_24_,
         u0_0_leon3x0_p0_iu_fe_npc_25_, u0_0_leon3x0_p0_iu_fe_npc_26_,
         u0_0_leon3x0_p0_iu_fe_npc_27_, u0_0_leon3x0_p0_iu_fe_npc_28_,
         u0_0_leon3x0_p0_iu_fe_npc_29_, u0_0_leon3x0_p0_iu_fe_npc_30_,
         u0_0_leon3x0_p0_iu_fe_npc_31_, u0_0_leon3x0_p0_iu_fe_pc_2_,
         u0_0_leon3x0_p0_iu_fe_pc_3_, u0_0_leon3x0_p0_iu_fe_pc_4_,
         u0_0_leon3x0_p0_iu_fe_pc_5_, u0_0_leon3x0_p0_iu_fe_pc_6_,
         u0_0_leon3x0_p0_iu_fe_pc_7_, u0_0_leon3x0_p0_iu_fe_pc_8_,
         u0_0_leon3x0_p0_iu_fe_pc_9_, u0_0_leon3x0_p0_iu_fe_pc_10_,
         u0_0_leon3x0_p0_iu_fe_pc_11_, u0_0_leon3x0_p0_iu_fe_pc_12_,
         u0_0_leon3x0_p0_iu_fe_pc_13_, u0_0_leon3x0_p0_iu_fe_pc_14_,
         u0_0_leon3x0_p0_iu_fe_pc_15_, u0_0_leon3x0_p0_iu_fe_pc_16_,
         u0_0_leon3x0_p0_iu_fe_pc_17_, u0_0_leon3x0_p0_iu_fe_pc_18_,
         u0_0_leon3x0_p0_iu_fe_pc_19_, u0_0_leon3x0_p0_iu_fe_pc_20_,
         u0_0_leon3x0_p0_iu_fe_pc_21_, u0_0_leon3x0_p0_iu_fe_pc_22_,
         u0_0_leon3x0_p0_iu_fe_pc_23_, u0_0_leon3x0_p0_iu_fe_pc_24_,
         u0_0_leon3x0_p0_iu_fe_pc_25_, u0_0_leon3x0_p0_iu_fe_pc_26_,
         u0_0_leon3x0_p0_iu_fe_pc_27_, u0_0_leon3x0_p0_iu_fe_pc_28_,
         u0_0_leon3x0_p0_iu_fe_pc_29_, u0_0_leon3x0_p0_iu_fe_pc_30_,
         u0_0_leon3x0_p0_iu_de_icc_0_, u0_0_leon3x0_p0_iu_de_icc_1_,
         u0_0_leon3x0_p0_iu_de_icc_2_, u0_0_leon3x0_p0_iu_de_icc_3_,
         u0_0_leon3x0_p0_iu_ex_jump_address_2_, u0_0_leon3x0_p0_iu_vp_ERROR_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__0_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__1_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__2_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__3_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__4_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__5_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__6_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__7_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__8_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__9_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__10_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__11_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__12_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__13_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__14_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__15_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__16_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__17_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__18_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__19_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__20_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__21_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__22_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__23_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__24_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__25_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__26_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__27_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__28_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__29_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__30_,
         u0_0_leon3x0_p0_iu_r_W__RESULT__31_, u0_0_leon3x0_p0_iu_r_W__S__Y__0_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__1_, u0_0_leon3x0_p0_iu_r_W__S__Y__2_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__3_, u0_0_leon3x0_p0_iu_r_W__S__Y__4_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__5_, u0_0_leon3x0_p0_iu_r_W__S__Y__6_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__7_, u0_0_leon3x0_p0_iu_r_W__S__Y__8_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__9_, u0_0_leon3x0_p0_iu_r_W__S__Y__10_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__11_, u0_0_leon3x0_p0_iu_r_W__S__Y__12_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__13_, u0_0_leon3x0_p0_iu_r_W__S__Y__14_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__15_, u0_0_leon3x0_p0_iu_r_W__S__Y__16_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__17_, u0_0_leon3x0_p0_iu_r_W__S__Y__18_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__19_, u0_0_leon3x0_p0_iu_r_W__S__Y__20_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__21_, u0_0_leon3x0_p0_iu_r_W__S__Y__22_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__23_, u0_0_leon3x0_p0_iu_r_W__S__Y__24_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__25_, u0_0_leon3x0_p0_iu_r_W__S__Y__26_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__27_, u0_0_leon3x0_p0_iu_r_W__S__Y__28_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__29_, u0_0_leon3x0_p0_iu_r_W__S__Y__30_,
         u0_0_leon3x0_p0_iu_r_W__S__Y__31_, u0_0_leon3x0_p0_iu_r_W__S__ET_,
         u0_0_leon3x0_p0_iu_r_W__S__PS_, u0_0_leon3x0_p0_iu_r_W__S__PIL__0_,
         u0_0_leon3x0_p0_iu_r_W__S__PIL__1_,
         u0_0_leon3x0_p0_iu_r_W__S__WIM__0_,
         u0_0_leon3x0_p0_iu_r_W__S__WIM__1_,
         u0_0_leon3x0_p0_iu_r_W__S__WIM__2_,
         u0_0_leon3x0_p0_iu_r_W__S__WIM__3_,
         u0_0_leon3x0_p0_iu_r_W__S__WIM__4_,
         u0_0_leon3x0_p0_iu_r_W__S__WIM__5_,
         u0_0_leon3x0_p0_iu_r_W__S__WIM__6_,
         u0_0_leon3x0_p0_iu_r_W__S__WIM__7_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__0_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__1_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__2_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__3_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__4_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__5_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__6_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__7_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__8_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__9_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__10_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__11_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__12_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__13_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__14_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__15_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__16_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__17_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__18_,
         u0_0_leon3x0_p0_iu_r_W__S__TBA__19_,
         u0_0_leon3x0_p0_iu_r_W__S__TT__4_, u0_0_leon3x0_p0_iu_r_W__S__TT__6_,
         u0_0_leon3x0_p0_iu_r_W__S__TT__7_, u0_0_leon3x0_p0_iu_r_W__S__ICC__0_,
         u0_0_leon3x0_p0_iu_r_W__S__ICC__1_,
         u0_0_leon3x0_p0_iu_r_W__S__ICC__2_,
         u0_0_leon3x0_p0_iu_r_W__S__ICC__3_,
         u0_0_leon3x0_p0_iu_r_W__S__CWP__0_,
         u0_0_leon3x0_p0_iu_r_W__S__CWP__1_,
         u0_0_leon3x0_p0_iu_r_W__S__CWP__2_, u0_0_leon3x0_p0_iu_r_X__NERROR_,
         u0_0_leon3x0_p0_iu_r_X__INTACK_, u0_0_leon3x0_p0_iu_r_X__NPC__0_,
         u0_0_leon3x0_p0_iu_r_X__NPC__1_, u0_0_leon3x0_p0_iu_r_X__NPC__2_,
         u0_0_leon3x0_p0_iu_r_X__LADDR__0_, u0_0_leon3x0_p0_iu_r_X__LADDR__1_,
         u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__0_,
         u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__1_,
         u0_0_leon3x0_p0_iu_r_X__DCI__SIGNED_, u0_0_leon3x0_p0_iu_r_X__MEXC_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__0_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__1_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__2_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__3_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__4_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__5_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__6_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__7_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__8_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__9_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__10_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__11_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__12_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__13_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__14_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__15_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__16_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__17_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__18_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__19_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__20_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__21_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__22_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__23_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__24_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__25_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__26_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__27_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__28_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__29_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__30_,
         u0_0_leon3x0_p0_iu_r_X__DATA__0__31_, u0_0_leon3x0_p0_iu_r_X__ICC__0_,
         u0_0_leon3x0_p0_iu_r_X__ICC__1_, u0_0_leon3x0_p0_iu_r_X__ICC__2_,
         u0_0_leon3x0_p0_iu_r_X__ICC__3_, u0_0_leon3x0_p0_iu_r_X__Y__8_,
         u0_0_leon3x0_p0_iu_r_X__Y__9_, u0_0_leon3x0_p0_iu_r_X__Y__10_,
         u0_0_leon3x0_p0_iu_r_X__Y__11_, u0_0_leon3x0_p0_iu_r_X__Y__12_,
         u0_0_leon3x0_p0_iu_r_X__Y__13_, u0_0_leon3x0_p0_iu_r_X__Y__14_,
         u0_0_leon3x0_p0_iu_r_X__Y__15_, u0_0_leon3x0_p0_iu_r_X__Y__16_,
         u0_0_leon3x0_p0_iu_r_X__Y__17_, u0_0_leon3x0_p0_iu_r_X__Y__18_,
         u0_0_leon3x0_p0_iu_r_X__Y__19_, u0_0_leon3x0_p0_iu_r_X__Y__20_,
         u0_0_leon3x0_p0_iu_r_X__Y__21_, u0_0_leon3x0_p0_iu_r_X__Y__22_,
         u0_0_leon3x0_p0_iu_r_X__Y__23_, u0_0_leon3x0_p0_iu_r_X__Y__24_,
         u0_0_leon3x0_p0_iu_r_X__Y__25_, u0_0_leon3x0_p0_iu_r_X__Y__26_,
         u0_0_leon3x0_p0_iu_r_X__Y__27_, u0_0_leon3x0_p0_iu_r_X__Y__28_,
         u0_0_leon3x0_p0_iu_r_X__Y__29_, u0_0_leon3x0_p0_iu_r_X__Y__30_,
         u0_0_leon3x0_p0_iu_r_X__Y__31_, u0_0_leon3x0_p0_iu_r_X__RESULT__0_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__1_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__2_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__3_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__4_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__5_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__6_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__7_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__8_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__9_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__10_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__11_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__12_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__13_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__14_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__15_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__16_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__17_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__18_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__19_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__20_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__21_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__22_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__23_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__24_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__25_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__26_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__27_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__28_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__29_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__30_,
         u0_0_leon3x0_p0_iu_r_X__RESULT__31_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RETT_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__LD_, u0_0_leon3x0_p0_iu_r_X__CTRL__WY_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__WREG_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__ANNUL_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__TRAP_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__TT__0_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__TT__1_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__TT__2_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__TT__3_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__TT__4_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__TT__5_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RD__0_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RD__1_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RD__2_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RD__3_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RD__4_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RD__5_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RD__6_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__RD__7_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__INST__19_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__INST__20_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__INST__25_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__INST__26_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__INST__27_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__INST__28_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__INST__29_,
         u0_0_leon3x0_p0_iu_r_X__CTRL__PC__2_, u0_0_leon3x0_p0_iu_r_M__CASA_,
         u0_0_leon3x0_p0_iu_r_M__MUL_, u0_0_leon3x0_p0_iu_r_M__DIVZ_,
         u0_0_leon3x0_p0_iu_r_M__IRQEN2_, u0_0_leon3x0_p0_iu_r_M__WCWP_,
         u0_0_leon3x0_p0_iu_r_M__NALIGN_, u0_0_leon3x0_p0_iu_r_M__CTRL__RETT_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__WICC_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__ANNUL_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__TRAP_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__TT__0_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__TT__1_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__TT__2_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__TT__3_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__TT__4_,
         u0_0_leon3x0_p0_iu_r_M__CTRL__TT__5_, u0_0_leon3x0_p0_iu_r_E__BP_,
         u0_0_leon3x0_p0_iu_r_E__MULSTEP_, u0_0_leon3x0_p0_iu_r_E__CWP__0_,
         u0_0_leon3x0_p0_iu_r_E__CWP__1_, u0_0_leon3x0_p0_iu_r_E__CWP__2_,
         u0_0_leon3x0_p0_iu_r_E__ET_, u0_0_leon3x0_p0_iu_r_E__JMPL_,
         u0_0_leon3x0_p0_iu_r_E__YMSB_, u0_0_leon3x0_p0_iu_r_E__SHLEFT_,
         u0_0_leon3x0_p0_iu_r_E__SARI_, u0_0_leon3x0_p0_iu_r_E__SHCNT__0_,
         u0_0_leon3x0_p0_iu_r_E__SHCNT__1_, u0_0_leon3x0_p0_iu_r_E__SHCNT__2_,
         u0_0_leon3x0_p0_iu_r_E__SHCNT__3_, u0_0_leon3x0_p0_iu_r_E__SHCNT__4_,
         u0_0_leon3x0_p0_iu_r_E__INVOP2_, u0_0_leon3x0_p0_iu_r_E__LDBP2_,
         u0_0_leon3x0_p0_iu_r_E__LDBP1_, u0_0_leon3x0_p0_iu_r_E__ALUCIN_,
         u0_0_leon3x0_p0_iu_r_E__ALUADD_, u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_,
         u0_0_leon3x0_p0_iu_r_E__ALUSEL__1_, u0_0_leon3x0_p0_iu_r_E__ALUOP__0_,
         u0_0_leon3x0_p0_iu_r_E__ALUOP__1_, u0_0_leon3x0_p0_iu_r_E__ALUOP__2_,
         u0_0_leon3x0_p0_iu_r_E__OP2__0_, u0_0_leon3x0_p0_iu_r_E__OP2__1_,
         u0_0_leon3x0_p0_iu_r_E__OP2__2_, u0_0_leon3x0_p0_iu_r_E__OP2__3_,
         u0_0_leon3x0_p0_iu_r_E__OP2__4_, u0_0_leon3x0_p0_iu_r_E__OP2__5_,
         u0_0_leon3x0_p0_iu_r_E__OP2__6_, u0_0_leon3x0_p0_iu_r_E__OP2__7_,
         u0_0_leon3x0_p0_iu_r_E__OP2__8_, u0_0_leon3x0_p0_iu_r_E__OP2__9_,
         u0_0_leon3x0_p0_iu_r_E__OP2__10_, u0_0_leon3x0_p0_iu_r_E__OP2__11_,
         u0_0_leon3x0_p0_iu_r_E__OP2__12_, u0_0_leon3x0_p0_iu_r_E__OP2__13_,
         u0_0_leon3x0_p0_iu_r_E__OP2__14_, u0_0_leon3x0_p0_iu_r_E__OP2__15_,
         u0_0_leon3x0_p0_iu_r_E__OP2__16_, u0_0_leon3x0_p0_iu_r_E__OP2__17_,
         u0_0_leon3x0_p0_iu_r_E__OP2__18_, u0_0_leon3x0_p0_iu_r_E__OP2__19_,
         u0_0_leon3x0_p0_iu_r_E__OP2__20_, u0_0_leon3x0_p0_iu_r_E__OP2__21_,
         u0_0_leon3x0_p0_iu_r_E__OP2__22_, u0_0_leon3x0_p0_iu_r_E__OP2__23_,
         u0_0_leon3x0_p0_iu_r_E__OP2__24_, u0_0_leon3x0_p0_iu_r_E__OP2__25_,
         u0_0_leon3x0_p0_iu_r_E__OP2__26_, u0_0_leon3x0_p0_iu_r_E__OP2__27_,
         u0_0_leon3x0_p0_iu_r_E__OP2__28_, u0_0_leon3x0_p0_iu_r_E__OP2__29_,
         u0_0_leon3x0_p0_iu_r_E__OP2__30_, u0_0_leon3x0_p0_iu_r_E__OP2__31_,
         u0_0_leon3x0_p0_iu_r_E__OP1__0_, u0_0_leon3x0_p0_iu_r_E__OP1__1_,
         u0_0_leon3x0_p0_iu_r_E__OP1__2_, u0_0_leon3x0_p0_iu_r_E__OP1__3_,
         u0_0_leon3x0_p0_iu_r_E__OP1__4_, u0_0_leon3x0_p0_iu_r_E__OP1__5_,
         u0_0_leon3x0_p0_iu_r_E__OP1__6_, u0_0_leon3x0_p0_iu_r_E__OP1__7_,
         u0_0_leon3x0_p0_iu_r_E__OP1__8_, u0_0_leon3x0_p0_iu_r_E__OP1__9_,
         u0_0_leon3x0_p0_iu_r_E__OP1__10_, u0_0_leon3x0_p0_iu_r_E__OP1__11_,
         u0_0_leon3x0_p0_iu_r_E__OP1__12_, u0_0_leon3x0_p0_iu_r_E__OP1__13_,
         u0_0_leon3x0_p0_iu_r_E__OP1__14_, u0_0_leon3x0_p0_iu_r_E__OP1__15_,
         u0_0_leon3x0_p0_iu_r_E__OP1__16_, u0_0_leon3x0_p0_iu_r_E__OP1__17_,
         u0_0_leon3x0_p0_iu_r_E__OP1__18_, u0_0_leon3x0_p0_iu_r_E__OP1__19_,
         u0_0_leon3x0_p0_iu_r_E__OP1__20_, u0_0_leon3x0_p0_iu_r_E__OP1__21_,
         u0_0_leon3x0_p0_iu_r_E__OP1__22_, u0_0_leon3x0_p0_iu_r_E__OP1__23_,
         u0_0_leon3x0_p0_iu_r_E__OP1__24_, u0_0_leon3x0_p0_iu_r_E__OP1__25_,
         u0_0_leon3x0_p0_iu_r_E__OP1__26_, u0_0_leon3x0_p0_iu_r_E__OP1__27_,
         u0_0_leon3x0_p0_iu_r_E__OP1__28_, u0_0_leon3x0_p0_iu_r_E__OP1__29_,
         u0_0_leon3x0_p0_iu_r_E__OP1__30_, u0_0_leon3x0_p0_iu_r_E__OP1__31_,
         u0_0_leon3x0_p0_iu_r_E__CTRL__RETT_,
         u0_0_leon3x0_p0_iu_r_E__CTRL__WICC_,
         u0_0_leon3x0_p0_iu_r_E__CTRL__WREG_,
         u0_0_leon3x0_p0_iu_r_E__CTRL__ANNUL_, u0_0_leon3x0_p0_iu_r_A__NOBP_,
         u0_0_leon3x0_p0_iu_r_A__BP_, u0_0_leon3x0_p0_iu_r_A__DIVSTART_,
         u0_0_leon3x0_p0_iu_r_A__MULSTART_, u0_0_leon3x0_p0_iu_r_A__JMPL_,
         u0_0_leon3x0_p0_iu_r_A__TICC_, u0_0_leon3x0_p0_iu_r_A__WUNF_,
         u0_0_leon3x0_p0_iu_r_A__WOVF_, u0_0_leon3x0_p0_iu_r_A__IMM__0_,
         u0_0_leon3x0_p0_iu_r_A__IMM__1_, u0_0_leon3x0_p0_iu_r_A__IMM__2_,
         u0_0_leon3x0_p0_iu_r_A__IMM__3_, u0_0_leon3x0_p0_iu_r_A__IMM__4_,
         u0_0_leon3x0_p0_iu_r_A__IMM__5_, u0_0_leon3x0_p0_iu_r_A__IMM__6_,
         u0_0_leon3x0_p0_iu_r_A__IMM__7_, u0_0_leon3x0_p0_iu_r_A__IMM__8_,
         u0_0_leon3x0_p0_iu_r_A__IMM__9_, u0_0_leon3x0_p0_iu_r_A__IMM__10_,
         u0_0_leon3x0_p0_iu_r_A__IMM__11_, u0_0_leon3x0_p0_iu_r_A__IMM__12_,
         u0_0_leon3x0_p0_iu_r_A__IMM__13_, u0_0_leon3x0_p0_iu_r_A__IMM__14_,
         u0_0_leon3x0_p0_iu_r_A__IMM__15_, u0_0_leon3x0_p0_iu_r_A__IMM__16_,
         u0_0_leon3x0_p0_iu_r_A__IMM__17_, u0_0_leon3x0_p0_iu_r_A__IMM__18_,
         u0_0_leon3x0_p0_iu_r_A__IMM__19_, u0_0_leon3x0_p0_iu_r_A__IMM__20_,
         u0_0_leon3x0_p0_iu_r_A__IMM__21_, u0_0_leon3x0_p0_iu_r_A__IMM__22_,
         u0_0_leon3x0_p0_iu_r_A__IMM__23_, u0_0_leon3x0_p0_iu_r_A__IMM__24_,
         u0_0_leon3x0_p0_iu_r_A__IMM__25_, u0_0_leon3x0_p0_iu_r_A__IMM__26_,
         u0_0_leon3x0_p0_iu_r_A__IMM__27_, u0_0_leon3x0_p0_iu_r_A__IMM__28_,
         u0_0_leon3x0_p0_iu_r_A__IMM__29_, u0_0_leon3x0_p0_iu_r_A__IMM__30_,
         u0_0_leon3x0_p0_iu_r_A__IMM__31_, u0_0_leon3x0_p0_iu_r_A__RSEL2__0_,
         u0_0_leon3x0_p0_iu_r_A__RSEL2__1_, u0_0_leon3x0_p0_iu_r_A__RSEL2__2_,
         u0_0_leon3x0_p0_iu_r_A__RSEL1__0_, u0_0_leon3x0_p0_iu_r_A__RSEL1__1_,
         u0_0_leon3x0_p0_iu_r_A__RSEL1__2_, u0_0_leon3x0_p0_iu_r_A__RFA2__0_,
         u0_0_leon3x0_p0_iu_r_A__RFA2__1_, u0_0_leon3x0_p0_iu_r_A__RFA2__2_,
         u0_0_leon3x0_p0_iu_r_A__RFA2__3_, u0_0_leon3x0_p0_iu_r_A__RFA2__4_,
         u0_0_leon3x0_p0_iu_r_A__RFA2__5_, u0_0_leon3x0_p0_iu_r_A__RFA2__6_,
         u0_0_leon3x0_p0_iu_r_A__RFA2__7_, u0_0_leon3x0_p0_iu_r_A__RFA1__0_,
         u0_0_leon3x0_p0_iu_r_A__RFA1__1_, u0_0_leon3x0_p0_iu_r_A__RFA1__2_,
         u0_0_leon3x0_p0_iu_r_A__RFA1__3_, u0_0_leon3x0_p0_iu_r_A__RFA1__4_,
         u0_0_leon3x0_p0_iu_r_A__RFA1__5_, u0_0_leon3x0_p0_iu_r_A__RFA1__6_,
         u0_0_leon3x0_p0_iu_r_A__RFA1__7_, u0_0_leon3x0_p0_iu_r_A__CTRL__RETT_,
         u0_0_leon3x0_p0_iu_r_A__CTRL__WICC_,
         u0_0_leon3x0_p0_iu_r_A__CTRL__WREG_,
         u0_0_leon3x0_p0_iu_r_A__CTRL__ANNUL_,
         u0_0_leon3x0_p0_iu_r_A__CTRL__TT__0_, u0_0_leon3x0_p0_iu_r_D__DIVRDY_,
         u0_0_leon3x0_p0_iu_r_D__INULL_, u0_0_leon3x0_p0_iu_r_D__ANNUL_,
         u0_0_leon3x0_p0_iu_r_D__PV_, u0_0_leon3x0_p0_iu_v_X__DCI__LOCK_,
         u0_0_leon3x0_p0_iu_v_X__DCI__SIGNED_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PV_, u0_0_leon3x0_p0_iu_v_X__CTRL__LD_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__WY_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__WREG_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__RD__0_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__RD__1_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__RD__2_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__RD__3_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__RD__4_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__RD__5_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__RD__6_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__RD__7_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__0_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__1_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__19_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__20_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__21_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__25_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__26_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__27_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__28_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__29_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__30_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__INST__31_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__2_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__3_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__4_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__5_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__6_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__7_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__8_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__9_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__10_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__11_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__12_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__13_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__14_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__15_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__16_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__17_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__18_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__19_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__20_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__21_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__22_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__23_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__24_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__25_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__26_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__27_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__28_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__29_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__30_,
         u0_0_leon3x0_p0_iu_v_X__CTRL__PC__31_, u0_0_leon3x0_p0_iu_v_M__MUL_,
         u0_0_leon3x0_p0_iu_v_M__IRQEN2_, u0_0_leon3x0_p0_iu_v_M__WERR_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PV_, u0_0_leon3x0_p0_iu_v_M__CTRL__LD_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__WY_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__TRAP_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__TT__0_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__TT__1_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__TT__2_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__TT__3_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__TT__4_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__TT__5_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__RD__0_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__RD__1_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__RD__2_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__RD__3_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__RD__4_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__RD__5_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__RD__6_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__RD__7_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__0_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__1_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__5_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__6_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__7_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__8_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__9_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__14_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__17_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__18_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__23_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__25_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__26_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__28_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__29_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__30_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__INST__31_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__2_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__3_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__4_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__5_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__6_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__7_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__8_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__9_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__10_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__11_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__12_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__13_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__14_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__15_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__16_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__17_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__18_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__19_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__20_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__21_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__22_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__23_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__24_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__25_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__26_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__27_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__28_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__29_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__30_,
         u0_0_leon3x0_p0_iu_v_M__CTRL__PC__31_, u0_0_leon3x0_p0_iu_v_E__RFE2_,
         u0_0_leon3x0_p0_iu_v_E__RFE1_, u0_0_leon3x0_p0_iu_v_E__CWP__0_,
         u0_0_leon3x0_p0_iu_v_E__CWP__1_, u0_0_leon3x0_p0_iu_v_E__CWP__2_,
         u0_0_leon3x0_p0_iu_v_E__ET_, u0_0_leon3x0_p0_iu_v_E__SU_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PV_, u0_0_leon3x0_p0_iu_v_E__CTRL__LD_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__WY_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__RD__0_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__RD__1_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__RD__2_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__RD__3_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__RD__4_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__RD__5_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__RD__6_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__RD__7_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__0_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__1_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__5_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__6_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__7_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__8_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__9_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__10_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__11_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__13_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__14_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__17_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__18_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__25_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__26_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__27_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__28_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__29_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__30_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__2_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__3_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__4_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__5_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__6_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__7_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__8_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__9_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__10_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__11_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__12_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__13_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__14_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__15_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__16_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__17_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__18_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__19_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__20_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__21_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__22_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__23_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__24_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__25_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__26_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__27_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__28_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__29_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__30_,
         u0_0_leon3x0_p0_iu_v_E__CTRL__PC__31_,
         u0_0_leon3x0_p0_iu_v_A__CWP__0_, u0_0_leon3x0_p0_iu_v_A__CWP__1_,
         u0_0_leon3x0_p0_iu_v_A__CWP__2_, u0_0_leon3x0_p0_iu_v_A__CTRL__TRAP_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__0_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__5_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__6_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__7_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__8_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__9_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__10_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__11_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__12_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__14_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__15_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__16_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__21_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__22_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__27_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__28_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__30_,
         u0_0_leon3x0_p0_iu_v_A__CTRL__INST__31_,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N59,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N57,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N54,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N53,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N52,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N51,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N50,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N49,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N48,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N47,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N46,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N42,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N29,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N28,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N27,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N26,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N25,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N21,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N20,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N18,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N16,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N14,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N13,
         u0_0_leon3x0_p0_mul0_m3232_dwm_N12, u0_0_leon3x0_p0_mul0_m3232_dwm_N8,
         u0_0_leon3x0_p0_div0_vaddsub, u0_0_leon3x0_p0_div0_addout_0_,
         u0_0_leon3x0_p0_div0_addout_1_, u0_0_leon3x0_p0_div0_addout_2_,
         u0_0_leon3x0_p0_div0_addout_3_, u0_0_leon3x0_p0_div0_addout_4_,
         u0_0_leon3x0_p0_div0_addout_5_, u0_0_leon3x0_p0_div0_addout_6_,
         u0_0_leon3x0_p0_div0_addout_7_, u0_0_leon3x0_p0_div0_addout_8_,
         u0_0_leon3x0_p0_div0_addout_9_, u0_0_leon3x0_p0_div0_addout_10_,
         u0_0_leon3x0_p0_div0_addout_11_, u0_0_leon3x0_p0_div0_addout_12_,
         u0_0_leon3x0_p0_div0_addout_13_, u0_0_leon3x0_p0_div0_addout_14_,
         u0_0_leon3x0_p0_div0_addout_15_, u0_0_leon3x0_p0_div0_addout_16_,
         u0_0_leon3x0_p0_div0_addout_17_, u0_0_leon3x0_p0_div0_addout_18_,
         u0_0_leon3x0_p0_div0_addout_19_, u0_0_leon3x0_p0_div0_addout_20_,
         u0_0_leon3x0_p0_div0_addout_21_, u0_0_leon3x0_p0_div0_addout_22_,
         u0_0_leon3x0_p0_div0_addout_23_, u0_0_leon3x0_p0_div0_addout_24_,
         u0_0_leon3x0_p0_div0_addout_25_, u0_0_leon3x0_p0_div0_addout_26_,
         u0_0_leon3x0_p0_div0_addout_27_, u0_0_leon3x0_p0_div0_addout_28_,
         u0_0_leon3x0_p0_div0_addout_29_, u0_0_leon3x0_p0_div0_addout_30_,
         u0_0_leon3x0_p0_div0_addout_31_, u0_0_leon3x0_p0_div0_addout_32_,
         u0_0_leon3x0_p0_div0_r_CNT__0_, u0_0_leon3x0_p0_div0_r_CNT__1_,
         u0_0_leon3x0_p0_div0_r_CNT__2_, u0_0_leon3x0_p0_div0_r_CNT__3_,
         u0_0_leon3x0_p0_div0_r_CNT__4_, u0_0_leon3x0_p0_div0_r_NEG_,
         u0_0_leon3x0_p0_div0_r_QMSB_, u0_0_leon3x0_p0_div0_r_ZERO2_,
         u0_0_leon3x0_p0_div0_r_X__0_, u0_0_leon3x0_p0_div0_r_X__1_,
         u0_0_leon3x0_p0_div0_r_X__2_, u0_0_leon3x0_p0_div0_r_X__3_,
         u0_0_leon3x0_p0_div0_r_X__4_, u0_0_leon3x0_p0_div0_r_X__5_,
         u0_0_leon3x0_p0_div0_r_X__6_, u0_0_leon3x0_p0_div0_r_X__7_,
         u0_0_leon3x0_p0_div0_r_X__8_, u0_0_leon3x0_p0_div0_r_X__9_,
         u0_0_leon3x0_p0_div0_r_X__10_, u0_0_leon3x0_p0_div0_r_X__11_,
         u0_0_leon3x0_p0_div0_r_X__12_, u0_0_leon3x0_p0_div0_r_X__13_,
         u0_0_leon3x0_p0_div0_r_X__14_, u0_0_leon3x0_p0_div0_r_X__15_,
         u0_0_leon3x0_p0_div0_r_X__16_, u0_0_leon3x0_p0_div0_r_X__17_,
         u0_0_leon3x0_p0_div0_r_X__18_, u0_0_leon3x0_p0_div0_r_X__19_,
         u0_0_leon3x0_p0_div0_r_X__20_, u0_0_leon3x0_p0_div0_r_X__21_,
         u0_0_leon3x0_p0_div0_r_X__22_, u0_0_leon3x0_p0_div0_r_X__23_,
         u0_0_leon3x0_p0_div0_r_X__24_, u0_0_leon3x0_p0_div0_r_X__25_,
         u0_0_leon3x0_p0_div0_r_X__26_, u0_0_leon3x0_p0_div0_r_X__27_,
         u0_0_leon3x0_p0_div0_r_X__28_, u0_0_leon3x0_p0_div0_r_X__29_,
         u0_0_leon3x0_p0_div0_r_X__30_, u0_0_leon3x0_p0_div0_r_X__31_,
         u0_0_leon3x0_p0_div0_v_ZERO2_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__0_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__1_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__2_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__3_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__4_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__5_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__6_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_HIT_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__0_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__1_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__2_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__3_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__4_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__5_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__6_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__7_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__2_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__4_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__5_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__6_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__7_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__8_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__9_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__10_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__11_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__12_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__13_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__14_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__15_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__16_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__17_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__18_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__19_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__20_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__21_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__22_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__23_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__24_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__25_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__26_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__27_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__28_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__29_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__30_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__31_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_UNDERRUN_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_OVERRUN_,
         u0_0_leon3x0_p0_c0mmu_icache0_r_BURST_,
         u0_0_leon3x0_p0_c0mmu_icache0_v_VADDRESS__3_,
         u0_0_leon3x0_p0_c0mmu_icache0_v_WADDRESS__2_,
         u0_0_leon3x0_p0_c0mmu_icache0_v_WADDRESS__4_,
         u0_0_leon3x0_p0_c0mmu_icache0_v_HOLDN_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_NOFLUSH_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_CCTRLWR_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_ASI__0_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__0_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__1_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__2_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__3_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__4_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__5_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__6_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__7_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__8_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__9_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__10_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__11_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__12_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__13_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__14_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__15_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__16_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__17_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__18_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__19_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__20_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__21_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__22_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__23_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__24_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__25_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__26_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__27_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__28_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__29_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__30_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__31_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_BMEXC_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_MEXC_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_FLUSH2_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_VALID_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__0_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__1_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__2_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__3_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__4_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__5_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_STPEND_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_NOMDS_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_RBURST_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__0_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__1_,
         u0_0_leon3x0_p0_c0mmu_dcache0_r_READ_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_CCTRL__DCS__0_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__2_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__3_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__4_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_FLUSH_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_FADDR__6_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_XADDRESS__2_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_HOLDN_,
         u0_0_leon3x0_p0_c0mmu_dcache0_v_REQ_,
         u0_0_leon3x0_p0_c0mmu_a0_r_NBO__0_,
         u0_0_leon3x0_p0_c0mmu_a0_r_NBO__1_, u0_0_leon3x0_p0_c0mmu_a0_r_NBA_,
         u0_0_leon3x0_p0_c0mmu_a0_r_HCACHE_,
         u0_0_leon3x0_p0_c0mmu_a0_r_HLOCKEN_,
         u0_0_leon3x0_p0_c0mmu_a0_r_BO__0_, u0_0_leon3x0_p0_c0mmu_a0_r_BG_,
         u0_0_leon3x0_p0_c0mmu_a0_v_BO__1_, sr1_sdi_HWRITE_, sr1_sdi_HSIZE__0_,
         sr1_sdi_HSIZE__1_, sr1_r_HBURST__0_, sr1_r_SRHSEL_, sr1_r_MCFG2__RMW_,
         sr1_r_MCFG2__RAMBANKSZ__0_, sr1_r_MCFG2__RAMBANKSZ__1_,
         sr1_r_MCFG2__RAMBANKSZ__3_, sr1_r_MCFG2__RAMWIDTH__0_,
         sr1_r_MCFG2__RAMWIDTH__1_, sr1_r_MCFG2__RAMWWS__0_,
         sr1_r_MCFG2__RAMWWS__1_, sr1_r_MCFG2__RAMRWS__0_,
         sr1_r_MCFG2__RAMRWS__1_, sr1_r_MCFG1__IOWIDTH__0_,
         sr1_r_MCFG1__IOWIDTH__1_, sr1_r_MCFG1__BRDYEN_, sr1_r_MCFG1__BEXCEN_,
         sr1_r_MCFG1__IOWS__0_, sr1_r_MCFG1__IOWS__1_, sr1_r_MCFG1__IOWS__2_,
         sr1_r_MCFG1__IOWS__3_, sr1_r_MCFG1__IOEN_, sr1_r_MCFG1__ROMWRITE_,
         sr1_r_MCFG1__ROMWIDTH__0_, sr1_r_MCFG1__ROMWIDTH__1_,
         sr1_r_MCFG1__ROMWWS__0_, sr1_r_MCFG1__ROMWWS__1_,
         sr1_r_MCFG1__ROMWWS__2_, sr1_r_MCFG1__ROMWWS__3_,
         sr1_r_MCFG1__ROMRWS__0_, sr1_r_MCFG1__ROMRWS__1_,
         sr1_r_MCFG1__ROMRWS__2_, sr1_r_MCFG1__ROMRWS__3_, sr1_r_AREA__0_,
         sr1_r_BSTATE__0_, sr1_r_BSTATE__1_, sr1_r_IOSN__1_, sr1_r_BUSW__0_,
         sr1_r_BUSW__1_, sr1_r_WS__0_, sr1_r_WS__2_, sr1_r_WS__3_,
         sr1_r_READY_, sr1_v_ADDRESS__0_, sr1_v_ADDRESS__1_, apb0_N1148,
         apb0_r_CFGSEL_, apb0_r_STATE__0_, apb0_r_PSEL_, uart1_scaler_1_,
         uart1_scaler_2_, uart1_scaler_3_, uart1_scaler_4_, uart1_scaler_9_,
         uart1_scaler_10_, uart1_scaler_11_, uart1_r_TCNT__0_,
         uart1_r_TCNT__1_, uart1_r_TCNT__2_, uart1_r_TCNT__3_,
         uart1_r_TCNT__4_, uart1_r_TCNT__5_, uart1_r_RCNT__0_,
         uart1_r_RCNT__1_, uart1_r_RCNT__2_, uart1_r_RCNT__3_,
         uart1_r_RCNT__4_, uart1_r_RCNT__5_, uart1_r_TWADDR__0_,
         uart1_r_TWADDR__1_, uart1_r_TWADDR__2_, uart1_r_TWADDR__4_,
         uart1_r_TRADDR__0_, uart1_r_TRADDR__1_, uart1_r_TRADDR__2_,
         uart1_r_TRADDR__3_, uart1_r_TRADDR__4_, uart1_r_RWADDR__0_,
         uart1_r_RWADDR__1_, uart1_r_RWADDR__2_, uart1_r_RWADDR__4_,
         uart1_r_IRQCNT__0_, uart1_r_IRQCNT__1_, uart1_r_IRQCNT__2_,
         uart1_r_IRQCNT__3_, uart1_r_IRQCNT__4_, uart1_r_IRQCNT__5_,
         uart1_r_TFIFOIRQEN_, uart1_r_RFIFOIRQEN_, uart1_r_RXF__1_,
         uart1_r_RXF__2_, uart1_r_RXF__3_, uart1_r_RXF__4_, uart1_r_BRATE__0_,
         uart1_r_BRATE__1_, uart1_r_BRATE__2_, uart1_r_BRATE__3_,
         uart1_r_BRATE__4_, uart1_r_BRATE__5_, uart1_r_BRATE__6_,
         uart1_r_BRATE__7_, uart1_r_BRATE__8_, uart1_r_BRATE__9_,
         uart1_r_BRATE__10_, uart1_r_BRATE__11_, uart1_r_TICK_,
         uart1_r_RXTICK_, uart1_r_DPAR_, uart1_r_RXDB__1_, uart1_r_RXCLK__0_,
         uart1_r_RXCLK__1_, uart1_r_RXSTATE__0_, uart1_r_RXSTATE__1_,
         uart1_r_TXCLK__0_, uart1_r_TXCLK__1_, uart1_r_TPAR_, uart1_r_IRQPEND_,
         uart1_r_THOLD__31__0_, uart1_r_THOLD__31__1_, uart1_r_THOLD__31__2_,
         uart1_r_THOLD__31__3_, uart1_r_THOLD__31__4_, uart1_r_THOLD__31__5_,
         uart1_r_THOLD__31__6_, uart1_r_THOLD__31__7_, uart1_r_THOLD__30__0_,
         uart1_r_THOLD__30__1_, uart1_r_THOLD__30__2_, uart1_r_THOLD__30__3_,
         uart1_r_THOLD__30__4_, uart1_r_THOLD__30__5_, uart1_r_THOLD__30__6_,
         uart1_r_THOLD__30__7_, uart1_r_THOLD__29__0_, uart1_r_THOLD__29__1_,
         uart1_r_THOLD__29__2_, uart1_r_THOLD__29__3_, uart1_r_THOLD__29__4_,
         uart1_r_THOLD__29__5_, uart1_r_THOLD__29__6_, uart1_r_THOLD__29__7_,
         uart1_r_THOLD__28__0_, uart1_r_THOLD__28__1_, uart1_r_THOLD__28__2_,
         uart1_r_THOLD__28__3_, uart1_r_THOLD__28__4_, uart1_r_THOLD__28__5_,
         uart1_r_THOLD__28__6_, uart1_r_THOLD__28__7_, uart1_r_THOLD__27__0_,
         uart1_r_THOLD__27__1_, uart1_r_THOLD__27__2_, uart1_r_THOLD__27__3_,
         uart1_r_THOLD__27__4_, uart1_r_THOLD__27__5_, uart1_r_THOLD__27__6_,
         uart1_r_THOLD__27__7_, uart1_r_THOLD__26__0_, uart1_r_THOLD__26__1_,
         uart1_r_THOLD__26__2_, uart1_r_THOLD__26__3_, uart1_r_THOLD__26__4_,
         uart1_r_THOLD__26__5_, uart1_r_THOLD__26__6_, uart1_r_THOLD__26__7_,
         uart1_r_THOLD__25__0_, uart1_r_THOLD__25__1_, uart1_r_THOLD__25__2_,
         uart1_r_THOLD__25__3_, uart1_r_THOLD__25__4_, uart1_r_THOLD__25__5_,
         uart1_r_THOLD__25__6_, uart1_r_THOLD__25__7_, uart1_r_THOLD__24__0_,
         uart1_r_THOLD__24__1_, uart1_r_THOLD__24__2_, uart1_r_THOLD__24__3_,
         uart1_r_THOLD__24__4_, uart1_r_THOLD__24__5_, uart1_r_THOLD__24__6_,
         uart1_r_THOLD__24__7_, uart1_r_THOLD__23__0_, uart1_r_THOLD__23__1_,
         uart1_r_THOLD__23__2_, uart1_r_THOLD__23__3_, uart1_r_THOLD__23__4_,
         uart1_r_THOLD__23__5_, uart1_r_THOLD__23__6_, uart1_r_THOLD__23__7_,
         uart1_r_THOLD__22__0_, uart1_r_THOLD__22__1_, uart1_r_THOLD__22__2_,
         uart1_r_THOLD__22__3_, uart1_r_THOLD__22__4_, uart1_r_THOLD__22__5_,
         uart1_r_THOLD__22__6_, uart1_r_THOLD__22__7_, uart1_r_THOLD__21__0_,
         uart1_r_THOLD__21__1_, uart1_r_THOLD__21__2_, uart1_r_THOLD__21__3_,
         uart1_r_THOLD__21__4_, uart1_r_THOLD__21__5_, uart1_r_THOLD__21__6_,
         uart1_r_THOLD__21__7_, uart1_r_THOLD__20__0_, uart1_r_THOLD__20__1_,
         uart1_r_THOLD__20__2_, uart1_r_THOLD__20__3_, uart1_r_THOLD__20__4_,
         uart1_r_THOLD__20__5_, uart1_r_THOLD__20__6_, uart1_r_THOLD__20__7_,
         uart1_r_THOLD__19__0_, uart1_r_THOLD__19__1_, uart1_r_THOLD__19__2_,
         uart1_r_THOLD__19__3_, uart1_r_THOLD__19__4_, uart1_r_THOLD__19__5_,
         uart1_r_THOLD__19__6_, uart1_r_THOLD__19__7_, uart1_r_THOLD__18__0_,
         uart1_r_THOLD__18__1_, uart1_r_THOLD__18__2_, uart1_r_THOLD__18__3_,
         uart1_r_THOLD__18__4_, uart1_r_THOLD__18__5_, uart1_r_THOLD__18__6_,
         uart1_r_THOLD__18__7_, uart1_r_THOLD__17__0_, uart1_r_THOLD__17__1_,
         uart1_r_THOLD__17__2_, uart1_r_THOLD__17__3_, uart1_r_THOLD__17__4_,
         uart1_r_THOLD__17__5_, uart1_r_THOLD__17__6_, uart1_r_THOLD__17__7_,
         uart1_r_THOLD__16__0_, uart1_r_THOLD__16__1_, uart1_r_THOLD__16__2_,
         uart1_r_THOLD__16__3_, uart1_r_THOLD__16__4_, uart1_r_THOLD__16__5_,
         uart1_r_THOLD__16__6_, uart1_r_THOLD__16__7_, uart1_r_THOLD__15__0_,
         uart1_r_THOLD__15__1_, uart1_r_THOLD__15__2_, uart1_r_THOLD__15__3_,
         uart1_r_THOLD__15__4_, uart1_r_THOLD__15__5_, uart1_r_THOLD__15__6_,
         uart1_r_THOLD__15__7_, uart1_r_THOLD__14__0_, uart1_r_THOLD__14__1_,
         uart1_r_THOLD__14__2_, uart1_r_THOLD__14__3_, uart1_r_THOLD__14__4_,
         uart1_r_THOLD__14__5_, uart1_r_THOLD__14__6_, uart1_r_THOLD__14__7_,
         uart1_r_THOLD__13__0_, uart1_r_THOLD__13__1_, uart1_r_THOLD__13__2_,
         uart1_r_THOLD__13__3_, uart1_r_THOLD__13__4_, uart1_r_THOLD__13__5_,
         uart1_r_THOLD__13__6_, uart1_r_THOLD__13__7_, uart1_r_THOLD__12__0_,
         uart1_r_THOLD__12__1_, uart1_r_THOLD__12__2_, uart1_r_THOLD__12__3_,
         uart1_r_THOLD__12__4_, uart1_r_THOLD__12__5_, uart1_r_THOLD__12__6_,
         uart1_r_THOLD__12__7_, uart1_r_THOLD__11__0_, uart1_r_THOLD__11__1_,
         uart1_r_THOLD__11__2_, uart1_r_THOLD__11__3_, uart1_r_THOLD__11__4_,
         uart1_r_THOLD__11__5_, uart1_r_THOLD__11__6_, uart1_r_THOLD__11__7_,
         uart1_r_THOLD__10__0_, uart1_r_THOLD__10__1_, uart1_r_THOLD__10__2_,
         uart1_r_THOLD__10__3_, uart1_r_THOLD__10__4_, uart1_r_THOLD__10__5_,
         uart1_r_THOLD__10__6_, uart1_r_THOLD__10__7_, uart1_r_THOLD__9__0_,
         uart1_r_THOLD__9__1_, uart1_r_THOLD__9__2_, uart1_r_THOLD__9__3_,
         uart1_r_THOLD__9__4_, uart1_r_THOLD__9__5_, uart1_r_THOLD__9__6_,
         uart1_r_THOLD__9__7_, uart1_r_THOLD__8__0_, uart1_r_THOLD__8__1_,
         uart1_r_THOLD__8__2_, uart1_r_THOLD__8__3_, uart1_r_THOLD__8__4_,
         uart1_r_THOLD__8__5_, uart1_r_THOLD__8__6_, uart1_r_THOLD__8__7_,
         uart1_r_THOLD__7__0_, uart1_r_THOLD__7__1_, uart1_r_THOLD__7__2_,
         uart1_r_THOLD__7__3_, uart1_r_THOLD__7__4_, uart1_r_THOLD__7__5_,
         uart1_r_THOLD__7__6_, uart1_r_THOLD__7__7_, uart1_r_THOLD__6__0_,
         uart1_r_THOLD__6__1_, uart1_r_THOLD__6__2_, uart1_r_THOLD__6__3_,
         uart1_r_THOLD__6__4_, uart1_r_THOLD__6__5_, uart1_r_THOLD__6__6_,
         uart1_r_THOLD__6__7_, uart1_r_THOLD__5__0_, uart1_r_THOLD__5__1_,
         uart1_r_THOLD__5__2_, uart1_r_THOLD__5__3_, uart1_r_THOLD__5__4_,
         uart1_r_THOLD__5__5_, uart1_r_THOLD__5__6_, uart1_r_THOLD__5__7_,
         uart1_r_THOLD__4__0_, uart1_r_THOLD__4__1_, uart1_r_THOLD__4__2_,
         uart1_r_THOLD__4__3_, uart1_r_THOLD__4__4_, uart1_r_THOLD__4__5_,
         uart1_r_THOLD__4__6_, uart1_r_THOLD__4__7_, uart1_r_THOLD__3__0_,
         uart1_r_THOLD__3__1_, uart1_r_THOLD__3__2_, uart1_r_THOLD__3__3_,
         uart1_r_THOLD__3__4_, uart1_r_THOLD__3__5_, uart1_r_THOLD__3__6_,
         uart1_r_THOLD__3__7_, uart1_r_THOLD__2__0_, uart1_r_THOLD__2__1_,
         uart1_r_THOLD__2__2_, uart1_r_THOLD__2__3_, uart1_r_THOLD__2__4_,
         uart1_r_THOLD__2__5_, uart1_r_THOLD__2__6_, uart1_r_THOLD__2__7_,
         uart1_r_THOLD__1__0_, uart1_r_THOLD__1__1_, uart1_r_THOLD__1__2_,
         uart1_r_THOLD__1__3_, uart1_r_THOLD__1__4_, uart1_r_THOLD__1__5_,
         uart1_r_THOLD__1__6_, uart1_r_THOLD__1__7_, uart1_r_THOLD__0__0_,
         uart1_r_THOLD__0__1_, uart1_r_THOLD__0__2_, uart1_r_THOLD__0__3_,
         uart1_r_THOLD__0__4_, uart1_r_THOLD__0__5_, uart1_r_THOLD__0__6_,
         uart1_r_THOLD__0__7_, uart1_r_TSHIFT__0_, uart1_r_TSHIFT__2_,
         uart1_r_TSHIFT__3_, uart1_r_TSHIFT__4_, uart1_r_TSHIFT__5_,
         uart1_r_TSHIFT__6_, uart1_r_TSHIFT__7_, uart1_r_TSHIFT__8_,
         uart1_r_TSHIFT__9_, uart1_r_RSHIFT__0_, uart1_r_RSHIFT__1_,
         uart1_r_RSHIFT__2_, uart1_r_RSHIFT__3_, uart1_r_RSHIFT__4_,
         uart1_r_RSHIFT__5_, uart1_r_RSHIFT__6_, uart1_r_RSHIFT__7_,
         uart1_r_RHOLD__31__0_, uart1_r_RHOLD__31__1_, uart1_r_RHOLD__31__2_,
         uart1_r_RHOLD__31__3_, uart1_r_RHOLD__31__4_, uart1_r_RHOLD__31__5_,
         uart1_r_RHOLD__31__6_, uart1_r_RHOLD__31__7_, uart1_r_RHOLD__30__0_,
         uart1_r_RHOLD__30__1_, uart1_r_RHOLD__30__2_, uart1_r_RHOLD__30__3_,
         uart1_r_RHOLD__30__4_, uart1_r_RHOLD__30__5_, uart1_r_RHOLD__30__6_,
         uart1_r_RHOLD__30__7_, uart1_r_RHOLD__29__0_, uart1_r_RHOLD__29__1_,
         uart1_r_RHOLD__29__2_, uart1_r_RHOLD__29__3_, uart1_r_RHOLD__29__4_,
         uart1_r_RHOLD__29__5_, uart1_r_RHOLD__29__6_, uart1_r_RHOLD__29__7_,
         uart1_r_RHOLD__28__0_, uart1_r_RHOLD__28__1_, uart1_r_RHOLD__28__2_,
         uart1_r_RHOLD__28__3_, uart1_r_RHOLD__28__4_, uart1_r_RHOLD__28__5_,
         uart1_r_RHOLD__28__6_, uart1_r_RHOLD__28__7_, uart1_r_RHOLD__27__0_,
         uart1_r_RHOLD__27__1_, uart1_r_RHOLD__27__2_, uart1_r_RHOLD__27__3_,
         uart1_r_RHOLD__27__4_, uart1_r_RHOLD__27__5_, uart1_r_RHOLD__27__6_,
         uart1_r_RHOLD__27__7_, uart1_r_RHOLD__26__0_, uart1_r_RHOLD__26__1_,
         uart1_r_RHOLD__26__2_, uart1_r_RHOLD__26__3_, uart1_r_RHOLD__26__4_,
         uart1_r_RHOLD__26__5_, uart1_r_RHOLD__26__6_, uart1_r_RHOLD__26__7_,
         uart1_r_RHOLD__25__0_, uart1_r_RHOLD__25__1_, uart1_r_RHOLD__25__2_,
         uart1_r_RHOLD__25__3_, uart1_r_RHOLD__25__4_, uart1_r_RHOLD__25__5_,
         uart1_r_RHOLD__25__6_, uart1_r_RHOLD__25__7_, uart1_r_RHOLD__24__0_,
         uart1_r_RHOLD__24__1_, uart1_r_RHOLD__24__2_, uart1_r_RHOLD__24__3_,
         uart1_r_RHOLD__24__4_, uart1_r_RHOLD__24__5_, uart1_r_RHOLD__24__6_,
         uart1_r_RHOLD__24__7_, uart1_r_RHOLD__23__0_, uart1_r_RHOLD__23__1_,
         uart1_r_RHOLD__23__2_, uart1_r_RHOLD__23__3_, uart1_r_RHOLD__23__4_,
         uart1_r_RHOLD__23__5_, uart1_r_RHOLD__23__6_, uart1_r_RHOLD__23__7_,
         uart1_r_RHOLD__22__0_, uart1_r_RHOLD__22__1_, uart1_r_RHOLD__22__2_,
         uart1_r_RHOLD__22__3_, uart1_r_RHOLD__22__4_, uart1_r_RHOLD__22__5_,
         uart1_r_RHOLD__22__6_, uart1_r_RHOLD__22__7_, uart1_r_RHOLD__21__0_,
         uart1_r_RHOLD__21__1_, uart1_r_RHOLD__21__2_, uart1_r_RHOLD__21__3_,
         uart1_r_RHOLD__21__4_, uart1_r_RHOLD__21__5_, uart1_r_RHOLD__21__6_,
         uart1_r_RHOLD__21__7_, uart1_r_RHOLD__20__0_, uart1_r_RHOLD__20__1_,
         uart1_r_RHOLD__20__2_, uart1_r_RHOLD__20__3_, uart1_r_RHOLD__20__4_,
         uart1_r_RHOLD__20__5_, uart1_r_RHOLD__20__6_, uart1_r_RHOLD__20__7_,
         uart1_r_RHOLD__19__0_, uart1_r_RHOLD__19__1_, uart1_r_RHOLD__19__2_,
         uart1_r_RHOLD__19__3_, uart1_r_RHOLD__19__4_, uart1_r_RHOLD__19__5_,
         uart1_r_RHOLD__19__6_, uart1_r_RHOLD__19__7_, uart1_r_RHOLD__18__0_,
         uart1_r_RHOLD__18__1_, uart1_r_RHOLD__18__2_, uart1_r_RHOLD__18__3_,
         uart1_r_RHOLD__18__4_, uart1_r_RHOLD__18__5_, uart1_r_RHOLD__18__6_,
         uart1_r_RHOLD__18__7_, uart1_r_RHOLD__17__0_, uart1_r_RHOLD__17__1_,
         uart1_r_RHOLD__17__2_, uart1_r_RHOLD__17__3_, uart1_r_RHOLD__17__4_,
         uart1_r_RHOLD__17__5_, uart1_r_RHOLD__17__6_, uart1_r_RHOLD__17__7_,
         uart1_r_RHOLD__16__0_, uart1_r_RHOLD__16__1_, uart1_r_RHOLD__16__2_,
         uart1_r_RHOLD__16__3_, uart1_r_RHOLD__16__4_, uart1_r_RHOLD__16__5_,
         uart1_r_RHOLD__16__6_, uart1_r_RHOLD__16__7_, uart1_r_RHOLD__15__0_,
         uart1_r_RHOLD__15__1_, uart1_r_RHOLD__15__2_, uart1_r_RHOLD__15__3_,
         uart1_r_RHOLD__15__4_, uart1_r_RHOLD__15__5_, uart1_r_RHOLD__15__6_,
         uart1_r_RHOLD__15__7_, uart1_r_RHOLD__14__0_, uart1_r_RHOLD__14__1_,
         uart1_r_RHOLD__14__2_, uart1_r_RHOLD__14__3_, uart1_r_RHOLD__14__4_,
         uart1_r_RHOLD__14__5_, uart1_r_RHOLD__14__6_, uart1_r_RHOLD__14__7_,
         uart1_r_RHOLD__13__0_, uart1_r_RHOLD__13__1_, uart1_r_RHOLD__13__2_,
         uart1_r_RHOLD__13__3_, uart1_r_RHOLD__13__4_, uart1_r_RHOLD__13__5_,
         uart1_r_RHOLD__13__6_, uart1_r_RHOLD__13__7_, uart1_r_RHOLD__12__0_,
         uart1_r_RHOLD__12__1_, uart1_r_RHOLD__12__2_, uart1_r_RHOLD__12__3_,
         uart1_r_RHOLD__12__4_, uart1_r_RHOLD__12__5_, uart1_r_RHOLD__12__6_,
         uart1_r_RHOLD__12__7_, uart1_r_RHOLD__11__0_, uart1_r_RHOLD__11__1_,
         uart1_r_RHOLD__11__2_, uart1_r_RHOLD__11__3_, uart1_r_RHOLD__11__4_,
         uart1_r_RHOLD__11__5_, uart1_r_RHOLD__11__6_, uart1_r_RHOLD__11__7_,
         uart1_r_RHOLD__10__0_, uart1_r_RHOLD__10__1_, uart1_r_RHOLD__10__2_,
         uart1_r_RHOLD__10__3_, uart1_r_RHOLD__10__4_, uart1_r_RHOLD__10__5_,
         uart1_r_RHOLD__10__6_, uart1_r_RHOLD__10__7_, uart1_r_RHOLD__9__0_,
         uart1_r_RHOLD__9__1_, uart1_r_RHOLD__9__2_, uart1_r_RHOLD__9__3_,
         uart1_r_RHOLD__9__4_, uart1_r_RHOLD__9__5_, uart1_r_RHOLD__9__6_,
         uart1_r_RHOLD__9__7_, uart1_r_RHOLD__8__0_, uart1_r_RHOLD__8__1_,
         uart1_r_RHOLD__8__2_, uart1_r_RHOLD__8__3_, uart1_r_RHOLD__8__4_,
         uart1_r_RHOLD__8__5_, uart1_r_RHOLD__8__6_, uart1_r_RHOLD__8__7_,
         uart1_r_RHOLD__7__0_, uart1_r_RHOLD__7__1_, uart1_r_RHOLD__7__2_,
         uart1_r_RHOLD__7__3_, uart1_r_RHOLD__7__4_, uart1_r_RHOLD__7__5_,
         uart1_r_RHOLD__7__6_, uart1_r_RHOLD__7__7_, uart1_r_RHOLD__6__0_,
         uart1_r_RHOLD__6__1_, uart1_r_RHOLD__6__2_, uart1_r_RHOLD__6__3_,
         uart1_r_RHOLD__6__4_, uart1_r_RHOLD__6__5_, uart1_r_RHOLD__6__6_,
         uart1_r_RHOLD__6__7_, uart1_r_RHOLD__5__0_, uart1_r_RHOLD__5__1_,
         uart1_r_RHOLD__5__2_, uart1_r_RHOLD__5__3_, uart1_r_RHOLD__5__4_,
         uart1_r_RHOLD__5__5_, uart1_r_RHOLD__5__6_, uart1_r_RHOLD__5__7_,
         uart1_r_RHOLD__4__0_, uart1_r_RHOLD__4__1_, uart1_r_RHOLD__4__2_,
         uart1_r_RHOLD__4__3_, uart1_r_RHOLD__4__4_, uart1_r_RHOLD__4__5_,
         uart1_r_RHOLD__4__6_, uart1_r_RHOLD__4__7_, uart1_r_RHOLD__3__0_,
         uart1_r_RHOLD__3__1_, uart1_r_RHOLD__3__2_, uart1_r_RHOLD__3__3_,
         uart1_r_RHOLD__3__4_, uart1_r_RHOLD__3__5_, uart1_r_RHOLD__3__6_,
         uart1_r_RHOLD__3__7_, uart1_r_RHOLD__2__0_, uart1_r_RHOLD__2__1_,
         uart1_r_RHOLD__2__2_, uart1_r_RHOLD__2__3_, uart1_r_RHOLD__2__4_,
         uart1_r_RHOLD__2__5_, uart1_r_RHOLD__2__6_, uart1_r_RHOLD__2__7_,
         uart1_r_RHOLD__1__0_, uart1_r_RHOLD__1__1_, uart1_r_RHOLD__1__2_,
         uart1_r_RHOLD__1__3_, uart1_r_RHOLD__1__4_, uart1_r_RHOLD__1__5_,
         uart1_r_RHOLD__1__6_, uart1_r_RHOLD__1__7_, uart1_r_RHOLD__0__0_,
         uart1_r_RHOLD__0__1_, uart1_r_RHOLD__0__2_, uart1_r_RHOLD__0__3_,
         uart1_r_RHOLD__0__4_, uart1_r_RHOLD__0__5_, uart1_r_RHOLD__0__6_,
         uart1_r_RHOLD__0__7_, uart1_r_EXTCLKEN_, uart1_r_FRAME_,
         uart1_r_PARERR_, uart1_r_OVF_, uart1_r_BREAKIRQEN_, uart1_r_BREAK_,
         uart1_r_TSEMPTYIRQEN_, uart1_r_TSEMPTY_, uart1_r_RSEMPTY_,
         uart1_r_LOOPB_, uart1_r_FLOW_, uart1_r_PAREN_, uart1_r_PARSEL_,
         uart1_r_TIRQEN_, uart1_r_RIRQEN_, uart1_v_RWADDR__3_, uart1_v_RXF__1_,
         uart1_v_SCALER__11_, uart1_v_RXDB__1_, uart1_v_RXCLK__2_,
         uart1_v_TXTICK_, uart1_v_TXCLK__2_, uart1_uarto_RXEN_,
         uart1_uarto_TXEN_, uart1_uarto_SCALER__0_, uart1_uarto_SCALER__1_,
         uart1_uarto_SCALER__2_, uart1_uarto_SCALER__3_,
         uart1_uarto_SCALER__4_, uart1_uarto_SCALER__5_,
         uart1_uarto_SCALER__6_, uart1_uarto_SCALER__7_,
         uart1_uarto_SCALER__8_, uart1_uarto_SCALER__9_,
         uart1_uarto_SCALER__10_, uart1_uarto_SCALER__11_,
         irqctrl0_r_IFORCE__0__1_, irqctrl0_r_IFORCE__0__2_,
         irqctrl0_r_IFORCE__0__3_, irqctrl0_r_IFORCE__0__4_,
         irqctrl0_r_IFORCE__0__5_, irqctrl0_r_IFORCE__0__6_,
         irqctrl0_r_IFORCE__0__7_, irqctrl0_r_IFORCE__0__8_,
         irqctrl0_r_IFORCE__0__9_, irqctrl0_r_IFORCE__0__10_,
         irqctrl0_r_IFORCE__0__11_, irqctrl0_r_IFORCE__0__12_,
         irqctrl0_r_IFORCE__0__13_, irqctrl0_r_IFORCE__0__14_,
         irqctrl0_r_IFORCE__0__15_, irqctrl0_r_IPEND__1_, irqctrl0_r_IPEND__2_,
         irqctrl0_r_IPEND__3_, irqctrl0_r_IPEND__4_, irqctrl0_r_IPEND__5_,
         irqctrl0_r_IPEND__6_, irqctrl0_r_IPEND__7_, irqctrl0_r_IPEND__8_,
         irqctrl0_r_IPEND__9_, irqctrl0_r_IPEND__10_, irqctrl0_r_IPEND__11_,
         irqctrl0_r_IPEND__12_, irqctrl0_r_IPEND__13_, irqctrl0_r_IPEND__14_,
         irqctrl0_r_IPEND__15_, irqctrl0_r_ILEVEL__1_, irqctrl0_r_ILEVEL__2_,
         irqctrl0_r_ILEVEL__3_, irqctrl0_r_ILEVEL__4_, irqctrl0_r_ILEVEL__5_,
         irqctrl0_r_ILEVEL__6_, irqctrl0_r_ILEVEL__8_, irqctrl0_r_ILEVEL__9_,
         irqctrl0_r_ILEVEL__10_, irqctrl0_r_ILEVEL__12_,
         irqctrl0_r_ILEVEL__13_, irqctrl0_r_ILEVEL__14_,
         irqctrl0_r_ILEVEL__15_, irqctrl0_r_IMASK__0__1_,
         irqctrl0_r_IMASK__0__2_, irqctrl0_r_IMASK__0__3_,
         irqctrl0_r_IMASK__0__4_, irqctrl0_r_IMASK__0__5_,
         irqctrl0_r_IMASK__0__6_, irqctrl0_r_IMASK__0__8_,
         irqctrl0_r_IMASK__0__9_, irqctrl0_r_IMASK__0__10_,
         irqctrl0_r_IMASK__0__12_, irqctrl0_r_IMASK__0__13_,
         irqctrl0_r_IMASK__0__14_, irqctrl0_r_IMASK__0__15_,
         irqctrl0_v_IRL__0__1_, irqctrl0_v_IRL__0__2_, irqctrl0_v_IRL__0__3_,
         timer0_res_1_, timer0_res_2_, timer0_res_3_, timer0_res_4_,
         timer0_res_5_, timer0_res_6_, timer0_res_7_, timer0_res_8_,
         timer0_res_9_, timer0_res_10_, timer0_res_11_, timer0_res_12_,
         timer0_res_13_, timer0_res_14_, timer0_res_15_, timer0_res_16_,
         timer0_res_17_, timer0_res_18_, timer0_res_19_, timer0_res_20_,
         timer0_res_21_, timer0_res_22_, timer0_res_23_, timer0_res_24_,
         timer0_res_25_, timer0_res_26_, timer0_res_27_, timer0_res_28_,
         timer0_res_29_, timer0_res_30_, timer0_res_31_, timer0_N91,
         timer0_N90, timer0_N89, timer0_N88, timer0_N87, timer0_N86,
         timer0_N85, timer0_N84, timer0_N83, timer0_N82, timer0_N81,
         timer0_N80, timer0_N79, timer0_N78, timer0_N77, timer0_N76,
         timer0_N75, timer0_N74, timer0_N73, timer0_N72, timer0_N71,
         timer0_N70, timer0_N69, timer0_N68, timer0_N67, timer0_N66,
         timer0_N65, timer0_N64, timer0_N63, timer0_N62, timer0_N61,
         timer0_N60, timer0_scaler_1_, timer0_scaler_2_, timer0_scaler_3_,
         timer0_scaler_4_, timer0_scaler_5_, timer0_scaler_6_,
         timer0_vtimers_1__RELOAD__0_, timer0_vtimers_1__RELOAD__1_,
         timer0_vtimers_1__RELOAD__2_, timer0_vtimers_1__RELOAD__3_,
         timer0_vtimers_1__RELOAD__4_, timer0_vtimers_1__RELOAD__5_,
         timer0_vtimers_1__RELOAD__6_, timer0_vtimers_1__RELOAD__7_,
         timer0_vtimers_1__RELOAD__8_, timer0_vtimers_1__RELOAD__9_,
         timer0_vtimers_1__RELOAD__10_, timer0_vtimers_1__RELOAD__11_,
         timer0_vtimers_1__RELOAD__12_, timer0_vtimers_1__RELOAD__13_,
         timer0_vtimers_1__RELOAD__14_, timer0_vtimers_1__RELOAD__15_,
         timer0_vtimers_1__RELOAD__16_, timer0_vtimers_1__RELOAD__17_,
         timer0_vtimers_1__RELOAD__18_, timer0_vtimers_1__RELOAD__19_,
         timer0_vtimers_1__RELOAD__20_, timer0_vtimers_1__RELOAD__21_,
         timer0_vtimers_1__RELOAD__22_, timer0_vtimers_1__RELOAD__23_,
         timer0_vtimers_1__RELOAD__24_, timer0_vtimers_1__RELOAD__25_,
         timer0_vtimers_1__RELOAD__26_, timer0_vtimers_1__RELOAD__27_,
         timer0_vtimers_1__RELOAD__28_, timer0_vtimers_1__RELOAD__29_,
         timer0_vtimers_1__RELOAD__30_, timer0_vtimers_1__RELOAD__31_,
         timer0_vtimers_1__IRQEN_, timer0_vtimers_1__IRQPEN_,
         timer0_vtimers_1__RESTART_, timer0_vtimers_1__LOAD_,
         timer0_vtimers_1__ENABLE_, timer0_r_DISHLT_, timer0_r_RELOAD__0_,
         timer0_r_RELOAD__1_, timer0_r_RELOAD__2_, timer0_r_RELOAD__3_,
         timer0_r_RELOAD__4_, timer0_r_RELOAD__5_, timer0_r_RELOAD__6_,
         timer0_r_RELOAD__7_, timer0_r_SCALER__0_, timer0_r_SCALER__1_,
         timer0_r_SCALER__2_, timer0_r_SCALER__3_, timer0_r_SCALER__4_,
         timer0_r_SCALER__5_, timer0_r_SCALER__6_, timer0_r_SCALER__7_,
         timer0_v_TIMERS__1__VALUE__0_, timer0_v_TIMERS__1__VALUE__1_,
         timer0_v_TIMERS__1__VALUE__2_, timer0_v_TIMERS__1__VALUE__3_,
         timer0_v_TIMERS__1__VALUE__4_, timer0_v_TIMERS__1__VALUE__5_,
         timer0_v_TIMERS__1__VALUE__6_, timer0_v_TIMERS__1__VALUE__7_,
         timer0_v_TIMERS__1__VALUE__8_, timer0_v_TIMERS__1__VALUE__9_,
         timer0_v_TIMERS__1__VALUE__10_, timer0_v_TIMERS__1__VALUE__11_,
         timer0_v_TIMERS__1__VALUE__12_, timer0_v_TIMERS__1__VALUE__13_,
         timer0_v_TIMERS__1__VALUE__14_, timer0_v_TIMERS__1__VALUE__15_,
         timer0_v_TIMERS__1__VALUE__16_, timer0_v_TIMERS__1__VALUE__17_,
         timer0_v_TIMERS__1__VALUE__18_, timer0_v_TIMERS__1__VALUE__19_,
         timer0_v_TIMERS__1__VALUE__20_, timer0_v_TIMERS__1__VALUE__21_,
         timer0_v_TIMERS__1__VALUE__22_, timer0_v_TIMERS__1__VALUE__23_,
         timer0_v_TIMERS__1__VALUE__24_, timer0_v_TIMERS__1__VALUE__25_,
         timer0_v_TIMERS__1__VALUE__26_, timer0_v_TIMERS__1__VALUE__27_,
         timer0_v_TIMERS__1__VALUE__28_, timer0_v_TIMERS__1__VALUE__29_,
         timer0_v_TIMERS__1__VALUE__30_, timer0_v_TIMERS__1__VALUE__31_,
         timer0_v_TICK_, timer0_gpto_TICK__1_, timer0_gpto_TICK__0_, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1643, n1645, n1647, n1649, n1651,
         n1653, n1655, n1657, n1659, n1661, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1786, n1788, n1789, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2238, n2239, n2240, n2241, n2242,
         n2243, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2278, n2279, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2295, n2297,
         n2299, n2301, n2302, n2304, n2306, n2307, n2308, n2309, n2310, n2312,
         n2313, n2314, n2316, n2318, n2319, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2333, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2355, n2356, n2357, n2358, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2369, n2372, n2374, n2376, n2378,
         n2380, n2382, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2465, n2466, n2467, n2469, n2471, n2473, n2475, n2477,
         n2479, n2481, n2482, n2483, n2485, n2486, n2488, n2490, n2492, n2493,
         n2494, n2496, n2498, n2500, n2502, n2504, n2506, n2508, n2509, n2510,
         n2512, n2513, n2515, n2517, n2521, n2523, n2525, n2527, n2529, n2531,
         n2533, n2535, n2536, n2537, n2539, n2540, n2542, n2543, n2544, n2546,
         n2548, n2550, n2552, n2554, n2556, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2567, n2569, n2570, n2571, n2572, n2574, n2576, n2578,
         n2580, n2582, n2584, n2586, n2587, n2588, n2590, n2591, n2592, n2593,
         n2595, n2597, n2599, n2601, n2603, n2605, n2607, n2608, n2609, n2611,
         n2612, n2614, n2615, n2616, n2617, n2619, n2621, n2623, n2625, n2627,
         n2629, n2631, n2632, n2633, n2634, n2635, n2636, n2638, n2639, n2640,
         n2641, n2643, n2645, n2647, n2649, n2651, n2653, n2655, n2656, n2657,
         n2659, n2660, n2662, n2663, n2664, n2665, n2667, n2669, n2671, n2673,
         n2675, n2677, n2679, n2680, n2681, n2682, n2683, n2684, n2686, n2687,
         n2688, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2703, n2705, n2706, n2708, n2710, n2712, n2714,
         n2716, n2718, n2720, n2722, n2724, n2725, n2727, n2728, n2730, n2731,
         n2733, n2735, n2736, n2737, n2739, n2740, n2742, n2744, n2745, n2747,
         n2749, n2751, n2753, n2755, n2757, n2758, n2760, n2762, n2764, n2766,
         n2767, n2769, n2770, n2772, n2774, n2776, n2778, n2780, n2782, n2784,
         n2786, n2788, n2790, n2792, n2794, n2796, n2798, n2800, n2802, n2804,
         n2806, n2808, n2810, n2811, n2812, n2813, n2815, n2816, n2818, n2820,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2931, n2932, n2933,
         n2935, n2936, n2937, n2938, n2939, n2940, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3004, n3005, n3006, n3008, n3009, n3011, n3012, n3013,
         n3015, n3016, n3017, n3018, n3019, n3020, n3022, n3023, n3024, n3025,
         n3027, n3028, n3030, n3031, n3033, n3034, n3035, n3036, n3037, n3038,
         n3040, n3041, n3042, n3044, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3065, n3066, n3067, n3068, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3079, n3081, n3083, n3085, n3087, n3089, n3091,
         n3093, n3095, n3097, n3099, n3101, n3103, n3105, n3107, n3109, n3111,
         n3113, n3115, n3117, n3119, n3121, n3123, n3125, n3127, n3129, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3154, n3156, n3158, n3160, n3162, n3164, n3166, n3168, n3170,
         n3172, n3174, n3176, n3178, n3180, n3182, n3184, n3186, n3188, n3190,
         n3192, n3194, n3196, n3198, n3200, n3202, n3204, n3206, n3208, n3210,
         n3212, n3214, n3216, n3218, n3220, n3222, n3224, n3226, n3228, n3230,
         n3232, n3234, n3236, n3238, n3240, n3242, n3244, n3246, n3248, n3250,
         n3252, n3254, n3256, n3258, n3260, n3262, n3264, n3266, n3268, n3270,
         n3272, n3274, n3276, n3278, n3280, n3282, n3284, n3286, n3288, n3290,
         n3292, n3294, n3296, n3298, n3300, n3302, n3304, n3306, n3308, n3310,
         n3312, n3313, n3314, n3316, n3318, n3320, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3332, n3334, n3336, n3338, n3340,
         n3342, n3344, n3346, n3348, n3350, n3352, n3354, n3356, n3358, n3360,
         n3362, n3364, n3366, n3369, n3372, n3374, n3376, n3379, n3381, n3383,
         n3385, n3387, n3389, n3390, n3392, n3394, n3396, n3398, n3400, n3402,
         n3404, n3406, n3408, n3410, n3412, n3414, n3416, n3418, n3420, n3422,
         n3424, n3426, n3428, n3430, n3432, n3434, n3436, n3438, n3440, n3442,
         n3444, n3446, n3448, n3450, n3452, n3454, n3456, n3458, n3460, n3462,
         n3464, n3466, n3468, n3470, n3472, n3474, n3476, n3478, n3480, n3482,
         n3484, n3486, n3488, n3490, n3493, n3495, n3497, n3499, n3501, n3503,
         n3505, n3507, n3509, n3512, n3514, n3516, n3518, n3522, n3524, n3526,
         n3528, n3530, n3532, n3534, n3536, n3538, n3540, n3542, n3544, n3546,
         n3548, n3550, n3552, n3554, n3556, n3558, n3560, n3562, n3564, n3566,
         n3568, n3570, n3572, n3574, n3576, n3578, n3580, n3582, n3584, n3586,
         n3588, n3590, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3602, n3604, n3606, n3614, n3616, n3621, n3636, n3640, n3642,
         n3645, n3648, n3651, n3653, n3655, n3657, n3660, n3662, n3664, n3666,
         n3669, n3671, n3673, n3675, n3678, n3680, n3682, n3684, n3687, n3689,
         n3691, n3694, n3696, n3698, n3700, n3702, n3703, n3704, n3705, n3707,
         n3709, n3711, n3713, n3715, n3717, n3719, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3730, n3731, n3733, n3735, n3737, n3739,
         n3741, n3743, n3745, n3747, n3750, n3752, n3754, n3756, n3758, n3760,
         n3762, n3764, n3766, n3769, n3771, n3773, n3775, n3778, n3780, n3782,
         n3784, n3786, n3788, n3790, n3792, n3794, n3796, n3798, n3800, n3802,
         n3804, n3806, n3808, n3810, n3812, n3814, n3816, n3818, n3820, n3822,
         n3824, n3826, n3828, n3830, n3832, n3834, n3836, n3838, n3840, n3842,
         n3844, n3846, n3848, n3850, n3852, n3854, n3856, n3858, n3860, n3862,
         n3864, n3867, n3869, n3871, n3873, n3875, n3878, n3879, n3880, n3881,
         n3883, n3885, n3887, n3889, n3891, n3894, n3895, n3896, n3897, n3899,
         n3900, n3901, n3904, n3905, n3906, n3907, n3908, n3910, n3912, n3913,
         n3914, n3916, n3917, n3919, n3920, n3922, n3924, n3926, n3928, n3929,
         n3930, n3932, n3934, n3936, n3938, n3940, n3942, n3944, n3946, n3948,
         n3949, n3951, n3953, n3955, n3957, n3959, n3961, n3963, n3965, n3967,
         n3969, n3971, n3973, n3974, n3976, n3978, n3980, n3982, n3984, n3986,
         n3988, n3990, n3991, n3993, n3995, n3997, n3998, n4000, n4002, n4004,
         n4006, n4008, n4010, n4012, n4014, n4016, n4018, n4020, n4022, n4024,
         n4026, n4028, n4031, n4032, n4033, n4034, n4035, n4036, n4038, n4040,
         n4042, n4044, n4045, n4047, n4049, n4051, n4053, n4055, n4057, n4059,
         n4061, n4063, n4065, n4067, n4070, n4071, n4072, n4074, n4076, n4079,
         n4081, n4082, n4083, n4084, n4085, n4087, n4089, n4091, n4093, n4095,
         n4097, n4099, n4101, n4103, n4105, n4107, n4109, n4111, n4113, n4115,
         n4117, n4119, n4121, n4123, n4125, n4127, n4129, n4131, n4133, n4135,
         n4137, n4139, n4141, n4143, n4145, n4147, n4149, n4151, n4153, n4155,
         n4157, n4159, n4161, n4163, n4165, n4167, n4169, n4171, n4173, n4175,
         n4177, n4179, n4181, n4183, n4185, n4187, n4189, n4191, n4193, n4195,
         n4197, n4199, n4201, n4203, n4205, n4207, n4209, n4211, n4213, n4215,
         n4217, n4219, n4221, n4223, n4225, n4227, n4229, n4231, n4233, n4235,
         n4237, n4239, n4241, n4243, n4245, n4247, n4249, n4251, n4253, n4255,
         n4257, n4259, n4261, n4263, n4265, n4267, n4269, n4271, n4273, n4275,
         n4277, n4279, n4281, n4283, n4285, n4287, n4289, n4291, n4293, n4295,
         n4297, n4299, n4301, n4303, n4305, n4307, n4309, n4311, n4313, n4316,
         n4317, n4318, n4319, n4321, n4322, n4324, n4325, n4326, n4328, n4330,
         n4332, n4334, n4336, n4338, n4340, n4341, n4343, n4344, n4346, n4348,
         n4350, n4353, n4354, n4355, n4356, n4357, n4358, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4376, n4378, n4379, n4380, n4382, n4383, n4384, n4385,
         n4386, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4396, n4397,
         n4399, n4400, n4402, n4404, n4406, n4408, n4410, n4413, n4414, n4415,
         n4416, n4417, n4418, n4420, n4421, n4423, n4425, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4438, n4440, n4441,
         n4443, n4445, n4447, n4449, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4461, n4463, n4465, n4467, n4469, n4471, n4473,
         n4474, n4475, n4476, n4477, n4478, n4480, n4481, n4483, n4485, n4488,
         n4490, n4492, n4493, n4496, n4497, n4498, n4499, n4500, n4501, n4503,
         n4505, n4507, n4508, n4509, n4511, n4512, n4513, n4515, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4551, n4553, n4554, n4555, n4557, n4558, n4559, n4560, n4561,
         n4562, n4564, n4565, n4567, n4569, n4572, n4573, n4574, n4575, n4576,
         n4577, n4579, n4581, n4583, n4585, n4586, n4587, n4589, n4590, n4592,
         n4594, n4595, n4596, n4597, n4599, n4601, n4602, n4604, n4605, n4607,
         n4609, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4629, n4634, n4635,
         n4636, n4637, n4638, n4639, n4641, n4642, n4643, n4644, n4645, n4646,
         n4648, n4649, n4650, n4651, n4652, n4654, n4656, n4657, n4658, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4675, n4676, n4677, n4679, n4681, n4683, n4684,
         n4685, n4686, n4687, n4688, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4698, n4699, n4700, n4701, n4702, n4703, n4705, n4707, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4719, n4722, n4723,
         n4724, n4725, n4726, n4727, n4729, n4730, n4731, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4751, n4752, n4753, n4754, n4755, n4756,
         n4758, n4759, n4760, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4818, n4821, n4824, n4827,
         n4828, n4832, n4838, n4927, n4928, n4929, n4930, n4948, n4949, n5014,
         n5061, n5590, n5591, n5592, n10972, n10988, n11260, n11537, n12995,
         n13499, n14803, n15074, n15075, n16599, n16838, n16969, n17066,
         n17243, n17251, n17252, n17270, n17271, n17273, n17278, n17284,
         n17285, n17288, n17422, n17443, n17444, n17445, n17450, n17455,
         n17456, n17457, n17458, n17459, n17717, n17722, n17778, n17785,
         n17802, n17804, n17805, n17812, n17853, n17857, n17885, n17886,
         n17887, n17889, n17890, n17903, n17904, n18045, n18047, n18049,
         n18051, n18053, n18089, n18090, n18096, n18100, n18101, n18102,
         n18168, n18171, n18172, n18174, n18175, n18176, n18209, n18210,
         n18211, n18212, n18213, n18248, n18252, n18276, n18277,
         add_x_746_n155, add_x_746_n153, add_x_746_n152, add_x_746_n151,
         add_x_746_n149, add_x_746_n148, add_x_746_n146, add_x_746_n145,
         add_x_746_n144, add_x_746_n143, add_x_746_n140, add_x_746_n139,
         add_x_746_n135, add_x_746_n134, add_x_746_n133, add_x_746_n131,
         add_x_746_n130, add_x_746_n129, add_x_746_n127, add_x_746_n126,
         add_x_746_n125, add_x_746_n124, add_x_746_n123, add_x_746_n121,
         add_x_746_n120, add_x_746_n116, add_x_746_n115, add_x_746_n114,
         add_x_746_n113, add_x_746_n110, add_x_746_n109, add_x_746_n108,
         add_x_746_n106, add_x_746_n104, add_x_746_n103, add_x_746_n102,
         add_x_746_n99, add_x_746_n98, add_x_746_n97, add_x_746_n96,
         add_x_746_n92, add_x_746_n91, add_x_746_n90, add_x_746_n89,
         add_x_746_n86, add_x_746_n85, add_x_746_n84, add_x_746_n78,
         add_x_746_n76, add_x_746_n75, add_x_746_n71, add_x_746_n70,
         add_x_746_n69, add_x_746_n68, add_x_746_n65, add_x_746_n64,
         add_x_746_n63, add_x_746_n61, add_x_746_n59, add_x_746_n58,
         add_x_746_n57, add_x_746_n56, add_x_746_n53, add_x_746_n52,
         add_x_746_n51, add_x_746_n47, add_x_746_n46, add_x_746_n45,
         add_x_746_n44, add_x_746_n41, add_x_746_n40, add_x_746_n39,
         add_x_746_n37, add_x_746_n36, add_x_746_n34, add_x_746_n33,
         add_x_746_n32, add_x_746_n29, add_x_746_n28, add_x_746_n27,
         add_x_746_n23, add_x_746_n22, add_x_746_n21, add_x_746_n20,
         add_x_746_n17, add_x_746_n16, add_x_746_n15, add_x_746_n13,
         add_x_746_n12, add_x_746_n10, add_x_746_n9, add_x_746_n8,
         add_x_746_n5, add_x_746_n4, add_x_746_n2, add_x_746_n1,
         DP_OP_5187J1_124_3275_n336, DP_OP_5187J1_124_3275_n335,
         DP_OP_5187J1_124_3275_n334, DP_OP_5187J1_124_3275_n332,
         DP_OP_5187J1_124_3275_n330, DP_OP_5187J1_124_3275_n329,
         DP_OP_5187J1_124_3275_n327, DP_OP_5187J1_124_3275_n326,
         DP_OP_5187J1_124_3275_n323, DP_OP_5187J1_124_3275_n322,
         DP_OP_5187J1_124_3275_n321, DP_OP_5187J1_124_3275_n320,
         DP_OP_5187J1_124_3275_n319, DP_OP_5187J1_124_3275_n318,
         DP_OP_5187J1_124_3275_n317, DP_OP_5187J1_124_3275_n316,
         DP_OP_5187J1_124_3275_n315, DP_OP_5187J1_124_3275_n314,
         DP_OP_5187J1_124_3275_n313, DP_OP_5187J1_124_3275_n312,
         DP_OP_5187J1_124_3275_n311, DP_OP_5187J1_124_3275_n310,
         DP_OP_5187J1_124_3275_n308, DP_OP_5187J1_124_3275_n306,
         DP_OP_5187J1_124_3275_n305, DP_OP_5187J1_124_3275_n304,
         DP_OP_5187J1_124_3275_n301, DP_OP_5187J1_124_3275_n300,
         DP_OP_5187J1_124_3275_n299, DP_OP_5187J1_124_3275_n298,
         DP_OP_5187J1_124_3275_n297, DP_OP_5187J1_124_3275_n296,
         DP_OP_5187J1_124_3275_n295, DP_OP_5187J1_124_3275_n294,
         DP_OP_5187J1_124_3275_n293, DP_OP_5187J1_124_3275_n292,
         DP_OP_5187J1_124_3275_n291, DP_OP_5187J1_124_3275_n290,
         DP_OP_5187J1_124_3275_n289, DP_OP_5187J1_124_3275_n288,
         DP_OP_5187J1_124_3275_n287, DP_OP_5187J1_124_3275_n286,
         DP_OP_5187J1_124_3275_n284, DP_OP_5187J1_124_3275_n283,
         DP_OP_5187J1_124_3275_n282, DP_OP_5187J1_124_3275_n279,
         DP_OP_5187J1_124_3275_n278, DP_OP_5187J1_124_3275_n277,
         DP_OP_5187J1_124_3275_n276, DP_OP_5187J1_124_3275_n274,
         DP_OP_5187J1_124_3275_n271, DP_OP_5187J1_124_3275_n270,
         DP_OP_5187J1_124_3275_n269, DP_OP_5187J1_124_3275_n268,
         DP_OP_5187J1_124_3275_n267, DP_OP_5187J1_124_3275_n266,
         DP_OP_5187J1_124_3275_n265, DP_OP_5187J1_124_3275_n264,
         DP_OP_5187J1_124_3275_n263, DP_OP_5187J1_124_3275_n262,
         DP_OP_5187J1_124_3275_n261, DP_OP_5187J1_124_3275_n259,
         DP_OP_5187J1_124_3275_n258, DP_OP_5187J1_124_3275_n257,
         DP_OP_5187J1_124_3275_n256, DP_OP_5187J1_124_3275_n255,
         DP_OP_5187J1_124_3275_n250, DP_OP_5187J1_124_3275_n249,
         DP_OP_5187J1_124_3275_n245, DP_OP_5187J1_124_3275_n244,
         DP_OP_5187J1_124_3275_n238, DP_OP_5187J1_124_3275_n237,
         DP_OP_5187J1_124_3275_n236, DP_OP_5187J1_124_3275_n235,
         DP_OP_5187J1_124_3275_n232, DP_OP_5187J1_124_3275_n231,
         DP_OP_5187J1_124_3275_n230, DP_OP_5187J1_124_3275_n229,
         DP_OP_5187J1_124_3275_n228, DP_OP_5187J1_124_3275_n227,
         DP_OP_5187J1_124_3275_n226, DP_OP_5187J1_124_3275_n225,
         DP_OP_5187J1_124_3275_n223, DP_OP_5187J1_124_3275_n222,
         DP_OP_5187J1_124_3275_n221, DP_OP_5187J1_124_3275_n220,
         DP_OP_5187J1_124_3275_n219, DP_OP_5187J1_124_3275_n214,
         DP_OP_5187J1_124_3275_n213, DP_OP_5187J1_124_3275_n209,
         DP_OP_5187J1_124_3275_n206, DP_OP_5187J1_124_3275_n200,
         DP_OP_5187J1_124_3275_n199, DP_OP_5187J1_124_3275_n198,
         DP_OP_5187J1_124_3275_n197, DP_OP_5187J1_124_3275_n196,
         DP_OP_5187J1_124_3275_n195, DP_OP_5187J1_124_3275_n194,
         DP_OP_5187J1_124_3275_n193, DP_OP_5187J1_124_3275_n191,
         DP_OP_5187J1_124_3275_n190, DP_OP_5187J1_124_3275_n189,
         DP_OP_5187J1_124_3275_n188, DP_OP_5187J1_124_3275_n187,
         DP_OP_5187J1_124_3275_n182, DP_OP_5187J1_124_3275_n181,
         DP_OP_5187J1_124_3275_n180, DP_OP_5187J1_124_3275_n179,
         DP_OP_5187J1_124_3275_n178, DP_OP_5187J1_124_3275_n177,
         DP_OP_5187J1_124_3275_n176, DP_OP_5187J1_124_3275_n175,
         DP_OP_5187J1_124_3275_n173, DP_OP_5187J1_124_3275_n172,
         DP_OP_5187J1_124_3275_n171, DP_OP_5187J1_124_3275_n170,
         DP_OP_5187J1_124_3275_n169, DP_OP_5187J1_124_3275_n168,
         DP_OP_5187J1_124_3275_n167, DP_OP_5187J1_124_3275_n164,
         DP_OP_5187J1_124_3275_n163, DP_OP_5187J1_124_3275_n162,
         DP_OP_5187J1_124_3275_n161, DP_OP_5187J1_124_3275_n160,
         DP_OP_5187J1_124_3275_n159, DP_OP_5187J1_124_3275_n158,
         DP_OP_5187J1_124_3275_n157, DP_OP_5187J1_124_3275_n155,
         DP_OP_5187J1_124_3275_n154, DP_OP_5187J1_124_3275_n153,
         DP_OP_5187J1_124_3275_n152, DP_OP_5187J1_124_3275_n151,
         DP_OP_5187J1_124_3275_n148, DP_OP_5187J1_124_3275_n147,
         DP_OP_5187J1_124_3275_n146, DP_OP_5187J1_124_3275_n145,
         DP_OP_5187J1_124_3275_n144, DP_OP_5187J1_124_3275_n143,
         DP_OP_5187J1_124_3275_n142, DP_OP_5187J1_124_3275_n141,
         DP_OP_5187J1_124_3275_n138, DP_OP_5187J1_124_3275_n137,
         DP_OP_5187J1_124_3275_n136, DP_OP_5187J1_124_3275_n135,
         DP_OP_5187J1_124_3275_n134, DP_OP_5187J1_124_3275_n133,
         DP_OP_5187J1_124_3275_n132, DP_OP_5187J1_124_3275_n131,
         DP_OP_5187J1_124_3275_n130, DP_OP_5187J1_124_3275_n129,
         DP_OP_5187J1_124_3275_n128, DP_OP_5187J1_124_3275_n127,
         DP_OP_5187J1_124_3275_n124, DP_OP_5187J1_124_3275_n123,
         DP_OP_5187J1_124_3275_n122, DP_OP_5187J1_124_3275_n121,
         DP_OP_5187J1_124_3275_n120, DP_OP_5187J1_124_3275_n119,
         DP_OP_5187J1_124_3275_n117, DP_OP_5187J1_124_3275_n116,
         DP_OP_5187J1_124_3275_n115, DP_OP_5187J1_124_3275_n114,
         DP_OP_5187J1_124_3275_n113, DP_OP_5187J1_124_3275_n110,
         DP_OP_5187J1_124_3275_n109, DP_OP_5187J1_124_3275_n108,
         DP_OP_5187J1_124_3275_n107, DP_OP_5187J1_124_3275_n106,
         DP_OP_5187J1_124_3275_n105, DP_OP_5187J1_124_3275_n104,
         DP_OP_5187J1_124_3275_n103, DP_OP_5187J1_124_3275_n100,
         DP_OP_5187J1_124_3275_n99, DP_OP_5187J1_124_3275_n98,
         DP_OP_5187J1_124_3275_n97, DP_OP_5187J1_124_3275_n96,
         DP_OP_5187J1_124_3275_n95, DP_OP_5187J1_124_3275_n94,
         DP_OP_5187J1_124_3275_n93, DP_OP_5187J1_124_3275_n92,
         DP_OP_5187J1_124_3275_n91, DP_OP_5187J1_124_3275_n88,
         DP_OP_5187J1_124_3275_n87, DP_OP_5187J1_124_3275_n86,
         DP_OP_5187J1_124_3275_n85, DP_OP_5187J1_124_3275_n84,
         DP_OP_5187J1_124_3275_n83, DP_OP_5187J1_124_3275_n80,
         DP_OP_5187J1_124_3275_n79, DP_OP_5187J1_124_3275_n78,
         DP_OP_5187J1_124_3275_n77, DP_OP_5187J1_124_3275_n76,
         DP_OP_5187J1_124_3275_n75, DP_OP_5187J1_124_3275_n74,
         DP_OP_5187J1_124_3275_n73, DP_OP_5187J1_124_3275_n72,
         DP_OP_5187J1_124_3275_n71, DP_OP_5187J1_124_3275_n70,
         DP_OP_5187J1_124_3275_n69, DP_OP_5187J1_124_3275_n68,
         DP_OP_5187J1_124_3275_n67, DP_OP_5187J1_124_3275_n66,
         DP_OP_5187J1_124_3275_n65, DP_OP_5187J1_124_3275_n64,
         DP_OP_5187J1_124_3275_n63, DP_OP_5187J1_124_3275_n62,
         DP_OP_5187J1_124_3275_n61, DP_OP_5187J1_124_3275_n60,
         DP_OP_5187J1_124_3275_n59, DP_OP_5187J1_124_3275_n58,
         DP_OP_5187J1_124_3275_n57, DP_OP_5187J1_124_3275_n56,
         DP_OP_5187J1_124_3275_n55, DP_OP_5187J1_124_3275_n54,
         DP_OP_5187J1_124_3275_n53, DP_OP_5187J1_124_3275_n52,
         DP_OP_5187J1_124_3275_n51, DP_OP_5187J1_124_3275_n50,
         DP_OP_5187J1_124_3275_n49, DP_OP_5187J1_124_3275_n48,
         DP_OP_5187J1_124_3275_n47, DP_OP_5187J1_124_3275_n46,
         DP_OP_5187J1_124_3275_n45, DP_OP_5187J1_124_3275_n44,
         DP_OP_5187J1_124_3275_n43, DP_OP_5187J1_124_3275_n42,
         DP_OP_5187J1_124_3275_n41, DP_OP_5187J1_124_3275_n36,
         DP_OP_5187J1_124_3275_n34, DP_OP_5187J1_124_3275_n32,
         DP_OP_5187J1_124_3275_n30, DP_OP_5187J1_124_3275_n27,
         DP_OP_5187J1_124_3275_n26, DP_OP_5187J1_124_3275_n23,
         DP_OP_5187J1_124_3275_n14, DP_OP_5187J1_124_3275_n13,
         DP_OP_5187J1_124_3275_n11, DP_OP_5187J1_124_3275_n8,
         DP_OP_5187J1_124_3275_n7, DP_OP_5187J1_124_3275_n6,
         DP_OP_5187J1_124_3275_n5, DP_OP_5187J1_124_3275_n4,
         DP_OP_5187J1_124_3275_n3, DP_OP_5187J1_124_3275_n2, add_x_735_A_32_,
         add_x_735_A_29_, add_x_735_A_26_, add_x_735_A_25_, add_x_735_A_24_,
         add_x_735_A_22_, add_x_735_A_20_, add_x_735_A_19_, add_x_735_A_16_,
         add_x_735_A_15_, add_x_735_A_14_, add_x_735_A_12_, add_x_735_A_10_,
         add_x_735_A_9_, add_x_735_A_4_, add_x_735_A_2_, add_x_735_n301,
         add_x_735_n299, add_x_735_n298, add_x_735_n297, add_x_735_n296,
         add_x_735_n295, add_x_735_n294, add_x_735_n293, add_x_735_n292,
         add_x_735_n291, add_x_735_n290, add_x_735_n289, add_x_735_n288,
         add_x_735_n287, add_x_735_n286, add_x_735_n285, add_x_735_n284,
         add_x_735_n283, add_x_735_n282, add_x_735_n281, add_x_735_n280,
         add_x_735_n279, add_x_735_n278, add_x_735_n276, add_x_735_n275,
         add_x_735_n274, add_x_735_n272, add_x_735_n270, add_x_735_n268,
         add_x_735_n267, add_x_735_n266, add_x_735_n265, add_x_735_n264,
         add_x_735_n263, add_x_735_n262, add_x_735_n261, add_x_735_n260,
         add_x_735_n259, add_x_735_n258, add_x_735_n257, add_x_735_n256,
         add_x_735_n255, add_x_735_n254, add_x_735_n253, add_x_735_n252,
         add_x_735_n251, add_x_735_n250, add_x_735_n249, add_x_735_n248,
         add_x_735_n247, add_x_735_n246, add_x_735_n245, add_x_735_n242,
         add_x_735_n241, add_x_735_n240, add_x_735_n238, add_x_735_n237,
         add_x_735_n236, add_x_735_n232, add_x_735_n231, add_x_735_n230,
         add_x_735_n229, add_x_735_n228, add_x_735_n225, add_x_735_n224,
         add_x_735_n223, add_x_735_n222, add_x_735_n221, add_x_735_n220,
         add_x_735_n219, add_x_735_n218, add_x_735_n217, add_x_735_n216,
         add_x_735_n215, add_x_735_n214, add_x_735_n213, add_x_735_n212,
         add_x_735_n211, add_x_735_n210, add_x_735_n209, add_x_735_n204,
         add_x_735_n203, add_x_735_n202, add_x_735_n201, add_x_735_n200,
         add_x_735_n199, add_x_735_n198, add_x_735_n197, add_x_735_n195,
         add_x_735_n194, add_x_735_n193, add_x_735_n192, add_x_735_n191,
         add_x_735_n190, add_x_735_n189, add_x_735_n186, add_x_735_n185,
         add_x_735_n184, add_x_735_n183, add_x_735_n182, add_x_735_n181,
         add_x_735_n180, add_x_735_n179, add_x_735_n177, add_x_735_n176,
         add_x_735_n175, add_x_735_n174, add_x_735_n173, add_x_735_n168,
         add_x_735_n167, add_x_735_n166, add_x_735_n165, add_x_735_n164,
         add_x_735_n163, add_x_735_n160, add_x_735_n159, add_x_735_n158,
         add_x_735_n157, add_x_735_n156, add_x_735_n155, add_x_735_n154,
         add_x_735_n153, add_x_735_n152, add_x_735_n151, add_x_735_n150,
         add_x_735_n149, add_x_735_n148, add_x_735_n147, add_x_735_n145,
         add_x_735_n144, add_x_735_n143, add_x_735_n142, add_x_735_n141,
         add_x_735_n136, add_x_735_n135, add_x_735_n134, add_x_735_n133,
         add_x_735_n132, add_x_735_n131, add_x_735_n130, add_x_735_n129,
         add_x_735_n127, add_x_735_n126, add_x_735_n125, add_x_735_n124,
         add_x_735_n123, add_x_735_n122, add_x_735_n121, add_x_735_n118,
         add_x_735_n117, add_x_735_n116, add_x_735_n115, add_x_735_n114,
         add_x_735_n113, add_x_735_n112, add_x_735_n111, add_x_735_n109,
         add_x_735_n108, add_x_735_n107, add_x_735_n106, add_x_735_n105,
         add_x_735_n102, add_x_735_n100, add_x_735_n99, add_x_735_n98,
         add_x_735_n97, add_x_735_n96, add_x_735_n95, add_x_735_n92,
         add_x_735_n91, add_x_735_n90, add_x_735_n89, add_x_735_n88,
         add_x_735_n87, add_x_735_n86, add_x_735_n85, add_x_735_n84,
         add_x_735_n83, add_x_735_n82, add_x_735_n81, add_x_735_n78,
         add_x_735_n77, add_x_735_n76, add_x_735_n75, add_x_735_n74,
         add_x_735_n73, add_x_735_n72, add_x_735_n71, add_x_735_n70,
         add_x_735_n69, add_x_735_n68, add_x_735_n67, add_x_735_n64,
         add_x_735_n62, add_x_735_n61, add_x_735_n60, add_x_735_n59,
         add_x_735_n58, add_x_735_n57, add_x_735_n54, add_x_735_n53,
         add_x_735_n52, add_x_735_n51, add_x_735_n50, add_x_735_n49,
         add_x_735_n48, add_x_735_n47, add_x_735_n46, add_x_735_n45,
         add_x_735_n40, add_x_735_n39, add_x_735_n38, add_x_735_n37,
         add_x_735_n32, add_x_735_n30, add_x_735_n29, add_x_735_n28,
         add_x_735_n27, add_x_735_n26, add_x_735_n25, add_x_735_n24,
         add_x_735_n23, add_x_735_n22, add_x_735_n21, add_x_735_n20,
         add_x_735_n19, add_x_735_n18, add_x_735_n17, add_x_735_n16,
         add_x_735_n15, add_x_735_n14, add_x_735_n13, add_x_735_n12,
         add_x_735_n11, add_x_735_n10, add_x_735_n9, add_x_735_n8,
         add_x_735_n7, add_x_735_n6, add_x_735_n5, add_x_735_n4, add_x_735_n3,
         add_x_735_n2, add_x_735_n1, mult_x_1196_n3330, mult_x_1196_n3329,
         mult_x_1196_n3327, mult_x_1196_n3323, mult_x_1196_n3320,
         mult_x_1196_n3317, mult_x_1196_n3316, mult_x_1196_n3280,
         mult_x_1196_n3279, mult_x_1196_n3278, mult_x_1196_n3277,
         mult_x_1196_n3276, mult_x_1196_n3275, mult_x_1196_n3274,
         mult_x_1196_n3273, mult_x_1196_n3272, mult_x_1196_n3271,
         mult_x_1196_n3270, mult_x_1196_n3269, mult_x_1196_n3268,
         mult_x_1196_n3267, mult_x_1196_n3266, mult_x_1196_n3265,
         mult_x_1196_n3264, mult_x_1196_n3263, mult_x_1196_n3262,
         mult_x_1196_n3261, mult_x_1196_n3260, mult_x_1196_n3259,
         mult_x_1196_n3257, mult_x_1196_n3256, mult_x_1196_n3255,
         mult_x_1196_n3254, mult_x_1196_n3253, mult_x_1196_n3252,
         mult_x_1196_n3251, mult_x_1196_n3250, mult_x_1196_n3249,
         mult_x_1196_n3248, mult_x_1196_n3247, mult_x_1196_n3245,
         mult_x_1196_n3244, mult_x_1196_n3243, mult_x_1196_n3242,
         mult_x_1196_n3241, mult_x_1196_n3240, mult_x_1196_n3239,
         mult_x_1196_n3238, mult_x_1196_n3237, mult_x_1196_n3236,
         mult_x_1196_n3235, mult_x_1196_n3234, mult_x_1196_n3233,
         mult_x_1196_n3232, mult_x_1196_n3231, mult_x_1196_n3230,
         mult_x_1196_n3229, mult_x_1196_n3228, mult_x_1196_n3227,
         mult_x_1196_n3226, mult_x_1196_n3225, mult_x_1196_n3224,
         mult_x_1196_n3223, mult_x_1196_n3222, mult_x_1196_n3221,
         mult_x_1196_n3220, mult_x_1196_n3219, mult_x_1196_n3218,
         mult_x_1196_n3217, mult_x_1196_n3216, mult_x_1196_n3215,
         mult_x_1196_n3214, mult_x_1196_n3213, mult_x_1196_n3212,
         mult_x_1196_n3211, mult_x_1196_n3210, mult_x_1196_n3209,
         mult_x_1196_n3208, mult_x_1196_n3207, mult_x_1196_n3206,
         mult_x_1196_n3205, mult_x_1196_n3204, mult_x_1196_n3203,
         mult_x_1196_n3202, mult_x_1196_n3201, mult_x_1196_n3200,
         mult_x_1196_n3199, mult_x_1196_n3198, mult_x_1196_n3197,
         mult_x_1196_n3196, mult_x_1196_n3195, mult_x_1196_n3194,
         mult_x_1196_n3193, mult_x_1196_n3192, mult_x_1196_n3191,
         mult_x_1196_n3190, mult_x_1196_n3189, mult_x_1196_n3188,
         mult_x_1196_n3187, mult_x_1196_n3186, mult_x_1196_n3185,
         mult_x_1196_n3184, mult_x_1196_n3183, mult_x_1196_n3182,
         mult_x_1196_n3181, mult_x_1196_n3180, mult_x_1196_n3179,
         mult_x_1196_n3178, mult_x_1196_n3177, mult_x_1196_n3176,
         mult_x_1196_n3175, mult_x_1196_n3174, mult_x_1196_n3173,
         mult_x_1196_n3172, mult_x_1196_n3171, mult_x_1196_n3170,
         mult_x_1196_n3169, mult_x_1196_n3168, mult_x_1196_n3167,
         mult_x_1196_n3166, mult_x_1196_n3165, mult_x_1196_n3163,
         mult_x_1196_n3162, mult_x_1196_n3161, mult_x_1196_n3160,
         mult_x_1196_n3159, mult_x_1196_n3158, mult_x_1196_n3157,
         mult_x_1196_n3156, mult_x_1196_n3155, mult_x_1196_n3154,
         mult_x_1196_n3153, mult_x_1196_n3152, mult_x_1196_n3151,
         mult_x_1196_n3150, mult_x_1196_n3149, mult_x_1196_n3148,
         mult_x_1196_n3147, mult_x_1196_n3146, mult_x_1196_n3145,
         mult_x_1196_n3144, mult_x_1196_n3143, mult_x_1196_n3142,
         mult_x_1196_n3141, mult_x_1196_n3140, mult_x_1196_n3139,
         mult_x_1196_n3138, mult_x_1196_n3137, mult_x_1196_n3136,
         mult_x_1196_n3135, mult_x_1196_n3134, mult_x_1196_n3133,
         mult_x_1196_n3132, mult_x_1196_n3131, mult_x_1196_n3130,
         mult_x_1196_n3128, mult_x_1196_n3127, mult_x_1196_n3126,
         mult_x_1196_n3125, mult_x_1196_n3124, mult_x_1196_n3123,
         mult_x_1196_n3122, mult_x_1196_n3121, mult_x_1196_n3120,
         mult_x_1196_n3119, mult_x_1196_n3118, mult_x_1196_n3117,
         mult_x_1196_n3116, mult_x_1196_n3115, mult_x_1196_n3114,
         mult_x_1196_n3113, mult_x_1196_n3112, mult_x_1196_n3111,
         mult_x_1196_n3110, mult_x_1196_n3109, mult_x_1196_n3108,
         mult_x_1196_n3107, mult_x_1196_n3106, mult_x_1196_n3105,
         mult_x_1196_n3104, mult_x_1196_n3103, mult_x_1196_n3102,
         mult_x_1196_n3101, mult_x_1196_n3100, mult_x_1196_n3099,
         mult_x_1196_n3098, mult_x_1196_n3097, mult_x_1196_n3095,
         mult_x_1196_n3094, mult_x_1196_n3093, mult_x_1196_n3092,
         mult_x_1196_n3091, mult_x_1196_n3090, mult_x_1196_n3089,
         mult_x_1196_n3088, mult_x_1196_n3087, mult_x_1196_n3086,
         mult_x_1196_n3085, mult_x_1196_n3084, mult_x_1196_n3083,
         mult_x_1196_n3082, mult_x_1196_n3081, mult_x_1196_n3080,
         mult_x_1196_n3079, mult_x_1196_n3078, mult_x_1196_n3077,
         mult_x_1196_n3076, mult_x_1196_n3075, mult_x_1196_n3074,
         mult_x_1196_n3073, mult_x_1196_n3072, mult_x_1196_n3071,
         mult_x_1196_n3070, mult_x_1196_n3069, mult_x_1196_n3068,
         mult_x_1196_n3067, mult_x_1196_n3066, mult_x_1196_n3065,
         mult_x_1196_n3064, mult_x_1196_n3063, mult_x_1196_n3062,
         mult_x_1196_n3061, mult_x_1196_n3060, mult_x_1196_n3059,
         mult_x_1196_n3058, mult_x_1196_n3057, mult_x_1196_n3056,
         mult_x_1196_n3055, mult_x_1196_n3054, mult_x_1196_n3053,
         mult_x_1196_n3052, mult_x_1196_n3051, mult_x_1196_n3050,
         mult_x_1196_n3049, mult_x_1196_n3048, mult_x_1196_n3047,
         mult_x_1196_n3046, mult_x_1196_n3045, mult_x_1196_n3044,
         mult_x_1196_n3043, mult_x_1196_n3042, mult_x_1196_n3041,
         mult_x_1196_n3039, mult_x_1196_n3038, mult_x_1196_n3037,
         mult_x_1196_n3036, mult_x_1196_n3035, mult_x_1196_n3034,
         mult_x_1196_n3033, mult_x_1196_n3032, mult_x_1196_n3031,
         mult_x_1196_n3030, mult_x_1196_n3029, mult_x_1196_n3028,
         mult_x_1196_n3027, mult_x_1196_n3026, mult_x_1196_n3025,
         mult_x_1196_n3024, mult_x_1196_n3023, mult_x_1196_n3022,
         mult_x_1196_n3021, mult_x_1196_n3020, mult_x_1196_n3019,
         mult_x_1196_n3018, mult_x_1196_n3017, mult_x_1196_n3016,
         mult_x_1196_n3015, mult_x_1196_n3014, mult_x_1196_n3013,
         mult_x_1196_n3012, mult_x_1196_n3011, mult_x_1196_n3010,
         mult_x_1196_n3009, mult_x_1196_n3008, mult_x_1196_n3007,
         mult_x_1196_n3006, mult_x_1196_n3005, mult_x_1196_n3004,
         mult_x_1196_n3003, mult_x_1196_n3002, mult_x_1196_n3001,
         mult_x_1196_n3000, mult_x_1196_n2999, mult_x_1196_n2998,
         mult_x_1196_n2997, mult_x_1196_n2996, mult_x_1196_n2995,
         mult_x_1196_n2994, mult_x_1196_n2993, mult_x_1196_n2992,
         mult_x_1196_n2991, mult_x_1196_n2990, mult_x_1196_n2989,
         mult_x_1196_n2988, mult_x_1196_n2987, mult_x_1196_n2986,
         mult_x_1196_n2985, mult_x_1196_n2984, mult_x_1196_n2983,
         mult_x_1196_n2982, mult_x_1196_n2981, mult_x_1196_n2980,
         mult_x_1196_n2979, mult_x_1196_n2978, mult_x_1196_n2977,
         mult_x_1196_n2976, mult_x_1196_n2975, mult_x_1196_n2973,
         mult_x_1196_n2972, mult_x_1196_n2971, mult_x_1196_n2970,
         mult_x_1196_n2969, mult_x_1196_n2968, mult_x_1196_n2967,
         mult_x_1196_n2966, mult_x_1196_n2965, mult_x_1196_n2964,
         mult_x_1196_n2963, mult_x_1196_n2962, mult_x_1196_n2961,
         mult_x_1196_n2960, mult_x_1196_n2959, mult_x_1196_n2958,
         mult_x_1196_n2957, mult_x_1196_n2956, mult_x_1196_n2955,
         mult_x_1196_n2954, mult_x_1196_n2953, mult_x_1196_n2952,
         mult_x_1196_n2951, mult_x_1196_n2950, mult_x_1196_n2949,
         mult_x_1196_n2948, mult_x_1196_n2947, mult_x_1196_n2946,
         mult_x_1196_n2945, mult_x_1196_n2944, mult_x_1196_n2943,
         mult_x_1196_n2942, mult_x_1196_n2941, mult_x_1196_n2939,
         mult_x_1196_n2938, mult_x_1196_n2936, mult_x_1196_n2935,
         mult_x_1196_n2934, mult_x_1196_n2933, mult_x_1196_n2932,
         mult_x_1196_n2931, mult_x_1196_n2930, mult_x_1196_n2929,
         mult_x_1196_n2928, mult_x_1196_n2927, mult_x_1196_n2926,
         mult_x_1196_n2925, mult_x_1196_n2924, mult_x_1196_n2923,
         mult_x_1196_n2922, mult_x_1196_n2921, mult_x_1196_n2920,
         mult_x_1196_n2919, mult_x_1196_n2918, mult_x_1196_n2917,
         mult_x_1196_n2916, mult_x_1196_n2915, mult_x_1196_n2914,
         mult_x_1196_n2913, mult_x_1196_n2912, mult_x_1196_n2911,
         mult_x_1196_n2910, mult_x_1196_n2909, mult_x_1196_n2908,
         mult_x_1196_n2907, mult_x_1196_n2906, mult_x_1196_n2905,
         mult_x_1196_n2904, mult_x_1196_n2903, mult_x_1196_n2902,
         mult_x_1196_n2901, mult_x_1196_n2900, mult_x_1196_n2899,
         mult_x_1196_n2898, mult_x_1196_n2897, mult_x_1196_n2896,
         mult_x_1196_n2895, mult_x_1196_n2894, mult_x_1196_n2893,
         mult_x_1196_n2892, mult_x_1196_n2891, mult_x_1196_n2890,
         mult_x_1196_n2889, mult_x_1196_n2888, mult_x_1196_n2887,
         mult_x_1196_n2886, mult_x_1196_n2885, mult_x_1196_n2884,
         mult_x_1196_n2882, mult_x_1196_n2881, mult_x_1196_n2880,
         mult_x_1196_n2879, mult_x_1196_n2878, mult_x_1196_n2877,
         mult_x_1196_n2876, mult_x_1196_n2875, mult_x_1196_n2874,
         mult_x_1196_n2873, mult_x_1196_n2872, mult_x_1196_n2871,
         mult_x_1196_n2870, mult_x_1196_n2868, mult_x_1196_n2867,
         mult_x_1196_n2866, mult_x_1196_n2865, mult_x_1196_n2864,
         mult_x_1196_n2863, mult_x_1196_n2862, mult_x_1196_n2861,
         mult_x_1196_n2859, mult_x_1196_n2858, mult_x_1196_n2857,
         mult_x_1196_n2856, mult_x_1196_n2855, mult_x_1196_n2854,
         mult_x_1196_n2853, mult_x_1196_n2852, mult_x_1196_n2851,
         mult_x_1196_n2850, mult_x_1196_n2849, mult_x_1196_n2848,
         mult_x_1196_n2847, mult_x_1196_n2846, mult_x_1196_n2845,
         mult_x_1196_n2844, mult_x_1196_n2843, mult_x_1196_n2842,
         mult_x_1196_n2841, mult_x_1196_n2840, mult_x_1196_n2839,
         mult_x_1196_n2838, mult_x_1196_n2836, mult_x_1196_n2835,
         mult_x_1196_n2834, mult_x_1196_n2833, mult_x_1196_n2832,
         mult_x_1196_n2831, mult_x_1196_n2830, mult_x_1196_n2829,
         mult_x_1196_n2828, mult_x_1196_n2826, mult_x_1196_n2824,
         mult_x_1196_n2823, mult_x_1196_n2822, mult_x_1196_n2821,
         mult_x_1196_n2820, mult_x_1196_n2819, mult_x_1196_n2818,
         mult_x_1196_n2817, mult_x_1196_n2816, mult_x_1196_n2815,
         mult_x_1196_n2814, mult_x_1196_n2813, mult_x_1196_n2812,
         mult_x_1196_n2811, mult_x_1196_n2810, mult_x_1196_n2809,
         mult_x_1196_n2808, mult_x_1196_n2807, mult_x_1196_n2806,
         mult_x_1196_n2805, mult_x_1196_n2804, mult_x_1196_n2803,
         mult_x_1196_n2802, mult_x_1196_n2801, mult_x_1196_n2800,
         mult_x_1196_n2798, mult_x_1196_n2797, mult_x_1196_n2796,
         mult_x_1196_n2795, mult_x_1196_n2794, mult_x_1196_n2793,
         mult_x_1196_n2792, mult_x_1196_n2791, mult_x_1196_n2790,
         mult_x_1196_n2789, mult_x_1196_n2788, mult_x_1196_n2787,
         mult_x_1196_n2786, mult_x_1196_n2785, mult_x_1196_n2784,
         mult_x_1196_n2783, mult_x_1196_n2782, mult_x_1196_n2781,
         mult_x_1196_n2780, mult_x_1196_n2779, mult_x_1196_n2778,
         mult_x_1196_n2777, mult_x_1196_n2776, mult_x_1196_n2775,
         mult_x_1196_n2774, mult_x_1196_n2773, mult_x_1196_n2772,
         mult_x_1196_n2771, mult_x_1196_n2770, mult_x_1196_n2769,
         mult_x_1196_n2768, mult_x_1196_n2767, mult_x_1196_n2765,
         mult_x_1196_n2764, mult_x_1196_n2763, mult_x_1196_n2762,
         mult_x_1196_n2761, mult_x_1196_n2760, mult_x_1196_n2759,
         mult_x_1196_n2758, mult_x_1196_n2757, mult_x_1196_n2756,
         mult_x_1196_n2755, mult_x_1196_n2754, mult_x_1196_n2753,
         mult_x_1196_n2752, mult_x_1196_n2751, mult_x_1196_n2750,
         mult_x_1196_n2749, mult_x_1196_n2747, mult_x_1196_n2746,
         mult_x_1196_n2745, mult_x_1196_n2744, mult_x_1196_n2743,
         mult_x_1196_n2742, mult_x_1196_n2741, mult_x_1196_n2740,
         mult_x_1196_n2739, mult_x_1196_n2738, mult_x_1196_n2737,
         mult_x_1196_n2736, mult_x_1196_n2734, mult_x_1196_n2733,
         mult_x_1196_n2732, mult_x_1196_n2731, mult_x_1196_n2730,
         mult_x_1196_n2729, mult_x_1196_n2728, mult_x_1196_n2727,
         mult_x_1196_n2726, mult_x_1196_n2725, mult_x_1196_n2724,
         mult_x_1196_n2723, mult_x_1196_n2722, mult_x_1196_n2718,
         mult_x_1196_n2717, mult_x_1196_n2710, mult_x_1196_n2708,
         mult_x_1196_n2703, mult_x_1196_n2702, mult_x_1196_n2701,
         mult_x_1196_n2700, mult_x_1196_n2699, mult_x_1196_n2698,
         mult_x_1196_n2693, mult_x_1196_n2692, mult_x_1196_n2690,
         mult_x_1196_n2689, mult_x_1196_n2688, mult_x_1196_n2687,
         mult_x_1196_n2686, mult_x_1196_n2684, mult_x_1196_n2679,
         mult_x_1196_n2677, mult_x_1196_n2675, mult_x_1196_n2674,
         mult_x_1196_n2673, mult_x_1196_n2670, mult_x_1196_n2669,
         mult_x_1196_n2668, mult_x_1196_n2666, mult_x_1196_n2665,
         mult_x_1196_n2664, mult_x_1196_n2663, mult_x_1196_n2662,
         mult_x_1196_n2658, mult_x_1196_n2657, mult_x_1196_n2655,
         mult_x_1196_n2653, mult_x_1196_n2652, mult_x_1196_n2651,
         mult_x_1196_n2650, mult_x_1196_n2649, mult_x_1196_n2647,
         mult_x_1196_n2646, mult_x_1196_n2645, mult_x_1196_n2644,
         mult_x_1196_n2642, mult_x_1196_n2640, mult_x_1196_n2638,
         mult_x_1196_n2637, mult_x_1196_n2636, mult_x_1196_n2635,
         mult_x_1196_n2633, mult_x_1196_n2632, mult_x_1196_n2631,
         mult_x_1196_n2630, mult_x_1196_n2629, mult_x_1196_n2628,
         mult_x_1196_n2627, mult_x_1196_n2625, mult_x_1196_n2624,
         mult_x_1196_n2623, mult_x_1196_n2622, mult_x_1196_n2619,
         mult_x_1196_n2615, mult_x_1196_n2614, mult_x_1196_n2613,
         mult_x_1196_n2611, mult_x_1196_n2609, mult_x_1196_n2608,
         mult_x_1196_n2607, mult_x_1196_n2606, mult_x_1196_n2605,
         mult_x_1196_n2604, mult_x_1196_n2602, mult_x_1196_n2599,
         mult_x_1196_n2596, mult_x_1196_n2595, mult_x_1196_n2594,
         mult_x_1196_n2589, mult_x_1196_n2588, mult_x_1196_n2587,
         mult_x_1196_n2585, mult_x_1196_n2584, mult_x_1196_n2583,
         mult_x_1196_n2581, mult_x_1196_n2580, mult_x_1196_n2578,
         mult_x_1196_n2577, mult_x_1196_n2576, mult_x_1196_n2574,
         mult_x_1196_n2573, mult_x_1196_n2571, mult_x_1196_n2570,
         mult_x_1196_n2569, mult_x_1196_n2568, mult_x_1196_n2566,
         mult_x_1196_n2565, mult_x_1196_n2564, mult_x_1196_n2563,
         mult_x_1196_n2562, mult_x_1196_n2561, mult_x_1196_n2560,
         mult_x_1196_n2559, mult_x_1196_n2558, mult_x_1196_n2555,
         mult_x_1196_n2554, mult_x_1196_n2552, mult_x_1196_n2551,
         mult_x_1196_n2550, mult_x_1196_n2549, mult_x_1196_n2548,
         mult_x_1196_n2547, mult_x_1196_n2545, mult_x_1196_n2544,
         mult_x_1196_n2540, mult_x_1196_n2539, mult_x_1196_n2538,
         mult_x_1196_n2537, mult_x_1196_n2535, mult_x_1196_n2534,
         mult_x_1196_n2531, mult_x_1196_n2529, mult_x_1196_n2528,
         mult_x_1196_n2527, mult_x_1196_n2526, mult_x_1196_n2521,
         mult_x_1196_n2520, mult_x_1196_n2519, mult_x_1196_n2516,
         mult_x_1196_n2515, mult_x_1196_n2514, mult_x_1196_n2513,
         mult_x_1196_n2512, mult_x_1196_n2510, mult_x_1196_n2509,
         mult_x_1196_n2508, mult_x_1196_n2507, mult_x_1196_n2506,
         mult_x_1196_n2504, mult_x_1196_n2503, mult_x_1196_n2501,
         mult_x_1196_n2498, mult_x_1196_n2496, mult_x_1196_n2495,
         mult_x_1196_n2493, mult_x_1196_n2492, mult_x_1196_n2491,
         mult_x_1196_n2490, mult_x_1196_n2485, mult_x_1196_n2483,
         mult_x_1196_n2481, mult_x_1196_n2480, mult_x_1196_n2478,
         mult_x_1196_n2476, mult_x_1196_n2475, mult_x_1196_n2474,
         mult_x_1196_n2473, mult_x_1196_n2472, mult_x_1196_n2471,
         mult_x_1196_n2470, mult_x_1196_n2468, mult_x_1196_n2467,
         mult_x_1196_n2466, mult_x_1196_n2465, mult_x_1196_n2461,
         mult_x_1196_n2457, mult_x_1196_n2456, mult_x_1196_n2455,
         mult_x_1196_n2454, mult_x_1196_n2453, mult_x_1196_n2452,
         mult_x_1196_n2451, mult_x_1196_n2450, mult_x_1196_n2449,
         mult_x_1196_n2447, mult_x_1196_n2446, mult_x_1196_n2445,
         mult_x_1196_n2444, mult_x_1196_n2443, mult_x_1196_n2440,
         mult_x_1196_n2439, mult_x_1196_n2437, mult_x_1196_n2436,
         mult_x_1196_n2433, mult_x_1196_n2430, mult_x_1196_n2429,
         mult_x_1196_n2426, mult_x_1196_n2422, mult_x_1196_n2419,
         mult_x_1196_n2418, mult_x_1196_n2417, mult_x_1196_n2410,
         mult_x_1196_n2409, mult_x_1196_n2408, mult_x_1196_n2407,
         mult_x_1196_n2406, mult_x_1196_n2405, mult_x_1196_n2404,
         mult_x_1196_n2402, mult_x_1196_n2401, mult_x_1196_n2400,
         mult_x_1196_n2399, mult_x_1196_n2398, mult_x_1196_n2397,
         mult_x_1196_n2396, mult_x_1196_n2395, mult_x_1196_n2394,
         mult_x_1196_n2393, mult_x_1196_n2392, mult_x_1196_n2391,
         mult_x_1196_n2390, mult_x_1196_n2389, mult_x_1196_n2388,
         mult_x_1196_n2387, mult_x_1196_n2386, mult_x_1196_n2385,
         mult_x_1196_n2383, mult_x_1196_n2381, mult_x_1196_n2380,
         mult_x_1196_n2379, mult_x_1196_n2378, mult_x_1196_n2377,
         mult_x_1196_n2376, mult_x_1196_n2375, mult_x_1196_n2374,
         mult_x_1196_n2372, mult_x_1196_n2371, mult_x_1196_n2370,
         mult_x_1196_n2369, mult_x_1196_n2368, mult_x_1196_n2367,
         mult_x_1196_n2365, mult_x_1196_n2364, mult_x_1196_n2363,
         mult_x_1196_n2362, mult_x_1196_n2361, mult_x_1196_n2360,
         mult_x_1196_n2359, mult_x_1196_n2358, mult_x_1196_n2357,
         mult_x_1196_n2356, mult_x_1196_n2355, mult_x_1196_n2354,
         mult_x_1196_n2353, mult_x_1196_n2352, mult_x_1196_n2351,
         mult_x_1196_n2350, mult_x_1196_n2349, mult_x_1196_n2347,
         mult_x_1196_n2345, mult_x_1196_n2344, mult_x_1196_n2343,
         mult_x_1196_n2342, mult_x_1196_n2341, mult_x_1196_n2340,
         mult_x_1196_n2339, mult_x_1196_n2338, mult_x_1196_n2337,
         mult_x_1196_n2336, mult_x_1196_n2335, mult_x_1196_n2334,
         mult_x_1196_n2333, mult_x_1196_n2330, mult_x_1196_n2328,
         mult_x_1196_n2327, mult_x_1196_n2326, mult_x_1196_n2325,
         mult_x_1196_n2324, mult_x_1196_n2323, mult_x_1196_n2319,
         mult_x_1196_n2318, mult_x_1196_n2315, mult_x_1196_n2313,
         mult_x_1196_n2312, mult_x_1196_n2308, mult_x_1196_n2306,
         mult_x_1196_n2305, mult_x_1196_n2302, mult_x_1196_n2301,
         mult_x_1196_n2300, mult_x_1196_n2299, mult_x_1196_n2298,
         mult_x_1196_n2295, mult_x_1196_n2294, mult_x_1196_n2292,
         mult_x_1196_n2290, mult_x_1196_n2289, mult_x_1196_n2288,
         mult_x_1196_n2286, mult_x_1196_n2284, mult_x_1196_n2282,
         mult_x_1196_n2281, mult_x_1196_n2280, mult_x_1196_n2279,
         mult_x_1196_n2278, mult_x_1196_n2277, mult_x_1196_n2275,
         mult_x_1196_n2273, mult_x_1196_n2272, mult_x_1196_n2269,
         mult_x_1196_n2268, mult_x_1196_n2266, mult_x_1196_n2264,
         mult_x_1196_n2262, mult_x_1196_n2258, mult_x_1196_n2257,
         mult_x_1196_n2256, mult_x_1196_n2255, mult_x_1196_n2254,
         mult_x_1196_n2253, mult_x_1196_n2252, mult_x_1196_n2251,
         mult_x_1196_n2250, mult_x_1196_n2249, mult_x_1196_n2247,
         mult_x_1196_n2246, mult_x_1196_n2245, mult_x_1196_n2244,
         mult_x_1196_n2242, mult_x_1196_n2241, mult_x_1196_n2239,
         mult_x_1196_n2238, mult_x_1196_n2235, mult_x_1196_n2233,
         mult_x_1196_n2232, mult_x_1196_n2231, mult_x_1196_n2230,
         mult_x_1196_n2229, mult_x_1196_n2228, mult_x_1196_n2227,
         mult_x_1196_n2226, mult_x_1196_n2225, mult_x_1196_n2223,
         mult_x_1196_n2222, mult_x_1196_n2220, mult_x_1196_n2219,
         mult_x_1196_n2218, mult_x_1196_n2213, mult_x_1196_n2211,
         mult_x_1196_n2210, mult_x_1196_n2209, mult_x_1196_n2207,
         mult_x_1196_n2206, mult_x_1196_n2199, mult_x_1196_n2197,
         mult_x_1196_n2196, mult_x_1196_n2195, mult_x_1196_n2194,
         mult_x_1196_n2190, mult_x_1196_n2186, mult_x_1196_n2185,
         mult_x_1196_n2183, mult_x_1196_n2182, mult_x_1196_n2181,
         mult_x_1196_n2180, mult_x_1196_n2178, mult_x_1196_n2177,
         mult_x_1196_n2173, mult_x_1196_n2172, mult_x_1196_n2171,
         mult_x_1196_n2170, mult_x_1196_n2169, mult_x_1196_n2168,
         mult_x_1196_n2167, mult_x_1196_n2166, mult_x_1196_n2165,
         mult_x_1196_n2164, mult_x_1196_n2163, mult_x_1196_n2162,
         mult_x_1196_n2161, mult_x_1196_n2160, mult_x_1196_n2158,
         mult_x_1196_n2157, mult_x_1196_n2156, mult_x_1196_n2155,
         mult_x_1196_n2154, mult_x_1196_n2153, mult_x_1196_n2152,
         mult_x_1196_n2151, mult_x_1196_n2150, mult_x_1196_n2149,
         mult_x_1196_n2148, mult_x_1196_n2146, mult_x_1196_n2143,
         mult_x_1196_n2142, mult_x_1196_n2141, mult_x_1196_n2140,
         mult_x_1196_n2139, mult_x_1196_n2138, mult_x_1196_n2137,
         mult_x_1196_n2136, mult_x_1196_n2135, mult_x_1196_n2134,
         mult_x_1196_n2133, mult_x_1196_n2132, mult_x_1196_n2130,
         mult_x_1196_n2129, mult_x_1196_n2128, mult_x_1196_n2127,
         mult_x_1196_n2091, mult_x_1196_n2090, mult_x_1196_n2089,
         mult_x_1196_n2088, mult_x_1196_n2087, mult_x_1196_n2086,
         mult_x_1196_n2084, mult_x_1196_n2083, mult_x_1196_n2082,
         mult_x_1196_n2080, mult_x_1196_n2078, mult_x_1196_n2077,
         mult_x_1196_n2075, mult_x_1196_n2071, mult_x_1196_n2070,
         mult_x_1196_n2069, mult_x_1196_n2068, mult_x_1196_n2067,
         mult_x_1196_n2065, mult_x_1196_n2064, mult_x_1196_n2063,
         mult_x_1196_n2062, mult_x_1196_n2061, mult_x_1196_n2060,
         mult_x_1196_n2059, mult_x_1196_n2058, mult_x_1196_n2057,
         mult_x_1196_n2055, mult_x_1196_n2054, mult_x_1196_n2053,
         mult_x_1196_n2052, mult_x_1196_n2051, mult_x_1196_n2050,
         mult_x_1196_n2049, mult_x_1196_n2048, mult_x_1196_n2046,
         mult_x_1196_n2045, mult_x_1196_n2044, mult_x_1196_n2043,
         mult_x_1196_n2040, mult_x_1196_n2037, mult_x_1196_n2035,
         mult_x_1196_n2034, mult_x_1196_n2031, mult_x_1196_n2030,
         mult_x_1196_n2029, mult_x_1196_n2027, mult_x_1196_n2024,
         mult_x_1196_n2022, mult_x_1196_n2018, mult_x_1196_n2013,
         mult_x_1196_n2012, mult_x_1196_n2010, mult_x_1196_n2009,
         mult_x_1196_n2008, mult_x_1196_n2006, mult_x_1196_n2005,
         mult_x_1196_n2004, mult_x_1196_n2002, mult_x_1196_n2001,
         mult_x_1196_n2000, mult_x_1196_n1995, mult_x_1196_n1994,
         mult_x_1196_n1991, mult_x_1196_n1989, mult_x_1196_n1985,
         mult_x_1196_n1984, mult_x_1196_n1983, mult_x_1196_n1982,
         mult_x_1196_n1981, mult_x_1196_n1979, mult_x_1196_n1976,
         mult_x_1196_n1975, mult_x_1196_n1974, mult_x_1196_n1973,
         mult_x_1196_n1972, mult_x_1196_n1969, mult_x_1196_n1968,
         mult_x_1196_n1967, mult_x_1196_n1966, mult_x_1196_n1965,
         mult_x_1196_n1964, mult_x_1196_n1963, mult_x_1196_n1962,
         mult_x_1196_n1961, mult_x_1196_n1959, mult_x_1196_n1957,
         mult_x_1196_n1956, mult_x_1196_n1955, mult_x_1196_n1954,
         mult_x_1196_n1949, mult_x_1196_n1948, mult_x_1196_n1946,
         mult_x_1196_n1945, mult_x_1196_n1944, mult_x_1196_n1943,
         mult_x_1196_n1940, mult_x_1196_n1937, mult_x_1196_n1936,
         mult_x_1196_n1934, mult_x_1196_n1932, mult_x_1196_n1931,
         mult_x_1196_n1929, mult_x_1196_n1928, mult_x_1196_n1927,
         mult_x_1196_n1924, mult_x_1196_n1922, mult_x_1196_n1921,
         mult_x_1196_n1918, mult_x_1196_n1916, mult_x_1196_n1913,
         mult_x_1196_n1912, mult_x_1196_n1911, mult_x_1196_n1906,
         mult_x_1196_n1905, mult_x_1196_n1904, mult_x_1196_n1903,
         mult_x_1196_n1902, mult_x_1196_n1901, mult_x_1196_n1900,
         mult_x_1196_n1899, mult_x_1196_n1891, mult_x_1196_n1889,
         mult_x_1196_n1887, mult_x_1196_n1884, mult_x_1196_n1883,
         mult_x_1196_n1882, mult_x_1196_n1879, mult_x_1196_n1877,
         mult_x_1196_n1876, mult_x_1196_n1872, mult_x_1196_n1870,
         mult_x_1196_n1869, mult_x_1196_n1868, mult_x_1196_n1866,
         mult_x_1196_n1864, mult_x_1196_n1863, mult_x_1196_n1862,
         mult_x_1196_n1860, mult_x_1196_n1859, mult_x_1196_n1858,
         mult_x_1196_n1852, mult_x_1196_n1847, mult_x_1196_n1846,
         mult_x_1196_n1845, mult_x_1196_n1844, mult_x_1196_n1840,
         mult_x_1196_n1839, mult_x_1196_n1838, mult_x_1196_n1837,
         mult_x_1196_n1836, mult_x_1196_n1835, mult_x_1196_n1834,
         mult_x_1196_n1833, mult_x_1196_n1832, mult_x_1196_n1830,
         mult_x_1196_n1828, mult_x_1196_n1825, mult_x_1196_n1822,
         mult_x_1196_n1820, mult_x_1196_n1819, mult_x_1196_n1818,
         mult_x_1196_n1817, mult_x_1196_n1814, mult_x_1196_n1813,
         mult_x_1196_n1812, mult_x_1196_n1811, mult_x_1196_n1810,
         mult_x_1196_n1809, mult_x_1196_n1807, mult_x_1196_n1806,
         mult_x_1196_n1805, mult_x_1196_n1802, mult_x_1196_n1801,
         mult_x_1196_n1797, mult_x_1196_n1796, mult_x_1196_n1794,
         mult_x_1196_n1793, mult_x_1196_n1792, mult_x_1196_n1791,
         mult_x_1196_n1790, mult_x_1196_n1789, mult_x_1196_n1788,
         mult_x_1196_n1787, mult_x_1196_n1783, mult_x_1196_n1781,
         mult_x_1196_n1780, mult_x_1196_n1777, mult_x_1196_n1775,
         mult_x_1196_n1772, mult_x_1196_n1771, mult_x_1196_n1767,
         mult_x_1196_n1766, mult_x_1196_n1765, mult_x_1196_n1763,
         mult_x_1196_n1762, mult_x_1196_n1760, mult_x_1196_n1757,
         mult_x_1196_n1756, mult_x_1196_n1755, mult_x_1196_n1754,
         mult_x_1196_n1753, mult_x_1196_n1751, mult_x_1196_n1750,
         mult_x_1196_n1749, mult_x_1196_n1748, mult_x_1196_n1747,
         mult_x_1196_n1745, mult_x_1196_n1744, mult_x_1196_n1739,
         mult_x_1196_n1738, mult_x_1196_n1737, mult_x_1196_n1736,
         mult_x_1196_n1735, mult_x_1196_n1734, mult_x_1196_n1733,
         mult_x_1196_n1732, mult_x_1196_n1730, mult_x_1196_n1727,
         mult_x_1196_n1721, mult_x_1196_n1719, mult_x_1196_n1718,
         mult_x_1196_n1712, mult_x_1196_n1711, mult_x_1196_n1709,
         mult_x_1196_n1708, mult_x_1196_n1707, mult_x_1196_n1706,
         mult_x_1196_n1705, mult_x_1196_n1704, mult_x_1196_n1703,
         mult_x_1196_n1699, mult_x_1196_n1697, mult_x_1196_n1696,
         mult_x_1196_n1695, mult_x_1196_n1694, mult_x_1196_n1691,
         mult_x_1196_n1690, mult_x_1196_n1689, mult_x_1196_n1686,
         mult_x_1196_n1685, mult_x_1196_n1684, mult_x_1196_n1681,
         mult_x_1196_n1678, mult_x_1196_n1677, mult_x_1196_n1676,
         mult_x_1196_n1675, mult_x_1196_n1674, mult_x_1196_n1672,
         mult_x_1196_n1671, mult_x_1196_n1670, mult_x_1196_n1669,
         mult_x_1196_n1668, mult_x_1196_n1666, mult_x_1196_n1665,
         mult_x_1196_n1662, mult_x_1196_n1661, mult_x_1196_n1660,
         mult_x_1196_n1659, mult_x_1196_n1658, mult_x_1196_n1653,
         mult_x_1196_n1650, mult_x_1196_n1648, mult_x_1196_n1643,
         mult_x_1196_n1642, mult_x_1196_n1641, mult_x_1196_n1640,
         mult_x_1196_n1639, mult_x_1196_n1638, mult_x_1196_n1637,
         mult_x_1196_n1636, mult_x_1196_n1633, mult_x_1196_n1630,
         mult_x_1196_n1629, mult_x_1196_n1627, mult_x_1196_n1625,
         mult_x_1196_n1624, mult_x_1196_n1620, mult_x_1196_n1619,
         mult_x_1196_n1614, mult_x_1196_n1613, mult_x_1196_n1612,
         mult_x_1196_n1611, mult_x_1196_n1610, mult_x_1196_n1609,
         mult_x_1196_n1606, mult_x_1196_n1605, mult_x_1196_n1604,
         mult_x_1196_n1603, mult_x_1196_n1602, mult_x_1196_n1599,
         mult_x_1196_n1597, mult_x_1196_n1596, mult_x_1196_n1593,
         mult_x_1196_n1591, mult_x_1196_n1586, mult_x_1196_n1583,
         mult_x_1196_n1581, mult_x_1196_n1580, mult_x_1196_n1579,
         mult_x_1196_n1578, mult_x_1196_n1577, mult_x_1196_n1574,
         mult_x_1196_n1572, mult_x_1196_n1571, mult_x_1196_n1570,
         mult_x_1196_n1569, mult_x_1196_n1568, mult_x_1196_n1567,
         mult_x_1196_n1566, mult_x_1196_n1565, mult_x_1196_n1563,
         mult_x_1196_n1561, mult_x_1196_n1559, mult_x_1196_n1557,
         mult_x_1196_n1556, mult_x_1196_n1554, mult_x_1196_n1553,
         mult_x_1196_n1552, mult_x_1196_n1548, mult_x_1196_n1544,
         mult_x_1196_n1542, mult_x_1196_n1538, mult_x_1196_n1537,
         mult_x_1196_n1536, mult_x_1196_n1535, mult_x_1196_n1534,
         mult_x_1196_n1532, mult_x_1196_n1531, mult_x_1196_n1528,
         mult_x_1196_n1527, mult_x_1196_n1526, mult_x_1196_n1525,
         mult_x_1196_n1524, mult_x_1196_n1522, mult_x_1196_n1520,
         mult_x_1196_n1517, mult_x_1196_n1516, mult_x_1196_n1512,
         mult_x_1196_n1510, mult_x_1196_n1509, mult_x_1196_n1504,
         mult_x_1196_n1501, mult_x_1196_n1500, mult_x_1196_n1497,
         mult_x_1196_n1496, mult_x_1196_n1495, mult_x_1196_n1494,
         mult_x_1196_n1493, mult_x_1196_n1490, mult_x_1196_n1488,
         mult_x_1196_n1487, mult_x_1196_n1486, mult_x_1196_n1484,
         mult_x_1196_n1483, mult_x_1196_n1480, mult_x_1196_n1479,
         mult_x_1196_n1477, mult_x_1196_n1476, mult_x_1196_n1475,
         mult_x_1196_n1474, mult_x_1196_n1473, mult_x_1196_n1472,
         mult_x_1196_n1471, mult_x_1196_n1467, mult_x_1196_n1463,
         mult_x_1196_n1460, mult_x_1196_n1459, mult_x_1196_n1455,
         mult_x_1196_n1454, mult_x_1196_n1452, mult_x_1196_n1448,
         mult_x_1196_n1447, mult_x_1196_n1446, mult_x_1196_n1443,
         mult_x_1196_n1442, mult_x_1196_n1441, mult_x_1196_n1440,
         mult_x_1196_n1439, mult_x_1196_n1438, mult_x_1196_n1435,
         mult_x_1196_n1434, mult_x_1196_n1433, mult_x_1196_n1427,
         mult_x_1196_n1426, mult_x_1196_n1425, mult_x_1196_n1424,
         mult_x_1196_n1423, mult_x_1196_n1422, mult_x_1196_n1421,
         mult_x_1196_n1420, mult_x_1196_n1419, mult_x_1196_n1418,
         mult_x_1196_n1417, mult_x_1196_n1416, mult_x_1196_n1415,
         mult_x_1196_n1411, mult_x_1196_n1409, mult_x_1196_n1408,
         mult_x_1196_n1407, mult_x_1196_n1406, mult_x_1196_n1405,
         mult_x_1196_n1404, mult_x_1196_n1400, mult_x_1196_n1397,
         mult_x_1196_n1395, mult_x_1196_n1394, mult_x_1196_n1392,
         mult_x_1196_n1391, mult_x_1196_n1387, mult_x_1196_n1386,
         mult_x_1196_n1385, mult_x_1196_n1383, mult_x_1196_n1381,
         mult_x_1196_n1380, mult_x_1196_n1379, mult_x_1196_n1378,
         mult_x_1196_n1376, mult_x_1196_n1374, mult_x_1196_n1373,
         mult_x_1196_n1372, mult_x_1196_n1371, mult_x_1196_n1369,
         mult_x_1196_n1368, mult_x_1196_n1367, mult_x_1196_n1365,
         mult_x_1196_n1364, mult_x_1196_n1363, mult_x_1196_n1362,
         mult_x_1196_n1361, mult_x_1196_n1359, mult_x_1196_n1358,
         mult_x_1196_n1357, mult_x_1196_n1355, mult_x_1196_n1353,
         mult_x_1196_n1352, mult_x_1196_n1351, mult_x_1196_n1350,
         mult_x_1196_n1349, mult_x_1196_n1348, mult_x_1196_n1346,
         mult_x_1196_n1345, mult_x_1196_n1344, mult_x_1196_n1341,
         mult_x_1196_n1340, mult_x_1196_n1336, mult_x_1196_n1334,
         mult_x_1196_n1331, mult_x_1196_n1329, mult_x_1196_n1328,
         mult_x_1196_n1327, mult_x_1196_n1323, mult_x_1196_n1322,
         mult_x_1196_n1321, mult_x_1196_n1320, mult_x_1196_n1318,
         mult_x_1196_n1317, mult_x_1196_n1316, mult_x_1196_n1315,
         mult_x_1196_n1314, mult_x_1196_n1312, mult_x_1196_n1310,
         mult_x_1196_n1308, mult_x_1196_n1305, mult_x_1196_n1299,
         mult_x_1196_n1298, mult_x_1196_n1297, mult_x_1196_n1295,
         mult_x_1196_n1294, mult_x_1196_n1288, mult_x_1196_n1286,
         mult_x_1196_n1285, mult_x_1196_n1284, mult_x_1196_n1283,
         mult_x_1196_n1282, mult_x_1196_n1281, mult_x_1196_n1280,
         mult_x_1196_n1279, mult_x_1196_n1274, mult_x_1196_n1273,
         mult_x_1196_n1271, mult_x_1196_n1270, mult_x_1196_n1269,
         mult_x_1196_n1268, mult_x_1196_n1267, mult_x_1196_n1265,
         mult_x_1196_n1264, mult_x_1196_n1263, mult_x_1196_n1262,
         mult_x_1196_n1260, mult_x_1196_n1259, mult_x_1196_n1255,
         mult_x_1196_n1253, mult_x_1196_n1252, mult_x_1196_n1251,
         mult_x_1196_n1250, mult_x_1196_n1249, mult_x_1196_n1248,
         mult_x_1196_n1247, mult_x_1196_n1246, mult_x_1196_n1245,
         mult_x_1196_n1243, mult_x_1196_n1242, mult_x_1196_n1240,
         mult_x_1196_n1239, mult_x_1196_n1237, mult_x_1196_n1235,
         mult_x_1196_n1234, mult_x_1196_n1230, mult_x_1196_n1229,
         mult_x_1196_n1225, mult_x_1196_n1223, mult_x_1196_n1222,
         mult_x_1196_n1221, mult_x_1196_n1220, mult_x_1196_n1219,
         mult_x_1196_n1218, mult_x_1196_n1217, mult_x_1196_n1216,
         mult_x_1196_n1214, mult_x_1196_n1212, mult_x_1196_n1210,
         mult_x_1196_n1209, mult_x_1196_n1204, mult_x_1196_n1203,
         mult_x_1196_n1202, mult_x_1196_n1200, mult_x_1196_n1198,
         mult_x_1196_n1197, mult_x_1196_n1196, mult_x_1196_n1194,
         mult_x_1196_n1191, mult_x_1196_n1190, mult_x_1196_n1188,
         mult_x_1196_n1187, mult_x_1196_n1186, mult_x_1196_n1185,
         mult_x_1196_n1184, mult_x_1196_n1183, mult_x_1196_n1178,
         mult_x_1196_n1177, mult_x_1196_n1175, mult_x_1196_n1173,
         mult_x_1196_n1172, mult_x_1196_n1169, mult_x_1196_n1168,
         mult_x_1196_n1167, mult_x_1196_n1166, mult_x_1196_n1163,
         mult_x_1196_n1162, mult_x_1196_n1161, mult_x_1196_n1160,
         mult_x_1196_n1159, mult_x_1196_n1158, mult_x_1196_n1156,
         mult_x_1196_n1154, mult_x_1196_n1153, mult_x_1196_n1152,
         mult_x_1196_n1148, mult_x_1196_n1147, mult_x_1196_n1145,
         mult_x_1196_n1144, mult_x_1196_n1142, mult_x_1196_n1141,
         mult_x_1196_n1140, mult_x_1196_n1139, mult_x_1196_n1136,
         mult_x_1196_n1135, mult_x_1196_n1134, mult_x_1196_n1133,
         mult_x_1196_n1131, mult_x_1196_n1130, mult_x_1196_n1129,
         mult_x_1196_n1128, mult_x_1196_n1127, mult_x_1196_n1126,
         mult_x_1196_n1125, mult_x_1196_n1124, mult_x_1196_n1122,
         mult_x_1196_n1119, mult_x_1196_n1117, mult_x_1196_n1113,
         mult_x_1196_n1112, mult_x_1196_n1110, mult_x_1196_n1105,
         mult_x_1196_n1104, mult_x_1196_n1103, mult_x_1196_n1102,
         mult_x_1196_n1101, mult_x_1196_n1100, mult_x_1196_n1099,
         mult_x_1196_n1098, mult_x_1196_n1097, mult_x_1196_n1096,
         mult_x_1196_n1095, mult_x_1196_n1094, mult_x_1196_n1093,
         mult_x_1196_n1092, mult_x_1196_n1091, mult_x_1196_n1090,
         mult_x_1196_n1089, mult_x_1196_n1088, mult_x_1196_n1086,
         mult_x_1196_n1084, mult_x_1196_n1083, mult_x_1196_n1081,
         mult_x_1196_n1080, mult_x_1196_n1078, mult_x_1196_n1077,
         mult_x_1196_n1076, mult_x_1196_n1075, mult_x_1196_n1074,
         mult_x_1196_n1072, mult_x_1196_n1069, mult_x_1196_n1068,
         mult_x_1196_n1067, mult_x_1196_n1066, mult_x_1196_n1064,
         mult_x_1196_n1063, mult_x_1196_n1062, mult_x_1196_n1061,
         mult_x_1196_n1059, mult_x_1196_n1058, mult_x_1196_n1057,
         mult_x_1196_n1055, mult_x_1196_n1054, mult_x_1196_n1053,
         mult_x_1196_n1052, mult_x_1196_n1050, mult_x_1196_n1049,
         mult_x_1196_n1048, mult_x_1196_n1047, mult_x_1196_n1046,
         mult_x_1196_n1045, mult_x_1196_n1044, mult_x_1196_n1043,
         mult_x_1196_n1042, mult_x_1196_n1039, mult_x_1196_n1037,
         mult_x_1196_n1036, mult_x_1196_n1034, mult_x_1196_n1033,
         mult_x_1196_n1032, mult_x_1196_n1029, mult_x_1196_n1028,
         mult_x_1196_n1027, mult_x_1196_n1025, mult_x_1196_n1023,
         mult_x_1196_n1022, mult_x_1196_n1021, mult_x_1196_n1020,
         mult_x_1196_n1017, mult_x_1196_n1016, mult_x_1196_n1015,
         mult_x_1196_n1014, mult_x_1196_n1013, mult_x_1196_n1011,
         mult_x_1196_n1010, mult_x_1196_n1009, mult_x_1196_n1006,
         mult_x_1196_n1005, mult_x_1196_n1004, mult_x_1196_n1002,
         mult_x_1196_n998, mult_x_1196_n997, mult_x_1196_n995,
         mult_x_1196_n994, mult_x_1196_n993, mult_x_1196_n992,
         mult_x_1196_n991, mult_x_1196_n990, mult_x_1196_n989,
         mult_x_1196_n987, mult_x_1196_n986, mult_x_1196_n984,
         mult_x_1196_n982, mult_x_1196_n981, mult_x_1196_n979,
         mult_x_1196_n978, mult_x_1196_n976, mult_x_1196_n975,
         mult_x_1196_n972, mult_x_1196_n971, mult_x_1196_n970,
         mult_x_1196_n969, mult_x_1196_n968, mult_x_1196_n967,
         mult_x_1196_n966, mult_x_1196_n965, mult_x_1196_n964,
         mult_x_1196_n963, mult_x_1196_n962, mult_x_1196_n960,
         mult_x_1196_n958, mult_x_1196_n957, mult_x_1196_n955,
         mult_x_1196_n954, mult_x_1196_n953, mult_x_1196_n952,
         mult_x_1196_n951, mult_x_1196_n949, mult_x_1196_n948,
         mult_x_1196_n947, mult_x_1196_n946, mult_x_1196_n945,
         mult_x_1196_n944, mult_x_1196_n943, mult_x_1196_n940,
         mult_x_1196_n937, mult_x_1196_n933, mult_x_1196_n932,
         mult_x_1196_n929, mult_x_1196_n928, mult_x_1196_n927,
         mult_x_1196_n926, mult_x_1196_n925, mult_x_1196_n924,
         mult_x_1196_n921, mult_x_1196_n918, mult_x_1196_n915,
         mult_x_1196_n913, mult_x_1196_n912, mult_x_1196_n911,
         mult_x_1196_n910, mult_x_1196_n907, mult_x_1196_n905,
         mult_x_1196_n904, mult_x_1196_n902, mult_x_1196_n901,
         mult_x_1196_n900, mult_x_1196_n899, mult_x_1196_n898,
         mult_x_1196_n897, mult_x_1196_n896, mult_x_1196_n894,
         mult_x_1196_n893, mult_x_1196_n891, mult_x_1196_n890,
         mult_x_1196_n889, mult_x_1196_n888, mult_x_1196_n887,
         mult_x_1196_n886, mult_x_1196_n885, mult_x_1196_n884,
         mult_x_1196_n883, mult_x_1196_n882, mult_x_1196_n881,
         mult_x_1196_n878, mult_x_1196_n877, mult_x_1196_n875,
         mult_x_1196_n874, mult_x_1196_n873, mult_x_1196_n872,
         mult_x_1196_n871, mult_x_1196_n870, mult_x_1196_n869,
         mult_x_1196_n867, mult_x_1196_n866, mult_x_1196_n865,
         mult_x_1196_n864, mult_x_1196_n863, mult_x_1196_n862,
         mult_x_1196_n861, mult_x_1196_n860, mult_x_1196_n859,
         mult_x_1196_n858, mult_x_1196_n856, mult_x_1196_n855,
         mult_x_1196_n854, mult_x_1196_n853, mult_x_1196_n852,
         mult_x_1196_n851, mult_x_1196_n850, mult_x_1196_n849,
         mult_x_1196_n848, mult_x_1196_n847, mult_x_1196_n844,
         mult_x_1196_n843, mult_x_1196_n842, mult_x_1196_n840,
         mult_x_1196_n839, mult_x_1196_n837, mult_x_1196_n829,
         mult_x_1196_n825, mult_x_1196_n824, mult_x_1196_n821,
         mult_x_1196_n820, mult_x_1196_n819, mult_x_1196_n818,
         mult_x_1196_n816, mult_x_1196_n815, mult_x_1196_n814,
         mult_x_1196_n813, mult_x_1196_n812, mult_x_1196_n810,
         mult_x_1196_n808, mult_x_1196_n807, mult_x_1196_n806,
         mult_x_1196_n805, mult_x_1196_n804, mult_x_1196_n803,
         mult_x_1196_n802, mult_x_1196_n801, mult_x_1196_n800,
         mult_x_1196_n799, mult_x_1196_n798, mult_x_1196_n796,
         mult_x_1196_n795, mult_x_1196_n794, mult_x_1196_n793,
         mult_x_1196_n792, mult_x_1196_n791, mult_x_1196_n788,
         mult_x_1196_n787, mult_x_1196_n785, mult_x_1196_n784,
         mult_x_1196_n781, mult_x_1196_n775, mult_x_1196_n771,
         mult_x_1196_n770, mult_x_1196_n766, mult_x_1196_n765,
         mult_x_1196_n764, mult_x_1196_n761, mult_x_1196_n760,
         mult_x_1196_n759, mult_x_1196_n758, mult_x_1196_n756,
         mult_x_1196_n753, mult_x_1196_n752, mult_x_1196_n750,
         mult_x_1196_n748, mult_x_1196_n747, mult_x_1196_n744,
         mult_x_1196_n735, mult_x_1196_n734, mult_x_1196_n732,
         mult_x_1196_n730, mult_x_1196_n729, mult_x_1196_n728,
         mult_x_1196_n726, mult_x_1196_n724, mult_x_1196_n723,
         mult_x_1196_n721, mult_x_1196_n719, mult_x_1196_n718,
         mult_x_1196_n717, mult_x_1196_n716, mult_x_1196_n715,
         mult_x_1196_n714, mult_x_1196_n713, mult_x_1196_n712,
         mult_x_1196_n710, mult_x_1196_n709, mult_x_1196_n708,
         mult_x_1196_n707, mult_x_1196_n706, mult_x_1196_n704,
         mult_x_1196_n702, mult_x_1196_n701, mult_x_1196_n699,
         mult_x_1196_n697, mult_x_1196_n696, mult_x_1196_n695,
         mult_x_1196_n693, mult_x_1196_n692, mult_x_1196_n691,
         mult_x_1196_n690, mult_x_1196_n689, mult_x_1196_n688,
         mult_x_1196_n687, mult_x_1196_n684, mult_x_1196_n683,
         mult_x_1196_n682, mult_x_1196_n680, mult_x_1196_n678,
         mult_x_1196_n677, mult_x_1196_n676, mult_x_1196_n675,
         mult_x_1196_n674, mult_x_1196_n672, mult_x_1196_n668,
         mult_x_1196_n667, mult_x_1196_n664, mult_x_1196_n661,
         mult_x_1196_n660, mult_x_1196_n657, mult_x_1196_n655,
         mult_x_1196_n654, mult_x_1196_n653, mult_x_1196_n652,
         mult_x_1196_n651, mult_x_1196_n648, mult_x_1196_n646,
         mult_x_1196_n645, mult_x_1196_n644, mult_x_1196_n642,
         mult_x_1196_n641, mult_x_1196_n640, mult_x_1196_n639,
         mult_x_1196_n638, mult_x_1196_n637, mult_x_1196_n636,
         mult_x_1196_n629, mult_x_1196_n626, mult_x_1196_n623,
         mult_x_1196_n622, mult_x_1196_n617, mult_x_1196_n616,
         mult_x_1196_n615, mult_x_1196_n614, mult_x_1196_n613,
         mult_x_1196_n612, mult_x_1196_n611, mult_x_1196_n607,
         mult_x_1196_n606, mult_x_1196_n604, mult_x_1196_n603,
         mult_x_1196_n602, mult_x_1196_n599, mult_x_1196_n597,
         mult_x_1196_n596, mult_x_1196_n595, mult_x_1196_n594,
         mult_x_1196_n591, mult_x_1196_n590, mult_x_1196_n589,
         mult_x_1196_n588, mult_x_1196_n587, mult_x_1196_n586,
         mult_x_1196_n584, mult_x_1196_n582, mult_x_1196_n580,
         mult_x_1196_n579, mult_x_1196_n578, mult_x_1196_n577,
         mult_x_1196_n575, mult_x_1196_n570, mult_x_1196_n568,
         mult_x_1196_n566, mult_x_1196_n565, mult_x_1196_n564,
         mult_x_1196_n563, mult_x_1196_n561, mult_x_1196_n560,
         mult_x_1196_n559, mult_x_1196_n558, mult_x_1196_n557,
         mult_x_1196_n556, mult_x_1196_n555, mult_x_1196_n552,
         mult_x_1196_n550, mult_x_1196_n549, mult_x_1196_n548,
         mult_x_1196_n547, mult_x_1196_n546, mult_x_1196_n545,
         mult_x_1196_n543, mult_x_1196_n542, mult_x_1196_n541,
         mult_x_1196_n540, mult_x_1196_n539, mult_x_1196_n535,
         mult_x_1196_n534, mult_x_1196_n533, mult_x_1196_n532,
         mult_x_1196_n531, mult_x_1196_n530, mult_x_1196_n529,
         mult_x_1196_n526, mult_x_1196_n525, mult_x_1196_n524,
         mult_x_1196_n520, mult_x_1196_n519, mult_x_1196_n518,
         mult_x_1196_n517, mult_x_1196_n516, mult_x_1196_n515,
         mult_x_1196_n514, mult_x_1196_n513, mult_x_1196_n507,
         mult_x_1196_n506, mult_x_1196_n505, mult_x_1196_n504,
         mult_x_1196_n496, mult_x_1196_n495, mult_x_1196_n494,
         mult_x_1196_n491, mult_x_1196_n489, mult_x_1196_n488,
         mult_x_1196_n487, mult_x_1196_n486, mult_x_1196_n485,
         mult_x_1196_n484, mult_x_1196_n483, mult_x_1196_n482,
         mult_x_1196_n481, mult_x_1196_n480, mult_x_1196_n478,
         mult_x_1196_n477, mult_x_1196_n476, mult_x_1196_n475,
         mult_x_1196_n474, mult_x_1196_n473, mult_x_1196_n472,
         mult_x_1196_n470, mult_x_1196_n467, mult_x_1196_n466,
         mult_x_1196_n465, mult_x_1196_n464, mult_x_1196_n460,
         mult_x_1196_n457, mult_x_1196_n456, mult_x_1196_n455,
         mult_x_1196_n454, mult_x_1196_n453, mult_x_1196_n452,
         mult_x_1196_n451, mult_x_1196_n449, mult_x_1196_n445,
         mult_x_1196_n444, mult_x_1196_n443, mult_x_1196_n442,
         mult_x_1196_n434, mult_x_1196_n432, mult_x_1196_n430,
         mult_x_1196_n429, mult_x_1196_n428, mult_x_1196_n425,
         mult_x_1196_n423, mult_x_1196_n421, mult_x_1196_n420,
         mult_x_1196_n418, mult_x_1196_n416, mult_x_1196_n411,
         mult_x_1196_n407, mult_x_1196_n405, mult_x_1196_n398,
         mult_x_1196_n396, mult_x_1196_n394, mult_x_1196_n393,
         mult_x_1196_n392, mult_x_1196_n391, mult_x_1196_n390,
         mult_x_1196_n387, mult_x_1196_n386, mult_x_1196_n385,
         mult_x_1196_n379, mult_x_1196_n378, mult_x_1196_n377,
         mult_x_1196_n375, mult_x_1196_n368, mult_x_1196_n366,
         mult_x_1196_n364, mult_x_1196_n361, mult_x_1196_n360,
         mult_x_1196_n359, mult_x_1196_n358, mult_x_1196_n357,
         mult_x_1196_n356, mult_x_1196_n355, mult_x_1196_n354,
         mult_x_1196_n350, mult_x_1196_n348, mult_x_1196_n347,
         mult_x_1196_n343, mult_x_1196_n339, mult_x_1196_n335,
         mult_x_1196_n334, mult_x_1196_n333, mult_x_1196_n331,
         mult_x_1196_n330, mult_x_1196_n328, mult_x_1196_n324,
         mult_x_1196_n323, mult_x_1196_n317, mult_x_1196_n316,
         mult_x_1196_n315, mult_x_1196_n313, mult_x_1196_n312,
         mult_x_1196_n308, mult_x_1196_n306, mult_x_1196_n302,
         mult_x_1196_n301, mult_x_1196_n299, mult_x_1196_n298,
         mult_x_1196_n297, mult_x_1196_n296, mult_x_1196_n295,
         mult_x_1196_n294, mult_x_1196_n288, mult_x_1196_n282,
         mult_x_1196_n278, mult_x_1196_n277, mult_x_1196_n276,
         mult_x_1196_n275, mult_x_1196_n274, mult_x_1196_n272,
         mult_x_1196_n271, mult_x_1196_n270, mult_x_1196_n269,
         mult_x_1196_n268, mult_x_1196_n267, mult_x_1196_n266,
         mult_x_1196_n265, mult_x_1196_n264, mult_x_1196_n263,
         mult_x_1196_n262, mult_x_1196_n261, mult_x_1196_n258,
         mult_x_1196_n257, mult_x_1196_n256, mult_x_1196_n255,
         mult_x_1196_n254, mult_x_1196_n253, mult_x_1196_n251,
         mult_x_1196_n250, mult_x_1196_n249, mult_x_1196_n248,
         mult_x_1196_n247, mult_x_1196_n246, mult_x_1196_n245,
         mult_x_1196_n244, mult_x_1196_n243, mult_x_1196_n242,
         mult_x_1196_n241, mult_x_1196_n240, mult_x_1196_n239,
         mult_x_1196_n238, mult_x_1196_n237, mult_x_1196_n236,
         mult_x_1196_n233, mult_x_1196_n231, mult_x_1196_n230,
         mult_x_1196_n229, mult_x_1196_n228, mult_x_1196_n227,
         mult_x_1196_n226, mult_x_1196_n225, mult_x_1196_n224,
         mult_x_1196_n223, mult_x_1196_n135, mult_x_1196_n126, mult_x_1196_n99,
         mult_x_1196_n96, mult_x_1196_n72, mult_x_1196_n60, mult_x_1196_n39,
         mult_x_1196_n9, mult_x_1196_n6, DP_OP_1196_128_7433_n480,
         DP_OP_1196_128_7433_n479, DP_OP_1196_128_7433_n478,
         DP_OP_1196_128_7433_n477, DP_OP_1196_128_7433_n476,
         DP_OP_1196_128_7433_n475, DP_OP_1196_128_7433_n474,
         DP_OP_1196_128_7433_n456, DP_OP_1196_128_7433_n455,
         DP_OP_1196_128_7433_n454, DP_OP_1196_128_7433_n453,
         DP_OP_1196_128_7433_n452, DP_OP_1196_128_7433_n386,
         DP_OP_1196_128_7433_n385, DP_OP_1196_128_7433_n380,
         DP_OP_1196_128_7433_n378, DP_OP_1196_128_7433_n376,
         DP_OP_1196_128_7433_n374, DP_OP_1196_128_7433_n372,
         DP_OP_1196_128_7433_n370, DP_OP_1196_128_7433_n368,
         DP_OP_1196_128_7433_n367, DP_OP_1196_128_7433_n365,
         DP_OP_1196_128_7433_n361, DP_OP_1196_128_7433_n357,
         DP_OP_1196_128_7433_n355, DP_OP_1196_128_7433_n354,
         DP_OP_1196_128_7433_n353, DP_OP_1196_128_7433_n352,
         DP_OP_1196_128_7433_n351, DP_OP_1196_128_7433_n350,
         DP_OP_1196_128_7433_n348, DP_OP_1196_128_7433_n347,
         DP_OP_1196_128_7433_n346, DP_OP_1196_128_7433_n345,
         DP_OP_1196_128_7433_n339, DP_OP_1196_128_7433_n338,
         DP_OP_1196_128_7433_n337, DP_OP_1196_128_7433_n336,
         DP_OP_1196_128_7433_n334, DP_OP_1196_128_7433_n330,
         DP_OP_1196_128_7433_n329, DP_OP_1196_128_7433_n328,
         DP_OP_1196_128_7433_n327, DP_OP_1196_128_7433_n325,
         DP_OP_1196_128_7433_n319, DP_OP_1196_128_7433_n318,
         DP_OP_1196_128_7433_n317, DP_OP_1196_128_7433_n316,
         DP_OP_1196_128_7433_n315, DP_OP_1196_128_7433_n314,
         DP_OP_1196_128_7433_n313, DP_OP_1196_128_7433_n310,
         DP_OP_1196_128_7433_n308, DP_OP_1196_128_7433_n307,
         DP_OP_1196_128_7433_n306, DP_OP_1196_128_7433_n305,
         DP_OP_1196_128_7433_n304, DP_OP_1196_128_7433_n303,
         DP_OP_1196_128_7433_n302, DP_OP_1196_128_7433_n301,
         DP_OP_1196_128_7433_n299, DP_OP_1196_128_7433_n297,
         DP_OP_1196_128_7433_n296, DP_OP_1196_128_7433_n291,
         DP_OP_1196_128_7433_n290, DP_OP_1196_128_7433_n289,
         DP_OP_1196_128_7433_n288, DP_OP_1196_128_7433_n285,
         DP_OP_1196_128_7433_n284, DP_OP_1196_128_7433_n283,
         DP_OP_1196_128_7433_n280, DP_OP_1196_128_7433_n278,
         DP_OP_1196_128_7433_n277, DP_OP_1196_128_7433_n276,
         DP_OP_1196_128_7433_n275, DP_OP_1196_128_7433_n274,
         DP_OP_1196_128_7433_n273, DP_OP_1196_128_7433_n272,
         DP_OP_1196_128_7433_n271, DP_OP_1196_128_7433_n269,
         DP_OP_1196_128_7433_n267, DP_OP_1196_128_7433_n266,
         DP_OP_1196_128_7433_n264, DP_OP_1196_128_7433_n263,
         DP_OP_1196_128_7433_n262, DP_OP_1196_128_7433_n261,
         DP_OP_1196_128_7433_n260, DP_OP_1196_128_7433_n259,
         DP_OP_1196_128_7433_n258, DP_OP_1196_128_7433_n257,
         DP_OP_1196_128_7433_n254, DP_OP_1196_128_7433_n252,
         DP_OP_1196_128_7433_n251, DP_OP_1196_128_7433_n250,
         DP_OP_1196_128_7433_n249, DP_OP_1196_128_7433_n248,
         DP_OP_1196_128_7433_n247, DP_OP_1196_128_7433_n246,
         DP_OP_1196_128_7433_n245, DP_OP_1196_128_7433_n243,
         DP_OP_1196_128_7433_n241, DP_OP_1196_128_7433_n240,
         DP_OP_1196_128_7433_n239, DP_OP_1196_128_7433_n238,
         DP_OP_1196_128_7433_n235, DP_OP_1196_128_7433_n234,
         DP_OP_1196_128_7433_n233, DP_OP_1196_128_7433_n232,
         DP_OP_1196_128_7433_n224, DP_OP_1196_128_7433_n222,
         DP_OP_1196_128_7433_n221, DP_OP_1196_128_7433_n220,
         DP_OP_1196_128_7433_n219, DP_OP_1196_128_7433_n218,
         DP_OP_1196_128_7433_n217, DP_OP_1196_128_7433_n216,
         DP_OP_1196_128_7433_n215, DP_OP_1196_128_7433_n213,
         DP_OP_1196_128_7433_n211, DP_OP_1196_128_7433_n210,
         DP_OP_1196_128_7433_n208, DP_OP_1196_128_7433_n207,
         DP_OP_1196_128_7433_n206, DP_OP_1196_128_7433_n205,
         DP_OP_1196_128_7433_n204, DP_OP_1196_128_7433_n203,
         DP_OP_1196_128_7433_n202, DP_OP_1196_128_7433_n201,
         DP_OP_1196_128_7433_n198, DP_OP_1196_128_7433_n196,
         DP_OP_1196_128_7433_n195, DP_OP_1196_128_7433_n194,
         DP_OP_1196_128_7433_n193, DP_OP_1196_128_7433_n192,
         DP_OP_1196_128_7433_n191, DP_OP_1196_128_7433_n190,
         DP_OP_1196_128_7433_n189, DP_OP_1196_128_7433_n187,
         DP_OP_1196_128_7433_n185, DP_OP_1196_128_7433_n184,
         DP_OP_1196_128_7433_n183, DP_OP_1196_128_7433_n180,
         DP_OP_1196_128_7433_n179, DP_OP_1196_128_7433_n178,
         DP_OP_1196_128_7433_n177, DP_OP_1196_128_7433_n176,
         DP_OP_1196_128_7433_n175, DP_OP_1196_128_7433_n174,
         DP_OP_1196_128_7433_n173, DP_OP_1196_128_7433_n168,
         DP_OP_1196_128_7433_n167, DP_OP_1196_128_7433_n166,
         DP_OP_1196_128_7433_n165, DP_OP_1196_128_7433_n164,
         DP_OP_1196_128_7433_n163, DP_OP_1196_128_7433_n162,
         DP_OP_1196_128_7433_n161, DP_OP_1196_128_7433_n157,
         DP_OP_1196_128_7433_n154, DP_OP_1196_128_7433_n153,
         DP_OP_1196_128_7433_n152, DP_OP_1196_128_7433_n151,
         DP_OP_1196_128_7433_n150, DP_OP_1196_128_7433_n149,
         DP_OP_1196_128_7433_n148, DP_OP_1196_128_7433_n147,
         DP_OP_1196_128_7433_n146, DP_OP_1196_128_7433_n145,
         DP_OP_1196_128_7433_n144, DP_OP_1196_128_7433_n143,
         DP_OP_1196_128_7433_n140, DP_OP_1196_128_7433_n139,
         DP_OP_1196_128_7433_n138, DP_OP_1196_128_7433_n137,
         DP_OP_1196_128_7433_n136, DP_OP_1196_128_7433_n135,
         DP_OP_1196_128_7433_n134, DP_OP_1196_128_7433_n131,
         DP_OP_1196_128_7433_n129, DP_OP_1196_128_7433_n128,
         DP_OP_1196_128_7433_n127, DP_OP_1196_128_7433_n126,
         DP_OP_1196_128_7433_n125, DP_OP_1196_128_7433_n124,
         DP_OP_1196_128_7433_n123, DP_OP_1196_128_7433_n122,
         DP_OP_1196_128_7433_n120, DP_OP_1196_128_7433_n118,
         DP_OP_1196_128_7433_n115, DP_OP_1196_128_7433_n114,
         DP_OP_1196_128_7433_n113, DP_OP_1196_128_7433_n112,
         DP_OP_1196_128_7433_n111, DP_OP_1196_128_7433_n110,
         DP_OP_1196_128_7433_n109, DP_OP_1196_128_7433_n108,
         DP_OP_1196_128_7433_n107, DP_OP_1196_128_7433_n106,
         DP_OP_1196_128_7433_n105, DP_OP_1196_128_7433_n104,
         DP_OP_1196_128_7433_n98, DP_OP_1196_128_7433_n97,
         DP_OP_1196_128_7433_n96, DP_OP_1196_128_7433_n95,
         DP_OP_1196_128_7433_n94, DP_OP_1196_128_7433_n93,
         DP_OP_1196_128_7433_n92, DP_OP_1196_128_7433_n91,
         DP_OP_1196_128_7433_n90, DP_OP_1196_128_7433_n87,
         DP_OP_1196_128_7433_n86, DP_OP_1196_128_7433_n85,
         DP_OP_1196_128_7433_n84, DP_OP_1196_128_7433_n80,
         DP_OP_1196_128_7433_n77, DP_OP_1196_128_7433_n76,
         DP_OP_1196_128_7433_n75, DP_OP_1196_128_7433_n74,
         DP_OP_1196_128_7433_n73, DP_OP_1196_128_7433_n72,
         DP_OP_1196_128_7433_n71, DP_OP_1196_128_7433_n70,
         DP_OP_1196_128_7433_n69, DP_OP_1196_128_7433_n68,
         DP_OP_1196_128_7433_n67, DP_OP_1196_128_7433_n66,
         DP_OP_1196_128_7433_n60, DP_OP_1196_128_7433_n57,
         DP_OP_1196_128_7433_n51, DP_OP_1196_128_7433_n50,
         DP_OP_1196_128_7433_n37, DP_OP_1196_128_7433_n36,
         DP_OP_1196_128_7433_n34, DP_OP_1196_128_7433_n33,
         DP_OP_1196_128_7433_n32, DP_OP_1196_128_7433_n31,
         DP_OP_1196_128_7433_n30, DP_OP_1196_128_7433_n29,
         DP_OP_1196_128_7433_n28, DP_OP_1196_128_7433_n27,
         DP_OP_1196_128_7433_n26, DP_OP_1196_128_7433_n24,
         DP_OP_1196_128_7433_n23, DP_OP_1196_128_7433_n22,
         DP_OP_1196_128_7433_n21, DP_OP_1196_128_7433_n20,
         DP_OP_1196_128_7433_n19, DP_OP_1196_128_7433_n18,
         DP_OP_1196_128_7433_n17, DP_OP_1196_128_7433_n16,
         DP_OP_1196_128_7433_n14, DP_OP_1196_128_7433_n12,
         DP_OP_1196_128_7433_n8, DP_OP_1196_128_7433_n7,
         DP_OP_1196_128_7433_n6, DP_OP_1196_128_7433_n4,
         DP_OP_1196_128_7433_n2, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24571, n24572, n24573, n24574, n24575, n24576,
         n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,
         n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,
         n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600,
         n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608,
         n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,
         n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624,
         n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
         n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640,
         n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648,
         n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,
         n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,
         n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672,
         n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680,
         n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,
         n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696,
         n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,
         n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,
         n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720,
         n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728,
         n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
         n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744,
         n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752,
         n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,
         n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,
         n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
         n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784,
         n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792,
         n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800,
         n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,
         n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816,
         n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824,
         n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,
         n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,
         n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848,
         n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856,
         n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864,
         n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
         n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,
         n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888,
         n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896,
         n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
         n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,
         n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,
         n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
         n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936,
         n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,
         n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,
         n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960,
         n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,
         n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
         n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
         n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
         n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
         n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,
         n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
         n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,
         n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032,
         n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,
         n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
         n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,
         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,
         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
         n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400,
         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,
         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512,
         n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,
         n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
         n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,
         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,
         n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
         n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
         n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
         n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,
         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
         n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
         n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,
         n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
         n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
         n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,
         n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
         n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,
         n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656,
         n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
         n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,
         n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
         n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704,
         n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
         n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,
         n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728,
         n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
         n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
         n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,
         n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
         n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
         n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776,
         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
         n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
         n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
         n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
         n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,
         n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
         n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
         n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848,
         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
         n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,
         n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
         n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,
         n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
         n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,
         n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
         n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
         n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920,
         n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
         n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,
         n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
         n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,
         n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
         n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,
         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
         n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,
         n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992,
         n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
         n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,
         n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016,
         n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024,
         n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
         n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
         n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,
         n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
         n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064,
         n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
         n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
         n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088,
         n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
         n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
         n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
         n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
         n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
         n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
         n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,
         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
         n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
         n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,
         n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
         n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
         n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
         n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
         n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
         n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240,
         n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
         n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256,
         n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264,
         n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,
         n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,
         n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
         n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,
         n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304,
         n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
         n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
         n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,
         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,
         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,
         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
         n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,
         n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,
         n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
         n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
         n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
         n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
         n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,
         n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
         n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,
         n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520,
         n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528,
         n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,
         n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544,
         n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
         n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
         n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,
         n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
         n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584,
         n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,
         n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600,
         n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
         n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616,
         n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,
         n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,
         n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,
         n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
         n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,
         n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664,
         n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672,
         n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
         n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688,
         n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696,
         n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
         n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712,
         n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
         n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,
         n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736,
         n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744,
         n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
         n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760,
         n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,
         n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,
         n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784,
         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
         n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,
         n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808,
         n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816,
         n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
         n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832,
         n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840,
         n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
         n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
         n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
         n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872,
         n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880,
         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
         n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
         n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904,
         n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912,
         n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
         n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928,
         n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
         n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,
         n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952,
         n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
         n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
         n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976,
         n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984,
         n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
         n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000,
         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
         n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,
         n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,
         n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
         n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
         n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048,
         n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056,
         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
         n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072,
         n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
         n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088,
         n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,
         n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
         n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
         n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120,
         n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
         n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
         n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144,
         n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
         n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
         n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168,
         n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
         n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192,
         n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200,
         n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,
         n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,
         n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224,
         n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232,
         n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240,
         n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
         n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256,
         n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264,
         n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272,
         n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,
         n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288,
         n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,
         n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
         n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,
         n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,
         n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328,
         n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,
         n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344,
         n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352,
         n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360,
         n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
         n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376,
         n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384,
         n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
         n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,
         n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408,
         n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416,
         n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
         n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
         n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,
         n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448,
         n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456,
         n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
         n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,
         n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,
         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,
         n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
         n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,
         n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,
         n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,
         n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528,
         n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536,
         n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544,
         n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552,
         n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560,
         n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568,
         n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576,
         n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584,
         n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592,
         n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600,
         n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608,
         n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
         n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624,
         n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632,
         n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640,
         n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648,
         n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656,
         n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664,
         n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672,
         n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680,
         n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688,
         n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696,
         n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704,
         n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712,
         n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720,
         n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728,
         n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736,
         n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744,
         n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752,
         n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760,
         n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768,
         n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776,
         n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784,
         n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792,
         n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800,
         n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808,
         n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816,
         n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824,
         n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832,
         n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840,
         n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848,
         n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856,
         n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864,
         n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872,
         n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880,
         n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888,
         n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896,
         n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904,
         n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912,
         n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920,
         n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928,
         n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936,
         n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944,
         n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952,
         n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960,
         n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968,
         n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976,
         n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984,
         n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992,
         n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000,
         n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008,
         n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016,
         n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024,
         n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032,
         n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040,
         n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048,
         n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056,
         n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064,
         n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072,
         n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080,
         n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088,
         n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096,
         n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104,
         n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112,
         n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120,
         n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128,
         n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136,
         n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144,
         n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152,
         n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160,
         n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168,
         n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176,
         n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184,
         n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192,
         n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200,
         n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208,
         n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216,
         n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224,
         n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232,
         n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240,
         n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248,
         n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256,
         n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264,
         n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272,
         n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280,
         n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288,
         n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296,
         n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304,
         n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312,
         n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320,
         n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328,
         n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336,
         n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344,
         n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352,
         n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360,
         n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368,
         n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376,
         n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
         n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392,
         n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400,
         n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408,
         n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416,
         n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424,
         n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432,
         n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440,
         n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448,
         n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
         n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464,
         n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472,
         n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480,
         n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488,
         n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496,
         n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504,
         n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512,
         n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520,
         n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528,
         n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536,
         n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544,
         n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552,
         n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560,
         n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568,
         n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576,
         n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584,
         n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
         n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600,
         n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608,
         n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616,
         n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624,
         n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632,
         n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640,
         n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648,
         n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656,
         n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
         n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672,
         n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680,
         n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688,
         n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696,
         n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704,
         n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712,
         n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720,
         n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728,
         n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
         n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744,
         n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752,
         n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760,
         n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768,
         n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776,
         n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784,
         n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792,
         n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800,
         n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808,
         n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816,
         n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824,
         n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832,
         n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840,
         n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848,
         n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856,
         n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864,
         n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872,
         n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
         n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888,
         n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896,
         n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904,
         n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912,
         n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920,
         n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928,
         n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936,
         n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
         n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952,
         n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960,
         n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968,
         n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976,
         n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
         n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992,
         n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000,
         n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008,
         n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016,
         n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024,
         n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032,
         n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040,
         n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048,
         n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056,
         n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064,
         n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072,
         n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
         n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088,
         n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096,
         n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104,
         n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112,
         n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120,
         n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128,
         n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136,
         n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144,
         n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
         n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160,
         n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168,
         n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176,
         n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184,
         n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192,
         n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200,
         n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208,
         n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216,
         n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224,
         n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232,
         n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240,
         n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248,
         n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256,
         n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264,
         n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272,
         n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280,
         n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288,
         n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
         n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304,
         n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
         n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320,
         n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328,
         n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336,
         n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344,
         n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352,
         n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360,
         n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368,
         n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376,
         n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384,
         n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392,
         n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400,
         n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408,
         n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416,
         n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424,
         n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432,
         n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
         n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448,
         n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456,
         n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464,
         n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472,
         n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480,
         n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488,
         n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496,
         n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
         n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
         n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520,
         n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528,
         n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536,
         n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544,
         n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552,
         n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560,
         n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568,
         n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576,
         n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
         n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592,
         n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600,
         n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608,
         n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616,
         n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624,
         n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632,
         n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640,
         n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648,
         n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656,
         n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664,
         n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672,
         n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680,
         n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688,
         n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696,
         n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704,
         n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712,
         n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720,
         n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
         n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736,
         n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744,
         n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752,
         n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760,
         n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768,
         n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776,
         n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784,
         n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792,
         n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
         n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808,
         n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816,
         n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824,
         n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832,
         n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840,
         n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848,
         n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856,
         n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864,
         n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
         n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880,
         n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888,
         n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896,
         n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904,
         n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912,
         n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920,
         n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928,
         n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936,
         n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
         n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952,
         n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960,
         n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968,
         n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976,
         n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984,
         n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992,
         n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000,
         n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008,
         n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
         n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024,
         n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032,
         n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040,
         n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048,
         n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056,
         n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064,
         n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072,
         n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080,
         n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088,
         n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096,
         n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104,
         n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112,
         n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120,
         n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128,
         n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136,
         n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144,
         n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152,
         n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
         n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168,
         n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176,
         n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184,
         n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192,
         n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200,
         n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208,
         n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216,
         n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224,
         n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
         n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240,
         n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248,
         n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256,
         n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264,
         n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272,
         n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280,
         n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288,
         n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296,
         n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
         n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312,
         n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320,
         n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328,
         n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336,
         n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344,
         n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352,
         n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360,
         n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368,
         n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
         n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384,
         n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
         n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400,
         n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408,
         n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416,
         n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424,
         n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432,
         n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440,
         n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448,
         n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456,
         n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464,
         n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472,
         n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480,
         n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488,
         n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496,
         n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504,
         n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512,
         n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520,
         n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528,
         n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536,
         n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544,
         n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552,
         n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560,
         n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568,
         n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576,
         n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584,
         n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592,
         n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600,
         n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608,
         n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616,
         n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624,
         n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632,
         n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640,
         n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648,
         n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656,
         n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664,
         n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672,
         n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680,
         n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688,
         n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696,
         n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704,
         n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712,
         n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720,
         n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728,
         n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736,
         n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744,
         n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752,
         n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760,
         n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768,
         n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776,
         n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784,
         n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792,
         n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800,
         n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808,
         n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816,
         n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824,
         n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832,
         n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840,
         n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848,
         n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856,
         n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864,
         n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872,
         n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880,
         n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888,
         n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896,
         n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904,
         n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912,
         n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920,
         n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928,
         n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936,
         n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944,
         n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952,
         n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960,
         n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968,
         n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976,
         n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984,
         n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992,
         n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000,
         n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008,
         n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016,
         n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024,
         n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032,
         n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040,
         n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048,
         n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056,
         n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064,
         n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072,
         n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080,
         n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088,
         n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096,
         n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104,
         n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112,
         n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
         n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128,
         n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136,
         n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
         n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152,
         n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160,
         n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168,
         n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176,
         n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
         n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192,
         n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200,
         n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208,
         n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216,
         n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224,
         n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232,
         n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240,
         n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248,
         n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256,
         n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264,
         n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272,
         n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280,
         n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288,
         n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296,
         n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304,
         n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312,
         n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320,
         n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328,
         n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336,
         n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344,
         n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352,
         n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360,
         n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368,
         n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376,
         n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384,
         n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392,
         n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400,
         n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408,
         n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416,
         n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424,
         n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432,
         n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440,
         n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448,
         n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456,
         n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464,
         n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472,
         n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480,
         n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488,
         n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496,
         n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504,
         n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512,
         n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520,
         n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528,
         n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536,
         n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544,
         n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552,
         n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560,
         n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568,
         n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576,
         n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584,
         n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592,
         n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600,
         n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608,
         n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
         n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624,
         n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632,
         n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640,
         n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648,
         n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656,
         n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664,
         n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672,
         n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680,
         n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688,
         n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696,
         n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704,
         n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712,
         n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720,
         n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728,
         n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736,
         n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744,
         n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752,
         n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760,
         n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768,
         n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776,
         n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784,
         n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792,
         n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800,
         n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808,
         n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816,
         n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824,
         n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832,
         n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840,
         n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848,
         n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856,
         n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864,
         n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872,
         n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880,
         n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888,
         n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896,
         n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904,
         n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912,
         n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920,
         n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928,
         n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936,
         n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944,
         n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952,
         n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960,
         n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968,
         n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976,
         n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984,
         n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992,
         n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000,
         n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008,
         n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016,
         n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024,
         n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032,
         n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040,
         n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048,
         n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056,
         n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064,
         n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072,
         n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080,
         n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088,
         n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096,
         n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104,
         n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112,
         n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120,
         n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128,
         n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136,
         n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144,
         n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152,
         n32153, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33061, n33062, n33063, n33064, n33065, n33066, n33067,
         n33068, n33069;
  wire   [1:0] irqo;
  wire   [46:0] apbi;
  wire   [33:0] u0_0_leon3x0_p0_divo;
  wire   [62:0] u0_0_leon3x0_p0_divi;
  wire   [63:0] u0_0_leon3x0_p0_mulo;
  wire   [48:0] u0_0_leon3x0_p0_muli;
  wire   [41:0] u0_0_leon3x0_p0_dci;
  wire   [89:0] u0_0_leon3x0_p0_ici;
  wire   [32:0] u0_0_leon3x0_p0_div0_b;
  wire   [32:0] u0_0_leon3x0_p0_div0_vaddin1;
  wire   [63:0] u0_0_leon3x0_p0_c0mmu_mcdi;
  wire   [31:0] u0_0_leon3x0_p0_c0mmu_mmudci;
  wire   [28:0] u0_0_leon3x0_p0_c0mmu_mcii;

  ASYNC_DFFHx1_ASAP7_75t_SL rst0_r_reg_0_ ( .D(n19002), .CLK(clk), .RESET(
        n18295), .SET(n4828), .QN(n4827) );
  ASYNC_DFFHx1_ASAP7_75t_SL rst0_r_reg_1_ ( .D(n4827), .CLK(clk), .RESET(n4828), .SET(n18295), .QN(rst0_r_1_) );
  ASYNC_DFFHx1_ASAP7_75t_SL rst0_r_reg_2_ ( .D(rst0_r_1_), .CLK(clk), .RESET(
        n18295), .SET(n4828), .QN(n4824) );
  ASYNC_DFFHx1_ASAP7_75t_SL rst0_r_reg_3_ ( .D(n4824), .CLK(clk), .RESET(n4828), .SET(n18295), .QN(rst0_r_3_) );
  ASYNC_DFFHx1_ASAP7_75t_SL rst0_r_reg_4_ ( .D(rst0_r_3_), .CLK(clk), .RESET(
        n18295), .SET(n4828), .QN(n4821) );
  ASYNC_DFFHx1_ASAP7_75t_SL rst0_rstoutl_reg ( .D(n11537), .CLK(clk), .RESET(
        n4828), .SET(n18295), .QN(rstn) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_rst_reg ( .D(n24694), .CLK(clk), .QN(
        n4818) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__0_ ( .D(n4816), .CLK(clk), .QN(
        ahbso_0__HRDATA__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__1_ ( .D(n4815), .CLK(clk), .QN(
        ahbso_0__HRDATA__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__2_ ( .D(n4814), .CLK(clk), .QN(
        ahbso_0__HRDATA__2_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__3_ ( .D(n4813), .CLK(clk), .QN(
        ahbso_0__HRDATA__3_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__4_ ( .D(n4812), .CLK(clk), .QN(
        ahbso_0__HRDATA__4_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__5_ ( .D(n4811), .CLK(clk), .QN(
        ahbso_0__HRDATA__5_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__6_ ( .D(n4810), .CLK(clk), .QN(
        ahbso_0__HRDATA__6_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__7_ ( .D(n4809), .CLK(clk), .QN(
        ahbso_0__HRDATA__7_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__8_ ( .D(n4808), .CLK(clk), .QN(
        ahbso_0__HRDATA__8_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__9_ ( .D(n4807), .CLK(clk), .QN(
        ahbso_0__HRDATA__9_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__10_ ( .D(n4806), .CLK(clk), .QN(
        ahbso_0__HRDATA__10_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__11_ ( .D(n4805), .CLK(clk), .QN(
        ahbso_0__HRDATA__11_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__12_ ( .D(n4804), .CLK(clk), .QN(
        ahbso_0__HRDATA__12_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__13_ ( .D(n4803), .CLK(clk), .QN(
        ahbso_0__HRDATA__13_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__14_ ( .D(n4802), .CLK(clk), .QN(
        ahbso_0__HRDATA__14_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__15_ ( .D(n4801), .CLK(clk), .QN(
        ahbso_0__HRDATA__15_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__16_ ( .D(n4800), .CLK(clk), .QN(
        ahbso_0__HRDATA__16_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__17_ ( .D(n4799), .CLK(clk), .QN(
        ahbso_0__HRDATA__17_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__18_ ( .D(n4798), .CLK(clk), .QN(
        ahbso_0__HRDATA__18_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__19_ ( .D(n4797), .CLK(clk), .QN(
        ahbso_0__HRDATA__19_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__20_ ( .D(n4796), .CLK(clk), .QN(
        ahbso_0__HRDATA__20_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__21_ ( .D(n4795), .CLK(clk), .QN(
        ahbso_0__HRDATA__21_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__22_ ( .D(n4794), .CLK(clk), .QN(
        ahbso_0__HRDATA__22_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__23_ ( .D(n4793), .CLK(clk), .QN(
        ahbso_0__HRDATA__23_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__24_ ( .D(n4792), .CLK(clk), .QN(
        ahbso_0__HRDATA__24_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__25_ ( .D(n4791), .CLK(clk), .QN(
        ahbso_0__HRDATA__25_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__26_ ( .D(n4790), .CLK(clk), .QN(
        ahbso_0__HRDATA__26_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__27_ ( .D(n4789), .CLK(clk), .QN(
        ahbso_0__HRDATA__27_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__28_ ( .D(n4788), .CLK(clk), .QN(
        ahbso_0__HRDATA__28_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__29_ ( .D(n4787), .CLK(clk), .QN(
        ahbso_0__HRDATA__29_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__30_ ( .D(n4786), .CLK(clk), .QN(
        ahbso_0__HRDATA__30_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_DATA__31_ ( .D(n4785), .CLK(clk), .QN(
        ahbso_0__HRDATA__31_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXF__0_ ( .D(n4784), .CLK(clk), .QN(
        uart1_v_RXF__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXF__1_ ( .D(n4783), .CLK(clk), .QN(
        uart1_r_RXF__1_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TICK_ ( .D(n33064), .CLK(clk), .QN(
        timer0_gpto_TICK__0_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_SCALER__7_ ( .D(n4780), .CLK(clk), .QN(
        timer0_r_SCALER__7_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__7_ ( .D(n4779), .CLK(clk), .QN(
        ahbso_1__HRDATA__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__7_ ( 
        .D(n4778), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__7_ ( 
        .D(n4777), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[11]) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__7_ ( .D(n17853), .CLK(clk), 
        .QN(n4775) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IRL__0__3_ ( .D(irqctrl0_v_IRL__0__3_), 
        .CLK(clk), .QN(n4774) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__31_ ( 
        .D(n4773), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__31_ ( 
        .D(n4772), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[35]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__31_ ( .D(n4771), .CLK(clk), .QN(
        apbi[31]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__31_ ( .D(
        timer0_v_TIMERS__1__VALUE__31_), .CLK(clk), .QN(n4770) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__IRQPEN_ ( .D(n4769), .CLK(clk), 
        .QN(timer0_vtimers_1__IRQPEN_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__4_ ( .D(n4768), .CLK(clk), .QN(
        ahbso_1__HRDATA__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__4_ ( 
        .D(n4767), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__4_ ( 
        .D(n4766), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[8]) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__4_ ( .D(n4764), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__4_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IRL__0__2_ ( .D(irqctrl0_v_IRL__0__2_), 
        .CLK(clk), .QN(n4763) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__TT__3_ ( .D(n4762), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__7_ ( .D(n4760), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[65]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__7_ ( .D(
        n4759), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[4]) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__7_ ( .D(n4758), .CLK(clk), .QN(
        ahb0_r_HADDR__7_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__5_ ( .D(n33066), .CLK(clk), .QN(
        ahb0_r_HRDATAS__5_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__12_ ( .D(n33066), .CLK(clk), .QN(
        ahb0_r_HRDATAS__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__12_ ( 
        .D(n4756), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__12_ ( 
        .D(n4755), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[16]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__12_ ( .D(n4754), .CLK(clk), .QN(
        apbi[12]) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__12_ ( .D(n4753), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__12_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IRL__0__1_ ( .D(irqctrl0_v_IRL__0__1_), 
        .CLK(clk), .QN(n4752) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__TT__1_ ( .D(n4751), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__5_ ( .D(n4749), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[63]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__5_ ( .D(
        n4748), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[2]) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__5_ ( .D(n4747), .CLK(clk), .QN(
        ahb0_r_HADDR__5_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAM__6_ ( .D(n4746), .CLK(clk), .QN(
        ahb0_r_HRDATAM__6_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAM__24_ ( .D(n4746), .CLK(clk), .QN(
        ahb0_r_HRDATAM__24_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAM__12_ ( .D(n4746), .CLK(clk), .QN(
        ahb0_r_HRDATAM__12_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAM__13_ ( .D(n4746), .CLK(clk), .QN(
        ahb0_r_HRDATAM__13_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAM__5_ ( .D(n4746), .CLK(clk), .QN(
        ahb0_r_HRDATAM__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__5_ ( 
        .D(n4745), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__5_ ( 
        .D(n4744), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[9]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__CHAIN_ ( .D(n17722), .CLK(clk), 
        .QN(n4742) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__30_ ( .D(
        timer0_v_TIMERS__1__VALUE__30_), .CLK(clk), .QN(n4741) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__30_ ( .D(n4740), .CLK(clk), .QN(
        ahbso_1__HRDATA__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__30_ ( 
        .D(n4739), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__30_ ( 
        .D(n4738), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[34]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__30_ ( .D(n4737), .CLK(clk), .QN(
        apbi[30]) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__14_ ( .D(n4736), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__14_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__14_ ( .D(n4735), .CLK(clk), .QN(
        irqctrl0_r_IPEND__14_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IRL__0__0_ ( .D(n4734), .CLK(clk), .QN(
        irqi_0__IRL__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__TT__0_ ( .D(n4733), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__4_ ( .D(n4731), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[62]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_BURST_ ( .D(n4730), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_BURST_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_HBURST__0_ ( .D(n4729), .CLK(clk), .QN(
        sr1_r_HBURST__0_) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_OEN_ ( .D(n4727), .CLK(clk), .RESET(
        n18295), .SET(n24695), .QN(oen) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_BSTATE__1_ ( .D(n4726), .CLK(clk), .QN(
        sr1_r_BSTATE__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WS__3_ ( .D(n4725), .CLK(clk), .QN(
        sr1_r_WS__3_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WS__1_ ( .D(n17422), .CLK(clk), .QN(n4724)
         );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WS__0_ ( .D(n4723), .CLK(clk), .QN(
        sr1_r_WS__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_READY_ ( .D(n4722), .CLK(clk), .QN(
        sr1_r_READY_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__19_ ( .D(n4719), .CLK(clk), .QN(
        apbi[45]) );
  SDFHx4_ASAP7_75t_SL apb0_r_reg_CFGSEL_ ( .D(n17251), .SI(n19002), .SE(n17252), .CLK(clk), .QN(apb0_r_CFGSEL_) );
  SDFHx4_ASAP7_75t_SL apb0_r_reg_PENABLE_ ( .D(apb0_N1148), .SI(n19002), .SE(
        n17243), .CLK(clk), .QN(apbi[46]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PSEL_ ( .D(n4716), .CLK(clk), .QN(
        apb0_r_PSEL_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RRADDR__4_ ( .D(n17455), .CLK(clk), .QN(
        n4715) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__6_ ( .D(n4714), .CLK(clk), .QN(
        ahbso_1__HRDATA__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__6_ ( 
        .D(n4713), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__6_ ( 
        .D(n4712), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[10]) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_FLOW_ ( .D(n4710), .CLK(clk), .QN(
        uart1_r_FLOW_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__9_ ( .D(n4709), .CLK(clk), .QN(
        uart1_r_TSHIFT__9_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__8_ ( .D(n24528), .CLK(clk), .QN(
        uart1_r_TSHIFT__8_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__7_ ( .D(n4707), .CLK(clk), .QN(
        uart1_r_TSHIFT__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__6_ ( .D(n24525), .CLK(clk), .QN(
        uart1_r_TSHIFT__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__5_ ( .D(n4705), .CLK(clk), .QN(
        uart1_r_TSHIFT__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__4_ ( .D(n24521), .CLK(clk), .QN(
        uart1_r_TSHIFT__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__3_ ( .D(n4703), .CLK(clk), .QN(
        uart1_r_TSHIFT__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__2_ ( .D(n4702), .CLK(clk), .QN(
        uart1_r_TSHIFT__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TPAR_ ( .D(n4700), .CLK(clk), .QN(
        uart1_r_TPAR_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSHIFT__0_ ( .D(n4699), .CLK(clk), .QN(
        uart1_r_TSHIFT__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXDB__0_ ( .D(n4698), .CLK(clk), .QN(
        uart1_v_RXDB__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXDB__1_ ( .D(n33065), .CLK(clk), .QN(
        uart1_r_RXDB__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSEMPTY_ ( .D(n4696), .CLK(clk), .QN(
        uart1_r_RSEMPTY_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__0__3_ ( .D(n4695), .CLK(clk), .QN(
        uart1_r_RHOLD__0__3_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__3_ ( .D(n4694), .CLK(clk), .QN(
        ahbso_1__HRDATA__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__3_ ( 
        .D(n4693), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__3_ ( 
        .D(n4692), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[7]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__IRQEN_ ( .D(n4690), .CLK(clk), 
        .QN(timer0_vtimers_1__IRQEN_) );
  SDFHx4_ASAP7_75t_SL irqctrl0_r_reg_IPEND__8_ ( .D(n15074), .SI(n19002), .SE(
        n15075), .CLK(clk), .QN(irqctrl0_r_IPEND__8_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__8_ ( .D(n4688), .CLK(clk), .QN(
        ahbso_1__HRDATA__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__8_ ( 
        .D(n4687), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__8_ ( 
        .D(n4686), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[12]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__8_ ( .D(n4685), .CLK(clk), .QN(
        apbi[8]) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_EXTCLKEN_ ( .D(n4684), .CLK(clk), .QN(
        uart1_r_EXTCLKEN_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TICK_ ( .D(n4683), .CLK(clk), .QN(
        uart1_r_TICK_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXF__2_ ( .D(n4681), .CLK(clk), .QN(
        uart1_r_RXF__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXF__3_ ( .D(n4679), .CLK(clk), .QN(
        uart1_r_RXF__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXF__4_ ( .D(n4677), .CLK(clk), .QN(
        uart1_r_RXF__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXTICK_ ( .D(n4676), .CLK(clk), .QN(
        uart1_r_RXTICK_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__0__2_ ( .D(n4675), .CLK(clk), .QN(
        uart1_r_RHOLD__0__2_) );
  SDFHx4_ASAP7_75t_SL apb0_r_reg_PRDATA__2_ ( .D(apb0_r_CFGSEL_), .SI(n19002), 
        .SE(n16838), .CLK(clk), .QN(ahbso_1__HRDATA__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__2_ ( 
        .D(n4673), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__2_ ( 
        .D(n4672), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[6]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__LOAD_ ( .D(n4670), .CLK(clk), 
        .QN(timer0_vtimers_1__LOAD_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__29_ ( .D(
        timer0_v_TIMERS__1__VALUE__29_), .CLK(clk), .QN(n4669) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__29_ ( .D(n4668), .CLK(clk), .QN(
        ahbso_1__HRDATA__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__29_ ( 
        .D(n4667), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__29_ ( 
        .D(n4666), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[33]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__29_ ( .D(n4665), .CLK(clk), .QN(
        apbi[29]) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__13_ ( .D(n4664), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__13_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__13_ ( .D(n4663), .CLK(clk), .QN(
        irqctrl0_r_IPEND__13_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__13_ ( .D(n4662), .CLK(clk), .QN(
        ahbso_1__HRDATA__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__13_ ( 
        .D(n4661), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__13_ ( .D(n4658), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__13_ ( .D(n4657), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__46_ ( .D(n4656), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[14]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__14_ ( .D(n4654), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__14_ ( .D(n4652), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[14]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__14_ ( 
        .D(n4651), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[47]) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_DEFSLV_ ( .D(n4650), .CLK(clk), .QN(
        ahb0_r_DEFSLV_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_WERR_ ( .D(n4649), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dco_WERR_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__TT__4_ ( .D(n4648), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__8_ ( .D(n4646), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[66]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__8_ ( .D(
        n4645), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[5]) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__8_ ( .D(n4644), .CLK(clk), .QN(
        ahb0_r_HADDR__8_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__17_ ( .D(n4643), .CLK(clk), .QN(
        ahb0_r_HRDATAS__17_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__16_ ( .D(n4643), .CLK(clk), .QN(
        ahb0_r_HRDATAS__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__16_ ( 
        .D(n4642), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__16_ ( .D(n4641), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__15_ ( 
        .D(n4638), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__15_ ( 
        .D(n4637), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[19]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__15_ ( .D(n4636), .CLK(clk), .QN(
        apbi[15]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__15_ ( .D(
        timer0_v_TIMERS__1__VALUE__15_), .CLK(clk), .QN(n4635) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__15_ ( .D(n4634), .CLK(clk), .QN(
        ahbso_1__HRDATA__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__15_ ( .D(n24437), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__25_ ( .D(n24509), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__25_ ( .D(n4629), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__25_ ( .D(n4627), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__25_ ( 
        .D(n4626), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[29]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__25_ ( .D(n4625), .CLK(clk), .QN(
        apbi[25]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__25_ ( .D(
        timer0_v_TIMERS__1__VALUE__25_), .CLK(clk), .QN(n4624) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__25_ ( .D(n4623), .CLK(clk), .QN(
        ahbso_1__HRDATA__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__25_ ( 
        .D(n4622), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__25_ ( .D(n4621), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__25_ ( .D(n4620), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__58_ ( .D(n4619), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[26]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__26_ ( .D(n4617), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__26_ ( 
        .D(n4616), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[30]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__26_ ( .D(n4615), .CLK(clk), .QN(
        apbi[26]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__26_ ( .D(
        timer0_v_TIMERS__1__VALUE__26_), .CLK(clk), .QN(n4614) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__26_ ( .D(n4613), .CLK(clk), .QN(
        ahbso_1__HRDATA__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__26_ ( 
        .D(n4612), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__26_ ( .D(n4609), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__26_ ( .D(n4607), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[57]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__25_ ( .D(n4605), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[56]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__57_ ( .D(n4604), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[25]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__25_ ( .D(n4602), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__13_ ( .D(n4601), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__25_ ( .D(n4599), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[83]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__25_ ( 
        .D(n31783), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[22]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__18_ ( .D(n4597), .CLK(clk), .QN(
        apbi[44]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__28_ ( .D(n4596), .CLK(clk), .QN(
        ahbso_1__HRDATA__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__28_ ( 
        .D(n4595), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__28_ ( .D(n4594), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__28_ ( .D(n4592), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__28_ ( .D(n4590), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[59]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__60_ ( .D(n4589), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[28]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__28_ ( .D(n4587), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__28_ ( .D(n4586), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__61_ ( .D(n4585), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[29]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__29_ ( .D(n4583), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__29_ ( .D(n4581), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__22_ ( .D(n4577), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__22_ ( 
        .D(n4576), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__22_ ( 
        .D(n4575), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[26]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__22_ ( .D(n4574), .CLK(clk), .QN(
        apbi[22]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__22_ ( .D(
        timer0_v_TIMERS__1__VALUE__22_), .CLK(clk), .QN(n4573) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__22_ ( .D(n4572), .CLK(clk), .QN(
        ahbso_1__HRDATA__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__WOVF_ ( .D(n4569), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__WOVF_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__TT__5_ ( .D(n4567), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__TT__5_ ( .D(n4565), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__TT__5_ ( .D(n4564), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__9_ ( .D(n4562), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[67]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__9_ ( .D(
        n4561), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[6]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__9_ ( .D(n4560), .CLK(clk), .QN(
        apbi[35]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__9_ ( .D(n4559), .CLK(clk), .QN(
        ahbso_1__HRDATA__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__9_ ( .D(n4557), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__9_ ( .D(n4555), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__9_ ( .D(n4554), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__42_ ( .D(n4553), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[10]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__10_ ( .D(n4551), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__10_ ( .D(n4549), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[10]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__10_ ( 
        .D(n4548), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__10_ ( 
        .D(n4547), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[43]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__10_ ( .D(n4546), .CLK(clk), .QN(
        apbi[36]) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXEN_ ( .D(n4545), .CLK(clk), .QN(
        uart1_uarto_RXEN_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSHIFT__7_ ( .D(n4544), .CLK(clk), .QN(
        uart1_r_RSHIFT__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSHIFT__6_ ( .D(n4543), .CLK(clk), .QN(
        uart1_r_RSHIFT__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSHIFT__5_ ( .D(n4542), .CLK(clk), .QN(
        uart1_r_RSHIFT__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSHIFT__4_ ( .D(n4541), .CLK(clk), .QN(
        uart1_r_RSHIFT__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSHIFT__3_ ( .D(n4540), .CLK(clk), .QN(
        uart1_r_RSHIFT__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSHIFT__2_ ( .D(n4539), .CLK(clk), .QN(
        uart1_r_RSHIFT__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSHIFT__1_ ( .D(n4538), .CLK(clk), .QN(
        uart1_r_RSHIFT__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__0__1_ ( .D(n4537), .CLK(clk), .QN(
        uart1_r_RHOLD__0__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__1_ ( 
        .D(n4535), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__1_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RESTART_ ( .D(n4532), .CLK(clk), .QN(timer0_vtimers_1__RESTART_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__27_ ( .D(
        timer0_v_TIMERS__1__VALUE__27_), .CLK(clk), .QN(n4531) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__27_ ( .D(n4530), .CLK(clk), .QN(
        ahbso_1__HRDATA__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__27_ ( 
        .D(n4529), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__27_ ( 
        .D(n4528), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[31]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__27_ ( .D(n4527), .CLK(clk), .QN(
        apbi[27]) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__11_ ( .D(n4526), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__11_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__11_ ( .D(n4525), .CLK(clk), .QN(
        irqctrl0_r_IPEND__11_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__11_ ( .D(n4524), .CLK(clk), .QN(
        ahbso_1__HRDATA__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__11_ ( 
        .D(n4523), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__11_ ( 
        .D(n4522), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[15]) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_DEBUG_ ( .D(n17804), .CLK(clk), .QN(n4520)
         );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TXTICK_ ( .D(uart1_v_TXTICK_), .CLK(clk), 
        .QN(n4519) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TXSTATE__0_ ( .D(n17444), .CLK(clk), .QN(
        n4518) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TXSTATE__1_ ( .D(n17445), .CLK(clk), .QN(
        n4517) );
  SDFHx4_ASAP7_75t_SL uart1_r_reg_TCNT__5_ ( .D(n5590), .SI(n19002), .SE(
        n24695), .CLK(clk), .QN(uart1_r_TCNT__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TCNT__2_ ( .D(n4515), .CLK(clk), .QN(
        uart1_r_TCNT__2_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__24_ ( .D(n4513), .CLK(clk), .QN(
        ahbso_1__HRDATA__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__24_ ( 
        .D(n4512), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__24_ ( .D(n4511), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_OVF_ ( .D(n4508), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_divo[31]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__63_ ( .D(n4507), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[33]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__31_ ( .D(n4505), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__ICC__0_ ( .D(n4503), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_de_icc_0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__20_ ( .D(n4501), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__20_ ( 
        .D(n4500), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__20_ ( 
        .D(n4499), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[24]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__20_ ( .D(n4498), .CLK(clk), .QN(
        apbi[20]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__20_ ( .D(
        timer0_v_TIMERS__1__VALUE__20_), .CLK(clk), .QN(n4497) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__20_ ( .D(n4496), .CLK(clk), .QN(
        ahbso_1__HRDATA__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PV_ ( .D(n4493), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_iu_r_D__PV_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__NPC__0_ ( .D(n4492), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__NPC__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__31_ ( .D(n4490), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__31_ ( .D(n4488), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__31_ ( .D(n26453), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[31]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__31_ ( 
        .D(n4485), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[63]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_BSTATE__0_ ( .D(n4483), .CLK(clk), .QN(
        sr1_r_BSTATE__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_HRESP__0_ ( .D(n33061), .CLK(clk), .QN(
        ahbso_0__HRESP__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_MEXC_ ( .D(n4481), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_MEXC_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__MEXC_ ( .D(n4480), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__MEXC_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__11_ ( .D(n4478), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[69]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__11_ ( 
        .D(n4477), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[8]) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_CFGA11_ ( .D(n4476), .CLK(clk), .QN(
        ahb0_r_CFGA11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__31_ ( .D(n4475), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__0_ ( .D(n4474), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__33_ ( .D(n4473), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[1]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__1_ ( .D(n4469), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__1_ ( .D(n4467), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[32]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__30_ ( .D(n4465), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__30_ ( .D(n4463), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__10_ ( .D(n4459), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__10_ ( 
        .D(n4458), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[14]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__10_ ( .D(n4457), .CLK(clk), .QN(
        apbi[10]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__10_ ( .D(
        timer0_v_TIMERS__1__VALUE__10_), .CLK(clk), .QN(n4456) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__10_ ( .D(n4455), .CLK(clk), .QN(
        ahbso_1__HRDATA__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__10_ ( 
        .D(n4454), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__10_ ( .D(n4453), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__10_ ( .D(n4452), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__43_ ( .D(n4451), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[11]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__11_ ( .D(n4449), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__11_ ( .D(n4447), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[42]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__10_ ( .D(n4445), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[41]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__9_ ( .D(n4443), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[40]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__8_ ( .D(n4441), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[39]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__40_ ( .D(n4440), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[8]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__8_ ( .D(n4438), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__8_ ( .D(n4436), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[8]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__8_ ( .D(
        n4435), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__8_ ( .D(
        n4434), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[41]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__8_ ( .D(n4433), .CLK(clk), .QN(
        apbi[34]) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__14_ ( .D(n4432), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__14_ ( 
        .D(n4430), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__14_ ( .D(n4429), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__14_ ( .D(n4428), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__47_ ( .D(n4427), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[15]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__14_ ( .D(n4425), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__23_ ( .D(n4423), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__23_ ( .D(n4421), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[54]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__55_ ( .D(n4420), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[23]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__23_ ( .D(n4418), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__23_ ( 
        .D(n4417), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__23_ ( 
        .D(n4416), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[27]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__23_ ( .D(n4415), .CLK(clk), .QN(
        apbi[23]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__23_ ( .D(
        timer0_v_TIMERS__1__VALUE__23_), .CLK(clk), .QN(n4414) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__23_ ( .D(n4413), .CLK(clk), .QN(
        ahbso_1__HRDATA__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__WICC_ ( .D(n4410), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__CTRL__WICC_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RSEL1__0_ ( .D(n4406), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RSEL1__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__27_ ( .D(n4404), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__27_ ( .D(n4402), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__27_ ( .D(n4400), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[58]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__59_ ( .D(n4399), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[27]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__27_ ( .D(n4397), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__15_ ( .D(n4396), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__27_ ( .D(n4394), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[85]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__27_ ( 
        .D(n4393), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[24]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HREADY_ ( .D(n4392), .CLK(clk), .QN(
        ahbso_1__HREADY_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HSLAVE__0_ ( .D(ahb0_v_HSLAVE__0_), .CLK(
        clk), .QN(n4391) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_BG_ ( .D(n4390), .CLK(
        clk), .QN(u0_0_leon3x0_p0_c0mmu_a0_r_BG_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_STATE__0_ ( .D(n4389), .CLK(clk), .QN(
        apb0_r_STATE__0_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__21_ ( .D(n4386), .CLK(clk), .QN(
        apbi[21]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__21_ ( .D(
        timer0_v_TIMERS__1__VALUE__21_), .CLK(clk), .QN(n4385) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__21_ ( .D(n4384), .CLK(clk), .QN(
        ahbso_1__HRDATA__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__21_ ( 
        .D(n4383), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__5_ ( .D(n4382), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__5_ ( .D(n4379), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__38_ ( .D(n4378), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[6]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__6_ ( .D(n4376), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__6_ ( .D(n4374), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[6]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__6_ ( .D(
        n4373), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__6_ ( .D(
        n4372), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[39]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__6_ ( .D(n17889), .CLK(clk), .QN(
        n4371) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_RELOAD__0_ ( .D(n4370), .CLK(clk), .QN(
        timer0_r_RELOAD__0_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_SCALER__0_ ( .D(n4369), .CLK(clk), .QN(
        timer0_r_SCALER__0_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__0_ ( .D(n4368), .CLK(clk), .QN(
        ahbso_1__HRDATA__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__0_ ( 
        .D(n4367), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__0_ ( 
        .D(n4366), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[4]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__ENABLE_ ( .D(n4364), .CLK(clk), 
        .QN(timer0_vtimers_1__ENABLE_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__19_ ( .D(
        timer0_v_TIMERS__1__VALUE__19_), .CLK(clk), .QN(n4363) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__19_ ( .D(n4362), .CLK(clk), .QN(
        ahbso_1__HRDATA__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__19_ ( 
        .D(n4361), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__19_ ( .D(n4360), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__18_ ( .D(n4358), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__18_ ( 
        .D(n4357), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__18_ ( 
        .D(n4356), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[22]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__18_ ( .D(n4355), .CLK(clk), .QN(
        apbi[18]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__18_ ( .D(
        timer0_v_TIMERS__1__VALUE__18_), .CLK(clk), .QN(n4354) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__18_ ( .D(n4353), .CLK(clk), .QN(
        ahbso_1__HRDATA__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__18_ ( .D(n24451), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RSEL1__1_ ( .D(n4350), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RSEL1__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__21_ ( .D(n4348), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__21_ ( .D(n4346), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__21_ ( .D(n4344), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[52]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__53_ ( .D(n4343), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[21]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__21_ ( .D(n4341), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__ICC__1_ ( .D(n4340), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__ICC__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__31_ ( .D(n4334), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[89]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__31_ ( .D(n4332), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[59]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__31_ ( .D(n4330), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__31_ ( .D(n4328), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__ICC__3_ ( .D(n4326), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_de_icc_3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_STATE__0_ ( .D(n18176), 
        .CLK(clk), .QN(n4325) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__62_ ( .D(n4324), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[30]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__30_ ( .D(n4322), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__18_ ( .D(n4321), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__30_ ( .D(n4319), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[88]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_HOLDN_ ( .D(
        u0_0_leon3x0_p0_c0mmu_icache0_v_HOLDN_), .CLK(clk), .QN(n4318) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_NOMDS_ ( .D(n4317), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_NOMDS_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_HOLDN_ ( .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_HOLDN_), .CLK(clk), .QN(n4316) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_ZERO_ ( .D(n4313), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_v_ZERO2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_ZERO2_ ( .D(n4311), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_ZERO2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__0_ ( .D(
        n4309), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[0]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__1_ ( .D(
        n4307), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[1]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__2_ ( .D(
        n4305), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[2]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__3_ ( .D(
        n4303), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[3]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__4_ ( .D(
        n4301), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[4]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__5_ ( .D(
        n4299), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[5]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__6_ ( .D(
        n4297), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[6]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__7_ ( .D(
        n4295), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[7]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__8_ ( .D(
        n4293), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[8]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__9_ ( .D(
        n4291), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[9]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__10_ ( .D(
        n4289), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[10]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__11_ ( .D(
        n4287), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[11]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__12_ ( .D(
        n4285), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[12]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__13_ ( .D(
        n4283), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[13]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__14_ ( .D(
        n4281), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[14]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__15_ ( .D(
        n4279), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[15]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__16_ ( .D(
        n4277), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[16]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__17_ ( .D(
        n4275), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[17]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__18_ ( .D(
        n4273), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[18]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__19_ ( .D(
        n4271), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[19]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__20_ ( .D(
        n4269), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[20]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__21_ ( .D(
        n4267), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[21]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__22_ ( .D(
        n4265), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[22]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__23_ ( .D(
        n4263), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[23]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__24_ ( .D(
        n4261), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[24]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__25_ ( .D(
        n4259), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[25]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__26_ ( .D(
        n4257), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[26]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__27_ ( .D(
        n4255), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[27]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__28_ ( .D(
        n4253), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[28]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__29_ ( .D(
        n4251), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[29]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__30_ ( .D(
        n4249), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[30]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__31_ ( .D(
        n4247), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[63]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__32_ ( .D(
        n4245), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[31]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__33_ ( .D(
        n4243), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[32]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__34_ ( .D(
        n4241), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[33]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__35_ ( .D(
        n4239), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[34]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__36_ ( .D(
        n4237), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[35]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__37_ ( .D(
        n4235), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[36]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__38_ ( .D(
        n4233), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[37]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__39_ ( .D(
        n4231), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[38]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__40_ ( .D(
        n4229), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[39]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__42_ ( .D(
        n4225), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[41]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__52_ ( .D(
        n4205), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[51]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__53_ ( .D(
        n4203), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[52]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__57_ ( .D(
        n4195), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[56]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__62_ ( .D(
        n4185), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[61]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__18_ ( .D(n4181), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__23_ ( .D(n4175), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__ANNUL_ ( .D(n4173), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_D__ANNUL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RSEL1__2_ ( .D(n4171), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RSEL1__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA1__0_ ( .D(n4169), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA1__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__CNT__0_ ( .D(n4167), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__CNT__0_ ( .D(n4163), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__CNT__1_ ( .D(n4161), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__18_ ( .D(n4159), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__20_ ( .D(n4157), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__22_ ( .D(n4155), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__23_ ( .D(n4153), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__31_ ( .D(n4151), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__1_ ( .D(n4149), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[1]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__5_ ( .D(n4147), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[5]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__9_ ( .D(n4145), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[9]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__11_ ( .D(n4143), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[11]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__12_ ( .D(n4141), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[12]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__13_ ( .D(n4139), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[13]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__16_ ( .D(n4137), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[16]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__19_ ( .D(n4135), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[19]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__20_ ( .D(n4133), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[20]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__21_ ( .D(n4131), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[21]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__22_ ( .D(n4129), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[22]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__23_ ( .D(n4127), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[23]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__24_ ( .D(n4125), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[24]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__25_ ( .D(n4123), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[25]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__26_ ( .D(n4121), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[26]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__27_ ( .D(n4119), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[27]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__28_ ( .D(n4117), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[28]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__29_ ( .D(n4115), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[29]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__30_ ( .D(n4113), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[30]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__CNT__0_ ( .D(n4111), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__CNT__1_ ( .D(n4109), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__20_ ( .D(n4107), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__23_ ( .D(n4103), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__20_ ( .D(n4101), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__22_ ( .D(n4099), .CLK(clk), .QN(u0_0_dbgo_OPTYPE__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__23_ ( .D(n4097), .CLK(clk), .QN(u0_0_dbgo_OPTYPE__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__31_ ( .D(n4095), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[28]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DIVZ_ ( .D(n4093), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_M__DIVZ_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__NALIGN_ ( .D(n4091), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_M__NALIGN_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__0_ ( .D(n4089), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[31]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__LADDR__1_ ( .D(n4087), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__LADDR__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__23_ ( .D(n4085), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CCTRL__DCS__1_ ( 
        .D(n4084), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DCS__1_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_BURST_ ( .D(n4083), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[1]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_REQ_ ( .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_REQ_), .CLK(clk), .QN(n4082) );
  SDFHx4_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_NBA_ ( .D(n22380), .SI(
        n19002), .SE(n10972), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_a0_r_NBA_)
         );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HWRITE_ ( .D(n4072), .CLK(clk), .QN(
        apbi[32]) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RCNT__5_ ( .D(n4071), .CLK(clk), .QN(
        uart1_r_RCNT__5_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__31_ ( .D(n4070), .CLK(clk), .QN(
        ahbso_1__HRDATA__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__31_ ( .D(n4067), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__31_ ( .D(n4065), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__31_ ( .D(n4063), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__31_ ( .D(n4061), .CLK(clk), .QN(u0_0_dbgo_OPTYPE__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RD__4_ ( .D(n4059), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RD__4_ ( .D(n4057), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RD__4_ ( .D(n4055), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RD__4_ ( .D(n4053), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RSEL2__1_ ( .D(n4051), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RSEL2__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__20_ ( .D(n4049), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__20_ ( .D(n4047), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[51]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__19_ ( .D(n4045), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[50]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__51_ ( .D(n4044), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[19]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__19_ ( .D(n4042), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__19_ ( .D(n4040), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__17_ ( .D(n4038), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[17]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__17_ ( .D(n4036), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__17_ ( 
        .D(n4035), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__17_ ( 
        .D(n4034), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[21]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__17_ ( .D(n4033), .CLK(clk), .QN(
        apbi[17]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__17_ ( .D(
        timer0_v_TIMERS__1__VALUE__17_), .CLK(clk), .QN(n4032) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__17_ ( .D(n4031), .CLK(clk), .QN(
        ahbso_1__HRDATA__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__17_ ( .D(n24440), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__17_ ( .D(n4028), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__17_ ( .D(n4026), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PV_ ( .D(n4024), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PV_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PV_ ( .D(n4022), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PV_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PV_ ( .D(n4020), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PV_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__CWP__2_ ( .D(n4018), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_A__CWP__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CWP__2_ ( .D(n4016), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_E__CWP__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CWP__2_ ( .D(n4014), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__CWP__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RD__6_ ( .D(n4012), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RD__6_ ( .D(n4010), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RD__6_ ( .D(n4008), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RD__6_ ( .D(n4006), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RSEL2__0_ ( .D(n4004), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RSEL2__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__18_ ( .D(n4002), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__18_ ( .D(n4000), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[18]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__18_ ( .D(n3998), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__18_ ( .D(n3997), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__18_ ( .D(n3995), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[49]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__17_ ( .D(n3993), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[48]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__16_ ( .D(n3991), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[47]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__48_ ( .D(n3990), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[16]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__16_ ( .D(n3988), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__16_ ( .D(n3986), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__15_ ( .D(n3984), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[15]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__15_ ( .D(n3982), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__15_ ( .D(n3980), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[46]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__14_ ( .D(n3978), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[45]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__13_ ( .D(n3976), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[44]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__12_ ( .D(n3974), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[43]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__44_ ( .D(n3973), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[12]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__12_ ( .D(n3971), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__12_ ( .D(n3969), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__7_ ( .D(n3967), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[7]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__7_ ( .D(n3965), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__4_ ( .D(n3963), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[4]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__3_ ( .D(n3957), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__2_ ( .D(n3955), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__2_ ( .D(n3953), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[2]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__2_ ( .D(n3951), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__2_ ( .D(n3949), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[33]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__34_ ( .D(n3948), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[2]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__2_ ( .D(n3946), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__6_ ( .D(n3944), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[64]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__6_ ( .D(n3942), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[34]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__6_ ( .D(n3940), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__6_ ( .D(n3938), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__6_ ( .D(n3936), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__6_ ( .D(n3934), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[3]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__6_ ( .D(n3932), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__6_ ( .D(n3930), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__6_ ( .D(n3929), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__39_ ( .D(n3928), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[7]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__7_ ( .D(n3926), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__7_ ( .D(n3924), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[38]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__6_ ( .D(n3922), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[37]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__5_ ( .D(n3920), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[36]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__37_ ( .D(n3919), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[5]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__5_ ( .D(n3917), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TT__5_ ( .D(n18053), 
        .CLK(clk), .QN(n3916) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__INTACK_ ( .D(n3914), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__INTACK_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CCTRL__ICS__1_ ( 
        .D(n3913), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__1_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__1_ ( .D(n3912), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__LADDR__0_ ( .D(n3908), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__LADDR__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CCTRL__ICS__0_ ( 
        .D(n3907), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__0_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_REQ_ ( .D(n3906), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[0]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_NBO__0_ ( .D(n3905), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_a0_r_NBO__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_BO__0_ ( .D(n3904), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_a0_r_BO__0_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HMASTERD_ ( .D(n3901), .CLK(clk), .QN(
        ahb0_r_HMASTERD_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HTRANS__1_ ( .D(n3900), .CLK(clk), .QN(
        ahb0_r_HTRANS__1_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HREADY_ ( .D(ahb0_v_HREADY_), .CLK(clk), 
        .QN(n4832) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_CFGSEL_ ( .D(ahb0_v_CFGSEL_), .CLK(clk), 
        .QN(n3899) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_BO__1_ ( .D(
        u0_0_leon3x0_p0_c0mmu_a0_v_BO__1_), .CLK(clk), .QN(n3897) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_HLOCKEN_ ( .D(n3896), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_a0_r_HLOCKEN_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_UNDERRUN_ ( .D(
        n3895), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_UNDERRUN_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_OVERRUN_ ( .D(
        n3894), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_OVERRUN_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__30_ ( .D(n3891), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__30_ ( .D(n3889), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__30_ ( .D(n3887), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__30_ ( .D(n3885), .CLK(clk), .QN(u0_0_dbgo_OPTYPE__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RETT_ ( .D(n3883), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__CTRL__RETT_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INULL_ ( .D(n3881), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_D__INULL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_ISTATE__0_ ( .D(
        n18248), .CLK(clk), .QN(n3880) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_ISTATE__1_ ( .D(
        n3879), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__1_ ( .D(n18212), 
        .CLK(clk), .QN(n4928) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__2_ ( .D(n18211), 
        .CLK(clk), .QN(n4929) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__3_ ( .D(n18210), 
        .CLK(clk), .QN(n4930) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__4_ ( .D(n18209), 
        .CLK(clk), .QN(n3878) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__21_ ( .D(n3875), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__21_ ( .D(n3873), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__21_ ( .D(n3871), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__21_ ( .D(n3869), .CLK(clk), .QN(u0_0_dbgo_OPTYPE__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__MULSTART_ ( .D(n3867), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__MULSTART_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__24_ ( .D(n3864), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__24_ ( .D(n3862), .CLK(clk), .QN(u0_0_leon3x0_p0_muli[8]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__24_ ( .D(n3860), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__24_ ( .D(n3858), .CLK(clk), .QN(u0_0_dbgo_OPTYPE__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__ICC__1_ ( .D(n3856), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__ICC__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__1_ ( .D(n3854), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__6_ ( .D(n3852), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__7_ ( .D(n3850), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__8_ ( .D(n3848), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__10_ ( .D(n3846), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__11_ ( .D(n3844), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__14_ ( .D(n3842), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__15_ ( .D(n3840), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__26_ ( .D(n3838), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__28_ ( .D(n3836), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__29_ ( .D(n3834), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__31_ ( .D(n3832), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__0_ ( .D(n3830), .CLK(
        clk), .QN(u0_0_leon3x0_p0_muli[0]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__1_ ( .D(n3828), .CLK(
        clk), .QN(u0_0_leon3x0_p0_muli[1]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__2_ ( .D(n3826), .CLK(
        clk), .QN(u0_0_leon3x0_p0_muli[2]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__5_ ( .D(n3824), .CLK(
        clk), .QN(u0_0_leon3x0_p0_muli[5]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__6_ ( .D(n3822), .CLK(
        clk), .QN(u0_0_leon3x0_p0_muli[6]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__7_ ( .D(n3820), .CLK(
        clk), .QN(u0_0_leon3x0_p0_muli[7]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__8_ ( .D(n3818), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__9_ ( .D(n3816), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__10_ ( .D(n3814), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__11_ ( .D(n3812), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__12_ ( .D(n3810), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__13_ ( .D(n3808), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__14_ ( .D(n3806), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__15_ ( .D(n3804), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__16_ ( .D(n3802), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__17_ ( .D(n3800), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__18_ ( .D(n3798), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__19_ ( .D(n3796), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__20_ ( .D(n3794), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__21_ ( .D(n3792), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__23_ ( .D(n3790), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__25_ ( .D(n3788), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__26_ ( .D(n3786), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__27_ ( .D(n3784), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__28_ ( .D(n3782), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__MUL_ ( .D(n3780), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__MUL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__MUL_ ( .D(n3778), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__MUL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__25_ ( .D(n24454), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__25_ ( .D(n3775), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__25_ ( .D(n3773), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__25_ ( .D(n3771), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__25_ ( .D(n3769), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__26_ ( .D(n24441), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__26_ ( .D(n3764), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__26_ ( .D(n3762), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__26_ ( .D(n3760), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA1__1_ ( .D(n3758), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA1__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RD__1_ ( .D(n3756), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RD__1_ ( .D(n3754), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RD__1_ ( .D(n3752), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RD__1_ ( .D(n3750), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__29_ ( .D(n24438), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__29_ ( .D(n3747), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__29_ ( .D(n3745), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__29_ ( .D(n3743), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__29_ ( .D(n3741), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__ANNUL_ ( .D(n3739), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__CTRL__ANNUL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__TRAP_ ( .D(n3737), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__TRAP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__TRAP_ ( .D(n3735), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__TRAP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__TRAP_ ( .D(n3733), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__TRAP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__ET_ ( .D(n3731), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__ET_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RSTATE__1_ ( .D(n18277), 
        .CLK(clk), .QN(n3730) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__ANNUL_ALL_ ( .D(n3728), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_muli[10]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_STATE__1_ ( .D(n18175), 
        .CLK(clk), .QN(n3727) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_CNT__4_ ( .D(n3726), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_CNT__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_STATE__2_ ( .D(n18174), 
        .CLK(clk), .QN(n3725) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_CNT__0_ ( .D(n3724), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_CNT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_CNT__1_ ( .D(n3723), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_CNT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_CNT__2_ ( .D(n3722), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_CNT__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_CNT__3_ ( .D(n3721), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_CNT__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_ZCORR_ ( .D(n18171), .CLK(
        clk), .QN(n4949) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__DIVRDY_ ( .D(n3719), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_D__DIVRDY_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__DIVSTART_ ( .D(n3717), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__DIVSTART_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__WICC_ ( .D(n3715), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__CTRL__WICC_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__WICC_ ( .D(n3713), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__WICC_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__ANNUL_ ( .D(n3709), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__CTRL__ANNUL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__ANNUL_ ( .D(n3707), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__ANNUL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__ANNUL_ ( .D(n3705), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__ANNUL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RSTATE__0_ ( .D(n18276), 
        .CLK(clk), .QN(n3704) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__NPC__1_ ( .D(n3703), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__NPC__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__MEXC_ ( .D(n3702), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__TRAP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__TT__0_ ( .D(n3700), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__CTRL__TT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RETT_ ( .D(n3698), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__CTRL__RETT_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RETT_ ( .D(n3696), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__RETT_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RETT_ ( .D(n3694), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RETT_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__5_ ( .D(n24457), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__5_ ( .D(n3691), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__5_ ( .D(n3689), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__5_ ( .D(n3687), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__6_ ( .D(n24455), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__6_ ( .D(n3684), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__6_ ( .D(n3682), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__ASI__1_ ( .D(n3680), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[38]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__6_ ( .D(n3678), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__7_ ( .D(n24443), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__7_ ( .D(n3675), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__7_ ( .D(n3673), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__ASI__2_ ( .D(n3671), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[39]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__7_ ( .D(n3669), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__8_ ( .D(n24434), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__8_ ( .D(n3666), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__8_ ( .D(n3664), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__ASI__3_ ( .D(n3662), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[40]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__8_ ( .D(n3660), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__9_ ( .D(n24445), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__9_ ( .D(n3657), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__9_ ( .D(n3655), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__ASI__4_ ( .D(n3653), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[41]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__9_ ( .D(n3651), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__10_ ( .D(n24435), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__10_ ( .D(n3648), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__11_ ( .D(n24433), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__11_ ( .D(n3645), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__12_ ( .D(n22217), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__22_ ( .D(n3642), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__15_ ( .D(n3640), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__16_ ( .D(n24508), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__17_ ( .D(n3636), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__18_ ( .D(n24507), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__19_ ( .D(n24506), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__20_ ( .D(n24505), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__21_ ( .D(n24504), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__30_ ( .D(n24497), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__31_ ( .D(n24499), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__13_ ( .D(n24458), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__13_ ( .D(n3621), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__23_ ( .D(n24500), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__14_ ( .D(n24444), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__14_ ( .D(n3616), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__14_ ( .D(n3614), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__24_ ( .D(n24503), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__16_ ( .D(n24436), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__26_ ( .D(n24502), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__19_ ( .D(n3602), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__19_ ( .D(n3600), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__2_ ( .D(n3599), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__3_ ( .D(n3598), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__9_ ( .D(n3597), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__11_ ( .D(n3596), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__14_ ( .D(n3595), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__16_ ( .D(n3594), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__17_ ( .D(n3593), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__19_ ( .D(n3592), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__SIZE__1_ ( .D(n3590), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[5]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DCI__SIZE__1_ ( .D(n3588), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__LOCK_ ( .D(n3586), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__DCI__LOCK_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__SIZE__0_ ( .D(n3584), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[4]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DCI__SIZE__0_ ( .D(n3582), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__SIGNED_ ( .D(n3580), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__DCI__SIGNED_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DCI__SIGNED_ ( .D(n3578), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DCI__SIGNED_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__WCWP_ ( .D(n3576), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_M__WCWP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__MULSTEP_ ( .D(n3574), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__MULSTEP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__SARI_ ( .D(n3572), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__SARI_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__ALUOP__2_ ( .D(n3570), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__ALUOP__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__SHLEFT_ ( .D(n3568), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__SHLEFT_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__SHCNT__1_ ( .D(n3566), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__SHCNT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__SHCNT__2_ ( .D(n3564), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__SHCNT__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__SHCNT__3_ ( .D(n3562), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__SHCNT__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__TICC_ ( .D(n3556), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__TICC_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__14_ ( .D(n3554), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA2__3_ ( .D(n3552), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA2__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA2__7_ ( .D(n3550), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA2__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__13_ ( .D(n3548), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__1_ ( .D(n3546), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__2_ ( .D(n3544), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__3_ ( .D(n3542), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA2__1_ ( .D(n3540), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA2__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__11_ ( .D(n3538), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA2__2_ ( .D(n3536), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA2__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__12_ ( .D(n3534), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RD__0_ ( .D(n3532), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RD__0_ ( .D(n3530), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RD__0_ ( .D(n3528), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RD__0_ ( .D(n3526), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__WUNF_ ( .D(n3524), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__WUNF_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__4_ ( .D(n3522), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__29_ ( .D(n24501), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__LD_ ( .D(n3518), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__LD_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__LD_ ( .D(n3516), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__LD_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__LD_ ( .D(n3514), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__LD_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__LD_ ( .D(n3512), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__LD_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__27_ ( .D(n24453), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__27_ ( .D(n3509), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__27_ ( .D(n3507), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__27_ ( .D(n3505), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__27_ ( .D(n3503), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA1__2_ ( .D(n3501), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA1__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RD__2_ ( .D(n3499), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RD__2_ ( .D(n3497), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RD__2_ ( .D(n3495), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RD__2_ ( .D(n3493), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__28_ ( .D(n24452), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__28_ ( .D(n3490), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__28_ ( .D(n3488), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__28_ ( .D(n3486), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__INST__28_ ( .D(n3484), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__DWT_ ( .D(n18252), 
        .CLK(clk), .QN(n4838) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RD__3_ ( .D(n3482), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RD__3_ ( .D(n3480), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RD__3_ ( .D(n3478), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RD__3_ ( .D(n3476), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__0_ ( .D(n18213), 
        .CLK(clk), .QN(n4927) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA2__0_ ( .D(n3474), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA2__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__10_ ( .D(n3472), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__0_ ( .D(n3470), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__4_ ( .D(n3468), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[32]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__4_ ( .D(n3466), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__4_ ( .D(n3464), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__4_ ( .D(n3462), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__4_ ( .D(n3460), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[1]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__5_ ( .D(n3458), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[33]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__5_ ( .D(n3456), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__5_ ( .D(n3454), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__5_ ( .D(n3452), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__5_ ( .D(n3450), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[2]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__7_ ( .D(n3448), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[35]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__7_ ( .D(n3446), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__7_ ( .D(n3444), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__7_ ( .D(n3442), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__7_ ( .D(n3440), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[4]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__8_ ( .D(n3438), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[36]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__8_ ( .D(n3436), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__8_ ( .D(n3434), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__8_ ( .D(n3432), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__8_ ( .D(n3430), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[5]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__9_ ( .D(n3428), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[37]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__9_ ( .D(n3426), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__9_ ( .D(n3424), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__9_ ( .D(n3422), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__9_ ( .D(n3420), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[6]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__11_ ( .D(n3418), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[39]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__11_ ( .D(n3416), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__11_ ( .D(n3414), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__11_ ( .D(n3412), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__11_ ( .D(n3410), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[8]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__25_ ( .D(n3408), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[53]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__25_ ( .D(n3406), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__25_ ( .D(n3404), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__25_ ( .D(n3402), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__25_ ( .D(n3400), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[22]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__27_ ( .D(n3398), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[55]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__27_ ( .D(n3396), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__27_ ( .D(n3394), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__27_ ( .D(n3392), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__27_ ( .D(n3390), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[24]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__NPC__2_ ( .D(n3389), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__NPC__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__1_ ( .D(n3387), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__IRQEN_ ( .D(n3385), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_M__IRQEN2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__IRQEN2_ ( .D(n3383), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_M__IRQEN2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__5_ ( .D(n3381), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__25_ ( .D(n3379), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__NERROR_ ( .D(n3376), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__NERROR_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__ET_ ( .D(n3374), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_iu_v_E__ET_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__ET_ ( .D(n3372), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_iu_r_E__ET_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__ASI__0_ ( .D(n3364), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[37]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__SU_ ( .D(n3362), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_iu_v_E__SU_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__SU_ ( .D(n3360), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_dci[0]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__TT__1_ ( .D(n3358), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__TT__1_ ( .D(n3356), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__TT__2_ ( .D(n3354), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__TT__2_ ( .D(n3352), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__TT__4_ ( .D(n3350), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__TT__4_ ( .D(n3348), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__TT__3_ ( .D(n3346), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__TT__3_ ( .D(n3344), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__TT__0_ ( .D(n3342), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__TT__0_ ( .D(n3340), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__WIM__1_ ( .D(n3338), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__WIM__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__WIM__2_ ( .D(n3336), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__WIM__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__WIM__5_ ( .D(n3334), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__WIM__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__WIM__6_ ( .D(n3332), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__WIM__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__WIM__7_ ( .D(n3330), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__WIM__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__PIL__0_ ( .D(n3329), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__PIL__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__PIL__2_ ( .D(n18089), 
        .CLK(clk), .QN(n3328) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__PIL__3_ ( .D(n18090), 
        .CLK(clk), .QN(n3327) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__TT__2_ ( .D(n3326), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TT__1_ ( .D(n18049), 
        .CLK(clk), .QN(n3325) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TT__6_ ( .D(n3324), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TT__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TT__7_ ( .D(n3323), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TT__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TT__2_ ( .D(n3322), 
        .CLK(clk), .QN(irqo[1]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__WRITE_ ( .D(n3320), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[1]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CASA_ ( .D(n3318), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_M__CASA_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__26_ ( .D(n3313), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__1_ ( .D(n3312), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__ALUSEL__0_ ( .D(n3310), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__ALUSEL__1_ ( .D(n3308), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__ALUSEL__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__ALUADD_ ( .D(n3306), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__ALUADD_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__ENADDR_ ( .D(n3304), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[3]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__NOBP_ ( .D(n3300), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__NOBP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__BP_ ( .D(n3298), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_iu_r_A__BP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__BRANCH_ ( .D(n3296), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[29]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__BP_ ( .D(n3294), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_iu_r_E__BP_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__29_ ( .D(n3292), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[87]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__29_ ( .D(n3290), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[57]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__29_ ( .D(n3288), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__29_ ( .D(n3286), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__29_ ( .D(n3284), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__29_ ( .D(n3282), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[26]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__28_ ( .D(n3280), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[86]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__28_ ( .D(n3278), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[56]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__28_ ( .D(n3276), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__28_ ( .D(n3274), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__28_ ( .D(n3272), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__28_ ( .D(n3270), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[25]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__28_ ( .D(n3268), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__26_ ( .D(n3266), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[84]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__26_ ( .D(n3264), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[54]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__26_ ( .D(n3262), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__26_ ( .D(n3260), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__26_ ( .D(n3258), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__26_ ( .D(n3256), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[23]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__26_ ( .D(n3254), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__23_ ( .D(n3252), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[81]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__23_ ( .D(n3250), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[51]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__23_ ( .D(n3248), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__23_ ( .D(n3246), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__23_ ( .D(n3244), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__23_ ( .D(n3242), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[20]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__21_ ( .D(n3240), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[79]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__21_ ( .D(n3238), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[49]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__21_ ( .D(n3236), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__21_ ( .D(n3234), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__21_ ( .D(n3232), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__21_ ( .D(n3230), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[18]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__15_ ( .D(n3228), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[73]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__15_ ( .D(n3226), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[43]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__15_ ( .D(n3224), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__15_ ( .D(n3222), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__15_ ( .D(n3220), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__15_ ( .D(n3218), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[12]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__14_ ( .D(n3216), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[72]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__14_ ( .D(n3214), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[42]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__14_ ( .D(n3212), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__14_ ( .D(n3210), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__14_ ( .D(n3208), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__14_ ( .D(n3206), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[11]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__14_ ( .D(n3204), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__2_ ( .D(n3200), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[30]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__2_ ( .D(n3198), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__2_ ( .D(n3196), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__2_ ( .D(n3194), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__2_ ( .D(n3192), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__PC__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__3_ ( .D(n3190), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[61]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__3_ ( .D(n3188), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[31]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__3_ ( .D(n3186), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__3_ ( .D(n3184), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__3_ ( .D(n3182), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__3_ ( .D(n3180), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[0]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__10_ ( .D(n3178), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[68]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__10_ ( .D(n3176), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[38]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__10_ ( .D(n3174), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__10_ ( .D(n3172), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__10_ ( .D(n3170), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__10_ ( .D(n3168), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[7]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__10_ ( .D(n3166), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__JMPL_ ( .D(n3164), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_A__JMPL_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA1__7_ ( .D(n3160), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA1__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__WY_ ( .D(n3158), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__WY_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__WY_ ( .D(n3156), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__WY_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__WY_ ( .D(n3154), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__WY_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__WY_ ( .D(n3152), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__WY_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__1_ ( .D(n3151), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__2_ ( .D(n3150), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__5_ ( .D(n3149), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__6_ ( .D(n3148), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__7_ ( .D(n3147), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__8_ ( .D(n3146), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__10_ ( .D(n3145), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__11_ ( .D(n3144), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__14_ ( .D(n3143), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__15_ ( .D(n3142), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__21_ ( .D(n3141), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__23_ ( .D(n3140), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__25_ ( .D(n3139), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__26_ ( .D(n3138), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__27_ ( .D(n3137), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__28_ ( .D(n3136), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FLUSH_ ( .D(n18096), .CLK(clk), .QN(n3135) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_DSTATE__2_ ( .D(
        n18101), .CLK(clk), .QN(n3134) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__4_ ( .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__4_), .CLK(clk), .QN(n3133)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_DSTATE__3_ ( .D(
        n18102), .CLK(clk), .QN(n3132) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CCTRLWR_ ( .D(
        n3131), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_CCTRLWR_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_SIZE__1_ ( .D(
        n3129), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_SIZE__0_ ( .D(
        n3127), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__31_ ( 
        .D(n3125), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__30_ ( 
        .D(n3123), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__29_ ( 
        .D(n3121), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__28_ ( 
        .D(n3119), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__27_ ( 
        .D(n3117), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__26_ ( 
        .D(n3115), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__25_ ( 
        .D(n3113), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__24_ ( 
        .D(n3111), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__23_ ( 
        .D(n3109), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__22_ ( 
        .D(n3107), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__21_ ( 
        .D(n3105), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__20_ ( 
        .D(n3103), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__19_ ( 
        .D(n3101), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__18_ ( 
        .D(n3099), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__17_ ( 
        .D(n3097), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__16_ ( 
        .D(n3095), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__15_ ( 
        .D(n3093), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__14_ ( 
        .D(n3091), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__13_ ( 
        .D(n3089), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__12_ ( 
        .D(n3087), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__4_ ( .D(
        n3085), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__3_ ( .D(
        n3083), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__1_ ( .D(
        n3081), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__0_ ( .D(
        n3079), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_ASI__0_ ( .D(n3077), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_ASI__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_READ_ ( .D(n3076), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_READ_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__5_ ( .D(
        n3075), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__7_ ( .D(
        n3074), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__9_ ( .D(
        n3073), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__11_ ( 
        .D(n3072), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_DSTATE__1_ ( .D(
        n18100), .CLK(clk), .QN(n3071) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_DSTATE__0_ ( .D(
        n3070), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_DIAGRDY_ ( .D(
        n14803), .CLK(clk), .QN(u0_0_leon3x0_p0_ico_DIAGRDY_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CACHE_ ( .D(n18047), .CLK(clk), .QN(n3068) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_XADDRESS__2_ ( .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_XADDRESS__2_), .CLK(clk), .QN(n3067)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FADDR__6_ ( .D(
        n3066), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FADDR__5_ ( .D(
        n3062), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FADDR__4_ ( .D(
        n3061), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FADDR__3_ ( .D(
        n3060), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FADDR__2_ ( .D(
        n3059), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FADDR__1_ ( .D(
        n3058), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FADDR__0_ ( .D(
        n3057), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_NOFLUSH_ ( .D(
        n3056), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_NOFLUSH_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FLUSH_ ( .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_FLUSH_), .CLK(clk), .QN(n3055) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FADDR__6_ ( .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_FADDR__6_), .CLK(clk), .QN(n3054) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FADDR__0_ ( .D(
        n3052), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FADDR__1_ ( .D(
        n3051), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FADDR__2_ ( .D(
        n3050), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FADDR__3_ ( .D(
        n3049), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FADDR__4_ ( .D(
        n3048), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FADDR__5_ ( .D(
        n3047), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CCTRL__DCS__0_ ( 
        .D(u0_0_leon3x0_p0_c0mmu_dcache0_v_CCTRL__DCS__0_), .CLK(clk), .QN(
        n3046) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_VALID_ ( .D(n3044), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_VALID_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_STPEND_ ( .D(n3042), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_STPEND_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__0_ ( .D(n3041), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__2_ ( .D(n3040), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__2_ ( .D(n3038), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__2_ ( .D(n3037), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__3_ ( .D(n3036), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__3_ ( .D(n3035), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__6_ ( .D(n3034), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__7_ ( .D(n3033), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__7_ ( .D(n3031), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__8_ ( .D(n3030), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__8_ ( .D(n3028), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__11_ ( .D(n3027), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__11_ ( .D(n3025), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__11_ ( .D(n3024), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__12_ ( .D(n3023), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__15_ ( .D(n3022), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__15_ ( .D(n3020), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__15_ ( .D(n3019), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__17_ ( .D(n3018), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__18_ ( .D(n3017), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__20_ ( .D(n3016), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__21_ ( .D(n3015), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__21_ ( .D(n3013), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__22_ ( .D(n3012), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__23_ ( .D(n3011), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__23_ ( .D(n3009), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__27_ ( .D(n3008), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__27_ ( .D(n3006), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__27_ ( .D(n3005), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__29_ ( .D(n3004), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__29_ ( .D(n3002), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__29_ ( .D(n3001), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__30_ ( .D(n3000), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_BMEXC_ ( .D(n2999), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_BMEXC_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__READ_ ( .D(
        n2998), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[0]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__SIZE__0_ ( .D(
        n2997), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[2]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__SIZE__1_ ( .D(
        n2996), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[3]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__5_ ( .D(
        n2995), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[38]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__5_ ( .D(n2994), .CLK(clk), .QN(
        apbi[33]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__7_ ( .D(
        n2993), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[40]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__7_ ( .D(n17890), .CLK(clk), .QN(
        n2992) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__9_ ( .D(
        n2991), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[42]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__11_ ( 
        .D(n2990), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[44]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__11_ ( .D(n2989), .CLK(clk), .QN(
        apbi[37]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__12_ ( 
        .D(n2988), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[45]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__13_ ( 
        .D(n2987), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[46]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__15_ ( 
        .D(n2986), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[48]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__16_ ( 
        .D(n2985), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[49]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__17_ ( 
        .D(n2984), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[50]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__19_ ( 
        .D(n2983), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[52]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__20_ ( 
        .D(n2982), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[53]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__21_ ( 
        .D(n2981), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[54]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__22_ ( 
        .D(n2980), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[55]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__23_ ( 
        .D(n2979), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[56]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__24_ ( 
        .D(n2978), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[57]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__25_ ( 
        .D(n2977), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[58]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__26_ ( 
        .D(n2976), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[59]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__27_ ( 
        .D(n2975), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[60]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__28_ ( 
        .D(n2974), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[61]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__29_ ( 
        .D(n2973), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[62]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__30_ ( 
        .D(n18045), .CLK(clk), .QN(n2972) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_RBURST_ ( .D(n2971), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_dcache0_r_RBURST_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__1_ ( .D(
        n2970), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[37]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_HIT_ ( .D(n2968), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dco_HIT_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CCTRL__IFRZ_ ( .D(
        n2967), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__IFRZ_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__4_ ( .D(n2966), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CCTRL__DFRZ_ ( .D(
        n2965), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DFRZ_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_CCTRL__BURST_ ( 
        .D(n2964), .CLK(clk), .QN(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__BURST_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__2_ ( .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__2_), .CLK(clk), .QN(n2963)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__3_ ( .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__3_), .CLK(clk), .QN(n2962)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__5_ ( .D(
        n2961), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__5_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__7_ ( .D(
        n2960), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__7_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__8_ ( .D(
        n2959), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__8_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__9_ ( .D(
        n2958), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__9_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__11_ ( 
        .D(n2957), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__11_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__25_ ( 
        .D(n32548), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__25_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__27_ ( 
        .D(n2955), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__10_ ( 
        .D(n2954), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__10_ ( 
        .D(n2953), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[7]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__14_ ( 
        .D(n2952), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__14_ ( 
        .D(n2951), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[11]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__14_ ( .D(n2950), .CLK(clk), .QN(
        apbi[40]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__15_ ( 
        .D(n2949), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__15_ ( 
        .D(n2948), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[12]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__15_ ( .D(n2947), .CLK(clk), .QN(
        apbi[41]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__21_ ( 
        .D(n2946), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__21_ ( 
        .D(n2945), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[18]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__23_ ( 
        .D(n32540), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__23_ ( 
        .D(n31762), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[20]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__26_ ( 
        .D(n32551), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__26_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__26_ ( 
        .D(n31779), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[23]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__28_ ( 
        .D(n2940), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__28_ ( 
        .D(n2939), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[25]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__29_ ( 
        .D(n2938), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__29_ ( 
        .D(n2937), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[26]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__2_ ( .D(
        n2936), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__2_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__3_ ( .D(
        u0_0_leon3x0_p0_c0mmu_icache0_v_VADDRESS__3_), .CLK(clk), .QN(n2935)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__4_ ( .D(
        n32685), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__4_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__2_ ( .D(
        u0_0_leon3x0_p0_c0mmu_icache0_v_WADDRESS__2_), .CLK(clk), .QN(n2933)
         );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__2_ ( .D(n2932), .CLK(clk), .QN(
        ahb0_r_HADDR__2_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__2_ ( .D(n17885), .CLK(clk), .QN(
        n2931) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__3_ ( .D(
        n30914), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[1]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__3_ ( .D(n17886), .CLK(clk), .QN(
        n2929) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__3_ ( .D(n2928), .CLK(clk), .QN(
        ahb0_r_HADDR__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__4_ ( .D(
        u0_0_leon3x0_p0_c0mmu_icache0_v_WADDRESS__4_), .CLK(clk), .QN(n2927)
         );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__4_ ( .D(ahb0_v_HADDR__4_), .CLK(clk), 
        .QN(n2926) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__4_ ( .D(n17887), .CLK(clk), .QN(
        n2925) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__BRDYEN_ ( .D(n2923), .CLK(clk), .QN(
        sr1_r_MCFG1__BRDYEN_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__BEXCEN_ ( .D(n2922), .CLK(clk), .QN(
        sr1_r_MCFG1__BEXCEN_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__IOWS__0_ ( .D(n2921), .CLK(clk), .QN(
        sr1_r_MCFG1__IOWS__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__IOWS__1_ ( .D(n2920), .CLK(clk), .QN(
        sr1_r_MCFG1__IOWS__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__IOWS__2_ ( .D(n2919), .CLK(clk), .QN(
        sr1_r_MCFG1__IOWS__2_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__IOWS__3_ ( .D(n2918), .CLK(clk), .QN(
        sr1_r_MCFG1__IOWS__3_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMWRITE_ ( .D(n2917), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMWRITE_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMWIDTH__0_ ( .D(n2916), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMWIDTH__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RMW_ ( .D(n2915), .CLK(clk), .QN(
        sr1_r_MCFG2__RMW_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMBANKSZ__1_ ( .D(n2914), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMBANKSZ__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMBANKSZ__3_ ( .D(n2913), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMBANKSZ__3_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMWIDTH__0_ ( .D(n2912), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMWIDTH__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMWIDTH__1_ ( .D(n2911), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMWIDTH__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMWWS__0_ ( .D(n2910), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMWWS__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMWWS__1_ ( .D(n2909), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMWWS__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMRWS__0_ ( .D(n2908), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMRWS__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMRWS__1_ ( .D(n2907), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMRWS__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__IOWIDTH__0_ ( .D(n2906), .CLK(clk), 
        .QN(sr1_r_MCFG1__IOWIDTH__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMWWS__0_ ( .D(n2905), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMWWS__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMWWS__1_ ( .D(n2904), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMWWS__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMWWS__2_ ( .D(n2903), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMWWS__2_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMWWS__3_ ( .D(n2902), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMWWS__3_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMRWS__0_ ( .D(n2901), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMRWS__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMRWS__1_ ( .D(n2900), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMRWS__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMRWS__2_ ( .D(n2899), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMRWS__2_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMRWS__3_ ( .D(n2898), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMRWS__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TCNT__0_ ( .D(n2896), .CLK(clk), .QN(
        uart1_r_TCNT__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TCNT__1_ ( .D(n2895), .CLK(clk), .QN(
        uart1_r_TCNT__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TXEN_ ( .D(n2894), .CLK(clk), .QN(
        uart1_uarto_TXEN_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__1_ ( .D(n2893), .CLK(clk), .QN(
        uart1_r_BRATE__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__2_ ( .D(n2892), .CLK(clk), .QN(
        uart1_r_BRATE__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__3_ ( .D(n2891), .CLK(clk), .QN(
        uart1_r_BRATE__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__4_ ( .D(n2890), .CLK(clk), .QN(
        uart1_r_BRATE__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__5_ ( .D(n2889), .CLK(clk), .QN(
        uart1_r_BRATE__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__6_ ( .D(n2888), .CLK(clk), .QN(
        uart1_r_BRATE__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__7_ ( .D(n2887), .CLK(clk), .QN(
        uart1_r_BRATE__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__8_ ( .D(n2886), .CLK(clk), .QN(
        uart1_r_BRATE__8_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__10_ ( .D(n2885), .CLK(clk), .QN(
        uart1_r_BRATE__10_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__11_ ( .D(n2884), .CLK(clk), .QN(
        uart1_r_BRATE__11_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__11_ ( .D(uart1_v_SCALER__11_), 
        .CLK(clk), .QN(n2883) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__8_ ( .D(n2882), .CLK(clk), .QN(
        uart1_uarto_SCALER__8_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__7_ ( .D(n2881), .CLK(clk), .QN(
        uart1_uarto_SCALER__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__6_ ( .D(n2880), .CLK(clk), .QN(
        uart1_uarto_SCALER__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__5_ ( .D(n2879), .CLK(clk), .QN(
        uart1_uarto_SCALER__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__4_ ( .D(n2878), .CLK(clk), .QN(
        uart1_uarto_SCALER__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__3_ ( .D(n2877), .CLK(clk), .QN(
        uart1_uarto_SCALER__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__2_ ( .D(n2876), .CLK(clk), .QN(
        uart1_uarto_SCALER__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__1_ ( .D(n2875), .CLK(clk), .QN(
        uart1_uarto_SCALER__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__10_ ( .D(n2874), .CLK(clk), .QN(
        uart1_uarto_SCALER__10_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__0_ ( .D(n2873), .CLK(clk), .QN(
        uart1_r_BRATE__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__0_ ( .D(n2872), .CLK(clk), .QN(
        uart1_uarto_SCALER__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RFIFOIRQEN_ ( .D(n2871), .CLK(clk), .QN(
        uart1_r_RFIFOIRQEN_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BREAKIRQEN_ ( .D(n2870), .CLK(clk), .QN(
        uart1_r_BREAKIRQEN_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_LOOPB_ ( .D(n2869), .CLK(clk), .QN(
        uart1_r_LOOPB_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_PAREN_ ( .D(n2868), .CLK(clk), .QN(
        uart1_r_PAREN_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXSTATE__2_ ( .D(n17450), .CLK(clk), .QN(
        n2867) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXSTATE__1_ ( .D(n2866), .CLK(clk), .QN(
        uart1_r_RXSTATE__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RSHIFT__0_ ( .D(n2865), .CLK(clk), .QN(
        uart1_r_RSHIFT__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXSTATE__0_ ( .D(n2864), .CLK(clk), .QN(
        uart1_r_RXSTATE__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXCLK__0_ ( .D(n2863), .CLK(clk), .QN(
        uart1_r_RXCLK__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXCLK__1_ ( .D(n2862), .CLK(clk), .QN(
        uart1_r_RXCLK__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RXCLK__2_ ( .D(uart1_v_RXCLK__2_), .CLK(
        clk), .QN(n2861) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_PARSEL_ ( .D(n2860), .CLK(clk), .QN(
        uart1_r_PARSEL_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_DPAR_ ( .D(n2859), .CLK(clk), .QN(
        uart1_r_DPAR_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TIRQEN_ ( .D(n2858), .CLK(clk), .QN(
        uart1_r_TIRQEN_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RIRQEN_ ( .D(n2857), .CLK(clk), .QN(
        uart1_r_RIRQEN_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__1_ ( .D(n2856), .CLK(clk), .QN(
        irqctrl0_r_ILEVEL__1_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__2_ ( .D(n2855), .CLK(clk), .QN(
        irqctrl0_r_ILEVEL__2_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__3_ ( .D(n2854), .CLK(clk), .QN(
        irqctrl0_r_ILEVEL__3_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__4_ ( .D(n2853), .CLK(clk), .QN(
        irqctrl0_r_ILEVEL__4_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__5_ ( .D(n2852), .CLK(clk), .QN(
        irqctrl0_r_ILEVEL__5_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__7_ ( .D(n17785), .CLK(clk), 
        .QN(n2851) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__10_ ( .D(n2850), .CLK(clk), 
        .QN(irqctrl0_r_ILEVEL__10_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__12_ ( .D(n2849), .CLK(clk), 
        .QN(irqctrl0_r_ILEVEL__12_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__15_ ( .D(n2848), .CLK(clk), 
        .QN(irqctrl0_r_ILEVEL__15_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__0_ ( .D(n2847), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__0_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__0_ ( .D(
        timer0_v_TIMERS__1__VALUE__0_), .CLK(clk), .QN(n2846) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__1_ ( .D(n2845), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__1_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__1_ ( .D(
        timer0_v_TIMERS__1__VALUE__1_), .CLK(clk), .QN(n2844) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__2_ ( .D(n2843), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__2_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__2_ ( .D(
        timer0_v_TIMERS__1__VALUE__2_), .CLK(clk), .QN(n2842) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__3_ ( .D(n2841), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__3_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__3_ ( .D(
        timer0_v_TIMERS__1__VALUE__3_), .CLK(clk), .QN(n2840) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__5_ ( .D(n2839), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__5_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__5_ ( .D(
        timer0_v_TIMERS__1__VALUE__5_), .CLK(clk), .QN(n2838) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__10_ ( .D(n2837), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__10_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__15_ ( .D(n2836), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__15_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__17_ ( .D(n2835), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__17_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__18_ ( .D(n2834), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__18_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__20_ ( .D(n2833), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__20_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__21_ ( .D(n2832), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__21_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__22_ ( .D(n2831), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__22_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__23_ ( .D(n2830), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__23_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__25_ ( .D(n2829), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__25_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__26_ ( .D(n2828), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__26_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__31_ ( .D(n2827), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__31_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__1_ ( .D(n2826), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__1_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__2_ ( .D(n2825), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__2_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__3_ ( .D(n2824), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__3_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__5_ ( .D(n2823), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__5_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__10_ ( .D(n2822), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RSEL2__2_ ( .D(n2820), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RSEL2__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__LDBP2_ ( .D(n2818), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__LDBP2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__31_ ( .D(n2816), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[62]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_NEG_ ( .D(n2815), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_div0_r_NEG_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__31_ ( .D(n2813), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__31_ ( .D(n2812), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_QCORR_ ( .D(n18172), .CLK(
        clk), .QN(n2811) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__32_ ( .D(n2810), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[0]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__0_ ( .D(n2808), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__CWP__0_ ( .D(n2806), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__CWP__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__CWP__1_ ( .D(n2804), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__CWP__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CWP__1_ ( .D(n2800), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_E__CWP__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CWP__1_ ( .D(n2798), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__CWP__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RD__5_ ( .D(n2796), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RD__5_ ( .D(n2794), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RD__5_ ( .D(n2792), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RD__5_ ( .D(n2790), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CWP__0_ ( .D(n2786), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_E__CWP__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CWP__0_ ( .D(n2784), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__CWP__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA2__5_ ( .D(n2782), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA2__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA2__6_ ( .D(n2780), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA2__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA1__4_ ( .D(n2778), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA1__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA2__4_ ( .D(n2776), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA2__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA1__6_ ( .D(n2774), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA1__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA1__5_ ( .D(n2772), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA1__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__0_ ( .D(n2770), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__0_ ( .D(n2769), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__WIM__0_ ( .D(n2767), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__WIM__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TT__0_ ( .D(n2766), 
        .CLK(clk), .QN(irqo[0]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__YMSB_ ( .D(n2764), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__YMSB_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__0_ ( .D(n2762), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__30_ ( .D(n2760), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[61]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__30_ ( .D(n2758), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__30_ ( .D(n2757), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__SHCNT__4_ ( .D(n2755), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__SHCNT__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__4_ ( .D(n2753), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__4_ ( .D(n2751), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[35]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__4_ ( .D(n2749), .CLK(
        clk), .QN(u0_0_leon3x0_p0_muli[4]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__3_ ( .D(n2747), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[34]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__3_ ( .D(n2745), .CLK(
        clk), .QN(u0_0_leon3x0_p0_muli[3]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__35_ ( .D(n2744), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[3]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__3_ ( .D(n2742), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__3_ ( .D(n2740), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__3_ ( .D(n2739), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__WIM__3_ ( .D(n2737), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__WIM__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TT__3_ ( .D(n18051), 
        .CLK(clk), .QN(n2736) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__36_ ( .D(n2735), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[4]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__4_ ( .D(n2733), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__4_ ( .D(n2731), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__4_ ( .D(n2730), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__4_ ( .D(n2728), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__4_ ( .D(n2727), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__WIM__4_ ( .D(n2725), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__WIM__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TT__4_ ( .D(n2724), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TT__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__RD__7_ ( .D(n2722), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__RD__7_ ( .D(n2720), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__RD__7_ ( .D(n2718), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__RD__7_ ( .D(n2716), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__WREG_ ( .D(n2714), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__CTRL__WREG_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__WREG_ ( .D(n2712), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__CTRL__WREG_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__WREG_ ( .D(n2710), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__WREG_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__WREG_ ( .D(n2708), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__WREG_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFE1_ ( .D(n2706), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_E__RFE1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__0_ ( .D(
        n2705), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[36]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__SHCNT__0_ ( .D(n2703), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__SHCNT__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__0_ ( .D(n2701), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__0_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__1_ ( .D(n2700), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__1_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__5_ ( .D(n2699), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__5_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__7_ ( .D(n2698), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__7_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__1_ ( .D(n2697), .CLK(clk), .QN(
        irqctrl0_r_IPEND__1_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__5_ ( .D(n2696), .CLK(clk), .QN(
        irqctrl0_r_IPEND__5_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__7_ ( .D(n2695), .CLK(clk), .QN(
        irqctrl0_r_IPEND__7_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__2_ ( .D(n2694), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__2_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__4_ ( .D(n2693), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__4_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__4_ ( .D(n2692), .CLK(clk), .QN(
        irqctrl0_r_IPEND__4_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__15_ ( .D(n2691), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__15_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__15_ ( .D(n2690), .CLK(clk), .QN(
        irqctrl0_r_IPEND__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__5_ ( .D(n2688), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__6_ ( .D(
        n2687), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__6_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__6_ ( .D(
        n2686), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[3]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__CWP__2_ ( .D(n2684), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__CWP__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__7_ ( .D(n2683), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__8_ ( .D(n2682), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_X__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__12_ ( .D(n2681), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__12_ ( .D(n2680), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__0_ ( .D(n2679), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__12_ ( .D(n2677), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[70]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__12_ ( .D(n2675), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[40]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__12_ ( .D(n2673), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__12_ ( .D(n2671), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__12_ ( .D(n2669), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__12_ ( .D(n2667), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[9]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__12_ ( .D(n2665), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__12_ ( 
        .D(n2664), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__12_ ( 
        .D(n2663), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[9]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__12_ ( .D(n2662), .CLK(clk), .QN(
        apbi[38]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__12_ ( .D(n2660), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__45_ ( .D(n2659), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[13]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__13_ ( .D(n2657), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__13_ ( .D(n2656), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__1_ ( .D(n2655), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__13_ ( .D(n2653), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[71]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__13_ ( .D(n2651), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[41]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__13_ ( .D(n2649), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__13_ ( .D(n2647), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__13_ ( .D(n2645), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__13_ ( .D(n2643), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[10]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__13_ ( .D(n2641), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__13_ ( 
        .D(n2640), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__13_ ( 
        .D(n2639), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[10]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__13_ ( .D(n2638), .CLK(clk), .QN(
        apbi[39]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__13_ ( .D(n2636), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__13_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__16_ ( .D(n2635), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__17_ ( .D(n2634), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__18_ ( .D(n2633), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__16_ ( .D(n2632), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__4_ ( .D(n2631), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__4_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__16_ ( .D(n2629), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[74]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__16_ ( .D(n2627), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[44]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__16_ ( .D(n2625), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__16_ ( .D(n2623), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__16_ ( .D(n2621), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__16_ ( .D(n2619), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[13]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__16_ ( .D(n2617), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__16_ ( 
        .D(n2616), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__16_ ( 
        .D(n2615), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[13]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__16_ ( .D(n2614), .CLK(clk), .QN(
        apbi[42]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__16_ ( .D(n2612), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__49_ ( .D(n2611), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[17]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__17_ ( .D(n2609), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__17_ ( .D(n2608), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__5_ ( .D(n2607), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__5_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__17_ ( .D(n2605), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[75]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__17_ ( .D(n2603), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[45]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__17_ ( .D(n2601), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__17_ ( .D(n2599), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__17_ ( .D(n2597), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__17_ ( .D(n2595), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[14]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__17_ ( .D(n2593), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__17_ ( 
        .D(n2592), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__17_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__17_ ( 
        .D(n2591), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[14]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_HADDR__17_ ( .D(n2590), .CLK(clk), .QN(
        apbi[43]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__50_ ( .D(n2587), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[18]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__6_ ( .D(n2586), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__6_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__18_ ( .D(n2584), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[76]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__18_ ( .D(n2582), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[46]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__18_ ( .D(n2580), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__18_ ( .D(n2578), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__18_ ( .D(n2576), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__18_ ( .D(n2574), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[15]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__18_ ( .D(n2572), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__18_ ( 
        .D(n2571), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__18_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__18_ ( 
        .D(n2570), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[15]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__ADDR__18_ ( 
        .D(n2569), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[51]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFA1__3_ ( .D(n2567), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__RFA1__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__27_ ( .D(n24498), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__27_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__19_ ( .D(n2564), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__20_ ( .D(n2563), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__21_ ( .D(n2562), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__21_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__22_ ( .D(n2561), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__23_ ( .D(n2560), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__23_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__19_ ( .D(n2559), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__7_ ( .D(n2558), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__7_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__19_ ( .D(n2556), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[77]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__19_ ( .D(n2554), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[47]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__19_ ( .D(n2552), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__19_ ( .D(n2550), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__19_ ( .D(n2548), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__19_ ( .D(n2546), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[16]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__19_ ( .D(n2544), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__19_ ( 
        .D(n2543), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__19_ ( 
        .D(n2542), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[16]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__19_ ( .D(n2540), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__19_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__52_ ( .D(n2539), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[20]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__20_ ( .D(n2537), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__20_ ( .D(n2536), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__8_ ( .D(n2535), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__20_ ( .D(n2533), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[78]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__20_ ( .D(n2531), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[48]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__20_ ( .D(n2529), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__20_ ( .D(n2527), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__20_ ( .D(n2525), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__20_ ( .D(n2523), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[17]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__20_ ( .D(n2521), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__20_ ( 
        .D(n32534), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__20_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__20_ ( 
        .D(n31769), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[17]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__22_ ( .D(n2517), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__22_ ( .D(n2515), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[53]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__22_ ( .D(n2513), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__54_ ( .D(n2512), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[22]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__22_ ( .D(n2510), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__22_ ( .D(n2509), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__10_ ( .D(n2508), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__22_ ( .D(n2506), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[80]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__22_ ( .D(n2504), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[50]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__22_ ( .D(n2502), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__22_ ( .D(n2500), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__22_ ( .D(n2498), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__22_ ( .D(n2496), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[19]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__22_ ( .D(n2494), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__22_ ( 
        .D(n2493), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__22_ ( 
        .D(n2492), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[19]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__24_ ( .D(n2490), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__24_ ( .D(n2488), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[55]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__24_ ( .D(n2486), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__56_ ( .D(n2485), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[24]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__24_ ( .D(n2483), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__24_ ( .D(n2482), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__TBA__12_ ( .D(n2481), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__TBA__12_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__24_ ( .D(n2479), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[82]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__24_ ( .D(n2477), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[52]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__24_ ( .D(n2475), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__24_ ( .D(n2473), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__24_ ( .D(n2471), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__24_ ( .D(n2469), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[21]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__24_ ( .D(n2467), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__24_ ( 
        .D(n2466), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__24_ ( 
        .D(n2465), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[21]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__RFE2_ ( .D(n2463), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_E__RFE2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RCNT__4_ ( .D(n2462), .CLK(clk), .QN(
        uart1_r_RCNT__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RCNT__0_ ( .D(n2461), .CLK(clk), .QN(
        uart1_r_RCNT__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RCNT__1_ ( .D(n2460), .CLK(clk), .QN(
        uart1_r_RCNT__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RCNT__2_ ( .D(n2459), .CLK(clk), .QN(
        uart1_r_RCNT__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RCNT__3_ ( .D(n2458), .CLK(clk), .QN(
        uart1_r_RCNT__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RWADDR__4_ ( .D(n2457), .CLK(clk), .QN(
        uart1_r_RWADDR__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RWADDR__3_ ( .D(uart1_v_RWADDR__3_), .CLK(
        clk), .QN(n2456) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RWADDR__2_ ( .D(n2455), .CLK(clk), .QN(
        uart1_r_RWADDR__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RWADDR__1_ ( .D(n2454), .CLK(clk), .QN(
        uart1_r_RWADDR__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RWADDR__0_ ( .D(n2453), .CLK(clk), .QN(
        uart1_r_RWADDR__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__15__0_ ( .D(n2452), .CLK(clk), .QN(
        uart1_r_RHOLD__15__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__15__1_ ( .D(n2451), .CLK(clk), .QN(
        uart1_r_RHOLD__15__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__7__0_ ( .D(n2450), .CLK(clk), .QN(
        uart1_r_RHOLD__7__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__7__1_ ( .D(n2449), .CLK(clk), .QN(
        uart1_r_RHOLD__7__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__0__0_ ( .D(n2448), .CLK(clk), .QN(
        uart1_r_RHOLD__0__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__31__0_ ( .D(n2447), .CLK(clk), .QN(
        uart1_r_RHOLD__31__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__31__1_ ( .D(n2446), .CLK(clk), .QN(
        uart1_r_RHOLD__31__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__30__0_ ( .D(n2445), .CLK(clk), .QN(
        uart1_r_RHOLD__30__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__30__1_ ( .D(n2444), .CLK(clk), .QN(
        uart1_r_RHOLD__30__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__29__0_ ( .D(n2443), .CLK(clk), .QN(
        uart1_r_RHOLD__29__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__29__1_ ( .D(n2442), .CLK(clk), .QN(
        uart1_r_RHOLD__29__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__28__0_ ( .D(n2441), .CLK(clk), .QN(
        uart1_r_RHOLD__28__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__28__1_ ( .D(n2440), .CLK(clk), .QN(
        uart1_r_RHOLD__28__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__27__0_ ( .D(n2439), .CLK(clk), .QN(
        uart1_r_RHOLD__27__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__27__1_ ( .D(n2438), .CLK(clk), .QN(
        uart1_r_RHOLD__27__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__26__0_ ( .D(n2437), .CLK(clk), .QN(
        uart1_r_RHOLD__26__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__26__1_ ( .D(n2436), .CLK(clk), .QN(
        uart1_r_RHOLD__26__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__25__0_ ( .D(n2435), .CLK(clk), .QN(
        uart1_r_RHOLD__25__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__25__1_ ( .D(n2434), .CLK(clk), .QN(
        uart1_r_RHOLD__25__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__24__0_ ( .D(n2433), .CLK(clk), .QN(
        uart1_r_RHOLD__24__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__24__1_ ( .D(n2432), .CLK(clk), .QN(
        uart1_r_RHOLD__24__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__23__0_ ( .D(n2431), .CLK(clk), .QN(
        uart1_r_RHOLD__23__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__23__1_ ( .D(n2430), .CLK(clk), .QN(
        uart1_r_RHOLD__23__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__22__0_ ( .D(n2429), .CLK(clk), .QN(
        uart1_r_RHOLD__22__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__22__1_ ( .D(n2428), .CLK(clk), .QN(
        uart1_r_RHOLD__22__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__21__0_ ( .D(n2427), .CLK(clk), .QN(
        uart1_r_RHOLD__21__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__21__1_ ( .D(n2426), .CLK(clk), .QN(
        uart1_r_RHOLD__21__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__20__0_ ( .D(n2425), .CLK(clk), .QN(
        uart1_r_RHOLD__20__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__20__1_ ( .D(n2424), .CLK(clk), .QN(
        uart1_r_RHOLD__20__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__19__0_ ( .D(n2423), .CLK(clk), .QN(
        uart1_r_RHOLD__19__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__19__1_ ( .D(n2422), .CLK(clk), .QN(
        uart1_r_RHOLD__19__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__18__0_ ( .D(n2421), .CLK(clk), .QN(
        uart1_r_RHOLD__18__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__18__1_ ( .D(n2420), .CLK(clk), .QN(
        uart1_r_RHOLD__18__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__17__0_ ( .D(n2419), .CLK(clk), .QN(
        uart1_r_RHOLD__17__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__17__1_ ( .D(n2418), .CLK(clk), .QN(
        uart1_r_RHOLD__17__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__16__0_ ( .D(n2417), .CLK(clk), .QN(
        uart1_r_RHOLD__16__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__16__1_ ( .D(n2416), .CLK(clk), .QN(
        uart1_r_RHOLD__16__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__14__0_ ( .D(n2415), .CLK(clk), .QN(
        uart1_r_RHOLD__14__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__14__1_ ( .D(n2414), .CLK(clk), .QN(
        uart1_r_RHOLD__14__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__13__0_ ( .D(n2413), .CLK(clk), .QN(
        uart1_r_RHOLD__13__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__13__1_ ( .D(n2412), .CLK(clk), .QN(
        uart1_r_RHOLD__13__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__12__0_ ( .D(n2411), .CLK(clk), .QN(
        uart1_r_RHOLD__12__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__12__1_ ( .D(n2410), .CLK(clk), .QN(
        uart1_r_RHOLD__12__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__11__0_ ( .D(n2409), .CLK(clk), .QN(
        uart1_r_RHOLD__11__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__11__1_ ( .D(n2408), .CLK(clk), .QN(
        uart1_r_RHOLD__11__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__10__0_ ( .D(n2407), .CLK(clk), .QN(
        uart1_r_RHOLD__10__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__10__1_ ( .D(n2406), .CLK(clk), .QN(
        uart1_r_RHOLD__10__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__9__0_ ( .D(n2405), .CLK(clk), .QN(
        uart1_r_RHOLD__9__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__9__1_ ( .D(n2404), .CLK(clk), .QN(
        uart1_r_RHOLD__9__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__8__0_ ( .D(n2403), .CLK(clk), .QN(
        uart1_r_RHOLD__8__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__8__1_ ( .D(n2402), .CLK(clk), .QN(
        uart1_r_RHOLD__8__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__6__0_ ( .D(n2401), .CLK(clk), .QN(
        uart1_r_RHOLD__6__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__6__1_ ( .D(n2400), .CLK(clk), .QN(
        uart1_r_RHOLD__6__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__5__0_ ( .D(n2399), .CLK(clk), .QN(
        uart1_r_RHOLD__5__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__5__1_ ( .D(n2398), .CLK(clk), .QN(
        uart1_r_RHOLD__5__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__4__0_ ( .D(n2397), .CLK(clk), .QN(
        uart1_r_RHOLD__4__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__4__1_ ( .D(n2396), .CLK(clk), .QN(
        uart1_r_RHOLD__4__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__3__0_ ( .D(n2395), .CLK(clk), .QN(
        uart1_r_RHOLD__3__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__3__1_ ( .D(n2394), .CLK(clk), .QN(
        uart1_r_RHOLD__3__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__2__0_ ( .D(n2393), .CLK(clk), .QN(
        uart1_r_RHOLD__2__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__2__1_ ( .D(n2392), .CLK(clk), .QN(
        uart1_r_RHOLD__2__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__1__0_ ( .D(n2391), .CLK(clk), .QN(
        uart1_r_RHOLD__1__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__1__1_ ( .D(n2390), .CLK(clk), .QN(
        uart1_r_RHOLD__1__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RRADDR__0_ ( .D(n17459), .CLK(clk), .QN(
        n2389) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RRADDR__1_ ( .D(n17458), .CLK(clk), .QN(
        n2388) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RRADDR__2_ ( .D(n17457), .CLK(clk), .QN(
        n2387) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RRADDR__3_ ( .D(n17456), .CLK(clk), .QN(
        n2386) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__10_ ( .D(n2385), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__10_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__10_ ( .D(n2384), .CLK(clk), .QN(
        irqctrl0_r_IPEND__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__PC__30_ ( .D(n2382), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[58]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__PC__30_ ( .D(n2380), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__PC__30_ ( .D(n2378), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__PC__30_ ( .D(n2376), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__PC__30_ ( .D(n2374), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_ici[27]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__30_ ( .D(n2372), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__30_ ( 
        .D(n32557), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__30_ ( 
        .D(n31998), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[27]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_QMSB_ ( .D(n2369), .CLK(clk), .QN(u0_0_leon3x0_p0_div0_r_QMSB_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__ICC__3_ ( .D(n2367), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__ICC__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__ICC__3_ ( .D(n2366), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__ICC__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VADDRESS__31_ ( 
        .D(n2365), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_WADDRESS__31_ ( 
        .D(n2364), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcii[28]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_HWRITE_ ( .D(n2363), .CLK(clk), .QN(
        sr1_sdi_HWRITE_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_SIZE__0_ ( .D(n2362), .CLK(clk), .QN(
        sr1_sdi_HSIZE__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_SIZE__1_ ( .D(n2361), .CLK(clk), .QN(
        sr1_sdi_HSIZE__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_SRHSEL_ ( .D(n2358), .CLK(clk), .QN(
        sr1_r_SRHSEL_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_BRMW_ ( .D(n17778), .CLK(clk), .QN(n2357) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_AREA__1_ ( .D(n17904), .CLK(clk), .QN(n2356)
         );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_AREA__0_ ( .D(n2355), .CLK(clk), .QN(
        sr1_r_AREA__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__IMM__28_ ( .D(n24496), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_A__IMM__28_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__19_ ( 
        .D(n2352), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[23]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__19_ ( .D(n2351), .CLK(clk), .QN(
        apbi[19]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__IOEN_ ( .D(n2350), .CLK(clk), .QN(
        sr1_r_MCFG1__IOEN_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__3_ ( .D(n2349), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__3_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__3_ ( .D(n2348), .CLK(clk), .QN(
        irqctrl0_r_IPEND__3_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__19_ ( .D(n2347), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__19_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__IRQ_ ( .D(n2346), .CLK(clk), 
        .QN(timer0_gpto_TICK__1_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__6_ ( .D(n2345), .CLK(clk), .QN(
        ahb0_r_HADDR__6_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__1_ ( .D(n33062), .CLK(clk), .QN(
        ahb0_r_HRDATAS__1_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__15_ ( .D(n2333), .CLK(clk), .QN(
        ahb0_r_HRDATAS__15_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__4_ ( .D(n33063), .CLK(clk), .QN(
        ahb0_r_HRDATAS__4_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__13_ ( .D(n2330), .CLK(clk), .QN(
        ahb0_r_HRDATAS__13_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__14_ ( .D(n2329), .CLK(clk), .QN(
        ahb0_r_HRDATAS__14_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__21_ ( 
        .D(n2328), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[25]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__14_ ( 
        .D(n2327), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[18]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__14_ ( .D(n2326), .CLK(clk), .QN(
        apbi[14]) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSEMPTYIRQEN_ ( .D(n2325), .CLK(clk), .QN(
        uart1_r_TSEMPTYIRQEN_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__14_ ( .D(n2324), .CLK(clk), 
        .QN(irqctrl0_r_ILEVEL__14_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__14_ ( .D(n2323), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__14_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__14_ ( .D(
        timer0_v_TIMERS__1__VALUE__14_), .CLK(clk), .QN(n2322) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__15_ ( .D(n2321), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__15_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__8_ ( .D(n2319), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__8_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__41_ ( .D(n2318), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[9]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__RESULT__9_ ( .D(n2316), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__RESULT__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__RESULT__9_ ( .D(n2314), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__RESULT__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__9_ ( .D(n2313), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__PIL__1_ ( .D(n2312), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__PIL__1_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__9_ ( .D(n2310), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__30_ ( .D(n2309), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__30_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__31_ ( .D(n2308), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__64_ ( .D(n18168), .CLK(
        clk), .QN(n2307) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_QZERO_ ( .D(n2306), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divo[32]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_IOSN__0_ ( .D(n2304), .CLK(clk), .RESET(
        n18295), .SET(n24695), .QN(iosn) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_IOSN__1_ ( .D(n2302), .CLK(clk), .RESET(
        n18295), .SET(n24695), .QN(sr1_r_IOSN__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEN_ ( .D(n2301), .CLK(clk), .QN(writen)
         );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_BDRIVE__0_ ( .D(n2299), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(datadir[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_BDRIVE__1_ ( .D(n2297), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(datadir[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_BDRIVE__2_ ( .D(n2295), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(datadir[2]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_BDRIVE__3_ ( .D(n2293), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(datadir[3]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_AREA__2_ ( .D(n17903), .CLK(clk), .QN(n2292)
         );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_BUSW__0_ ( .D(n2291), .CLK(clk), .QN(
        sr1_r_BUSW__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_HCACHE_ ( .D(n2290), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_a0_r_HCACHE_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_HIT_ ( .D(n2289), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_HIT_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VALID__0__4_ ( .D(
        n2288), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__4_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VALID__0__0_ ( .D(
        n2287), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__0_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VALID__0__1_ ( .D(
        n2286), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__1_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VALID__0__2_ ( .D(
        n2285), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__2_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VALID__0__3_ ( .D(
        n2284), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__3_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VALID__0__5_ ( .D(
        n2283), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__5_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VALID__0__6_ ( .D(
        n2282), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__6_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_VALID__0__7_ ( .D(
        n2281), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__7_)
         );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__ICC__0_ ( .D(n2279), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__ICC__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__ICC__0_ ( .D(n2278), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__ICC__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__ALUCIN_ ( .D(n2276), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__ALUCIN_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_div0_r_reg_X__24_ ( .D(n2275), .CLK(
        clk), .QN(u0_0_leon3x0_p0_div0_r_X__24_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__24_ ( 
        .D(n2274), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[28]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__24_ ( .D(n2273), .CLK(clk), .QN(
        apbi[24]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__24_ ( .D(n2272), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__24_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__24_ ( .D(
        timer0_v_TIMERS__1__VALUE__24_), .CLK(clk), .QN(n2271) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TWADDR__0_ ( .D(n2270), .CLK(clk), .QN(
        uart1_r_TWADDR__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TWADDR__1_ ( .D(n2269), .CLK(clk), .QN(
        uart1_r_TWADDR__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TWADDR__2_ ( .D(n2268), .CLK(clk), .QN(
        uart1_r_TWADDR__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TWADDR__3_ ( .D(n17717), .CLK(clk), .QN(
        n2267) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TWADDR__4_ ( .D(n2266), .CLK(clk), .QN(
        uart1_r_TWADDR__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__24__0_ ( .D(n2265), .CLK(clk), .QN(
        uart1_r_THOLD__24__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__22__0_ ( .D(n2264), .CLK(clk), .QN(
        uart1_r_THOLD__22__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__21__0_ ( .D(n2263), .CLK(clk), .QN(
        uart1_r_THOLD__21__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__19__0_ ( .D(n2262), .CLK(clk), .QN(
        uart1_r_THOLD__19__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__16__0_ ( .D(n2261), .CLK(clk), .QN(
        uart1_r_THOLD__16__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__14__0_ ( .D(n2260), .CLK(clk), .QN(
        uart1_r_THOLD__14__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__13__0_ ( .D(n2259), .CLK(clk), .QN(
        uart1_r_THOLD__13__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__12__0_ ( .D(n2258), .CLK(clk), .QN(
        uart1_r_THOLD__12__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__11__0_ ( .D(n2257), .CLK(clk), .QN(
        uart1_r_THOLD__11__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__10__0_ ( .D(n2256), .CLK(clk), .QN(
        uart1_r_THOLD__10__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__9__0_ ( .D(n2255), .CLK(clk), .QN(
        uart1_r_THOLD__9__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__8__0_ ( .D(n2254), .CLK(clk), .QN(
        uart1_r_THOLD__8__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__6__0_ ( .D(n2253), .CLK(clk), .QN(
        uart1_r_THOLD__6__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__5__0_ ( .D(n2252), .CLK(clk), .QN(
        uart1_r_THOLD__5__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__4__0_ ( .D(n2251), .CLK(clk), .QN(
        uart1_r_THOLD__4__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__3__0_ ( .D(n2250), .CLK(clk), .QN(
        uart1_r_THOLD__3__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__2__0_ ( .D(n2249), .CLK(clk), .QN(
        uart1_r_THOLD__2__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__1__0_ ( .D(n2248), .CLK(clk), .QN(
        uart1_r_THOLD__1__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__0__0_ ( .D(n2247), .CLK(clk), .QN(
        uart1_r_THOLD__0__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TXCLK__0_ ( .D(n2246), .CLK(clk), .QN(
        uart1_r_TXCLK__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TXCLK__1_ ( .D(n2245), .CLK(clk), .QN(
        uart1_r_TXCLK__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TXCLK__2_ ( .D(uart1_v_TXCLK__2_), .CLK(
        clk), .QN(n5014) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TSEMPTY_ ( .D(n2243), .CLK(clk), .QN(
        uart1_r_TSEMPTY_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TRADDR__4_ ( .D(n2242), .CLK(clk), .QN(
        uart1_r_TRADDR__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TRADDR__3_ ( .D(n2241), .CLK(clk), .QN(
        uart1_r_TRADDR__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TRADDR__2_ ( .D(n2240), .CLK(clk), .QN(
        uart1_r_TRADDR__2_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__11_ ( .D(n17802), .CLK(clk), 
        .QN(n2236) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__11_ ( .D(n17857), .CLK(clk), 
        .QN(n2235) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__11_ ( .D(n2234), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__11_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__11_ ( .D(
        timer0_v_TIMERS__1__VALUE__11_), .CLK(clk), .QN(n2233) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__27_ ( .D(n2232), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__27_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_RELOAD__1_ ( .D(n2231), .CLK(clk), .QN(
        timer0_r_RELOAD__1_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_SCALER__1_ ( .D(n2230), .CLK(clk), .QN(
        timer0_r_SCALER__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__31__2_ ( .D(n2229), .CLK(clk), .QN(
        uart1_r_RHOLD__31__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__30__2_ ( .D(n2228), .CLK(clk), .QN(
        uart1_r_RHOLD__30__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__29__2_ ( .D(n2227), .CLK(clk), .QN(
        uart1_r_RHOLD__29__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__28__2_ ( .D(n2226), .CLK(clk), .QN(
        uart1_r_RHOLD__28__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__27__2_ ( .D(n2225), .CLK(clk), .QN(
        uart1_r_RHOLD__27__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__26__2_ ( .D(n2224), .CLK(clk), .QN(
        uart1_r_RHOLD__26__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__25__2_ ( .D(n2223), .CLK(clk), .QN(
        uart1_r_RHOLD__25__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__24__2_ ( .D(n2222), .CLK(clk), .QN(
        uart1_r_RHOLD__24__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__23__2_ ( .D(n2221), .CLK(clk), .QN(
        uart1_r_RHOLD__23__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__22__2_ ( .D(n2220), .CLK(clk), .QN(
        uart1_r_RHOLD__22__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__21__2_ ( .D(n2219), .CLK(clk), .QN(
        uart1_r_RHOLD__21__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__20__2_ ( .D(n2218), .CLK(clk), .QN(
        uart1_r_RHOLD__20__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__19__2_ ( .D(n2217), .CLK(clk), .QN(
        uart1_r_RHOLD__19__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__18__2_ ( .D(n2216), .CLK(clk), .QN(
        uart1_r_RHOLD__18__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__17__2_ ( .D(n2215), .CLK(clk), .QN(
        uart1_r_RHOLD__17__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__16__2_ ( .D(n2214), .CLK(clk), .QN(
        uart1_r_RHOLD__16__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__15__2_ ( .D(n2213), .CLK(clk), .QN(
        uart1_r_RHOLD__15__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__14__2_ ( .D(n2212), .CLK(clk), .QN(
        uart1_r_RHOLD__14__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__13__2_ ( .D(n2211), .CLK(clk), .QN(
        uart1_r_RHOLD__13__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__12__2_ ( .D(n2210), .CLK(clk), .QN(
        uart1_r_RHOLD__12__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__11__2_ ( .D(n2209), .CLK(clk), .QN(
        uart1_r_RHOLD__11__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__10__2_ ( .D(n2208), .CLK(clk), .QN(
        uart1_r_RHOLD__10__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__9__2_ ( .D(n2207), .CLK(clk), .QN(
        uart1_r_RHOLD__9__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__8__2_ ( .D(n2206), .CLK(clk), .QN(
        uart1_r_RHOLD__8__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__7__2_ ( .D(n2205), .CLK(clk), .QN(
        uart1_r_RHOLD__7__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__6__2_ ( .D(n2204), .CLK(clk), .QN(
        uart1_r_RHOLD__6__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__5__2_ ( .D(n2203), .CLK(clk), .QN(
        uart1_r_RHOLD__5__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__4__2_ ( .D(n2202), .CLK(clk), .QN(
        uart1_r_RHOLD__4__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__3__2_ ( .D(n2201), .CLK(clk), .QN(
        uart1_r_RHOLD__3__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__2__2_ ( .D(n2200), .CLK(clk), .QN(
        uart1_r_RHOLD__2__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__1__2_ ( .D(n2199), .CLK(clk), .QN(
        uart1_r_RHOLD__1__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__31__3_ ( .D(n2198), .CLK(clk), .QN(
        uart1_r_RHOLD__31__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__30__3_ ( .D(n2197), .CLK(clk), .QN(
        uart1_r_RHOLD__30__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__29__3_ ( .D(n2196), .CLK(clk), .QN(
        uart1_r_RHOLD__29__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__28__3_ ( .D(n2195), .CLK(clk), .QN(
        uart1_r_RHOLD__28__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__27__3_ ( .D(n2194), .CLK(clk), .QN(
        uart1_r_RHOLD__27__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__26__3_ ( .D(n2193), .CLK(clk), .QN(
        uart1_r_RHOLD__26__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__25__3_ ( .D(n2192), .CLK(clk), .QN(
        uart1_r_RHOLD__25__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__24__3_ ( .D(n2191), .CLK(clk), .QN(
        uart1_r_RHOLD__24__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__23__3_ ( .D(n2190), .CLK(clk), .QN(
        uart1_r_RHOLD__23__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__22__3_ ( .D(n2189), .CLK(clk), .QN(
        uart1_r_RHOLD__22__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__21__3_ ( .D(n2188), .CLK(clk), .QN(
        uart1_r_RHOLD__21__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__20__3_ ( .D(n2187), .CLK(clk), .QN(
        uart1_r_RHOLD__20__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__19__3_ ( .D(n2186), .CLK(clk), .QN(
        uart1_r_RHOLD__19__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__18__3_ ( .D(n2185), .CLK(clk), .QN(
        uart1_r_RHOLD__18__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__17__3_ ( .D(n2184), .CLK(clk), .QN(
        uart1_r_RHOLD__17__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__16__3_ ( .D(n2183), .CLK(clk), .QN(
        uart1_r_RHOLD__16__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__15__3_ ( .D(n2182), .CLK(clk), .QN(
        uart1_r_RHOLD__15__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__14__3_ ( .D(n2181), .CLK(clk), .QN(
        uart1_r_RHOLD__14__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__13__3_ ( .D(n2180), .CLK(clk), .QN(
        uart1_r_RHOLD__13__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__12__3_ ( .D(n2179), .CLK(clk), .QN(
        uart1_r_RHOLD__12__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__11__3_ ( .D(n2178), .CLK(clk), .QN(
        uart1_r_RHOLD__11__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__10__3_ ( .D(n2177), .CLK(clk), .QN(
        uart1_r_RHOLD__10__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__9__3_ ( .D(n2176), .CLK(clk), .QN(
        uart1_r_RHOLD__9__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__8__3_ ( .D(n2175), .CLK(clk), .QN(
        uart1_r_RHOLD__8__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__7__3_ ( .D(n2174), .CLK(clk), .QN(
        uart1_r_RHOLD__7__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__6__3_ ( .D(n2173), .CLK(clk), .QN(
        uart1_r_RHOLD__6__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__5__3_ ( .D(n2172), .CLK(clk), .QN(
        uart1_r_RHOLD__5__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__4__3_ ( .D(n2171), .CLK(clk), .QN(
        uart1_r_RHOLD__4__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__3__3_ ( .D(n2170), .CLK(clk), .QN(
        uart1_r_RHOLD__3__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__2__3_ ( .D(n2169), .CLK(clk), .QN(
        uart1_r_RHOLD__2__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__1__3_ ( .D(n2168), .CLK(clk), .QN(
        uart1_r_RHOLD__1__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__31__4_ ( .D(n2167), .CLK(clk), .QN(
        uart1_r_RHOLD__31__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__30__4_ ( .D(n2166), .CLK(clk), .QN(
        uart1_r_RHOLD__30__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__29__4_ ( .D(n2165), .CLK(clk), .QN(
        uart1_r_RHOLD__29__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__28__4_ ( .D(n2164), .CLK(clk), .QN(
        uart1_r_RHOLD__28__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__27__4_ ( .D(n2163), .CLK(clk), .QN(
        uart1_r_RHOLD__27__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__26__4_ ( .D(n2162), .CLK(clk), .QN(
        uart1_r_RHOLD__26__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__25__4_ ( .D(n2161), .CLK(clk), .QN(
        uart1_r_RHOLD__25__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__24__4_ ( .D(n2160), .CLK(clk), .QN(
        uart1_r_RHOLD__24__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__23__4_ ( .D(n2159), .CLK(clk), .QN(
        uart1_r_RHOLD__23__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__22__4_ ( .D(n2158), .CLK(clk), .QN(
        uart1_r_RHOLD__22__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__21__4_ ( .D(n2157), .CLK(clk), .QN(
        uart1_r_RHOLD__21__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__20__4_ ( .D(n2156), .CLK(clk), .QN(
        uart1_r_RHOLD__20__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__19__4_ ( .D(n2155), .CLK(clk), .QN(
        uart1_r_RHOLD__19__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__18__4_ ( .D(n2154), .CLK(clk), .QN(
        uart1_r_RHOLD__18__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__17__4_ ( .D(n2153), .CLK(clk), .QN(
        uart1_r_RHOLD__17__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__16__4_ ( .D(n2152), .CLK(clk), .QN(
        uart1_r_RHOLD__16__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__15__4_ ( .D(n2151), .CLK(clk), .QN(
        uart1_r_RHOLD__15__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__14__4_ ( .D(n2150), .CLK(clk), .QN(
        uart1_r_RHOLD__14__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__13__4_ ( .D(n2149), .CLK(clk), .QN(
        uart1_r_RHOLD__13__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__12__4_ ( .D(n2148), .CLK(clk), .QN(
        uart1_r_RHOLD__12__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__11__4_ ( .D(n2147), .CLK(clk), .QN(
        uart1_r_RHOLD__11__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__10__4_ ( .D(n2146), .CLK(clk), .QN(
        uart1_r_RHOLD__10__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__9__4_ ( .D(n2145), .CLK(clk), .QN(
        uart1_r_RHOLD__9__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__8__4_ ( .D(n2144), .CLK(clk), .QN(
        uart1_r_RHOLD__8__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__7__4_ ( .D(n2143), .CLK(clk), .QN(
        uart1_r_RHOLD__7__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__6__4_ ( .D(n2142), .CLK(clk), .QN(
        uart1_r_RHOLD__6__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__5__4_ ( .D(n2141), .CLK(clk), .QN(
        uart1_r_RHOLD__5__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__4__4_ ( .D(n2140), .CLK(clk), .QN(
        uart1_r_RHOLD__4__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__3__4_ ( .D(n2139), .CLK(clk), .QN(
        uart1_r_RHOLD__3__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__2__4_ ( .D(n2138), .CLK(clk), .QN(
        uart1_r_RHOLD__2__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__1__4_ ( .D(n2137), .CLK(clk), .QN(
        uart1_r_RHOLD__1__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__31__5_ ( .D(n2136), .CLK(clk), .QN(
        uart1_r_RHOLD__31__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__30__5_ ( .D(n2135), .CLK(clk), .QN(
        uart1_r_RHOLD__30__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__29__5_ ( .D(n2134), .CLK(clk), .QN(
        uart1_r_RHOLD__29__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__28__5_ ( .D(n2133), .CLK(clk), .QN(
        uart1_r_RHOLD__28__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__27__5_ ( .D(n2132), .CLK(clk), .QN(
        uart1_r_RHOLD__27__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__26__5_ ( .D(n2131), .CLK(clk), .QN(
        uart1_r_RHOLD__26__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__25__5_ ( .D(n2130), .CLK(clk), .QN(
        uart1_r_RHOLD__25__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__24__5_ ( .D(n2129), .CLK(clk), .QN(
        uart1_r_RHOLD__24__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__23__5_ ( .D(n2128), .CLK(clk), .QN(
        uart1_r_RHOLD__23__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__22__5_ ( .D(n2127), .CLK(clk), .QN(
        uart1_r_RHOLD__22__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__21__5_ ( .D(n2126), .CLK(clk), .QN(
        uart1_r_RHOLD__21__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__20__5_ ( .D(n2125), .CLK(clk), .QN(
        uart1_r_RHOLD__20__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__19__5_ ( .D(n2124), .CLK(clk), .QN(
        uart1_r_RHOLD__19__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__18__5_ ( .D(n2123), .CLK(clk), .QN(
        uart1_r_RHOLD__18__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__17__5_ ( .D(n2122), .CLK(clk), .QN(
        uart1_r_RHOLD__17__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__16__5_ ( .D(n2121), .CLK(clk), .QN(
        uart1_r_RHOLD__16__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__15__5_ ( .D(n2120), .CLK(clk), .QN(
        uart1_r_RHOLD__15__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__14__5_ ( .D(n2119), .CLK(clk), .QN(
        uart1_r_RHOLD__14__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__13__5_ ( .D(n2118), .CLK(clk), .QN(
        uart1_r_RHOLD__13__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__12__5_ ( .D(n2117), .CLK(clk), .QN(
        uart1_r_RHOLD__12__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__11__5_ ( .D(n2116), .CLK(clk), .QN(
        uart1_r_RHOLD__11__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__10__5_ ( .D(n2115), .CLK(clk), .QN(
        uart1_r_RHOLD__10__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__9__5_ ( .D(n2114), .CLK(clk), .QN(
        uart1_r_RHOLD__9__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__8__5_ ( .D(n2113), .CLK(clk), .QN(
        uart1_r_RHOLD__8__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__7__5_ ( .D(n2112), .CLK(clk), .QN(
        uart1_r_RHOLD__7__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__6__5_ ( .D(n2111), .CLK(clk), .QN(
        uart1_r_RHOLD__6__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__5__5_ ( .D(n2110), .CLK(clk), .QN(
        uart1_r_RHOLD__5__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__4__5_ ( .D(n2109), .CLK(clk), .QN(
        uart1_r_RHOLD__4__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__3__5_ ( .D(n2108), .CLK(clk), .QN(
        uart1_r_RHOLD__3__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__2__5_ ( .D(n2107), .CLK(clk), .QN(
        uart1_r_RHOLD__2__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__1__5_ ( .D(n2106), .CLK(clk), .QN(
        uart1_r_RHOLD__1__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__31__6_ ( .D(n2105), .CLK(clk), .QN(
        uart1_r_RHOLD__31__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__30__6_ ( .D(n2104), .CLK(clk), .QN(
        uart1_r_RHOLD__30__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__29__6_ ( .D(n2103), .CLK(clk), .QN(
        uart1_r_RHOLD__29__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__28__6_ ( .D(n2102), .CLK(clk), .QN(
        uart1_r_RHOLD__28__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__27__6_ ( .D(n2101), .CLK(clk), .QN(
        uart1_r_RHOLD__27__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__26__6_ ( .D(n2100), .CLK(clk), .QN(
        uart1_r_RHOLD__26__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__25__6_ ( .D(n2099), .CLK(clk), .QN(
        uart1_r_RHOLD__25__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__24__6_ ( .D(n2098), .CLK(clk), .QN(
        uart1_r_RHOLD__24__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__23__6_ ( .D(n2097), .CLK(clk), .QN(
        uart1_r_RHOLD__23__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__22__6_ ( .D(n2096), .CLK(clk), .QN(
        uart1_r_RHOLD__22__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__21__6_ ( .D(n2095), .CLK(clk), .QN(
        uart1_r_RHOLD__21__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__20__6_ ( .D(n2094), .CLK(clk), .QN(
        uart1_r_RHOLD__20__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__19__6_ ( .D(n2093), .CLK(clk), .QN(
        uart1_r_RHOLD__19__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__18__6_ ( .D(n2092), .CLK(clk), .QN(
        uart1_r_RHOLD__18__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__17__6_ ( .D(n2091), .CLK(clk), .QN(
        uart1_r_RHOLD__17__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__16__6_ ( .D(n2090), .CLK(clk), .QN(
        uart1_r_RHOLD__16__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__15__6_ ( .D(n2089), .CLK(clk), .QN(
        uart1_r_RHOLD__15__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__14__6_ ( .D(n2088), .CLK(clk), .QN(
        uart1_r_RHOLD__14__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__13__6_ ( .D(n2087), .CLK(clk), .QN(
        uart1_r_RHOLD__13__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__12__6_ ( .D(n2086), .CLK(clk), .QN(
        uart1_r_RHOLD__12__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__11__6_ ( .D(n2085), .CLK(clk), .QN(
        uart1_r_RHOLD__11__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__10__6_ ( .D(n2084), .CLK(clk), .QN(
        uart1_r_RHOLD__10__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__9__6_ ( .D(n2083), .CLK(clk), .QN(
        uart1_r_RHOLD__9__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__8__6_ ( .D(n2082), .CLK(clk), .QN(
        uart1_r_RHOLD__8__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__7__6_ ( .D(n2081), .CLK(clk), .QN(
        uart1_r_RHOLD__7__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__6__6_ ( .D(n2080), .CLK(clk), .QN(
        uart1_r_RHOLD__6__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__5__6_ ( .D(n2079), .CLK(clk), .QN(
        uart1_r_RHOLD__5__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__4__6_ ( .D(n2078), .CLK(clk), .QN(
        uart1_r_RHOLD__4__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__3__6_ ( .D(n2077), .CLK(clk), .QN(
        uart1_r_RHOLD__3__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__2__6_ ( .D(n2076), .CLK(clk), .QN(
        uart1_r_RHOLD__2__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__1__6_ ( .D(n2075), .CLK(clk), .QN(
        uart1_r_RHOLD__1__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__31__7_ ( .D(n2074), .CLK(clk), .QN(
        uart1_r_RHOLD__31__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__30__7_ ( .D(n2073), .CLK(clk), .QN(
        uart1_r_RHOLD__30__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__29__7_ ( .D(n2072), .CLK(clk), .QN(
        uart1_r_RHOLD__29__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__28__7_ ( .D(n2071), .CLK(clk), .QN(
        uart1_r_RHOLD__28__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__27__7_ ( .D(n2070), .CLK(clk), .QN(
        uart1_r_RHOLD__27__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__26__7_ ( .D(n2069), .CLK(clk), .QN(
        uart1_r_RHOLD__26__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__25__7_ ( .D(n2068), .CLK(clk), .QN(
        uart1_r_RHOLD__25__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__24__7_ ( .D(n2067), .CLK(clk), .QN(
        uart1_r_RHOLD__24__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__23__7_ ( .D(n2066), .CLK(clk), .QN(
        uart1_r_RHOLD__23__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__22__7_ ( .D(n2065), .CLK(clk), .QN(
        uart1_r_RHOLD__22__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__21__7_ ( .D(n2064), .CLK(clk), .QN(
        uart1_r_RHOLD__21__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__20__7_ ( .D(n2063), .CLK(clk), .QN(
        uart1_r_RHOLD__20__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__19__7_ ( .D(n2062), .CLK(clk), .QN(
        uart1_r_RHOLD__19__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__18__7_ ( .D(n2061), .CLK(clk), .QN(
        uart1_r_RHOLD__18__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__17__7_ ( .D(n2060), .CLK(clk), .QN(
        uart1_r_RHOLD__17__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__16__7_ ( .D(n2059), .CLK(clk), .QN(
        uart1_r_RHOLD__16__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__15__7_ ( .D(n2058), .CLK(clk), .QN(
        uart1_r_RHOLD__15__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__14__7_ ( .D(n2057), .CLK(clk), .QN(
        uart1_r_RHOLD__14__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__13__7_ ( .D(n2056), .CLK(clk), .QN(
        uart1_r_RHOLD__13__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__12__7_ ( .D(n2055), .CLK(clk), .QN(
        uart1_r_RHOLD__12__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__11__7_ ( .D(n2054), .CLK(clk), .QN(
        uart1_r_RHOLD__11__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__10__7_ ( .D(n2053), .CLK(clk), .QN(
        uart1_r_RHOLD__10__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__9__7_ ( .D(n2052), .CLK(clk), .QN(
        uart1_r_RHOLD__9__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__8__7_ ( .D(n2051), .CLK(clk), .QN(
        uart1_r_RHOLD__8__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__7__7_ ( .D(n2050), .CLK(clk), .QN(
        uart1_r_RHOLD__7__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__6__7_ ( .D(n2049), .CLK(clk), .QN(
        uart1_r_RHOLD__6__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__5__7_ ( .D(n2048), .CLK(clk), .QN(
        uart1_r_RHOLD__5__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__4__7_ ( .D(n2047), .CLK(clk), .QN(
        uart1_r_RHOLD__4__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__3__7_ ( .D(n2046), .CLK(clk), .QN(
        uart1_r_RHOLD__3__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__2__7_ ( .D(n2045), .CLK(clk), .QN(
        uart1_r_RHOLD__2__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__1__7_ ( .D(n2044), .CLK(clk), .QN(
        uart1_r_RHOLD__1__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__31__0_ ( .D(n2043), .CLK(clk), .QN(
        uart1_r_THOLD__31__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__31__1_ ( .D(n2042), .CLK(clk), .QN(
        uart1_r_THOLD__31__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__31__2_ ( .D(n2041), .CLK(clk), .QN(
        uart1_r_THOLD__31__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__31__3_ ( .D(n2040), .CLK(clk), .QN(
        uart1_r_THOLD__31__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__31__4_ ( .D(n2039), .CLK(clk), .QN(
        uart1_r_THOLD__31__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__31__5_ ( .D(n2038), .CLK(clk), .QN(
        uart1_r_THOLD__31__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__31__6_ ( .D(n2037), .CLK(clk), .QN(
        uart1_r_THOLD__31__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__31__7_ ( .D(n2036), .CLK(clk), .QN(
        uart1_r_THOLD__31__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__30__0_ ( .D(n2035), .CLK(clk), .QN(
        uart1_r_THOLD__30__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__30__1_ ( .D(n2034), .CLK(clk), .QN(
        uart1_r_THOLD__30__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__24__1_ ( .D(n2033), .CLK(clk), .QN(
        uart1_r_THOLD__24__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__22__1_ ( .D(n2032), .CLK(clk), .QN(
        uart1_r_THOLD__22__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__21__1_ ( .D(n2031), .CLK(clk), .QN(
        uart1_r_THOLD__21__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__19__1_ ( .D(n2030), .CLK(clk), .QN(
        uart1_r_THOLD__19__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__16__1_ ( .D(n2029), .CLK(clk), .QN(
        uart1_r_THOLD__16__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__14__1_ ( .D(n2028), .CLK(clk), .QN(
        uart1_r_THOLD__14__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__13__1_ ( .D(n2027), .CLK(clk), .QN(
        uart1_r_THOLD__13__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__12__1_ ( .D(n2026), .CLK(clk), .QN(
        uart1_r_THOLD__12__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__11__1_ ( .D(n2025), .CLK(clk), .QN(
        uart1_r_THOLD__11__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__10__1_ ( .D(n2024), .CLK(clk), .QN(
        uart1_r_THOLD__10__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__9__1_ ( .D(n2023), .CLK(clk), .QN(
        uart1_r_THOLD__9__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__8__1_ ( .D(n2022), .CLK(clk), .QN(
        uart1_r_THOLD__8__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__6__1_ ( .D(n2021), .CLK(clk), .QN(
        uart1_r_THOLD__6__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__5__1_ ( .D(n2020), .CLK(clk), .QN(
        uart1_r_THOLD__5__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__4__1_ ( .D(n2019), .CLK(clk), .QN(
        uart1_r_THOLD__4__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__3__1_ ( .D(n2018), .CLK(clk), .QN(
        uart1_r_THOLD__3__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__2__1_ ( .D(n2017), .CLK(clk), .QN(
        uart1_r_THOLD__2__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__1__1_ ( .D(n2016), .CLK(clk), .QN(
        uart1_r_THOLD__1__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__0__1_ ( .D(n2015), .CLK(clk), .QN(
        uart1_r_THOLD__0__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__30__2_ ( .D(n2014), .CLK(clk), .QN(
        uart1_r_THOLD__30__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__24__2_ ( .D(n2013), .CLK(clk), .QN(
        uart1_r_THOLD__24__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__22__2_ ( .D(n2012), .CLK(clk), .QN(
        uart1_r_THOLD__22__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__21__2_ ( .D(n2011), .CLK(clk), .QN(
        uart1_r_THOLD__21__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__19__2_ ( .D(n2010), .CLK(clk), .QN(
        uart1_r_THOLD__19__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__16__2_ ( .D(n2009), .CLK(clk), .QN(
        uart1_r_THOLD__16__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__14__2_ ( .D(n2008), .CLK(clk), .QN(
        uart1_r_THOLD__14__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__13__2_ ( .D(n2007), .CLK(clk), .QN(
        uart1_r_THOLD__13__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__12__2_ ( .D(n2006), .CLK(clk), .QN(
        uart1_r_THOLD__12__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__11__2_ ( .D(n2005), .CLK(clk), .QN(
        uart1_r_THOLD__11__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__10__2_ ( .D(n2004), .CLK(clk), .QN(
        uart1_r_THOLD__10__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__9__2_ ( .D(n2003), .CLK(clk), .QN(
        uart1_r_THOLD__9__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__8__2_ ( .D(n2002), .CLK(clk), .QN(
        uart1_r_THOLD__8__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__6__2_ ( .D(n2001), .CLK(clk), .QN(
        uart1_r_THOLD__6__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__5__2_ ( .D(n2000), .CLK(clk), .QN(
        uart1_r_THOLD__5__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__4__2_ ( .D(n1999), .CLK(clk), .QN(
        uart1_r_THOLD__4__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__3__2_ ( .D(n1998), .CLK(clk), .QN(
        uart1_r_THOLD__3__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__2__2_ ( .D(n1997), .CLK(clk), .QN(
        uart1_r_THOLD__2__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__1__2_ ( .D(n1996), .CLK(clk), .QN(
        uart1_r_THOLD__1__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__0__2_ ( .D(n1995), .CLK(clk), .QN(
        uart1_r_THOLD__0__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__30__3_ ( .D(n1994), .CLK(clk), .QN(
        uart1_r_THOLD__30__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__24__3_ ( .D(n1993), .CLK(clk), .QN(
        uart1_r_THOLD__24__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__22__3_ ( .D(n1992), .CLK(clk), .QN(
        uart1_r_THOLD__22__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__21__3_ ( .D(n1991), .CLK(clk), .QN(
        uart1_r_THOLD__21__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__19__3_ ( .D(n1990), .CLK(clk), .QN(
        uart1_r_THOLD__19__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__16__3_ ( .D(n1989), .CLK(clk), .QN(
        uart1_r_THOLD__16__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__14__3_ ( .D(n1988), .CLK(clk), .QN(
        uart1_r_THOLD__14__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__13__3_ ( .D(n1987), .CLK(clk), .QN(
        uart1_r_THOLD__13__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__12__3_ ( .D(n1986), .CLK(clk), .QN(
        uart1_r_THOLD__12__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__11__3_ ( .D(n1985), .CLK(clk), .QN(
        uart1_r_THOLD__11__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__10__3_ ( .D(n1984), .CLK(clk), .QN(
        uart1_r_THOLD__10__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__9__3_ ( .D(n1983), .CLK(clk), .QN(
        uart1_r_THOLD__9__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__8__3_ ( .D(n1982), .CLK(clk), .QN(
        uart1_r_THOLD__8__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__6__3_ ( .D(n1981), .CLK(clk), .QN(
        uart1_r_THOLD__6__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__5__3_ ( .D(n1980), .CLK(clk), .QN(
        uart1_r_THOLD__5__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__4__3_ ( .D(n1979), .CLK(clk), .QN(
        uart1_r_THOLD__4__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__3__3_ ( .D(n1978), .CLK(clk), .QN(
        uart1_r_THOLD__3__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__2__3_ ( .D(n1977), .CLK(clk), .QN(
        uart1_r_THOLD__2__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__1__3_ ( .D(n1976), .CLK(clk), .QN(
        uart1_r_THOLD__1__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__0__3_ ( .D(n1975), .CLK(clk), .QN(
        uart1_r_THOLD__0__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__30__4_ ( .D(n1974), .CLK(clk), .QN(
        uart1_r_THOLD__30__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__24__4_ ( .D(n1973), .CLK(clk), .QN(
        uart1_r_THOLD__24__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__22__4_ ( .D(n1972), .CLK(clk), .QN(
        uart1_r_THOLD__22__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__21__4_ ( .D(n1971), .CLK(clk), .QN(
        uart1_r_THOLD__21__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__19__4_ ( .D(n1970), .CLK(clk), .QN(
        uart1_r_THOLD__19__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__16__4_ ( .D(n1969), .CLK(clk), .QN(
        uart1_r_THOLD__16__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__14__4_ ( .D(n1968), .CLK(clk), .QN(
        uart1_r_THOLD__14__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__13__4_ ( .D(n1967), .CLK(clk), .QN(
        uart1_r_THOLD__13__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__12__4_ ( .D(n1966), .CLK(clk), .QN(
        uart1_r_THOLD__12__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__11__4_ ( .D(n1965), .CLK(clk), .QN(
        uart1_r_THOLD__11__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__10__4_ ( .D(n1964), .CLK(clk), .QN(
        uart1_r_THOLD__10__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__9__4_ ( .D(n1963), .CLK(clk), .QN(
        uart1_r_THOLD__9__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__8__4_ ( .D(n1962), .CLK(clk), .QN(
        uart1_r_THOLD__8__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__6__4_ ( .D(n1961), .CLK(clk), .QN(
        uart1_r_THOLD__6__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__5__4_ ( .D(n1960), .CLK(clk), .QN(
        uart1_r_THOLD__5__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__4__4_ ( .D(n1959), .CLK(clk), .QN(
        uart1_r_THOLD__4__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__3__4_ ( .D(n1958), .CLK(clk), .QN(
        uart1_r_THOLD__3__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__2__4_ ( .D(n1957), .CLK(clk), .QN(
        uart1_r_THOLD__2__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__1__4_ ( .D(n1956), .CLK(clk), .QN(
        uart1_r_THOLD__1__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__0__4_ ( .D(n1955), .CLK(clk), .QN(
        uart1_r_THOLD__0__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__30__5_ ( .D(n1954), .CLK(clk), .QN(
        uart1_r_THOLD__30__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__24__5_ ( .D(n1953), .CLK(clk), .QN(
        uart1_r_THOLD__24__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__22__5_ ( .D(n1952), .CLK(clk), .QN(
        uart1_r_THOLD__22__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__21__5_ ( .D(n1951), .CLK(clk), .QN(
        uart1_r_THOLD__21__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__19__5_ ( .D(n1950), .CLK(clk), .QN(
        uart1_r_THOLD__19__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__16__5_ ( .D(n1949), .CLK(clk), .QN(
        uart1_r_THOLD__16__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__14__5_ ( .D(n1948), .CLK(clk), .QN(
        uart1_r_THOLD__14__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__13__5_ ( .D(n1947), .CLK(clk), .QN(
        uart1_r_THOLD__13__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__12__5_ ( .D(n1946), .CLK(clk), .QN(
        uart1_r_THOLD__12__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__11__5_ ( .D(n1945), .CLK(clk), .QN(
        uart1_r_THOLD__11__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__10__5_ ( .D(n1944), .CLK(clk), .QN(
        uart1_r_THOLD__10__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__9__5_ ( .D(n1943), .CLK(clk), .QN(
        uart1_r_THOLD__9__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__8__5_ ( .D(n1942), .CLK(clk), .QN(
        uart1_r_THOLD__8__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__6__5_ ( .D(n1941), .CLK(clk), .QN(
        uart1_r_THOLD__6__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__5__5_ ( .D(n1940), .CLK(clk), .QN(
        uart1_r_THOLD__5__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__4__5_ ( .D(n1939), .CLK(clk), .QN(
        uart1_r_THOLD__4__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__3__5_ ( .D(n1938), .CLK(clk), .QN(
        uart1_r_THOLD__3__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__2__5_ ( .D(n1937), .CLK(clk), .QN(
        uart1_r_THOLD__2__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__1__5_ ( .D(n1936), .CLK(clk), .QN(
        uart1_r_THOLD__1__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__0__5_ ( .D(n1935), .CLK(clk), .QN(
        uart1_r_THOLD__0__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__30__6_ ( .D(n1934), .CLK(clk), .QN(
        uart1_r_THOLD__30__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__24__6_ ( .D(n1933), .CLK(clk), .QN(
        uart1_r_THOLD__24__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__22__6_ ( .D(n1932), .CLK(clk), .QN(
        uart1_r_THOLD__22__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__21__6_ ( .D(n1931), .CLK(clk), .QN(
        uart1_r_THOLD__21__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__19__6_ ( .D(n1930), .CLK(clk), .QN(
        uart1_r_THOLD__19__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__16__6_ ( .D(n1929), .CLK(clk), .QN(
        uart1_r_THOLD__16__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__14__6_ ( .D(n1928), .CLK(clk), .QN(
        uart1_r_THOLD__14__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__13__6_ ( .D(n1927), .CLK(clk), .QN(
        uart1_r_THOLD__13__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__12__6_ ( .D(n1926), .CLK(clk), .QN(
        uart1_r_THOLD__12__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__11__6_ ( .D(n1925), .CLK(clk), .QN(
        uart1_r_THOLD__11__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__10__6_ ( .D(n1924), .CLK(clk), .QN(
        uart1_r_THOLD__10__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__9__6_ ( .D(n1923), .CLK(clk), .QN(
        uart1_r_THOLD__9__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__8__6_ ( .D(n1922), .CLK(clk), .QN(
        uart1_r_THOLD__8__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__6__6_ ( .D(n1921), .CLK(clk), .QN(
        uart1_r_THOLD__6__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__5__6_ ( .D(n1920), .CLK(clk), .QN(
        uart1_r_THOLD__5__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__4__6_ ( .D(n1919), .CLK(clk), .QN(
        uart1_r_THOLD__4__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__3__6_ ( .D(n1918), .CLK(clk), .QN(
        uart1_r_THOLD__3__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__2__6_ ( .D(n1917), .CLK(clk), .QN(
        uart1_r_THOLD__2__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__1__6_ ( .D(n1916), .CLK(clk), .QN(
        uart1_r_THOLD__1__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__0__6_ ( .D(n1915), .CLK(clk), .QN(
        uart1_r_THOLD__0__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__30__7_ ( .D(n1914), .CLK(clk), .QN(
        uart1_r_THOLD__30__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__24__7_ ( .D(n1913), .CLK(clk), .QN(
        uart1_r_THOLD__24__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__22__7_ ( .D(n1912), .CLK(clk), .QN(
        uart1_r_THOLD__22__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__21__7_ ( .D(n1911), .CLK(clk), .QN(
        uart1_r_THOLD__21__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__19__7_ ( .D(n1910), .CLK(clk), .QN(
        uart1_r_THOLD__19__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__16__7_ ( .D(n1909), .CLK(clk), .QN(
        uart1_r_THOLD__16__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__14__7_ ( .D(n1908), .CLK(clk), .QN(
        uart1_r_THOLD__14__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__13__7_ ( .D(n1907), .CLK(clk), .QN(
        uart1_r_THOLD__13__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__12__7_ ( .D(n1906), .CLK(clk), .QN(
        uart1_r_THOLD__12__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__11__7_ ( .D(n1905), .CLK(clk), .QN(
        uart1_r_THOLD__11__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__10__7_ ( .D(n1904), .CLK(clk), .QN(
        uart1_r_THOLD__10__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__9__7_ ( .D(n1903), .CLK(clk), .QN(
        uart1_r_THOLD__9__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__8__7_ ( .D(n1902), .CLK(clk), .QN(
        uart1_r_THOLD__8__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__6__7_ ( .D(n1901), .CLK(clk), .QN(
        uart1_r_THOLD__6__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__5__7_ ( .D(n1900), .CLK(clk), .QN(
        uart1_r_THOLD__5__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__4__7_ ( .D(n1899), .CLK(clk), .QN(
        uart1_r_THOLD__4__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__3__7_ ( .D(n1898), .CLK(clk), .QN(
        uart1_r_THOLD__3__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__2__7_ ( .D(n1897), .CLK(clk), .QN(
        uart1_r_THOLD__2__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__1__7_ ( .D(n1896), .CLK(clk), .QN(
        uart1_r_THOLD__1__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__0__7_ ( .D(n1895), .CLK(clk), .QN(
        uart1_r_THOLD__0__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__29__0_ ( .D(n1894), .CLK(clk), .QN(
        uart1_r_THOLD__29__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__29__1_ ( .D(n1893), .CLK(clk), .QN(
        uart1_r_THOLD__29__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__29__2_ ( .D(n1892), .CLK(clk), .QN(
        uart1_r_THOLD__29__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__29__3_ ( .D(n1891), .CLK(clk), .QN(
        uart1_r_THOLD__29__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__29__4_ ( .D(n1890), .CLK(clk), .QN(
        uart1_r_THOLD__29__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__29__5_ ( .D(n1889), .CLK(clk), .QN(
        uart1_r_THOLD__29__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__29__6_ ( .D(n1888), .CLK(clk), .QN(
        uart1_r_THOLD__29__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__29__7_ ( .D(n1887), .CLK(clk), .QN(
        uart1_r_THOLD__29__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__28__0_ ( .D(n1886), .CLK(clk), .QN(
        uart1_r_THOLD__28__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__28__1_ ( .D(n1885), .CLK(clk), .QN(
        uart1_r_THOLD__28__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__28__2_ ( .D(n1884), .CLK(clk), .QN(
        uart1_r_THOLD__28__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__28__3_ ( .D(n1883), .CLK(clk), .QN(
        uart1_r_THOLD__28__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__28__4_ ( .D(n1882), .CLK(clk), .QN(
        uart1_r_THOLD__28__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__28__5_ ( .D(n1881), .CLK(clk), .QN(
        uart1_r_THOLD__28__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__28__6_ ( .D(n1880), .CLK(clk), .QN(
        uart1_r_THOLD__28__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__28__7_ ( .D(n1879), .CLK(clk), .QN(
        uart1_r_THOLD__28__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__27__0_ ( .D(n1878), .CLK(clk), .QN(
        uart1_r_THOLD__27__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__27__1_ ( .D(n1877), .CLK(clk), .QN(
        uart1_r_THOLD__27__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__27__2_ ( .D(n1876), .CLK(clk), .QN(
        uart1_r_THOLD__27__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__27__3_ ( .D(n1875), .CLK(clk), .QN(
        uart1_r_THOLD__27__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__27__4_ ( .D(n1874), .CLK(clk), .QN(
        uart1_r_THOLD__27__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__27__5_ ( .D(n1873), .CLK(clk), .QN(
        uart1_r_THOLD__27__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__27__6_ ( .D(n1872), .CLK(clk), .QN(
        uart1_r_THOLD__27__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__27__7_ ( .D(n1871), .CLK(clk), .QN(
        uart1_r_THOLD__27__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__26__0_ ( .D(n1870), .CLK(clk), .QN(
        uart1_r_THOLD__26__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__26__1_ ( .D(n1869), .CLK(clk), .QN(
        uart1_r_THOLD__26__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__26__2_ ( .D(n1868), .CLK(clk), .QN(
        uart1_r_THOLD__26__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__26__3_ ( .D(n1867), .CLK(clk), .QN(
        uart1_r_THOLD__26__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__26__4_ ( .D(n1866), .CLK(clk), .QN(
        uart1_r_THOLD__26__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__26__5_ ( .D(n1865), .CLK(clk), .QN(
        uart1_r_THOLD__26__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__26__6_ ( .D(n1864), .CLK(clk), .QN(
        uart1_r_THOLD__26__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__26__7_ ( .D(n1863), .CLK(clk), .QN(
        uart1_r_THOLD__26__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__25__0_ ( .D(n1862), .CLK(clk), .QN(
        uart1_r_THOLD__25__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__25__1_ ( .D(n1861), .CLK(clk), .QN(
        uart1_r_THOLD__25__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__25__2_ ( .D(n1860), .CLK(clk), .QN(
        uart1_r_THOLD__25__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__25__3_ ( .D(n1859), .CLK(clk), .QN(
        uart1_r_THOLD__25__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__25__4_ ( .D(n1858), .CLK(clk), .QN(
        uart1_r_THOLD__25__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__25__5_ ( .D(n1857), .CLK(clk), .QN(
        uart1_r_THOLD__25__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__25__6_ ( .D(n1856), .CLK(clk), .QN(
        uart1_r_THOLD__25__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__25__7_ ( .D(n1855), .CLK(clk), .QN(
        uart1_r_THOLD__25__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__23__0_ ( .D(n1854), .CLK(clk), .QN(
        uart1_r_THOLD__23__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__23__1_ ( .D(n1853), .CLK(clk), .QN(
        uart1_r_THOLD__23__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__23__2_ ( .D(n1852), .CLK(clk), .QN(
        uart1_r_THOLD__23__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__23__3_ ( .D(n1851), .CLK(clk), .QN(
        uart1_r_THOLD__23__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__23__4_ ( .D(n1850), .CLK(clk), .QN(
        uart1_r_THOLD__23__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__23__5_ ( .D(n1849), .CLK(clk), .QN(
        uart1_r_THOLD__23__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__23__6_ ( .D(n1848), .CLK(clk), .QN(
        uart1_r_THOLD__23__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__23__7_ ( .D(n1847), .CLK(clk), .QN(
        uart1_r_THOLD__23__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__20__0_ ( .D(n1846), .CLK(clk), .QN(
        uart1_r_THOLD__20__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__20__1_ ( .D(n1845), .CLK(clk), .QN(
        uart1_r_THOLD__20__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__20__2_ ( .D(n1844), .CLK(clk), .QN(
        uart1_r_THOLD__20__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__20__3_ ( .D(n1843), .CLK(clk), .QN(
        uart1_r_THOLD__20__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__20__4_ ( .D(n1842), .CLK(clk), .QN(
        uart1_r_THOLD__20__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__20__5_ ( .D(n1841), .CLK(clk), .QN(
        uart1_r_THOLD__20__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__20__6_ ( .D(n1840), .CLK(clk), .QN(
        uart1_r_THOLD__20__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__20__7_ ( .D(n1839), .CLK(clk), .QN(
        uart1_r_THOLD__20__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__18__0_ ( .D(n1838), .CLK(clk), .QN(
        uart1_r_THOLD__18__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__18__1_ ( .D(n1837), .CLK(clk), .QN(
        uart1_r_THOLD__18__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__18__2_ ( .D(n1836), .CLK(clk), .QN(
        uart1_r_THOLD__18__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__18__3_ ( .D(n1835), .CLK(clk), .QN(
        uart1_r_THOLD__18__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__18__4_ ( .D(n1834), .CLK(clk), .QN(
        uart1_r_THOLD__18__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__18__5_ ( .D(n1833), .CLK(clk), .QN(
        uart1_r_THOLD__18__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__18__6_ ( .D(n1832), .CLK(clk), .QN(
        uart1_r_THOLD__18__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__18__7_ ( .D(n1831), .CLK(clk), .QN(
        uart1_r_THOLD__18__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__17__0_ ( .D(n1830), .CLK(clk), .QN(
        uart1_r_THOLD__17__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__17__1_ ( .D(n1829), .CLK(clk), .QN(
        uart1_r_THOLD__17__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__17__2_ ( .D(n1828), .CLK(clk), .QN(
        uart1_r_THOLD__17__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__17__3_ ( .D(n1827), .CLK(clk), .QN(
        uart1_r_THOLD__17__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__17__4_ ( .D(n1826), .CLK(clk), .QN(
        uart1_r_THOLD__17__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__17__5_ ( .D(n1825), .CLK(clk), .QN(
        uart1_r_THOLD__17__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__17__6_ ( .D(n1824), .CLK(clk), .QN(
        uart1_r_THOLD__17__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__17__7_ ( .D(n1823), .CLK(clk), .QN(
        uart1_r_THOLD__17__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__15__0_ ( .D(n1822), .CLK(clk), .QN(
        uart1_r_THOLD__15__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__15__1_ ( .D(n1821), .CLK(clk), .QN(
        uart1_r_THOLD__15__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__15__2_ ( .D(n1820), .CLK(clk), .QN(
        uart1_r_THOLD__15__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__15__3_ ( .D(n1819), .CLK(clk), .QN(
        uart1_r_THOLD__15__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__15__4_ ( .D(n1818), .CLK(clk), .QN(
        uart1_r_THOLD__15__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__15__5_ ( .D(n1817), .CLK(clk), .QN(
        uart1_r_THOLD__15__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__15__6_ ( .D(n1816), .CLK(clk), .QN(
        uart1_r_THOLD__15__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__15__7_ ( .D(n1815), .CLK(clk), .QN(
        uart1_r_THOLD__15__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__7__0_ ( .D(n1814), .CLK(clk), .QN(
        uart1_r_THOLD__7__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__7__1_ ( .D(n1813), .CLK(clk), .QN(
        uart1_r_THOLD__7__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__7__2_ ( .D(n1812), .CLK(clk), .QN(
        uart1_r_THOLD__7__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__7__3_ ( .D(n1811), .CLK(clk), .QN(
        uart1_r_THOLD__7__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__7__4_ ( .D(n1810), .CLK(clk), .QN(
        uart1_r_THOLD__7__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__7__5_ ( .D(n1809), .CLK(clk), .QN(
        uart1_r_THOLD__7__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__7__6_ ( .D(n1808), .CLK(clk), .QN(
        uart1_r_THOLD__7__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_THOLD__7__7_ ( .D(n1807), .CLK(clk), .QN(
        uart1_r_THOLD__7__7_) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__10_ ( .D(n1806), .CLK(clk), .QN(
        ahb0_r_HADDR__10_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__9_ ( 
        .D(n1805), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[13]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__9_ ( .D(n1804), .CLK(clk), .QN(
        apbi[9]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMBANKSZ__0_ ( .D(n1803), .CLK(clk), 
        .QN(sr1_r_MCFG2__RAMBANKSZ__0_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__ROMWIDTH__1_ ( .D(n1802), .CLK(clk), 
        .QN(sr1_r_MCFG1__ROMWIDTH__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TFIFOIRQEN_ ( .D(n1801), .CLK(clk), .QN(
        uart1_r_TFIFOIRQEN_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BRATE__9_ ( .D(n1800), .CLK(clk), .QN(
        uart1_r_BRATE__9_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_SCALER__9_ ( .D(n1799), .CLK(clk), .QN(
        uart1_uarto_SCALER__9_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__9_ ( .D(n1798), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__9_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__9_ ( .D(n1797), .CLK(clk), .QN(
        irqctrl0_r_IPEND__9_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__9_ ( .D(n1796), .CLK(clk), .QN(
        irqctrl0_r_ILEVEL__9_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__9_ ( .D(n1795), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__9_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_DISHLT_ ( .D(n1794), .CLK(clk), .QN(
        timer0_r_DISHLT_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__9_ ( .D(n1793), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__9_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__9_ ( .D(
        timer0_v_TIMERS__1__VALUE__9_), .CLK(clk), .QN(n1792) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HADDR__9_ ( .D(n1791), .CLK(clk), .QN(
        ahb0_r_HADDR__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__ICC__2_ ( .D(n1789), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__ICC__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__ICC__2_ ( .D(n1788), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__ICC__2_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__Y__29_ ( .D(n1786), .CLK(
        clk), .QN(u0_0_leon3x0_p0_divi[60]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__Y__29_ ( .D(n1784), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_X__Y__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_W__S__Y__29_ ( .D(n1783), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__Y__29_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__28_ ( 
        .D(n1782), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[32]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__28_ ( .D(n1781), .CLK(clk), .QN(
        apbi[28]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_MCFG1__IOWIDTH__1_ ( .D(n1780), .CLK(clk), 
        .QN(sr1_r_MCFG1__IOWIDTH__1_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_BUSW__1_ ( .D(n1779), .CLK(clk), .QN(
        sr1_r_BUSW__1_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__12_ ( .D(n1778), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__12_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__12_ ( .D(n1777), .CLK(clk), .QN(
        irqctrl0_r_IPEND__12_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__28_ ( .D(n1776), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__28_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__28_ ( .D(
        timer0_v_TIMERS__1__VALUE__28_), .CLK(clk), .QN(n1775) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__16_ ( 
        .D(n1774), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[20]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__16_ ( .D(n1773), .CLK(clk), .QN(
        apbi[16]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__16_ ( .D(n1772), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__16_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__16_ ( .D(
        timer0_v_TIMERS__1__VALUE__16_), .CLK(clk), .QN(n1771) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__16_ ( .D(n1770), .CLK(clk), .QN(
        ahbso_1__HRDATA__16_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__13_ ( 
        .D(n1767), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[17]) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__13_ ( .D(n1766), .CLK(clk), .QN(
        apbi[13]) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_DELAYIRQEN_ ( .D(n17812), .CLK(clk), .QN(
        n1765) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_IRQCNT__0_ ( .D(n1764), .CLK(clk), .QN(
        uart1_r_IRQCNT__0_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_IRQCNT__1_ ( .D(n1763), .CLK(clk), .QN(
        uart1_r_IRQCNT__1_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_IRQCNT__2_ ( .D(n1762), .CLK(clk), .QN(
        uart1_r_IRQCNT__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_IRQCNT__3_ ( .D(n1761), .CLK(clk), .QN(
        uart1_r_IRQCNT__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_IRQCNT__4_ ( .D(n1760), .CLK(clk), .QN(
        uart1_r_IRQCNT__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_IRQCNT__5_ ( .D(n1759), .CLK(clk), .QN(
        uart1_r_IRQCNT__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_IRQPEND_ ( .D(n1758), .CLK(clk), .QN(
        uart1_r_IRQPEND_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_IRQ_ ( .D(n1757), .CLK(clk), .QN(
        apbo_1__PIRQ__2_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__2_ ( .D(n1756), .CLK(clk), .QN(
        irqctrl0_r_IPEND__2_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__13_ ( .D(n1755), .CLK(clk), 
        .QN(irqctrl0_r_ILEVEL__13_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__13_ ( .D(n1754), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__13_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__13_ ( .D(n1753), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__13_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__13_ ( .D(
        timer0_v_TIMERS__1__VALUE__13_), .CLK(clk), .QN(n1752) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__29_ ( .D(n1751), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__29_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_RELOAD__2_ ( .D(n1750), .CLK(clk), .QN(
        timer0_r_RELOAD__2_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_SCALER__2_ ( .D(n1749), .CLK(clk), .QN(
        timer0_r_SCALER__2_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_PARERR_ ( .D(n1748), .CLK(clk), .QN(
        uart1_r_PARERR_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_FRAME_ ( .D(n1747), .CLK(clk), .QN(
        uart1_r_FRAME_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_BREAK_ ( .D(n1746), .CLK(clk), .QN(
        uart1_r_BREAK_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__8_ ( .D(n1745), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__8_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__8_ ( .D(n1744), .CLK(clk), .QN(
        irqctrl0_r_ILEVEL__8_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__8_ ( .D(n1743), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__8_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__8_ ( .D(n1742), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__8_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__8_ ( .D(
        timer0_v_TIMERS__1__VALUE__8_), .CLK(clk), .QN(n1741) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_RELOAD__3_ ( .D(n1740), .CLK(clk), .QN(
        timer0_r_RELOAD__3_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_SCALER__3_ ( .D(n1739), .CLK(clk), .QN(
        timer0_r_SCALER__3_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__0__4_ ( .D(n1738), .CLK(clk), .QN(
        uart1_r_RHOLD__0__4_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__0__5_ ( .D(n1737), .CLK(clk), .QN(
        uart1_r_RHOLD__0__5_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__0__6_ ( .D(n1736), .CLK(clk), .QN(
        uart1_r_RHOLD__0__6_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_RHOLD__0__7_ ( .D(n1735), .CLK(clk), .QN(
        uart1_r_RHOLD__0__7_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_OVF_ ( .D(n1734), .CLK(clk), .QN(
        uart1_r_OVF_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IFORCE__0__6_ ( .D(n1733), .CLK(clk), 
        .QN(irqctrl0_r_IFORCE__0__6_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IPEND__6_ ( .D(n1732), .CLK(clk), .QN(
        irqctrl0_r_IPEND__6_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_ILEVEL__6_ ( .D(n1731), .CLK(clk), .QN(
        irqctrl0_r_ILEVEL__6_) );
  DFFHQNx1_ASAP7_75t_SL irqctrl0_r_reg_IMASK__0__6_ ( .D(n1730), .CLK(clk), 
        .QN(irqctrl0_r_IMASK__0__6_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__6_ ( .D(n1729), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__6_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__6_ ( .D(
        timer0_v_TIMERS__1__VALUE__6_), .CLK(clk), .QN(n1728) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_RELOAD__6_ ( .D(n1727), .CLK(clk), .QN(
        timer0_r_RELOAD__6_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_SCALER__6_ ( .D(n1726), .CLK(clk), .QN(
        timer0_r_SCALER__6_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WS__2_ ( .D(n1725), .CLK(clk), .QN(
        sr1_r_WS__2_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__0_ ( .D(sr1_v_ADDRESS__0_), .CLK(
        clk), .QN(n1724) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__1_ ( .D(sr1_v_ADDRESS__1_), .CLK(
        clk), .QN(n1723) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRN__0_ ( .D(n1722), .CLK(clk), .QN(rwen[0])
         );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRN__1_ ( .D(n1721), .CLK(clk), .QN(rwen[1])
         );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRN__2_ ( .D(n1720), .CLK(clk), .QN(rwen[2])
         );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRN__3_ ( .D(n1719), .CLK(clk), .QN(rwen[3])
         );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__0_ ( .D(n1718), .CLK(clk), .QN(
        dataout[0]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__1_ ( .D(n1717), .CLK(clk), .QN(
        dataout[1]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__2_ ( .D(n1716), .CLK(clk), .QN(
        dataout[2]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__3_ ( .D(n1715), .CLK(clk), .QN(
        dataout[3]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__4_ ( .D(n1714), .CLK(clk), .QN(
        dataout[4]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__5_ ( .D(n1713), .CLK(clk), .QN(
        dataout[5]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__6_ ( .D(n1712), .CLK(clk), .QN(
        dataout[6]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__7_ ( .D(n1711), .CLK(clk), .QN(
        dataout[7]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__8_ ( .D(n1710), .CLK(clk), .QN(
        dataout[8]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__9_ ( .D(n1709), .CLK(clk), .QN(
        dataout[9]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__10_ ( .D(n1708), .CLK(clk), .QN(
        dataout[10]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__11_ ( .D(n1707), .CLK(clk), .QN(
        dataout[11]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__12_ ( .D(n1706), .CLK(clk), .QN(
        dataout[12]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__13_ ( .D(n1705), .CLK(clk), .QN(
        dataout[13]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__14_ ( .D(n1704), .CLK(clk), .QN(
        dataout[14]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__15_ ( .D(n1703), .CLK(clk), .QN(
        dataout[15]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__16_ ( .D(n1702), .CLK(clk), .QN(
        dataout[16]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__17_ ( .D(n1701), .CLK(clk), .QN(
        dataout[17]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__18_ ( .D(n1700), .CLK(clk), .QN(
        dataout[18]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__19_ ( .D(n1699), .CLK(clk), .QN(
        dataout[19]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__20_ ( .D(n1698), .CLK(clk), .QN(
        dataout[20]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__21_ ( .D(n1697), .CLK(clk), .QN(
        dataout[21]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__22_ ( .D(n1696), .CLK(clk), .QN(
        dataout[22]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__23_ ( .D(n1695), .CLK(clk), .QN(
        dataout[23]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__24_ ( .D(n1694), .CLK(clk), .QN(
        dataout[24]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__25_ ( .D(n1693), .CLK(clk), .QN(
        dataout[25]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__26_ ( .D(n1692), .CLK(clk), .QN(
        dataout[26]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__27_ ( .D(n1691), .CLK(clk), .QN(
        dataout[27]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__28_ ( .D(n1690), .CLK(clk), .QN(
        dataout[28]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__29_ ( .D(n1689), .CLK(clk), .QN(
        dataout[29]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__30_ ( .D(n1688), .CLK(clk), .QN(
        dataout[30]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_WRITEDATA__31_ ( .D(n1687), .CLK(clk), .QN(
        dataout[31]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__2_ ( .D(n1686), .CLK(clk), .QN(
        address[2]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__3_ ( .D(n1685), .CLK(clk), .QN(
        address[3]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__4_ ( .D(n1684), .CLK(clk), .QN(
        address[4]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__6_ ( .D(n1683), .CLK(clk), .QN(
        address[6]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__8_ ( .D(n1682), .CLK(clk), .QN(
        address[8]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__9_ ( .D(n1681), .CLK(clk), .QN(
        address[9]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__10_ ( .D(n1680), .CLK(clk), .QN(
        address[10]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__11_ ( .D(n1679), .CLK(clk), .QN(
        address[11]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__12_ ( .D(n1678), .CLK(clk), .QN(
        address[12]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__13_ ( .D(n1677), .CLK(clk), .QN(
        address[13]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__14_ ( .D(n1676), .CLK(clk), .QN(
        address[14]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__15_ ( .D(n1675), .CLK(clk), .QN(
        address[15]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__16_ ( .D(n1674), .CLK(clk), .QN(
        address[16]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__17_ ( .D(n1673), .CLK(clk), .QN(
        address[17]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__18_ ( .D(n1672), .CLK(clk), .QN(
        address[18]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__19_ ( .D(n1671), .CLK(clk), .QN(
        address[19]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__20_ ( .D(n1670), .CLK(clk), .QN(
        address[20]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__21_ ( .D(n1669), .CLK(clk), .QN(
        address[21]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__22_ ( .D(n1668), .CLK(clk), .QN(
        address[22]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__23_ ( .D(n1667), .CLK(clk), .QN(
        address[23]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__24_ ( .D(n1666), .CLK(clk), .QN(
        address[24]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__25_ ( .D(n1665), .CLK(clk), .QN(
        address[25]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__26_ ( .D(n1664), .CLK(clk), .QN(
        address[26]) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__27_ ( .D(n1663), .CLK(clk), .QN(
        address[27]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_ROMSN__0_ ( .D(n1661), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(romsn[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_ROMSN__1_ ( .D(n1659), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(romsn[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_RAMSN__0_ ( .D(n1657), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(ramsn[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_RAMOEN__0_ ( .D(n1655), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(ramoen[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_RAMSN__1_ ( .D(n1653), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(ramsn[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_RAMOEN__1_ ( .D(n1651), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(ramoen[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_RAMSN__2_ ( .D(n1649), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(ramsn[2]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_RAMOEN__2_ ( .D(n1647), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(ramoen[2]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_RAMSN__3_ ( .D(n1645), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(ramsn[3]) );
  ASYNC_DFFHx1_ASAP7_75t_SL sr1_r_reg_RAMOEN__3_ ( .D(n1643), .CLK(clk), 
        .RESET(n18295), .SET(n24695), .QN(ramoen[3]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__30_ ( .D(n1640), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__30_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_RELOAD__5_ ( .D(n1639), .CLK(clk), .QN(
        timer0_r_RELOAD__5_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_SCALER__5_ ( .D(n1638), .CLK(clk), .QN(
        timer0_r_SCALER__5_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__5_ ( .D(n1636), .CLK(clk), .QN(
        address[5]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__12_ ( .D(n1635), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__12_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__12_ ( .D(
        timer0_v_TIMERS__1__VALUE__12_), .CLK(clk), .QN(n1634) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PRDATA__12_ ( .D(n1633), .CLK(clk), .QN(
        ahbso_1__HRDATA__12_) );
  DFFHQNx1_ASAP7_75t_SL sr1_r_reg_ADDRESS__7_ ( .D(n1632), .CLK(clk), .QN(
        address[7]) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__4_ ( .D(n1631), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__4_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__4_ ( .D(
        timer0_v_TIMERS__1__VALUE__4_), .CLK(clk), .QN(n1630) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_RELOAD__4_ ( .D(n1629), .CLK(clk), .QN(
        timer0_r_RELOAD__4_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_SCALER__4_ ( .D(n1628), .CLK(clk), .QN(
        timer0_r_SCALER__4_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__RELOAD__7_ ( .D(n1627), .CLK(
        clk), .QN(timer0_vtimers_1__RELOAD__7_) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_TIMERS__1__VALUE__7_ ( .D(
        timer0_v_TIMERS__1__VALUE__7_), .CLK(clk), .QN(n1626) );
  DFFHQNx1_ASAP7_75t_SL timer0_r_reg_RELOAD__7_ ( .D(n1625), .CLK(clk), .QN(
        timer0_r_RELOAD__7_) );
  XNOR2xp5_ASAP7_75t_SL add_x_746_U180 ( .A(u0_0_leon3x0_p0_iu_fe_pc_2_), .B(
        add_x_746_n155), .Y(u0_0_leon3x0_p0_iu_fe_npc_3_) );
  XNOR2xp5_ASAP7_75t_SL add_x_746_U176 ( .A(add_x_746_n151), .B(add_x_746_n152), .Y(u0_0_leon3x0_p0_iu_fe_npc_4_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U170 ( .A(add_x_746_n148), .B(add_x_746_n149), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_5_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U165 ( .A(add_x_746_n143), .B(add_x_746_n144), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_6_) );
  XNOR2xp5_ASAP7_75t_SL add_x_746_U158 ( .A(add_x_746_n139), .B(add_x_746_n140), .Y(u0_0_leon3x0_p0_iu_fe_npc_7_) );
  XNOR2xp5_ASAP7_75t_SL add_x_746_U153 ( .A(add_x_746_n133), .B(add_x_746_n134), .Y(u0_0_leon3x0_p0_iu_fe_npc_8_) );
  XNOR2xp5_ASAP7_75t_SL add_x_746_U146 ( .A(add_x_746_n129), .B(add_x_746_n130), .Y(u0_0_leon3x0_p0_iu_fe_npc_9_) );
  XNOR2xp5_ASAP7_75t_SL add_x_746_U142 ( .A(add_x_746_n123), .B(add_x_746_n124), .Y(u0_0_leon3x0_p0_iu_fe_npc_10_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U134 ( .A(add_x_746_n120), .B(add_x_746_n121), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_11_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U128 ( .A(add_x_746_n113), .B(add_x_746_n114), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_12_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U120 ( .A(add_x_746_n108), .B(add_x_746_n109), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_13_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U114 ( .A(add_x_746_n99), .B(add_x_746_n102), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_14_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U106 ( .A(add_x_746_n96), .B(add_x_746_n97), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_15_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U100 ( .A(add_x_746_n89), .B(add_x_746_n90), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_16_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U93 ( .A(add_x_746_n84), .B(add_x_746_n85), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_17_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U81 ( .A(add_x_746_n75), .B(add_x_746_n76), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_19_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U75 ( .A(add_x_746_n68), .B(add_x_746_n69), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_20_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U67 ( .A(add_x_746_n63), .B(add_x_746_n64), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_21_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U61 ( .A(add_x_746_n56), .B(add_x_746_n57), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_22_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U53 ( .A(add_x_746_n51), .B(add_x_746_n52), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_23_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U47 ( .A(add_x_746_n44), .B(add_x_746_n45), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_24_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U39 ( .A(add_x_746_n39), .B(add_x_746_n40), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_25_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U33 ( .A(add_x_746_n32), .B(add_x_746_n33), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_26_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U25 ( .A(add_x_746_n27), .B(add_x_746_n28), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_27_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U19 ( .A(add_x_746_n20), .B(add_x_746_n21), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_28_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U11 ( .A(add_x_746_n15), .B(add_x_746_n16), 
        .Y(u0_0_leon3x0_p0_iu_fe_npc_29_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U5 ( .A(add_x_746_n8), .B(add_x_746_n9), .Y(
        u0_0_leon3x0_p0_iu_fe_npc_30_) );
  XOR2xp5_ASAP7_75t_SL add_x_746_U3 ( .A(n24493), .B(add_x_746_n4), .Y(
        u0_0_leon3x0_p0_iu_fe_npc_31_) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PWDATA__7_ ( .D(n4776), .CLK(clk), .QN(
        apbi[7]) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PWDATA__4_ ( .D(n4765), .CLK(clk), .QN(
        apbi[4]) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PWDATA__5_ ( .D(n4743), .CLK(clk), .QN(
        apbi[5]) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PWDATA__6_ ( .D(n4711), .CLK(clk), .QN(
        apbi[6]) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PWDATA__3_ ( .D(n4691), .CLK(clk), .QN(
        apbi[3]) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PWDATA__2_ ( .D(n4671), .CLK(clk), .QN(
        apbi[2]) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PWDATA__1_ ( .D(n4533), .CLK(clk), .QN(
        apbi[1]) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__20_ ( .D(n24449), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__23_ ( .D(n24448), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PWDATA__0_ ( .D(n4365), .CLK(clk), .QN(
        apbi[0]) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__CNT__0_ ( .D(n4336), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__0_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__20_ ( .D(n4179), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__22_ ( .D(n4177), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__CTRL__INST__22_ ( .D(n4105), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__24_ ( .D(n24456), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__CTRL__WICC_ ( .D(n3711), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__19_ ( .D(n3606), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__ALUOP__0_ ( .D(n3560), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__ALUOP__1_ ( .D(n3558), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__DCI__READ_ ( .D(n3302), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_dci[2]) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__JMPL_ ( .D(n3162), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__JMPL_) );
  DFFHQNx2_ASAP7_75t_SL sr1_r_reg_MCFG2__RAMBANKSZ__2_ ( .D(n17805), .CLK(clk), 
        .QN(n2924) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__CWP__1_ ( .D(n2802), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_A__CWP__1_) );
  DFFHQx4_ASAP7_75t_SL timer0_r_reg_TSEL_ ( .D(n24554), .CLK(clk), .Q(n5061)
         );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_PWDATA__11_ ( .D(n4521), .CLK(clk), .QN(
        apbi[11]) );
  SDFHx1_ASAP7_75t_SL apb0_r_reg_PRDATA__1_ ( .D(n16969), .SI(n4536), .SE(
        apb0_r_CFGSEL_), .CLK(clk), .QN(ahbso_1__HRDATA__1_) );
  DFFHQNx1_ASAP7_75t_SRAM uart1_r_reg_TSHIFT__1_ ( .D(n17443), .CLK(clk), .QN(
        n4701) );
  SDFHx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__9_ ( .D(n17271), .SI(n19002), .SE(
        n17270), .CLK(clk), .QN(ahb0_r_HRDATAS__9_) );
  SDFHx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__10_ ( .D(n17271), .SI(n19002), .SE(
        n17270), .CLK(clk), .QN(ahb0_r_HRDATAS__10_) );
  SDFHx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__8_ ( .D(n17271), .SI(n19002), .SE(
        n17270), .CLK(clk), .QN(ahb0_r_HRDATAS__8_) );
  SDFHx1_ASAP7_75t_SRAM u0_0_leon3x0_p0_iu_r_reg_W__S__PS_ ( .D(n3369), .SI(
        n18295), .SE(n22380), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_W__S__PS_)
         );
  SDFHx1_ASAP7_75t_SL apb0_r_reg_PRDATA__14_ ( .D(n17066), .SI(n4431), .SE(
        apb0_r_CFGSEL_), .CLK(clk), .QN(ahbso_1__HRDATA__14_) );
  SDFHx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__24_ ( .D(n17271), .SI(n19002), .SE(
        n17278), .CLK(clk), .QN(ahb0_r_HRDATAS__24_) );
  SDFHx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__29_ ( .D(ahb0_r_HADDR__3_), .SI(
        n19002), .SE(n17288), .CLK(clk), .QN(ahb0_r_HRDATAS__29_) );
  SDFHx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__26_ ( .D(n17284), .SI(n19002), .SE(
        n17285), .CLK(clk), .QN(ahb0_r_HRDATAS__26_) );
  DFFHQNx1_ASAP7_75t_SL uart1_r_reg_TRADDR__1_ ( .D(n2239), .CLK(clk), .QN(
        uart1_r_TRADDR__1_) );
  SDFHx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_FLUSH2_ ( .D(n24684), 
        .SI(n18295), .SE(n33067), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FLUSH2_) );
  SDFHx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__7_ ( .D(n17271), .SI(n19002), .SE(
        n17270), .CLK(clk), .QN(ahb0_r_HRDATAS__7_) );
  SDFHx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__31_ ( .D(n17271), .SI(n19002), .SE(
        n17270), .CLK(clk), .QN(ahb0_r_HRDATAS__31_) );
  SDFHx1_ASAP7_75t_SRAM u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_ICENABLE_ ( .D(
        u0_0_leon3x0_p0_ico_DIAGRDY_), .SI(n19002), .SE(n13499), .CLK(clk), 
        .QN(u0_0_leon3x0_p0_dco_ICDIAG__ENABLE_) );
  SDFHx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_a0_r_reg_NBO__1_ ( .D(n22380), 
        .SI(n19002), .SE(n10988), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_a0_r_NBO__1_) );
  SDFHx1_ASAP7_75t_SL uart1_r_reg_TCNT__4_ ( .D(n5591), .SI(n19002), .SE(
        n24695), .CLK(clk), .QN(uart1_r_TCNT__4_) );
  SDFHx1_ASAP7_75t_SL uart1_r_reg_TCNT__3_ ( .D(n5592), .SI(n19002), .SE(
        n24695), .CLK(clk), .QN(uart1_r_TCNT__3_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__3_ ( .D(n3959), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[3]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__RESULT__0_ ( .D(n3910), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mmudci[0]) );
  SDFHx1_ASAP7_75t_SRAM u0_0_leon3x0_p0_c0mmu_a0_r_reg_BA_ ( .D(n4079), .SI(
        n18295), .SE(n22380), .CLK(clk), .QN(n4081) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U130 ( .A(add_x_746_n113), .B(add_x_746_n116), .Y(add_x_746_n110) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U108 ( .A(add_x_746_n92), .B(add_x_746_n104), 
        .Y(add_x_746_n91) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U55 ( .A(add_x_746_n47), .B(add_x_746_n59), 
        .Y(add_x_746_n46) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U43 ( .A(add_x_746_n37), .B(add_x_746_n47), 
        .Y(add_x_746_n36) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U27 ( .A(add_x_746_n23), .B(add_x_746_n2), 
        .Y(add_x_746_n22) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U63 ( .A(add_x_746_n56), .B(add_x_746_n59), 
        .Y(add_x_746_n53) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U159 ( .A(add_x_746_n135), .B(add_x_746_n144), .Y(add_x_746_n134) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U154 ( .A(add_x_746_n144), .B(add_x_746_n131), .Y(add_x_746_n130) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U166 ( .A(add_x_746_n143), .B(add_x_746_n144), .Y(add_x_746_n140) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U35 ( .A(add_x_746_n32), .B(add_x_746_n2), 
        .Y(add_x_746_n29) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U116 ( .A(add_x_746_n99), .B(add_x_746_n104), 
        .Y(add_x_746_n98) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U77 ( .A(add_x_746_n68), .B(add_x_746_n71), 
        .Y(add_x_746_n65) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U172 ( .A(add_x_746_n153), .B(add_x_746_n146), .Y(add_x_746_n145) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U149 ( .A(add_x_746_n127), .B(add_x_746_n135), .Y(add_x_746_n126) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U124 ( .A(add_x_746_n116), .B(add_x_746_n106), .Y(add_x_746_n103) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U71 ( .A(add_x_746_n61), .B(add_x_746_n71), 
        .Y(add_x_746_n58) );
  NOR2xp33_ASAP7_75t_SL add_x_746_U15 ( .A(add_x_746_n13), .B(add_x_746_n23), 
        .Y(add_x_746_n12) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__INVOP2_ ( .D(n3316), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__INVOP2_) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U44 ( .A(
        DP_OP_5187J1_124_3275_n69), .B(DP_OP_5187J1_124_3275_n6), .Y(
        DP_OP_5187J1_124_3275_n67) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U58 ( .A(
        DP_OP_5187J1_124_3275_n80), .B(DP_OP_5187J1_124_3275_n6), .Y(
        DP_OP_5187J1_124_3275_n78) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U84 ( .A(
        DP_OP_5187J1_124_3275_n100), .B(DP_OP_5187J1_124_3275_n109), .Y(
        DP_OP_5187J1_124_3275_n98) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U30 ( .A(
        DP_OP_5187J1_124_3275_n58), .B(DP_OP_5187J1_124_3275_n6), .Y(
        DP_OP_5187J1_124_3275_n56) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U174 ( .A(
        DP_OP_5187J1_124_3275_n169), .B(DP_OP_5187J1_124_3275_n176), .Y(
        DP_OP_5187J1_124_3275_n167) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U178 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[19]), .B(u0_0_leon3x0_p0_div0_b[19]), .Y(
        DP_OP_5187J1_124_3275_n169) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U164 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[20]), .B(u0_0_leon3x0_p0_div0_b[20]), .Y(
        DP_OP_5187J1_124_3275_n158) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U140 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[22]), .B(u0_0_leon3x0_p0_div0_b[22]), .Y(
        DP_OP_5187J1_124_3275_n138) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U128 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[23]), .B(u0_0_leon3x0_p0_div0_b[23]), .Y(
        DP_OP_5187J1_124_3275_n131) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U16 ( .A(
        DP_OP_5187J1_124_3275_n47), .B(DP_OP_5187J1_124_3275_n6), .Y(
        DP_OP_5187J1_124_3275_n45) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U100 ( .A(
        DP_OP_5187J1_124_3275_n113), .B(DP_OP_5187J1_124_3275_n120), .Y(
        DP_OP_5187J1_124_3275_n107) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U114 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[24]), .B(u0_0_leon3x0_p0_div0_b[24]), .Y(
        DP_OP_5187J1_124_3275_n120) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U104 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[25]), .B(u0_0_leon3x0_p0_div0_b[25]), .Y(
        DP_OP_5187J1_124_3275_n113) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U74 ( .A(
        DP_OP_5187J1_124_3275_n93), .B(DP_OP_5187J1_124_3275_n100), .Y(
        DP_OP_5187J1_124_3275_n91) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U90 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[26]), .B(u0_0_leon3x0_p0_div0_b[26]), .Y(
        DP_OP_5187J1_124_3275_n100) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U78 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[27]), .B(u0_0_leon3x0_p0_div0_b[27]), .Y(
        DP_OP_5187J1_124_3275_n93) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U48 ( .A(
        DP_OP_5187J1_124_3275_n73), .B(DP_OP_5187J1_124_3275_n80), .Y(
        DP_OP_5187J1_124_3275_n71) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U64 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[28]), .B(u0_0_leon3x0_p0_div0_b[28]), .Y(
        DP_OP_5187J1_124_3275_n80) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U52 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[29]), .B(u0_0_leon3x0_p0_div0_b[29]), .Y(
        DP_OP_5187J1_124_3275_n73) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U38 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[30]), .B(u0_0_leon3x0_p0_div0_b[30]), .Y(
        DP_OP_5187J1_124_3275_n62) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U24 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[31]), .B(u0_0_leon3x0_p0_div0_b[31]), .Y(
        DP_OP_5187J1_124_3275_n51) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U198 ( .A(
        DP_OP_5187J1_124_3275_n187), .B(DP_OP_5187J1_124_3275_n190), .Y(
        DP_OP_5187J1_124_3275_n181) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U188 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[18]), .B(u0_0_leon3x0_p0_div0_b[18]), .Y(
        DP_OP_5187J1_124_3275_n176) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U329 ( .A(
        DP_OP_5187J1_124_3275_n282), .B(DP_OP_5187J1_124_3275_n287), .Y(
        DP_OP_5187J1_124_3275_n276) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U341 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[4]), .B(u0_0_leon3x0_p0_div0_b[4]), .Y(
        DP_OP_5187J1_124_3275_n287) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U311 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[7]), .B(u0_0_leon3x0_p0_div0_b[7]), .Y(
        DP_OP_5187J1_124_3275_n266) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U363 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[1]), .B(u0_0_leon3x0_p0_div0_b[1]), .Y(
        DP_OP_5187J1_124_3275_n300) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U346 ( .A(
        DP_OP_5187J1_124_3275_n293), .B(DP_OP_5187J1_124_3275_n296), .Y(
        DP_OP_5187J1_124_3275_n291) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U356 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[2]), .B(u0_0_leon3x0_p0_div0_b[2]), .Y(
        DP_OP_5187J1_124_3275_n296) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U350 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[3]), .B(u0_0_leon3x0_p0_div0_b[3]), .Y(
        DP_OP_5187J1_124_3275_n293) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U212 ( .A(
        DP_OP_5187J1_124_3275_n195), .B(DP_OP_5187J1_124_3275_n229), .Y(
        DP_OP_5187J1_124_3275_n193) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U280 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[10]), .B(u0_0_leon3x0_p0_div0_b[10]), .Y(
        DP_OP_5187J1_124_3275_n244) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U270 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[11]), .B(u0_0_leon3x0_p0_div0_b[11]), .Y(
        DP_OP_5187J1_124_3275_n237) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U256 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[12]), .B(u0_0_leon3x0_p0_div0_b[12]), .Y(
        DP_OP_5187J1_124_3275_n226) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U216 ( .A(
        DP_OP_5187J1_124_3275_n199), .B(DP_OP_5187J1_124_3275_n206), .Y(
        DP_OP_5187J1_124_3275_n197) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U220 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[15]), .B(u0_0_leon3x0_p0_div0_b[15]), .Y(
        DP_OP_5187J1_124_3275_n199) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U208 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[16]), .B(u0_0_leon3x0_p0_div0_b[16]), .Y(
        DP_OP_5187J1_124_3275_n190) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U202 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[17]), .B(u0_0_leon3x0_p0_div0_b[17]), .Y(
        DP_OP_5187J1_124_3275_n187) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U20 ( .A(
        DP_OP_5187J1_124_3275_n51), .B(DP_OP_5187J1_124_3275_n62), .Y(
        DP_OP_5187J1_124_3275_n49) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U134 ( .A(
        DP_OP_5187J1_124_3275_n138), .B(DP_OP_5187J1_124_3275_n147), .Y(
        DP_OP_5187J1_124_3275_n136) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U315 ( .A(
        DP_OP_5187J1_124_3275_n271), .B(DP_OP_5187J1_124_3275_n278), .Y(
        DP_OP_5187J1_124_3275_n269) );
  NOR2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U370 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[0]), .B(u0_0_leon3x0_p0_div0_vaddsub), 
        .Y(DP_OP_5187J1_124_3275_n304) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U343 ( .A(
        DP_OP_5187J1_124_3275_n36), .B(DP_OP_5187J1_124_3275_n295), .Y(
        u0_0_leon3x0_p0_div0_addout_3_) );
  XOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U323 ( .A(
        DP_OP_5187J1_124_3275_n34), .B(DP_OP_5187J1_124_3275_n284), .Y(
        u0_0_leon3x0_p0_div0_addout_5_) );
  XOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U302 ( .A(
        DP_OP_5187J1_124_3275_n32), .B(DP_OP_5187J1_124_3275_n268), .Y(
        u0_0_leon3x0_p0_div0_addout_7_) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U282 ( .A(
        DP_OP_5187J1_124_3275_n30), .B(DP_OP_5187J1_124_3275_n257), .Y(
        u0_0_leon3x0_p0_div0_addout_9_) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U248 ( .A(
        DP_OP_5187J1_124_3275_n27), .B(DP_OP_5187J1_124_3275_n228), .Y(
        u0_0_leon3x0_p0_div0_addout_12_) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U234 ( .A(
        DP_OP_5187J1_124_3275_n26), .B(DP_OP_5187J1_124_3275_n221), .Y(
        u0_0_leon3x0_p0_div0_addout_13_) );
  XOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U204 ( .A(
        DP_OP_5187J1_124_3275_n23), .B(n22225), .Y(
        u0_0_leon3x0_p0_div0_addout_16_) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U92 ( .A(
        DP_OP_5187J1_124_3275_n14), .B(DP_OP_5187J1_124_3275_n115), .Y(
        u0_0_leon3x0_p0_div0_addout_25_) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U80 ( .A(
        DP_OP_5187J1_124_3275_n13), .B(DP_OP_5187J1_124_3275_n104), .Y(
        u0_0_leon3x0_p0_div0_addout_26_) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U54 ( .A(
        DP_OP_5187J1_124_3275_n11), .B(DP_OP_5187J1_124_3275_n84), .Y(
        u0_0_leon3x0_p0_div0_addout_28_) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U12 ( .A(
        DP_OP_5187J1_124_3275_n8), .B(DP_OP_5187J1_124_3275_n53), .Y(
        u0_0_leon3x0_p0_div0_addout_31_) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U49 ( .A(add_x_735_n8), .B(add_x_735_n76), 
        .Y(u0_0_leon3x0_p0_dci[32]) );
  XOR2xp5_ASAP7_75t_SL add_x_735_U295 ( .A(add_x_735_n30), .B(add_x_735_n252), 
        .Y(u0_0_leon3x0_p0_dci[10]) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U286 ( .A(add_x_735_n29), .B(add_x_735_n249), 
        .Y(u0_0_leon3x0_p0_dci[11]) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U191 ( .A(add_x_735_n20), .B(add_x_735_n182), 
        .Y(u0_0_leon3x0_p0_dci[20]) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U17 ( .A(add_x_735_n54), .B(add_x_735_n47), 
        .Y(add_x_735_n45) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U35 ( .A(add_x_735_n7), .B(add_x_735_n69), 
        .Y(u0_0_leon3x0_p0_dci[33]) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U67 ( .A(add_x_735_n92), .B(add_x_735_n85), 
        .Y(add_x_735_n83) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U33 ( .A(n22968), .B(
        u0_0_leon3x0_p0_divi[28]), .Y(add_x_735_n54) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U73 ( .A(add_x_735_n10), .B(add_x_735_n96), 
        .Y(u0_0_leon3x0_p0_dci[30]) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U83 ( .A(n18606), .B(
        u0_0_leon3x0_p0_divi[24]), .Y(add_x_735_n92) );
  NAND2xp33_ASAP7_75t_SRAM add_x_735_U84 ( .A(n18606), .B(
        u0_0_leon3x0_p0_divi[24]), .Y(add_x_735_n95) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U109 ( .A(add_x_735_n13), .B(add_x_735_n125), 
        .Y(u0_0_leon3x0_p0_dci[27]) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U99 ( .A(add_x_735_n12), .B(add_x_735_n114), 
        .Y(u0_0_leon3x0_p0_dci[28]) );
  NAND2xp33_ASAP7_75t_SRAM add_x_735_U108 ( .A(n18296), .B(
        u0_0_leon3x0_p0_divi[22]), .Y(add_x_735_n113) );
  NAND2xp33_ASAP7_75t_SRAM add_x_735_U152 ( .A(n24231), .B(
        u0_0_leon3x0_p0_divi[18]), .Y(add_x_735_n145) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U159 ( .A(add_x_735_n160), .B(add_x_735_n153), .Y(add_x_735_n151) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U163 ( .A(add_x_735_A_19_), .B(
        u0_0_leon3x0_p0_divi[17]), .Y(add_x_735_n153) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U117 ( .A(add_x_735_n130), .B(add_x_735_n123), .Y(add_x_735_n121) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U141 ( .A(add_x_735_n144), .B(add_x_735_n141), .Y(add_x_735_n135) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U151 ( .A(n24231), .B(
        u0_0_leon3x0_p0_divi[18]), .Y(add_x_735_n144) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U107 ( .A(n18296), .B(
        u0_0_leon3x0_p0_divi[22]), .Y(add_x_735_n112) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U97 ( .A(n23002), .B(
        u0_0_leon3x0_p0_divi[23]), .Y(add_x_735_n105) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U165 ( .A(add_x_735_n18), .B(add_x_735_n164), 
        .Y(u0_0_leon3x0_p0_dci[22]) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U175 ( .A(n23965), .B(
        u0_0_leon3x0_p0_divi[16]), .Y(add_x_735_n160) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U177 ( .A(add_x_735_n19), .B(add_x_735_n175), 
        .Y(u0_0_leon3x0_p0_dci[21]) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U215 ( .A(add_x_735_n22), .B(add_x_735_n200), 
        .Y(u0_0_leon3x0_p0_dci[18]) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U284 ( .A(n18588), .B(
        u0_0_leon3x0_p0_divi[6]), .Y(add_x_735_n241) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U250 ( .A(add_x_735_n225), .B(add_x_735_n220), .Y(add_x_735_n218) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U310 ( .A(add_x_735_n262), .B(add_x_735_n259), .Y(add_x_735_n257) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U306 ( .A(u0_0_leon3x0_p0_muli[41]), .B(
        u0_0_leon3x0_p0_divi[3]), .Y(add_x_735_n254) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U289 ( .A(add_x_735_n247), .B(add_x_735_n250), .Y(add_x_735_n245) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U299 ( .A(n23958), .B(
        u0_0_leon3x0_p0_divi[4]), .Y(add_x_735_n250) );
  NAND2xp33_ASAP7_75t_SRAM add_x_735_U8 ( .A(add_x_735_A_32_), .B(
        u0_0_leon3x0_p0_divi[30]), .Y(add_x_735_n37) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U308 ( .A(add_x_735_n32), .B(add_x_735_n261), 
        .Y(u0_0_leon3x0_p0_dci[8]) );
  XOR2xp5_ASAP7_75t_SL add_x_735_U239 ( .A(add_x_735_n24), .B(add_x_735_n214), 
        .Y(u0_0_leon3x0_p0_dci[16]) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U169 ( .A(n18888), .B(n18898), .Y(
        add_x_735_n158) );
  NOR2xp33_ASAP7_75t_SL add_x_735_U258 ( .A(add_x_735_n225), .B(add_x_735_n232), .Y(add_x_735_n223) );
  XNOR2xp5_ASAP7_75t_SL add_x_735_U153 ( .A(add_x_735_n17), .B(add_x_735_n155), 
        .Y(u0_0_leon3x0_p0_dci[23]) );
  XOR2xp5_ASAP7_75t_SL add_x_735_U147 ( .A(add_x_735_n16), .B(n22228), .Y(
        u0_0_leon3x0_p0_dci[24]) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U864 ( .A(mult_x_1196_n282), .B(
        mult_x_1196_n759), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N8) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U828 ( .A(n23889), .B(mult_x_1196_n278), 
        .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N12) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U820 ( .A(mult_x_1196_n729), .B(
        mult_x_1196_n277), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N13) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U782 ( .A(mult_x_1196_n701), .B(n24310), 
        .Y(mult_x_1196_n272) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U771 ( .A(mult_x_1196_n693), .B(
        mult_x_1196_n821), .Y(mult_x_1196_n271) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U756 ( .A(mult_x_1196_n684), .B(
        mult_x_1196_n819), .Y(mult_x_1196_n269) );
  AOI21xp33_ASAP7_75t_SRAM mult_x_1196_U745 ( .A1(n23886), .A2(
        mult_x_1196_n676), .B(n18923), .Y(mult_x_1196_n675) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U684 ( .A(mult_x_1196_n636), .B(n24304), 
        .Y(mult_x_1196_n261) );
  OAI21xp33_ASAP7_75t_SRAM mult_x_1196_U621 ( .A1(mult_x_1196_n591), .A2(
        mult_x_1196_n599), .B(n22503), .Y(mult_x_1196_n590) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U614 ( .A(mult_x_1196_n587), .B(
        mult_x_1196_n804), .Y(mult_x_1196_n254) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U709 ( .A(mult_x_1196_n814), .B(
        mult_x_1196_n652), .Y(mult_x_1196_n264) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U603 ( .A(mult_x_1196_n579), .B(
        mult_x_1196_n803), .Y(mult_x_1196_n253) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U511 ( .A(mult_x_1196_n507), .B(
        mult_x_1196_n795), .Y(mult_x_1196_n245) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U653 ( .A(mult_x_1196_n614), .B(
        mult_x_1196_n808), .Y(mult_x_1196_n258) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U573 ( .A(mult_x_1196_n558), .B(
        mult_x_1196_n800), .Y(mult_x_1196_n250) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U549 ( .A(mult_x_1196_n540), .B(
        mult_x_1196_n798), .Y(mult_x_1196_n248) );
  AOI21xp33_ASAP7_75t_SRAM mult_x_1196_U542 ( .A1(mult_x_1196_n552), .A2(
        n22264), .B(n18914), .Y(mult_x_1196_n532) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1946 ( .A1(mult_x_1196_n2841), .A2(
        n24031), .B1(n24030), .B2(mult_x_1196_n2840), .Y(mult_x_1196_n2275) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1739 ( .A1(mult_x_1196_n2745), .A2(
        n24041), .B1(n24040), .B2(mult_x_1196_n2744), .Y(mult_x_1196_n2182) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1738 ( .A1(mult_x_1196_n2744), .A2(
        n24041), .B1(n24040), .B2(mult_x_1196_n2743), .Y(mult_x_1196_n2181) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1737 ( .A1(mult_x_1196_n2743), .A2(
        n24041), .B1(n24040), .B2(mult_x_1196_n2742), .Y(mult_x_1196_n2180) );
  NOR2xp33_ASAP7_75t_SL mult_x_1196_U247 ( .A(mult_x_1196_n851), .B(
        mult_x_1196_n848), .Y(mult_x_1196_n301) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1700 ( .A(n18615), .B(n22642), .Y(
        mult_x_1196_n2708) );
  AO21x1_ASAP7_75t_SL mult_x_1196_U1873 ( .A1(n18402), .A2(n24034), .B(
        mult_x_1196_n2805), .Y(mult_x_1196_n2239) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1735 ( .A1(mult_x_1196_n2741), .A2(
        n18364), .B1(n24040), .B2(mult_x_1196_n2740), .Y(mult_x_1196_n2178) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1770 ( .A(n24048), .B(n23976), .Y(
        mult_x_1196_n2741) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1804 ( .A1(mult_x_1196_n2773), .A2(
        n22509), .B1(mult_x_1196_n2772), .B2(n22481), .Y(mult_x_1196_n2210) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1803 ( .A1(n22481), .A2(
        mult_x_1196_n2771), .B1(mult_x_1196_n2772), .B2(n22412), .Y(
        mult_x_1196_n2209) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1734 ( .A1(mult_x_1196_n2740), .A2(
        n24041), .B1(n24040), .B2(mult_x_1196_n2739), .Y(mult_x_1196_n2177) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1768 ( .A(n24046), .B(n23976), .Y(
        mult_x_1196_n2739) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1769 ( .A(n24047), .B(n23976), .Y(
        mult_x_1196_n2740) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U2537 ( .A1(mult_x_1196_n3136), .A2(
        n23999), .B1(n23996), .B2(mult_x_1196_n3135), .Y(mult_x_1196_n2560) );
  XOR2xp5_ASAP7_75t_SL mult_x_1196_U1589 ( .A(mult_x_1196_n2529), .B(
        mult_x_1196_n2689), .Y(mult_x_1196_n1985) );
  NOR2xp33_ASAP7_75t_SL mult_x_1196_U877 ( .A(mult_x_1196_n2091), .B(
        mult_x_1196_n2088), .Y(mult_x_1196_n760) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2505 ( .A(n24073), .B(n23091), .Y(
        mult_x_1196_n3106) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2506 ( .A(n24074), .B(n23091), .Y(
        mult_x_1196_n3107) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2507 ( .A(n24075), .B(n23091), .Y(
        mult_x_1196_n3108) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2504 ( .A(n24072), .B(n23091), .Y(
        mult_x_1196_n3105) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2503 ( .A(n24071), .B(n23091), .Y(
        mult_x_1196_n3104) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2502 ( .A(n24070), .B(n23091), .Y(
        mult_x_1196_n3103) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2771 ( .A(n24055), .B(n23955), .Y(
        mult_x_1196_n3224) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2770 ( .A(n24054), .B(n23955), .Y(
        mult_x_1196_n3223) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2354 ( .A(n24064), .B(n23964), .Y(
        mult_x_1196_n3029) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2355 ( .A(n24065), .B(n23964), .Y(
        mult_x_1196_n3030) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2010 ( .A(n24075), .B(n23971), .Y(
        mult_x_1196_n2870) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2699 ( .A(n24054), .B(n23957), .Y(
        mult_x_1196_n3189) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2630 ( .A(n24056), .B(n23960), .Y(
        mult_x_1196_n3157) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2007 ( .A(n18306), .B(n23971), .Y(
        mult_x_1196_n2867) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2283 ( .A(n24064), .B(n23965), .Y(
        mult_x_1196_n2995) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2284 ( .A(n24065), .B(n23965), .Y(
        mult_x_1196_n2996) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2628 ( .A(n24054), .B(n23960), .Y(
        mult_x_1196_n3155) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2629 ( .A(n24055), .B(n23960), .Y(
        mult_x_1196_n3156) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2767 ( .A(n24051), .B(n23955), .Y(
        mult_x_1196_n3220) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2076 ( .A(n24070), .B(n23089), .Y(
        mult_x_1196_n2899) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2766 ( .A(n24050), .B(n22449), .Y(
        mult_x_1196_n3219) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2695 ( .A(n24050), .B(n23957), .Y(
        mult_x_1196_n3185) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1936 ( .A(n24072), .B(n22395), .Y(
        mult_x_1196_n2833) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2626 ( .A(n24052), .B(n23960), .Y(
        mult_x_1196_n3153) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2281 ( .A(n24062), .B(n23965), .Y(
        mult_x_1196_n2993) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2074 ( .A(n24068), .B(n23089), .Y(
        mult_x_1196_n2897) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2764 ( .A(n24048), .B(n23955), .Y(
        mult_x_1196_n3217) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2073 ( .A(n24067), .B(n23089), .Y(
        mult_x_1196_n2896) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2142 ( .A(n24065), .B(n23969), .Y(
        mult_x_1196_n2928) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2625 ( .A(n24051), .B(n23960), .Y(
        mult_x_1196_n3152) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2486 ( .A(n24054), .B(n22394), .Y(
        mult_x_1196_n3087) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2348 ( .A(n24058), .B(n23964), .Y(
        mult_x_1196_n3023) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2278 ( .A(u0_0_leon3x0_p0_muli[25]), .B(
        n23965), .Y(mult_x_1196_n2990) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1934 ( .A(n24070), .B(n22395), .Y(
        mult_x_1196_n2831) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2760 ( .A(n23955), .B(n24044), .Y(
        mult_x_1196_n3213) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2416 ( .A(n24055), .B(n24081), .Y(
        mult_x_1196_n3054) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2622 ( .A(n24048), .B(n23960), .Y(
        mult_x_1196_n3149) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2277 ( .A(n24058), .B(n23965), .Y(
        mult_x_1196_n2989) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2139 ( .A(n24062), .B(n23969), .Y(
        mult_x_1196_n2925) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2485 ( .A(n24053), .B(n22394), .Y(
        mult_x_1196_n3086) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2001 ( .A(n24066), .B(n23971), .Y(
        mult_x_1196_n2861) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2621 ( .A(n24047), .B(n23960), .Y(
        mult_x_1196_n3148) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2276 ( .A(n24057), .B(n23965), .Y(
        mult_x_1196_n2988) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1999 ( .A(n24064), .B(n23971), .Y(
        mult_x_1196_n2859) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U2306 ( .A1(mult_x_1196_n3016), .A2(
        n22815), .B1(mult_x_1196_n3015), .B2(n23442), .Y(mult_x_1196_n2444) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2483 ( .A(n24051), .B(n22394), .Y(
        mult_x_1196_n3084) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2411 ( .A(n24050), .B(n24081), .Y(
        mult_x_1196_n3049) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2134 ( .A(n24057), .B(n23969), .Y(
        mult_x_1196_n2920) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2409 ( .A(n24048), .B(n24081), .Y(
        mult_x_1196_n3047) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2408 ( .A(n24047), .B(n23396), .Y(
        mult_x_1196_n3046) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2339 ( .A(n24049), .B(n23964), .Y(
        mult_x_1196_n3014) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2271 ( .A(n24052), .B(n23965), .Y(
        mult_x_1196_n2983) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1787 ( .A(n24065), .B(n23975), .Y(
        mult_x_1196_n2758) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2479 ( .A(u0_0_leon3x0_p0_muli[35]), .B(
        n22394), .Y(mult_x_1196_n3080) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U2167 ( .A1(mult_x_1196_n2951), .A2(
        n23141), .B1(n24017), .B2(mult_x_1196_n2950), .Y(mult_x_1196_n2379) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1995 ( .A(n24060), .B(n23971), .Y(
        mult_x_1196_n2855) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2338 ( .A(n24048), .B(n23964), .Y(
        mult_x_1196_n3013) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1993 ( .A(n24058), .B(n23971), .Y(
        mult_x_1196_n2853) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1786 ( .A(n24064), .B(n23975), .Y(
        mult_x_1196_n2757) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2337 ( .A(n24047), .B(n23964), .Y(
        mult_x_1196_n3012) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1886 ( .A1(mult_x_1196_n2818), .A2(
        n24035), .B1(n22251), .B2(mult_x_1196_n2817), .Y(mult_x_1196_n2252) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1816 ( .A1(mult_x_1196_n2785), .A2(
        n24039), .B1(mult_x_1196_n2784), .B2(n22936), .Y(mult_x_1196_n2219) );
  AO21x1_ASAP7_75t_SL mult_x_1196_U2299 ( .A1(n22540), .A2(n22815), .B(
        mult_x_1196_n3009), .Y(mult_x_1196_n2437) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1990 ( .A(n24055), .B(n23971), .Y(
        mult_x_1196_n2850) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1991 ( .A(n24056), .B(n23971), .Y(
        mult_x_1196_n2851) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2058 ( .A(n24052), .B(n23089), .Y(
        mult_x_1196_n2881) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U2016 ( .A1(n24025), .A2(
        mult_x_1196_n2873), .B1(mult_x_1196_n2874), .B2(n24026), .Y(
        mult_x_1196_n2308) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1810 ( .A1(mult_x_1196_n2779), .A2(
        n22412), .B1(mult_x_1196_n2778), .B2(n22481), .Y(mult_x_1196_n2213) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1948 ( .A1(mult_x_1196_n2843), .A2(
        n24031), .B1(n24030), .B2(mult_x_1196_n2842), .Y(mult_x_1196_n2277) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U1950 ( .A1(mult_x_1196_n2845), .A2(
        n24031), .B1(n24030), .B2(mult_x_1196_n2844), .Y(mult_x_1196_n2279) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1839 ( .A(n24046), .B(n22968), .Y(
        mult_x_1196_n2773) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2481 ( .A(n24049), .B(n22394), .Y(
        mult_x_1196_n3082) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1997 ( .A(n24062), .B(n23971), .Y(
        mult_x_1196_n2857) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2478 ( .A(n24046), .B(n22394), .Y(
        mult_x_1196_n3079) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1716 ( .A(n24065), .B(n22642), .Y(
        mult_x_1196_n2724) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1785 ( .A(n24063), .B(n23975), .Y(
        mult_x_1196_n2756) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U2543 ( .A1(mult_x_1196_n3142), .A2(
        n18397), .B1(n23996), .B2(mult_x_1196_n3141), .Y(mult_x_1196_n2566) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2341 ( .A(n24051), .B(n23964), .Y(
        mult_x_1196_n3016) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2336 ( .A(n24046), .B(n23964), .Y(
        mult_x_1196_n3011) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2129 ( .A(n24052), .B(n23969), .Y(
        mult_x_1196_n2915) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1983 ( .A(n24048), .B(n23971), .Y(
        mult_x_1196_n2843) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2646 ( .A(n24072), .B(n23960), .Y(
        mult_x_1196_n3173) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2705 ( .A(n24060), .B(n23957), .Y(
        mult_x_1196_n3195) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U816 ( .A(mult_x_1196_n723), .B(n24307), 
        .Y(mult_x_1196_n276) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U805 ( .A(mult_x_1196_n715), .B(
        mult_x_1196_n825), .Y(mult_x_1196_n275) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2852 ( .A(n24065), .B(n18927), .Y(
        mult_x_1196_n3268) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2710 ( .A(n24065), .B(n23957), .Y(
        mult_x_1196_n3200) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2708 ( .A(n24063), .B(n23957), .Y(
        mult_x_1196_n3198) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2702 ( .A(n24057), .B(n23957), .Y(
        mult_x_1196_n3192) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2698 ( .A(n24053), .B(n23957), .Y(
        mult_x_1196_n3188) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2274 ( .A(n24055), .B(n23050), .Y(
        mult_x_1196_n2986) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1982 ( .A(n24047), .B(n23971), .Y(
        mult_x_1196_n2842) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2703 ( .A(n24058), .B(n23957), .Y(
        mult_x_1196_n3193) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1981 ( .A(n24046), .B(n23971), .Y(
        mult_x_1196_n2841) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2696 ( .A(n24051), .B(n23957), .Y(
        mult_x_1196_n3186) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2694 ( .A(n24049), .B(n23957), .Y(
        mult_x_1196_n3184) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2405 ( .A(n23396), .B(n24044), .Y(
        mult_x_1196_n3043) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2334 ( .A(n23964), .B(n24044), .Y(
        mult_x_1196_n3009) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1843 ( .A(n24050), .B(n22968), .Y(
        mult_x_1196_n2777) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1979 ( .A(n23971), .B(n24044), .Y(
        mult_x_1196_n2839) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1837 ( .A(n22968), .B(n18541), .Y(
        mult_x_1196_n2771) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U2828 ( .A1(mult_x_1196_n3279), .A2(
        n23982), .B1(n23980), .B2(mult_x_1196_n3278), .Y(mult_x_1196_n2703) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2476 ( .A(n22394), .B(
        u0_0_leon3x0_p0_muli[37]), .Y(mult_x_1196_n3077) );
  OAI22xp33_ASAP7_75t_SRAM mult_x_1196_U2795 ( .A1(n22389), .A2(
        mult_x_1196_n3280), .B1(n18614), .B2(n23981), .Y(mult_x_1196_n2143) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U833 ( .A(mult_x_1196_n734), .B(n24290), 
        .Y(mult_x_1196_n278) );
  NAND2xp33_ASAP7_75t_SRAM mult_x_1196_U824 ( .A(mult_x_1196_n728), .B(n24276), 
        .Y(mult_x_1196_n277) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U2367 ( .A(n22227), .B(n18299), .Y(
        mult_x_1196_n3042) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U2580 ( .A(n22227), .B(n23643), .Y(
        mult_x_1196_n3144) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U2864 ( .A(n22227), .B(n18614), .Y(
        mult_x_1196_n3280) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U2687 ( .A(n22227), .B(n23986), .Y(
        mult_x_1196_n2636) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U2651 ( .A(n22227), .B(n18414), .Y(
        mult_x_1196_n3178) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U2722 ( .A(n22227), .B(n23956), .Y(
        mult_x_1196_n3212) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U2403 ( .A(n22227), .B(n24004), .Y(
        mult_x_1196_n2504) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U2474 ( .A(n22227), .B(n24001), .Y(
        mult_x_1196_n2534) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U2296 ( .A(n22227), .B(n22216), .Y(
        mult_x_1196_n3008) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U2119 ( .A(n22227), .B(n18563), .Y(
        mult_x_1196_n2368) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U2048 ( .A(n22227), .B(n18536), .Y(
        mult_x_1196_n2334) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U2083 ( .A(n22227), .B(n18604), .Y(
        mult_x_1196_n2906) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U2012 ( .A(n22227), .B(n24691), .Y(
        mult_x_1196_n2872) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U1941 ( .A(n22227), .B(n22918), .Y(
        mult_x_1196_n2838) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U1799 ( .A(n22227), .B(n23974), .Y(
        mult_x_1196_n2770) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U1870 ( .A(n22227), .B(n23479), .Y(
        mult_x_1196_n2804) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U1764 ( .A(n22227), .B(n18339), .Y(
        mult_x_1196_n2207) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U1694 ( .A(n22227), .B(n24042), .Y(
        mult_x_1196_n2173) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2851 ( .A(n24064), .B(n18927), .Y(
        mult_x_1196_n3267) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2850 ( .A(n24063), .B(n18927), .Y(
        mult_x_1196_n3266) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2849 ( .A(n24062), .B(n18927), .Y(
        mult_x_1196_n3265) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2848 ( .A(n24061), .B(add_x_735_A_2_), 
        .Y(mult_x_1196_n3264) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2840 ( .A(n24053), .B(n18927), .Y(
        mult_x_1196_n3256) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2838 ( .A(n24051), .B(n18926), .Y(
        mult_x_1196_n3254) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2837 ( .A(n24050), .B(n18927), .Y(
        mult_x_1196_n3253) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2836 ( .A(n24049), .B(n18927), .Y(
        mult_x_1196_n3252) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2787 ( .A(n24071), .B(n23955), .Y(
        mult_x_1196_n3240) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2786 ( .A(n24070), .B(n23955), .Y(
        mult_x_1196_n3239) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2785 ( .A(n24069), .B(n23955), .Y(
        mult_x_1196_n3238) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2784 ( .A(n24068), .B(n23955), .Y(
        mult_x_1196_n3237) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2783 ( .A(n24067), .B(n23955), .Y(
        mult_x_1196_n3236) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2772 ( .A(n24056), .B(n23955), .Y(
        mult_x_1196_n3225) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2769 ( .A(n24053), .B(n23955), .Y(
        mult_x_1196_n3222) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2768 ( .A(n24052), .B(n23955), .Y(
        mult_x_1196_n3221) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2763 ( .A(n24047), .B(n23955), .Y(
        mult_x_1196_n3216) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2762 ( .A(n24046), .B(n23955), .Y(
        mult_x_1196_n3215) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2721 ( .A(n23957), .B(n22227), .Y(
        mult_x_1196_n3211) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2691 ( .A(n24046), .B(n23957), .Y(
        mult_x_1196_n3181) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2650 ( .A(n22227), .B(n23960), .Y(
        mult_x_1196_n3177) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2649 ( .A(n24075), .B(n23960), .Y(
        mult_x_1196_n3176) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2648 ( .A(n24074), .B(n23960), .Y(
        mult_x_1196_n3175) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2647 ( .A(n24073), .B(n23960), .Y(
        mult_x_1196_n3174) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2645 ( .A(n24071), .B(n23960), .Y(
        mult_x_1196_n3172) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2644 ( .A(n24070), .B(n23960), .Y(
        mult_x_1196_n3171) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2643 ( .A(n24069), .B(n23960), .Y(
        mult_x_1196_n3170) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2642 ( .A(n24068), .B(n23960), .Y(
        mult_x_1196_n3169) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2641 ( .A(n24067), .B(n23960), .Y(
        mult_x_1196_n3168) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2627 ( .A(n24053), .B(n23960), .Y(
        mult_x_1196_n3154) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2579 ( .A(n22227), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3143) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2578 ( .A(n24075), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3142) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2577 ( .A(n24074), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3141) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2574 ( .A(n24071), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3138) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2573 ( .A(n24070), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3137) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2572 ( .A(n24069), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3136) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2571 ( .A(n24068), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3135) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2569 ( .A(n24066), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3133) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2568 ( .A(n24065), .B(n23658), .Y(
        mult_x_1196_n3132) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2567 ( .A(n24064), .B(n23658), .Y(
        mult_x_1196_n3131) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2566 ( .A(n24063), .B(n23658), .Y(
        mult_x_1196_n3130) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2564 ( .A(n24061), .B(n22448), .Y(
        mult_x_1196_n3128) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2563 ( .A(n24060), .B(n23658), .Y(
        mult_x_1196_n3127) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2560 ( .A(n22442), .B(n23658), .Y(
        mult_x_1196_n3124) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2508 ( .A(n22394), .B(n22227), .Y(
        mult_x_1196_n3109) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2501 ( .A(n24069), .B(n23091), .Y(
        mult_x_1196_n3102) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2496 ( .A(n24064), .B(n22394), .Y(
        mult_x_1196_n3097) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2494 ( .A(n24062), .B(n22394), .Y(
        mult_x_1196_n3095) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2493 ( .A(n24061), .B(n22394), .Y(
        mult_x_1196_n3094) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2492 ( .A(n24060), .B(n22394), .Y(
        mult_x_1196_n3093) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2488 ( .A(n24056), .B(n22394), .Y(
        mult_x_1196_n3089) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2437 ( .A(n22227), .B(n23396), .Y(
        mult_x_1196_n3075) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2435 ( .A(n24074), .B(n24081), .Y(
        mult_x_1196_n3073) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2434 ( .A(n24081), .B(n24073), .Y(
        mult_x_1196_n3072) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2433 ( .A(n24072), .B(n23396), .Y(
        mult_x_1196_n3071) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2432 ( .A(n24071), .B(n24081), .Y(
        mult_x_1196_n3070) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2430 ( .A(n24069), .B(n24081), .Y(
        mult_x_1196_n3068) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2427 ( .A(n24066), .B(n24081), .Y(
        mult_x_1196_n3065) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2424 ( .A(n24063), .B(n24081), .Y(
        mult_x_1196_n3062) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2422 ( .A(n24061), .B(n24081), .Y(
        mult_x_1196_n3060) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2421 ( .A(n24060), .B(n23396), .Y(
        mult_x_1196_n3059) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2420 ( .A(n24059), .B(n23396), .Y(
        mult_x_1196_n3058) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2419 ( .A(n24058), .B(n23396), .Y(
        mult_x_1196_n3057) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2415 ( .A(n24054), .B(n23396), .Y(
        mult_x_1196_n3053) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2410 ( .A(n18615), .B(n23396), .Y(
        mult_x_1196_n3048) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2353 ( .A(n24063), .B(n23964), .Y(
        mult_x_1196_n3028) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2352 ( .A(n24062), .B(n23964), .Y(
        mult_x_1196_n3027) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2350 ( .A(n24060), .B(n23964), .Y(
        mult_x_1196_n3025) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2343 ( .A(n24053), .B(n23964), .Y(
        mult_x_1196_n3018) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2340 ( .A(n24050), .B(n23964), .Y(
        mult_x_1196_n3015) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2295 ( .A(n22227), .B(n23965), .Y(
        mult_x_1196_n3007) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2294 ( .A(n24075), .B(n23965), .Y(
        mult_x_1196_n3006) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2291 ( .A(n24072), .B(n23965), .Y(
        mult_x_1196_n3003) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2290 ( .A(n24071), .B(n23965), .Y(
        mult_x_1196_n3002) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2288 ( .A(n24069), .B(n23965), .Y(
        mult_x_1196_n3000) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2286 ( .A(n24067), .B(n23965), .Y(
        mult_x_1196_n2998) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2285 ( .A(n24066), .B(n23965), .Y(
        mult_x_1196_n2997) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2280 ( .A(n24061), .B(n23965), .Y(
        mult_x_1196_n2992) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2273 ( .A(n24054), .B(n23050), .Y(
        mult_x_1196_n2985) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2272 ( .A(n24053), .B(n23050), .Y(
        mult_x_1196_n2984) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2270 ( .A(n24051), .B(n23050), .Y(
        mult_x_1196_n2982) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2269 ( .A(n18788), .B(n23050), .Y(
        mult_x_1196_n2981) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2268 ( .A(n24049), .B(n23050), .Y(
        mult_x_1196_n2980) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2267 ( .A(n24048), .B(n23050), .Y(
        mult_x_1196_n2979) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2266 ( .A(n24047), .B(n23050), .Y(
        mult_x_1196_n2978) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2265 ( .A(n24046), .B(n23050), .Y(
        mult_x_1196_n2977) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2264 ( .A(n24045), .B(n23050), .Y(
        mult_x_1196_n2976) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2263 ( .A(n23050), .B(n24044), .Y(
        mult_x_1196_n2975) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2213 ( .A(n24065), .B(n23967), .Y(
        mult_x_1196_n2962) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2212 ( .A(n24064), .B(n23967), .Y(
        mult_x_1196_n2961) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2210 ( .A(n24062), .B(n24231), .Y(
        mult_x_1196_n2959) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2209 ( .A(n24061), .B(n23967), .Y(
        mult_x_1196_n2958) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2208 ( .A(n24060), .B(n23967), .Y(
        mult_x_1196_n2957) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2207 ( .A(n24059), .B(n23967), .Y(
        mult_x_1196_n2956) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2203 ( .A(n24055), .B(n24231), .Y(
        mult_x_1196_n2952) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2202 ( .A(n24054), .B(n23967), .Y(
        mult_x_1196_n2951) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2201 ( .A(n24053), .B(n24231), .Y(
        mult_x_1196_n2950) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2199 ( .A(n24051), .B(n23967), .Y(
        mult_x_1196_n2948) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2198 ( .A(n24050), .B(n24231), .Y(
        mult_x_1196_n2947) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2197 ( .A(n18615), .B(n24231), .Y(
        mult_x_1196_n2946) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2196 ( .A(n24048), .B(n24231), .Y(
        mult_x_1196_n2945) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2195 ( .A(n24047), .B(n24231), .Y(
        mult_x_1196_n2944) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2194 ( .A(n24046), .B(n24231), .Y(
        mult_x_1196_n2943) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2193 ( .A(n24045), .B(n24231), .Y(
        mult_x_1196_n2942) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2192 ( .A(n24231), .B(n18541), .Y(
        mult_x_1196_n2941) );
  AO21x1_ASAP7_75t_SL mult_x_1196_U2157 ( .A1(n22694), .A2(n22779), .B(
        mult_x_1196_n2941), .Y(mult_x_1196_n2369) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2153 ( .A(n22227), .B(n23969), .Y(
        mult_x_1196_n2939) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2152 ( .A(n24075), .B(n23969), .Y(
        mult_x_1196_n2938) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2150 ( .A(n24073), .B(n23969), .Y(
        mult_x_1196_n2936) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2149 ( .A(n24072), .B(n23969), .Y(
        mult_x_1196_n2935) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2148 ( .A(n24071), .B(n23969), .Y(
        mult_x_1196_n2934) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2147 ( .A(n24070), .B(n23969), .Y(
        mult_x_1196_n2933) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2146 ( .A(n24069), .B(n23969), .Y(
        mult_x_1196_n2932) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2145 ( .A(n24068), .B(n23969), .Y(
        mult_x_1196_n2931) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2144 ( .A(n24067), .B(n23969), .Y(
        mult_x_1196_n2930) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2143 ( .A(n24066), .B(n23969), .Y(
        mult_x_1196_n2929) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2082 ( .A(n22227), .B(n23089), .Y(
        mult_x_1196_n2905) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2081 ( .A(n24075), .B(n23089), .Y(
        mult_x_1196_n2904) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2077 ( .A(n24071), .B(n23089), .Y(
        mult_x_1196_n2900) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2070 ( .A(n24064), .B(n23089), .Y(
        mult_x_1196_n2893) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2069 ( .A(n24063), .B(n23089), .Y(
        mult_x_1196_n2892) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2066 ( .A(n24060), .B(n23089), .Y(
        mult_x_1196_n2889) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2064 ( .A(n24058), .B(n23089), .Y(
        mult_x_1196_n2887) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2062 ( .A(n24056), .B(n23089), .Y(
        mult_x_1196_n2885) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2061 ( .A(n24055), .B(n23089), .Y(
        mult_x_1196_n2884) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2057 ( .A(n24051), .B(n23089), .Y(
        mult_x_1196_n2880) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2056 ( .A(n24050), .B(n23089), .Y(
        mult_x_1196_n2879) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2055 ( .A(n24049), .B(n23089), .Y(
        mult_x_1196_n2878) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2053 ( .A(n24047), .B(n23089), .Y(
        mult_x_1196_n2876) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2052 ( .A(n24046), .B(n23089), .Y(
        mult_x_1196_n2875) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2051 ( .A(n24045), .B(n23089), .Y(
        mult_x_1196_n2874) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2050 ( .A(n23089), .B(n24044), .Y(
        mult_x_1196_n2873) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2011 ( .A(n22227), .B(n23971), .Y(
        mult_x_1196_n2871) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2006 ( .A(n24071), .B(n23971), .Y(
        mult_x_1196_n2866) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2005 ( .A(n24070), .B(n23971), .Y(
        mult_x_1196_n2865) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1996 ( .A(n24061), .B(n23971), .Y(
        mult_x_1196_n2856) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1989 ( .A(n24054), .B(n23971), .Y(
        mult_x_1196_n2849) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1988 ( .A(n24053), .B(n23971), .Y(
        mult_x_1196_n2848) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1987 ( .A(n18556), .B(n23971), .Y(
        mult_x_1196_n2847) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1986 ( .A(n24051), .B(n22897), .Y(
        mult_x_1196_n2846) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1985 ( .A(n24050), .B(n23971), .Y(
        mult_x_1196_n2845) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1984 ( .A(n24049), .B(n23971), .Y(
        mult_x_1196_n2844) );
  AO21x1_ASAP7_75t_SL mult_x_1196_U1944 ( .A1(n22743), .A2(n18309), .B(
        mult_x_1196_n2839), .Y(mult_x_1196_n2273) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1939 ( .A(n24075), .B(n22395), .Y(
        mult_x_1196_n2836) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1938 ( .A(n24074), .B(n22395), .Y(
        mult_x_1196_n2835) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1935 ( .A(n24071), .B(n22395), .Y(
        mult_x_1196_n2832) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1932 ( .A(n24068), .B(n22395), .Y(
        mult_x_1196_n2829) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1927 ( .A(n24063), .B(n22395), .Y(
        mult_x_1196_n2824) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1926 ( .A(n24062), .B(n22395), .Y(
        mult_x_1196_n2823) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1925 ( .A(n24061), .B(n22395), .Y(
        mult_x_1196_n2822) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1924 ( .A(n24060), .B(n22395), .Y(
        mult_x_1196_n2821) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1920 ( .A(n24056), .B(n22395), .Y(
        mult_x_1196_n2817) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1916 ( .A(n24052), .B(n22395), .Y(
        mult_x_1196_n2813) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1912 ( .A(n24048), .B(n18307), .Y(
        mult_x_1196_n2809) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1910 ( .A(n24046), .B(n22395), .Y(
        mult_x_1196_n2807) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1849 ( .A(n24056), .B(n22968), .Y(
        mult_x_1196_n2783) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1848 ( .A(n24055), .B(n22968), .Y(
        mult_x_1196_n2782) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1846 ( .A(n24053), .B(n22968), .Y(
        mult_x_1196_n2780) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1844 ( .A(n24051), .B(n22968), .Y(
        mult_x_1196_n2778) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1842 ( .A(n18615), .B(n22968), .Y(
        mult_x_1196_n2776) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1841 ( .A(n24048), .B(n22968), .Y(
        mult_x_1196_n2775) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1840 ( .A(n24047), .B(n22968), .Y(
        mult_x_1196_n2774) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1798 ( .A(n22227), .B(n22926), .Y(
        mult_x_1196_n2769) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1797 ( .A(n24075), .B(n22926), .Y(
        mult_x_1196_n2768) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1794 ( .A(n24072), .B(n22926), .Y(
        mult_x_1196_n2765) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1793 ( .A(n24071), .B(n22926), .Y(
        mult_x_1196_n2764) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1792 ( .A(n24070), .B(n22926), .Y(
        mult_x_1196_n2763) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1790 ( .A(n24068), .B(n22926), .Y(
        mult_x_1196_n2761) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1789 ( .A(n24067), .B(n22926), .Y(
        mult_x_1196_n2760) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1788 ( .A(n24066), .B(n22926), .Y(
        mult_x_1196_n2759) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1784 ( .A(n24062), .B(n23975), .Y(
        mult_x_1196_n2755) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1782 ( .A(n24060), .B(n23975), .Y(
        mult_x_1196_n2753) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1780 ( .A(n24058), .B(n23975), .Y(
        mult_x_1196_n2751) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1779 ( .A(n22442), .B(n23975), .Y(
        mult_x_1196_n2750) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1778 ( .A(n24056), .B(n23976), .Y(
        mult_x_1196_n2749) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1776 ( .A(n24054), .B(n23976), .Y(
        mult_x_1196_n2747) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1775 ( .A(n24053), .B(n23976), .Y(
        mult_x_1196_n2746) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1774 ( .A(n24052), .B(n22926), .Y(
        mult_x_1196_n2745) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1773 ( .A(n24051), .B(n23976), .Y(
        mult_x_1196_n2744) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1772 ( .A(n24050), .B(n23976), .Y(
        mult_x_1196_n2743) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1771 ( .A(n18615), .B(n23976), .Y(
        mult_x_1196_n2742) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1766 ( .A(n23976), .B(n18541), .Y(
        mult_x_1196_n2737) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1726 ( .A(n24075), .B(n23978), .Y(
        mult_x_1196_n2734) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1725 ( .A(n24074), .B(n23978), .Y(
        mult_x_1196_n2733) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1724 ( .A(n24073), .B(n23978), .Y(
        mult_x_1196_n2732) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1723 ( .A(n24072), .B(n23978), .Y(
        mult_x_1196_n2731) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1722 ( .A(n24071), .B(n23978), .Y(
        mult_x_1196_n2730) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1721 ( .A(n24070), .B(n23978), .Y(
        mult_x_1196_n2729) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1720 ( .A(n24069), .B(n23978), .Y(
        mult_x_1196_n2728) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1719 ( .A(n24068), .B(n23978), .Y(
        mult_x_1196_n2727) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1718 ( .A(n24067), .B(n23978), .Y(
        mult_x_1196_n2726) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1717 ( .A(n24066), .B(n23978), .Y(
        mult_x_1196_n2725) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1715 ( .A(n24064), .B(n22642), .Y(
        mult_x_1196_n2723) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1714 ( .A(n24063), .B(n22642), .Y(
        mult_x_1196_n2722) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1709 ( .A(n24058), .B(n22642), .Y(
        mult_x_1196_n2717) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1702 ( .A(n24051), .B(n23978), .Y(
        mult_x_1196_n2710) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U1661 ( .A(mult_x_1196_n2669), .B(
        mult_x_1196_n2701), .Y(mult_x_1196_n2091) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U1488 ( .A(mult_x_1196_n2521), .B(n23932), 
        .Y(mult_x_1196_n1818) );
  XOR2xp5_ASAP7_75t_SL mult_x_1196_U809 ( .A(mult_x_1196_n276), .B(
        mult_x_1196_n724), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N14) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U794 ( .A(mult_x_1196_n274), .B(
        mult_x_1196_n713), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N16) );
  XOR2xp5_ASAP7_75t_SL mult_x_1196_U775 ( .A(mult_x_1196_n272), .B(
        mult_x_1196_n702), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N18) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U760 ( .A(mult_x_1196_n270), .B(
        mult_x_1196_n691), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N20) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U752 ( .A(mult_x_1196_n269), .B(n23886), 
        .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N21) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U713 ( .A(mult_x_1196_n265), .B(
        mult_x_1196_n660), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N25) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U704 ( .A(mult_x_1196_n264), .B(
        mult_x_1196_n653), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N26) );
  XOR2xp5_ASAP7_75t_SL mult_x_1196_U688 ( .A(mult_x_1196_n262), .B(
        mult_x_1196_n642), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N28) );
  XOR2xp5_ASAP7_75t_SL mult_x_1196_U677 ( .A(mult_x_1196_n261), .B(
        mult_x_1196_n637), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N29) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U539 ( .A(mult_x_1196_n248), .B(
        mult_x_1196_n541), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N42) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U491 ( .A(mult_x_1196_n244), .B(
        mult_x_1196_n505), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N46) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U477 ( .A(mult_x_1196_n243), .B(
        mult_x_1196_n494), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N47) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U467 ( .A(mult_x_1196_n242), .B(
        mult_x_1196_n483), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N48) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U425 ( .A(mult_x_1196_n239), .B(
        mult_x_1196_n452), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N51) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U407 ( .A(mult_x_1196_n238), .B(
        mult_x_1196_n443), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N52) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U393 ( .A(mult_x_1196_n237), .B(
        mult_x_1196_n428), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N53) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U333 ( .A(mult_x_1196_n233), .B(
        mult_x_1196_n378), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N57) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U307 ( .A(mult_x_1196_n231), .B(
        mult_x_1196_n356), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N59) );
  XOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U406 ( .A(DP_OP_1196_128_7433_n357), 
        .B(DP_OP_1196_128_7433_n37), .Y(u0_0_leon3x0_p0_iu_N5467) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U48 ( .A(DP_OP_1196_128_7433_n70), 
        .B(DP_OP_1196_128_7433_n77), .Y(DP_OP_1196_128_7433_n68) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U38 ( .A(u0_0_leon3x0_p0_ici[57]), 
        .B(DP_OP_1196_128_7433_n479), .Y(DP_OP_1196_128_7433_n57) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U124 ( .A(DP_OP_1196_128_7433_n128), .B(DP_OP_1196_128_7433_n139), .Y(DP_OP_1196_128_7433_n126) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U172 ( .A(DP_OP_1196_128_7433_n167), .B(DP_OP_1196_128_7433_n178), .Y(DP_OP_1196_128_7433_n165) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U58 ( .A(DP_OP_1196_128_7433_n77), 
        .B(DP_OP_1196_128_7433_n86), .Y(DP_OP_1196_128_7433_n75) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U74 ( .A(DP_OP_1196_128_7433_n90), 
        .B(DP_OP_1196_128_7433_n97), .Y(DP_OP_1196_128_7433_n84) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U78 ( .A(u0_0_leon3x0_p0_ici[54]), 
        .B(DP_OP_1196_128_7433_n476), .Y(DP_OP_1196_128_7433_n90) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U64 ( .A(u0_0_leon3x0_p0_ici[55]), 
        .B(DP_OP_1196_128_7433_n477), .Y(DP_OP_1196_128_7433_n77) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U52 ( .A(u0_0_leon3x0_p0_ici[56]), 
        .B(DP_OP_1196_128_7433_n478), .Y(DP_OP_1196_128_7433_n70) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U94 ( .A(DP_OP_1196_128_7433_n104), 
        .B(DP_OP_1196_128_7433_n338), .Y(DP_OP_1196_128_7433_n8) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U98 ( .A(DP_OP_1196_128_7433_n115), 
        .B(DP_OP_1196_128_7433_n108), .Y(DP_OP_1196_128_7433_n106) );
  NAND2xp33_ASAP7_75t_SRAM DP_OP_1196_128_7433_U119 ( .A(
        u0_0_leon3x0_p0_ici[51]), .B(n18842), .Y(DP_OP_1196_128_7433_n122) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U142 ( .A(DP_OP_1196_128_7433_n232), .B(DP_OP_1196_128_7433_n143), .Y(DP_OP_1196_128_7433_n137) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U146 ( .A(DP_OP_1196_128_7433_n147), .B(DP_OP_1196_128_7433_n154), .Y(DP_OP_1196_128_7433_n145) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U180 ( .A(u0_0_leon3x0_p0_ici[47]), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_), .Y(
        DP_OP_1196_128_7433_n167) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U192 ( .A(DP_OP_1196_128_7433_n184), .B(DP_OP_1196_128_7433_n210), .Y(DP_OP_1196_128_7433_n180) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U132 ( .A(u0_0_leon3x0_p0_ici[50]), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), .Y(
        DP_OP_1196_128_7433_n128) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U102 ( .A(u0_0_leon3x0_p0_ici[52]), 
        .B(DP_OP_1196_128_7433_n474), .Y(DP_OP_1196_128_7433_n108) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U214 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__15_), .B(u0_0_leon3x0_p0_ici[45]), 
        .Y(DP_OP_1196_128_7433_n195) );
  NAND2xp33_ASAP7_75t_SRAM DP_OP_1196_128_7433_U269 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__12_), .B(u0_0_leon3x0_p0_ici[42]), 
        .Y(DP_OP_1196_128_7433_n245) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U260 ( .A(DP_OP_1196_128_7433_n240), .B(DP_OP_1196_128_7433_n266), .Y(DP_OP_1196_128_7433_n238) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U246 ( .A(u0_0_leon3x0_p0_ici[43]), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_), .Y(
        DP_OP_1196_128_7433_n221) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U328 ( .A(DP_OP_1196_128_7433_n296), .B(DP_OP_1196_128_7433_n318), .Y(DP_OP_1196_128_7433_n290) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U350 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__7_), .B(u0_0_leon3x0_p0_ici[37]), 
        .Y(DP_OP_1196_128_7433_n307) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U314 ( .A(u0_0_leon3x0_p0_ici[39]), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__9_), .Y(
        DP_OP_1196_128_7433_n277) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U282 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__11_), .B(u0_0_leon3x0_p0_ici[41]), 
        .Y(DP_OP_1196_128_7433_n251) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U108 ( .A(DP_OP_1196_128_7433_n115), .B(DP_OP_1196_128_7433_n139), .Y(DP_OP_1196_128_7433_n113) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U274 ( .A(DP_OP_1196_128_7433_n251), .B(DP_OP_1196_128_7433_n262), .Y(DP_OP_1196_128_7433_n249) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U238 ( .A(DP_OP_1196_128_7433_n221), .B(DP_OP_1196_128_7433_n232), .Y(DP_OP_1196_128_7433_n219) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U156 ( .A(DP_OP_1196_128_7433_n154), .B(DP_OP_1196_128_7433_n178), .Y(DP_OP_1196_128_7433_n152) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U306 ( .A(DP_OP_1196_128_7433_n277), .B(DP_OP_1196_128_7433_n288), .Y(DP_OP_1196_128_7433_n275) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U206 ( .A(DP_OP_1196_128_7433_n195), .B(DP_OP_1196_128_7433_n206), .Y(DP_OP_1196_128_7433_n193) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U26 ( .A(u0_0_leon3x0_p0_ici[58]), 
        .B(DP_OP_1196_128_7433_n480), .Y(DP_OP_1196_128_7433_n50) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U88 ( .A(u0_0_leon3x0_p0_ici[53]), 
        .B(DP_OP_1196_128_7433_n475), .Y(DP_OP_1196_128_7433_n97) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U411 ( .A(u0_0_leon3x0_p0_ici[31]), 
        .B(DP_OP_1196_128_7433_n453), .Y(DP_OP_1196_128_7433_n354) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U394 ( .A(DP_OP_1196_128_7433_n350), .B(DP_OP_1196_128_7433_n347), .Y(DP_OP_1196_128_7433_n345) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U398 ( .A(u0_0_leon3x0_p0_ici[33]), 
        .B(DP_OP_1196_128_7433_n455), .Y(DP_OP_1196_128_7433_n347) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U404 ( .A(u0_0_leon3x0_p0_ici[32]), 
        .B(DP_OP_1196_128_7433_n454), .Y(DP_OP_1196_128_7433_n350) );
  XOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U400 ( .A(DP_OP_1196_128_7433_n36), 
        .B(DP_OP_1196_128_7433_n352), .Y(u0_0_leon3x0_p0_iu_N5468) );
  XOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U382 ( .A(DP_OP_1196_128_7433_n34), 
        .B(n23941), .Y(u0_0_leon3x0_p0_iu_N5470) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U370 ( .A(DP_OP_1196_128_7433_n33), 
        .B(DP_OP_1196_128_7433_n337), .Y(u0_0_leon3x0_p0_iu_N5471) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U352 ( .A(DP_OP_1196_128_7433_n32), 
        .B(DP_OP_1196_128_7433_n328), .Y(u0_0_leon3x0_p0_iu_N5472) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U338 ( .A(DP_OP_1196_128_7433_n31), 
        .B(DP_OP_1196_128_7433_n313), .Y(u0_0_leon3x0_p0_iu_N5473) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U316 ( .A(DP_OP_1196_128_7433_n30), 
        .B(DP_OP_1196_128_7433_n302), .Y(u0_0_leon3x0_p0_iu_N5474) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U302 ( .A(DP_OP_1196_128_7433_n29), 
        .B(DP_OP_1196_128_7433_n283), .Y(u0_0_leon3x0_p0_iu_N5475) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U284 ( .A(DP_OP_1196_128_7433_n28), 
        .B(DP_OP_1196_128_7433_n272), .Y(u0_0_leon3x0_p0_iu_N5476) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U270 ( .A(DP_OP_1196_128_7433_n27), 
        .B(DP_OP_1196_128_7433_n257), .Y(u0_0_leon3x0_p0_iu_N5477) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U248 ( .A(DP_OP_1196_128_7433_n26), 
        .B(DP_OP_1196_128_7433_n246), .Y(u0_0_leon3x0_p0_iu_N5478) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U216 ( .A(DP_OP_1196_128_7433_n24), 
        .B(DP_OP_1196_128_7433_n216), .Y(u0_0_leon3x0_p0_iu_N5480) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U202 ( .A(DP_OP_1196_128_7433_n23), 
        .B(DP_OP_1196_128_7433_n201), .Y(u0_0_leon3x0_p0_iu_N5481) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U182 ( .A(DP_OP_1196_128_7433_n22), 
        .B(DP_OP_1196_128_7433_n190), .Y(u0_0_leon3x0_p0_iu_N5482) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U168 ( .A(DP_OP_1196_128_7433_n21), 
        .B(DP_OP_1196_128_7433_n173), .Y(u0_0_leon3x0_p0_iu_N5483) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U152 ( .A(DP_OP_1196_128_7433_n20), 
        .B(DP_OP_1196_128_7433_n162), .Y(u0_0_leon3x0_p0_iu_N5484) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U134 ( .A(DP_OP_1196_128_7433_n19), 
        .B(DP_OP_1196_128_7433_n149), .Y(u0_0_leon3x0_p0_iu_N5485) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U120 ( .A(DP_OP_1196_128_7433_n18), 
        .B(DP_OP_1196_128_7433_n134), .Y(u0_0_leon3x0_p0_iu_N5486) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U104 ( .A(DP_OP_1196_128_7433_n17), 
        .B(DP_OP_1196_128_7433_n123), .Y(u0_0_leon3x0_p0_iu_N5487) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U90 ( .A(DP_OP_1196_128_7433_n16), 
        .B(DP_OP_1196_128_7433_n110), .Y(u0_0_leon3x0_p0_iu_N5488) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U66 ( .A(DP_OP_1196_128_7433_n14), 
        .B(DP_OP_1196_128_7433_n92), .Y(u0_0_leon3x0_p0_iu_N5490) );
  XNOR2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U40 ( .A(DP_OP_1196_128_7433_n12), 
        .B(DP_OP_1196_128_7433_n72), .Y(u0_0_leon3x0_p0_iu_N5492) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_F__PC__2_ ( .D(n3202), .CLK(
        clk), .QN(u0_0_leon3x0_p0_ici[60]) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__30_ ( .D(n24439), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__30_) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U1900 ( .A1(mult_x_1196_n2832), .A2(n24034), .B1(n22251), .B2(mult_x_1196_n2831), .Y(mult_x_1196_n2266) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2447 ( .A1(mult_x_1196_n3083), .A2(n18919), .B1(mult_x_1196_n3082), .B2(n24003), .Y(mult_x_1196_n2509) );
  OAI21xp5_ASAP7_75t_SL mult_x_1196_U408 ( .A1(mult_x_1196_n429), .A2(n22533), 
        .B(mult_x_1196_n430), .Y(mult_x_1196_n428) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__43_ ( .D(
        n4223), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[42]) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U1876 ( .A1(mult_x_1196_n2808), .A2(n24034), .B1(n22251), .B2(mult_x_1196_n2807), .Y(mult_x_1196_n2242) );
  FAx1_ASAP7_75t_SL mult_x_1196_U911 ( .A(mult_x_1196_n856), .B(
        mult_x_1196_n2177), .CI(mult_x_1196_n2209), .CON(mult_x_1196_n853), 
        .SN(mult_x_1196_n854) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2309 ( .A1(mult_x_1196_n3019), .A2(n24009), .B1(mult_x_1196_n3018), .B2(n23442), .Y(mult_x_1196_n2447) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2730 ( .A1(n24082), .A2(mult_x_1196_n3218), .B1(mult_x_1196_n3217), .B2(n23984), .Y(mult_x_1196_n2642) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2443 ( .A1(mult_x_1196_n3079), .A2(n18920), .B1(mult_x_1196_n3078), .B2(n24002), .Y(mult_x_1196_n2507) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2301 ( .A1(mult_x_1196_n3011), .A2(n22815), .B1(mult_x_1196_n3010), .B2(n23442), .Y(mult_x_1196_n2439) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2442 ( .A1(n22756), .A2(mult_x_1196_n3077), .B1(mult_x_1196_n3078), .B2(n18920), .Y(mult_x_1196_n2506) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2298 ( .A1(n23442), .A2(mult_x_1196_n3042), .B1(n18299), .B2(n22563), .Y(mult_x_1196_n2136) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2813 ( .A1(mult_x_1196_n3264), .A2(n23982), .B1(n22389), .B2(mult_x_1196_n3263), .Y(mult_x_1196_n2688) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2023 ( .A1(mult_x_1196_n2881), .A2(n22464), .B1(mult_x_1196_n2880), .B2(n24025), .Y(mult_x_1196_n2312) );
  OAI22x1_ASAP7_75t_SL mult_x_1196_U2328 ( .A1(mult_x_1196_n3038), .A2(n22815), 
        .B1(mult_x_1196_n3037), .B2(n22540), .Y(mult_x_1196_n2466) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2382 ( .A1(mult_x_1196_n3055), .A2(n24007), .B1(n24005), .B2(mult_x_1196_n3054), .Y(mult_x_1196_n2483) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2308 ( .A1(mult_x_1196_n3018), .A2(n22815), .B1(mult_x_1196_n3017), .B2(n23442), .Y(mult_x_1196_n2446) );
  XNOR2x1_ASAP7_75t_SL mult_x_1196_U2555 ( .A(n24052), .B(add_x_735_A_10_), 
        .Y(mult_x_1196_n3119) );
  OAI21xp5_ASAP7_75t_SL mult_x_1196_U438 ( .A1(mult_x_1196_n453), .A2(n22258), 
        .B(mult_x_1196_n454), .Y(mult_x_1196_n452) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2390 ( .A1(mult_x_1196_n3063), .A2(n24007), .B1(n24005), .B2(mult_x_1196_n3062), .Y(mult_x_1196_n2491) );
  NOR2x1_ASAP7_75t_SL mult_x_1196_U585 ( .A(mult_x_1196_n1391), .B(
        mult_x_1196_n1358), .Y(mult_x_1196_n564) );
  FAx1_ASAP7_75t_SL mult_x_1196_U918 ( .A(mult_x_1196_n2210), .B(
        mult_x_1196_n875), .CI(mult_x_1196_n2178), .CON(mult_x_1196_n864), 
        .SN(mult_x_1196_n865) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2538 ( .A1(mult_x_1196_n3137), .A2(n23999), .B1(n23996), .B2(mult_x_1196_n3136), .Y(mult_x_1196_n2561) );
  OAI22x1_ASAP7_75t_SL mult_x_1196_U2535 ( .A1(mult_x_1196_n3134), .A2(n18397), 
        .B1(n23997), .B2(mult_x_1196_n3133), .Y(mult_x_1196_n2558) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2182 ( .A1(mult_x_1196_n2966), .A2(n22779), .B1(n22694), .B2(mult_x_1196_n2965), .Y(mult_x_1196_n2394) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U1878 ( .A1(mult_x_1196_n2810), .A2(n24034), .B1(n22251), .B2(mult_x_1196_n2809), .Y(mult_x_1196_n2244) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U1801 ( .A1(n22391), .A2(mult_x_1196_n2804), .B1(n23076), .B2(n24039), .Y(mult_x_1196_n2129) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2384 ( .A1(n24007), .A2(mult_x_1196_n3057), .B1(n24005), .B2(mult_x_1196_n3056), .Y(mult_x_1196_n2485) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U1806 ( .A1(mult_x_1196_n2775), .A2(n22412), .B1(mult_x_1196_n2774), .B2(n22481), .Y(mult_x_1196_n2211) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U1747 ( .A1(mult_x_1196_n2753), .A2(n24041), .B1(n24040), .B2(mult_x_1196_n2752), .Y(mult_x_1196_n2190) );
  NOR2x1_ASAP7_75t_SL mult_x_1196_U315 ( .A(mult_x_1196_n888), .B(
        mult_x_1196_n887), .Y(mult_x_1196_n354) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2380 ( .A1(mult_x_1196_n3053), .A2(n23637), .B1(n24005), .B2(mult_x_1196_n3052), .Y(mult_x_1196_n2481) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__44_ ( .D(
        n4221), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[43]) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__47_ ( .D(
        n4215), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[46]) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2817 ( .A1(mult_x_1196_n3268), .A2(n23981), .B1(n23980), .B2(mult_x_1196_n3267), .Y(mult_x_1196_n2692) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__45_ ( .D(
        n4219), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[44]) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2610 ( .A1(mult_x_1196_n3172), .A2(n23994), .B1(n23992), .B2(mult_x_1196_n3171), .Y(mult_x_1196_n2596) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2761 ( .A(n24045), .B(n23955), .Y(
        mult_x_1196_n3214) );
  NOR2x1_ASAP7_75t_SL mult_x_1196_U773 ( .A(mult_x_1196_n1949), .B(n22330), 
        .Y(mult_x_1196_n692) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U473 ( .A(mult_x_1196_n482), .B(
        mult_x_1196_n792), .Y(mult_x_1196_n242) );
  NAND2xp5_ASAP7_75t_SRAM mult_x_1196_U487 ( .A(n18422), .B(mult_x_1196_n793), 
        .Y(mult_x_1196_n243) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__46_ ( .D(
        n4217), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[45]) );
  OAI21xp5_ASAP7_75t_SL mult_x_1196_U468 ( .A1(mult_x_1196_n477), .A2(n22533), 
        .B(mult_x_1196_n478), .Y(mult_x_1196_n476) );
  XNOR2x1_ASAP7_75t_SL mult_x_1196_U2623 ( .A(n24049), .B(n23960), .Y(
        mult_x_1196_n3150) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2293 ( .A(n23965), .B(
        u0_0_leon3x0_p0_muli[13]), .Y(mult_x_1196_n3005) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2287 ( .A(n24068), .B(n23965), .Y(
        mult_x_1196_n2999) );
  NOR2x1_ASAP7_75t_SL mult_x_1196_U489 ( .A(n22353), .B(mult_x_1196_n1105), 
        .Y(mult_x_1196_n488) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2497 ( .A(n24065), .B(n22394), .Y(
        mult_x_1196_n3098) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__59_ ( .D(
        n4191), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[58]) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U368 ( .A(mult_x_1196_n947), .B(
        mult_x_1196_n933), .Y(mult_x_1196_n398) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U240 ( .A1(add_x_735_n212), .A2(
        add_x_735_n214), .B(add_x_735_n213), .Y(add_x_735_n211) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U226 ( .A1(add_x_735_n201), .A2(
        add_x_735_n214), .B(add_x_735_n202), .Y(add_x_735_n200) );
  NOR2x1_ASAP7_75t_SL mult_x_1196_U807 ( .A(n22334), .B(n23888), .Y(
        mult_x_1196_n714) );
  XNOR2x1_ASAP7_75t_SL mult_x_1196_U2618 ( .A(n23960), .B(n24044), .Y(
        mult_x_1196_n3145) );
  NOR2x1_ASAP7_75t_SL mult_x_1196_U513 ( .A(mult_x_1196_n1163), .B(
        mult_x_1196_n1162), .Y(mult_x_1196_n506) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U878 ( .A(mult_x_1196_n2091), .B(
        mult_x_1196_n2088), .Y(mult_x_1196_n761) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2414 ( .A(n24053), .B(n23396), .Y(
        mult_x_1196_n3052) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2689 ( .A(u0_0_leon3x0_p0_muli[37]), .B(
        n23958), .Y(mult_x_1196_n3179) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2690 ( .A(n24045), .B(n23957), .Y(
        mult_x_1196_n3180) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__48_ ( .D(
        n4213), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[47]) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__50_ ( .D(
        n4209), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[49]) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__54_ ( .D(
        n4201), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[53]) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77145 ( .A(uart1_uarto_SCALER__9_), .Y(
        n24600) );
  INVxp67_ASAP7_75t_SL sub_x_2325__cell_77154 ( .A(uart1_uarto_SCALER__0_), 
        .Y(n24609) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U315 ( .A(u0_0_leon3x0_p0_ici[39]), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__9_), .Y(DP_OP_1196_128_7433_n278) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U337 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__8_), .B(u0_0_leon3x0_p0_ici[38]), 
        .Y(DP_OP_1196_128_7433_n301) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U351 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__7_), .B(u0_0_leon3x0_p0_ici[37]), 
        .Y(DP_OP_1196_128_7433_n308) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U369 ( .A(u0_0_leon3x0_p0_ici[36]), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__6_), .Y(DP_OP_1196_128_7433_n327) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77148 ( .A(uart1_uarto_SCALER__6_), .Y(
        n24603) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77151 ( .A(uart1_uarto_SCALER__3_), .Y(
        n24606) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77149 ( .A(uart1_uarto_SCALER__5_), .Y(
        n24604) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77150 ( .A(uart1_uarto_SCALER__4_), .Y(
        n24605) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77152 ( .A(uart1_uarto_SCALER__2_), .Y(
        n24607) );
  INVxp67_ASAP7_75t_SL sub_x_2654__cell_77086 ( .A(timer0_r_SCALER__1_), .Y(
        n24627) );
  INVx1_ASAP7_75t_SL sub_x_2654__cell_77085 ( .A(timer0_r_SCALER__2_), .Y(
        n24626) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U283 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__11_), .B(u0_0_leon3x0_p0_ici[41]), 
        .Y(DP_OP_1196_128_7433_n252) );
  INVxp67_ASAP7_75t_SL sub_x_2654__cell_77082 ( .A(timer0_r_SCALER__5_), .Y(
        n24623) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U201 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__16_), .B(u0_0_leon3x0_p0_ici[46]), 
        .Y(DP_OP_1196_128_7433_n189) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U215 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__15_), .B(u0_0_leon3x0_p0_ici[45]), 
        .Y(DP_OP_1196_128_7433_n196) );
  INVx1_ASAP7_75t_SL sub_x_2654__cell_77087 ( .A(timer0_r_SCALER__0_), .Y(
        n24628) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U233 ( .A(u0_0_leon3x0_p0_ici[44]), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__14_), .Y(DP_OP_1196_128_7433_n215) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U133 ( .A(u0_0_leon3x0_p0_ici[50]), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), .Y(DP_OP_1196_128_7433_n129) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U167 ( .A(u0_0_leon3x0_p0_ici[48]), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_), .Y(DP_OP_1196_128_7433_n161) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U247 ( .A(u0_0_leon3x0_p0_ici[43]), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_), .Y(DP_OP_1196_128_7433_n222) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U181 ( .A(u0_0_leon3x0_p0_ici[47]), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_), .Y(DP_OP_1196_128_7433_n168) );
  INVx1_ASAP7_75t_SL sub_x_2654__cell_77081 ( .A(timer0_r_SCALER__6_), .Y(
        n24622) );
  INVx1_ASAP7_75t_SL sub_x_2654__cell_77084 ( .A(timer0_r_SCALER__3_), .Y(
        n24625) );
  INVxp33_ASAP7_75t_SL sub_x_2325__cell_77144 ( .A(uart1_uarto_SCALER__10_), 
        .Y(n24599) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U301 ( .A(u0_0_leon3x0_p0_ici[40]), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__10_), .Y(DP_OP_1196_128_7433_n271) );
  INVxp67_ASAP7_75t_SL sub_x_2654__cell_77083 ( .A(timer0_r_SCALER__4_), .Y(
        n24624) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U362 ( .A(n23950), .B(n23949), .Y(
        DP_OP_1196_128_7433_n318) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U334 ( .A(
        DP_OP_1196_128_7433_n301), .B(n23948), .Y(DP_OP_1196_128_7433_n30) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U230 ( .A(DP_OP_1196_128_7433_n215), .B(n23943), .Y(DP_OP_1196_128_7433_n24) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U198 ( .A(DP_OP_1196_128_7433_n189), .B(n23944), .Y(DP_OP_1196_128_7433_n22) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U266 ( .A(
        DP_OP_1196_128_7433_n245), .B(n23946), .Y(DP_OP_1196_128_7433_n26) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U164 ( .A(DP_OP_1196_128_7433_n161), .B(n23947), .Y(DP_OP_1196_128_7433_n20) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U298 ( .A(DP_OP_1196_128_7433_n271), .B(n23945), .Y(DP_OP_1196_128_7433_n28) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U294 ( .A(n23945), .B(
        DP_OP_1196_128_7433_n378), .Y(DP_OP_1196_128_7433_n266) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U295 ( .A1(n23945), .A2(
        DP_OP_1196_128_7433_n280), .B(DP_OP_1196_128_7433_n269), .Y(
        DP_OP_1196_128_7433_n267) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U262 ( .A(n23946), .B(
        DP_OP_1196_128_7433_n376), .Y(DP_OP_1196_128_7433_n240) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U148 ( .A(DP_OP_1196_128_7433_n148), .B(DP_OP_1196_128_7433_n368), .Y(DP_OP_1196_128_7433_n19) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U263 ( .A1(n23946), .A2(
        DP_OP_1196_128_7433_n254), .B(DP_OP_1196_128_7433_n243), .Y(
        DP_OP_1196_128_7433_n241) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U178 ( .A(DP_OP_1196_128_7433_n168), .B(DP_OP_1196_128_7433_n370), .Y(DP_OP_1196_128_7433_n21) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U112 ( .A(n23942), .B(
        DP_OP_1196_128_7433_n367), .Y(DP_OP_1196_128_7433_n115) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U212 ( .A(DP_OP_1196_128_7433_n196), .B(DP_OP_1196_128_7433_n372), .Y(DP_OP_1196_128_7433_n23) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U348 ( .A(
        DP_OP_1196_128_7433_n308), .B(DP_OP_1196_128_7433_n380), .Y(
        DP_OP_1196_128_7433_n31) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U280 ( .A(DP_OP_1196_128_7433_n252), .B(DP_OP_1196_128_7433_n376), .Y(DP_OP_1196_128_7433_n27) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U194 ( .A(n23944), .B(
        DP_OP_1196_128_7433_n372), .Y(DP_OP_1196_128_7433_n184) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U113 ( .A1(n23942), .A2(
        DP_OP_1196_128_7433_n131), .B(DP_OP_1196_128_7433_n120), .Y(
        DP_OP_1196_128_7433_n118) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U227 ( .A1(n23943), .A2(
        DP_OP_1196_128_7433_n224), .B(DP_OP_1196_128_7433_n213), .Y(
        DP_OP_1196_128_7433_n211) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U130 ( .A(DP_OP_1196_128_7433_n129), .B(DP_OP_1196_128_7433_n367), .Y(DP_OP_1196_128_7433_n18) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U160 ( .A(n23947), .B(
        DP_OP_1196_128_7433_n370), .Y(DP_OP_1196_128_7433_n154) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U363 ( .A1(n23949), .A2(
        DP_OP_1196_128_7433_n334), .B(DP_OP_1196_128_7433_n325), .Y(
        DP_OP_1196_128_7433_n319) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U330 ( .A(n23948), .B(
        DP_OP_1196_128_7433_n380), .Y(DP_OP_1196_128_7433_n296) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U226 ( .A(n23943), .B(
        DP_OP_1196_128_7433_n374), .Y(DP_OP_1196_128_7433_n210) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U27 ( .A(u0_0_leon3x0_p0_ici[58]), 
        .B(DP_OP_1196_128_7433_n480), .Y(DP_OP_1196_128_7433_n51) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U39 ( .A(u0_0_leon3x0_p0_ici[57]), 
        .B(DP_OP_1196_128_7433_n479), .Y(DP_OP_1196_128_7433_n60) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U53 ( .A(u0_0_leon3x0_p0_ici[56]), 
        .B(DP_OP_1196_128_7433_n478), .Y(DP_OP_1196_128_7433_n71) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U103 ( .A(u0_0_leon3x0_p0_ici[52]), .B(DP_OP_1196_128_7433_n474), .Y(DP_OP_1196_128_7433_n109) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U329 ( .A1(
        DP_OP_1196_128_7433_n319), .A2(DP_OP_1196_128_7433_n296), .B(
        DP_OP_1196_128_7433_n297), .Y(DP_OP_1196_128_7433_n291) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U147 ( .A1(
        DP_OP_1196_128_7433_n147), .A2(DP_OP_1196_128_7433_n157), .B(
        DP_OP_1196_128_7433_n148), .Y(DP_OP_1196_128_7433_n146) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U193 ( .A1(
        DP_OP_1196_128_7433_n211), .A2(DP_OP_1196_128_7433_n184), .B(
        DP_OP_1196_128_7433_n185), .Y(DP_OP_1196_128_7433_n183) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U343 ( .A1(
        DP_OP_1196_128_7433_n307), .A2(DP_OP_1196_128_7433_n319), .B(
        DP_OP_1196_128_7433_n308), .Y(DP_OP_1196_128_7433_n306) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U89 ( .A(u0_0_leon3x0_p0_ici[53]), 
        .B(DP_OP_1196_128_7433_n475), .Y(DP_OP_1196_128_7433_n98) );
  INVxp33_ASAP7_75t_SL sub_x_2655__cell_77050 ( .A(timer0_N63), .Y(n24390) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77064 ( .A(timer0_N77), .Y(n24403) );
  INVxp67_ASAP7_75t_SL sub_x_2655__cell_77054 ( .A(timer0_N67), .Y(n24393) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77061 ( .A(timer0_N74), .Y(n24400) );
  INVxp33_ASAP7_75t_SL sub_x_2655__cell_77048 ( .A(timer0_N61), .Y(n24388) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77053 ( .A(timer0_N66), .Y(n24392) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77063 ( .A(timer0_N76), .Y(n24402) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77060 ( .A(timer0_N73), .Y(n24399) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77057 ( .A(timer0_N70), .Y(n24396) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77055 ( .A(timer0_N68), .Y(n24394) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77049 ( .A(timer0_N62), .Y(n24389) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U65 ( .A(u0_0_leon3x0_p0_ici[55]), 
        .B(DP_OP_1196_128_7433_n477), .Y(DP_OP_1196_128_7433_n80) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77068 ( .A(timer0_N81), .Y(n24407) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77067 ( .A(timer0_N80), .Y(n24406) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U290 ( .A(
        DP_OP_1196_128_7433_n264), .B(DP_OP_1196_128_7433_n290), .Y(
        DP_OP_1196_128_7433_n262) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U49 ( .A1(DP_OP_1196_128_7433_n80), .A2(DP_OP_1196_128_7433_n70), .B(DP_OP_1196_128_7433_n71), .Y(
        DP_OP_1196_128_7433_n69) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U99 ( .A1(
        DP_OP_1196_128_7433_n118), .A2(DP_OP_1196_128_7433_n108), .B(
        DP_OP_1196_128_7433_n109), .Y(DP_OP_1196_128_7433_n107) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U145 ( .A1(
        DP_OP_1196_128_7433_n145), .A2(DP_OP_1196_128_7433_n183), .B(
        DP_OP_1196_128_7433_n146), .Y(DP_OP_1196_128_7433_n144) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U144 ( .A(DP_OP_1196_128_7433_n180), .B(DP_OP_1196_128_7433_n145), .Y(DP_OP_1196_128_7433_n143) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U259 ( .A1(
        DP_OP_1196_128_7433_n238), .A2(DP_OP_1196_128_7433_n291), .B(
        DP_OP_1196_128_7433_n239), .Y(DP_OP_1196_128_7433_n233) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U258 ( .A(DP_OP_1196_128_7433_n238), .B(DP_OP_1196_128_7433_n290), .Y(DP_OP_1196_128_7433_n232) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U47 ( .A1(DP_OP_1196_128_7433_n68), 
        .A2(DP_OP_1196_128_7433_n85), .B(DP_OP_1196_128_7433_n69), .Y(
        DP_OP_1196_128_7433_n67) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U307 ( .A(u0_0_leon3x0_p0_muli[41]), .B(
        u0_0_leon3x0_p0_divi[3]), .Y(add_x_735_n255) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U46 ( .A(DP_OP_1196_128_7433_n68), 
        .B(DP_OP_1196_128_7433_n84), .Y(DP_OP_1196_128_7433_n66) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U239 ( .A1(
        DP_OP_1196_128_7433_n221), .A2(DP_OP_1196_128_7433_n233), .B(
        DP_OP_1196_128_7433_n222), .Y(DP_OP_1196_128_7433_n220) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U2487 ( .A(n24055), .B(n23091), .Y(
        mult_x_1196_n3088) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U307 ( .A1(
        DP_OP_1196_128_7433_n277), .A2(DP_OP_1196_128_7433_n289), .B(
        DP_OP_1196_128_7433_n278), .Y(DP_OP_1196_128_7433_n276) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U143 ( .A1(
        DP_OP_1196_128_7433_n233), .A2(DP_OP_1196_128_7433_n143), .B(
        DP_OP_1196_128_7433_n144), .Y(DP_OP_1196_128_7433_n138) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U100 ( .A(DP_OP_1196_128_7433_n109), .B(DP_OP_1196_128_7433_n365), .Y(DP_OP_1196_128_7433_n16) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U275 ( .A1(
        DP_OP_1196_128_7433_n251), .A2(DP_OP_1196_128_7433_n263), .B(
        DP_OP_1196_128_7433_n252), .Y(DP_OP_1196_128_7433_n250) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U50 ( .A(DP_OP_1196_128_7433_n71), 
        .B(DP_OP_1196_128_7433_n361), .Y(DP_OP_1196_128_7433_n12) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U412 ( .A(u0_0_leon3x0_p0_ici[31]), 
        .B(DP_OP_1196_128_7433_n453), .Y(DP_OP_1196_128_7433_n355) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U405 ( .A(u0_0_leon3x0_p0_ici[32]), .B(DP_OP_1196_128_7433_n454), .Y(DP_OP_1196_128_7433_n351) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U391 ( .A(u0_0_leon3x0_p0_ici[34]), 
        .B(DP_OP_1196_128_7433_n456), .Y(DP_OP_1196_128_7433_n339) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U399 ( .A(u0_0_leon3x0_p0_ici[33]), 
        .B(DP_OP_1196_128_7433_n455), .Y(DP_OP_1196_128_7433_n348) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U222 ( .A(DP_OP_1196_128_7433_n208), .B(DP_OP_1196_128_7433_n234), .Y(DP_OP_1196_128_7433_n206) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U189 ( .A1(
        DP_OP_1196_128_7433_n235), .A2(DP_OP_1196_128_7433_n180), .B(
        DP_OP_1196_128_7433_n183), .Y(DP_OP_1196_128_7433_n179) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U188 ( .A(DP_OP_1196_128_7433_n180), .B(DP_OP_1196_128_7433_n234), .Y(DP_OP_1196_128_7433_n178) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U1931 ( .A(n24067), .B(n22395), .Y(
        mult_x_1196_n2828) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U59 ( .A1(DP_OP_1196_128_7433_n77), .A2(DP_OP_1196_128_7433_n87), .B(DP_OP_1196_128_7433_n80), .Y(
        DP_OP_1196_128_7433_n76) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U395 ( .A1(
        DP_OP_1196_128_7433_n351), .A2(DP_OP_1196_128_7433_n347), .B(
        DP_OP_1196_128_7433_n348), .Y(DP_OP_1196_128_7433_n346) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U97 ( .A1(
        DP_OP_1196_128_7433_n106), .A2(DP_OP_1196_128_7433_n138), .B(
        DP_OP_1196_128_7433_n107), .Y(DP_OP_1196_128_7433_n105) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U96 ( .A(DP_OP_1196_128_7433_n106), 
        .B(DP_OP_1196_128_7433_n137), .Y(DP_OP_1196_128_7433_n104) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U95 ( .A1(DP_OP_1196_128_7433_n104), .A2(DP_OP_1196_128_7433_n339), .B(DP_OP_1196_128_7433_n105), .Y(
        DP_OP_1196_128_7433_n7) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U272 ( .A(
        DP_OP_1196_128_7433_n249), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n247) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U157 ( .A1(
        DP_OP_1196_128_7433_n154), .A2(DP_OP_1196_128_7433_n179), .B(
        DP_OP_1196_128_7433_n157), .Y(DP_OP_1196_128_7433_n153) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U125 ( .A1(
        DP_OP_1196_128_7433_n128), .A2(DP_OP_1196_128_7433_n140), .B(
        DP_OP_1196_128_7433_n129), .Y(DP_OP_1196_128_7433_n127) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U236 ( .A(
        DP_OP_1196_128_7433_n219), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n217) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U207 ( .A1(
        DP_OP_1196_128_7433_n195), .A2(DP_OP_1196_128_7433_n207), .B(
        DP_OP_1196_128_7433_n196), .Y(DP_OP_1196_128_7433_n194) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U173 ( .A1(
        DP_OP_1196_128_7433_n167), .A2(DP_OP_1196_128_7433_n179), .B(
        DP_OP_1196_128_7433_n168), .Y(DP_OP_1196_128_7433_n166) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U137 ( .A1(DP_OP_1196_128_7433_n4), .A2(DP_OP_1196_128_7433_n137), .B(DP_OP_1196_128_7433_n138), .Y(
        DP_OP_1196_128_7433_n136) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U136 ( .A(
        DP_OP_1196_128_7433_n137), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n135) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U109 ( .A1(
        DP_OP_1196_128_7433_n115), .A2(DP_OP_1196_128_7433_n140), .B(
        DP_OP_1196_128_7433_n118), .Y(DP_OP_1196_128_7433_n114) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U304 ( .A(
        DP_OP_1196_128_7433_n275), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n273) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U286 ( .A(
        DP_OP_1196_128_7433_n260), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n258) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U373 ( .A1(DP_OP_1196_128_7433_n4), .A2(n23950), .B(DP_OP_1196_128_7433_n334), .Y(DP_OP_1196_128_7433_n330) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U402 ( .A(
        DP_OP_1196_128_7433_n351), .B(DP_OP_1196_128_7433_n385), .Y(
        DP_OP_1196_128_7433_n36) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U409 ( .A(
        DP_OP_1196_128_7433_n355), .B(DP_OP_1196_128_7433_n386), .Y(
        DP_OP_1196_128_7433_n37) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U318 ( .A(
        DP_OP_1196_128_7433_n290), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n284) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U388 ( .A(
        DP_OP_1196_128_7433_n339), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n34) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U319 ( .A1(DP_OP_1196_128_7433_n4), .A2(DP_OP_1196_128_7433_n290), .B(DP_OP_1196_128_7433_n291), .Y(
        DP_OP_1196_128_7433_n285) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U132 ( .A(n23969), .B(
        u0_0_leon3x0_p0_divi[20]), .Y(add_x_735_n131) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U372 ( .A(n23950), .B(
        DP_OP_1196_128_7433_n6), .Y(DP_OP_1196_128_7433_n329) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U354 ( .A(
        DP_OP_1196_128_7433_n316), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n314) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U34 ( .A(n22968), .B(
        u0_0_leon3x0_p0_divi[28]), .Y(add_x_735_n57) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U355 ( .A1(DP_OP_1196_128_7433_n4), .A2(DP_OP_1196_128_7433_n316), .B(DP_OP_1196_128_7433_n317), .Y(
        DP_OP_1196_128_7433_n315) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U277 ( .A(add_x_735_A_9_), .B(
        u0_0_leon3x0_p0_divi[7]), .Y(add_x_735_n237) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U341 ( .A1(DP_OP_1196_128_7433_n4), .A2(DP_OP_1196_128_7433_n305), .B(DP_OP_1196_128_7433_n306), .Y(
        DP_OP_1196_128_7433_n304) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U340 ( .A(
        DP_OP_1196_128_7433_n305), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n303) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U238 ( .A(u0_0_leon3x0_p0_muli[45]), .B(
        u0_0_leon3x0_p0_divi[11]), .Y(add_x_735_n210) );
  OAI21xp33_ASAP7_75t_SL add_x_735_U68 ( .A1(add_x_735_n95), .A2(add_x_735_n85), .B(add_x_735_n86), .Y(add_x_735_n84) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U122 ( .A(
        DP_OP_1196_128_7433_n126), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n124) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U82 ( .A(DP_OP_1196_128_7433_n95), 
        .B(DP_OP_1196_128_7433_n8), .Y(DP_OP_1196_128_7433_n93) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U83 ( .A1(DP_OP_1196_128_7433_n7), 
        .A2(DP_OP_1196_128_7433_n95), .B(DP_OP_1196_128_7433_n96), .Y(
        DP_OP_1196_128_7433_n94) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U56 ( .A(DP_OP_1196_128_7433_n75), 
        .B(DP_OP_1196_128_7433_n8), .Y(DP_OP_1196_128_7433_n73) );
  AOI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U57 ( .A1(DP_OP_1196_128_7433_n7), 
        .A2(DP_OP_1196_128_7433_n75), .B(DP_OP_1196_128_7433_n76), .Y(
        DP_OP_1196_128_7433_n74) );
  OAI21xp33_ASAP7_75t_SL add_x_735_U118 ( .A1(add_x_735_n131), .A2(
        add_x_735_n123), .B(add_x_735_n124), .Y(add_x_735_n122) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U154 ( .A(
        DP_OP_1196_128_7433_n152), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n150) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U170 ( .A(
        DP_OP_1196_128_7433_n165), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n163) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U184 ( .A(
        DP_OP_1196_128_7433_n176), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n174) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U204 ( .A(
        DP_OP_1196_128_7433_n193), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n191) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U218 ( .A(
        DP_OP_1196_128_7433_n204), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n202) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U106 ( .A(
        DP_OP_1196_128_7433_n113), .B(DP_OP_1196_128_7433_n6), .Y(
        DP_OP_1196_128_7433_n111) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U353 ( .A1(
        DP_OP_1196_128_7433_n314), .A2(n23941), .B(DP_OP_1196_128_7433_n315), 
        .Y(DP_OP_1196_128_7433_n313) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U187 ( .A(add_x_735_n174), .B(add_x_735_n288), .Y(add_x_735_n19) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U252 ( .A(add_x_735_n221), .B(
        add_x_735_n294), .Y(add_x_735_n25) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U339 ( .A1(
        DP_OP_1196_128_7433_n303), .A2(n23941), .B(DP_OP_1196_128_7433_n304), 
        .Y(DP_OP_1196_128_7433_n302) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U317 ( .A1(
        DP_OP_1196_128_7433_n284), .A2(n23941), .B(DP_OP_1196_128_7433_n285), 
        .Y(DP_OP_1196_128_7433_n283) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U271 ( .A1(
        DP_OP_1196_128_7433_n247), .A2(n23941), .B(DP_OP_1196_128_7433_n248), 
        .Y(DP_OP_1196_128_7433_n246) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U221 ( .A(add_x_735_n199), .B(
        add_x_735_n291), .Y(add_x_735_n22) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U153 ( .A1(
        DP_OP_1196_128_7433_n150), .A2(n23941), .B(DP_OP_1196_128_7433_n151), 
        .Y(DP_OP_1196_128_7433_n149) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U121 ( .A1(
        DP_OP_1196_128_7433_n124), .A2(n23941), .B(DP_OP_1196_128_7433_n125), 
        .Y(DP_OP_1196_128_7433_n123) );
  AOI21xp33_ASAP7_75t_SL add_x_735_U218 ( .A1(add_x_735_n204), .A2(
        add_x_735_n291), .B(add_x_735_n197), .Y(add_x_735_n195) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U217 ( .A(add_x_735_n291), .B(
        add_x_735_n203), .Y(add_x_735_n194) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U81 ( .A1(DP_OP_1196_128_7433_n93), 
        .A2(n23941), .B(DP_OP_1196_128_7433_n94), .Y(DP_OP_1196_128_7433_n92)
         );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U55 ( .A1(DP_OP_1196_128_7433_n73), 
        .A2(n23941), .B(DP_OP_1196_128_7433_n74), .Y(DP_OP_1196_128_7433_n72)
         );
  NAND2xp33_ASAP7_75t_SL add_x_735_U149 ( .A(n18889), .B(add_x_735_n285), .Y(
        add_x_735_n16) );
  AOI21xp33_ASAP7_75t_SL add_x_735_U66 ( .A1(add_x_735_n83), .A2(
        add_x_735_n100), .B(add_x_735_n84), .Y(add_x_735_n82) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U65 ( .A(add_x_735_n99), .B(add_x_735_n83), 
        .Y(add_x_735_n81) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U5 ( .A(add_x_735_n37), .B(n24313), .Y(
        add_x_735_n4) );
  AOI21xp33_ASAP7_75t_SL add_x_735_U126 ( .A1(add_x_735_n136), .A2(
        add_x_735_n283), .B(add_x_735_n129), .Y(add_x_735_n127) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U125 ( .A(add_x_735_n283), .B(
        add_x_735_n135), .Y(add_x_735_n126) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U119 ( .A(add_x_735_n124), .B(add_x_735_n282), .Y(add_x_735_n13) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U105 ( .A(add_x_735_n113), .B(
        add_x_735_n281), .Y(add_x_735_n12) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U95 ( .A(add_x_735_n106), .B(add_x_735_n280), 
        .Y(add_x_735_n11) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U143 ( .A(add_x_735_n142), .B(add_x_735_n284), .Y(add_x_735_n15) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U31 ( .A(add_x_735_n57), .B(add_x_735_n275), 
        .Y(add_x_735_n6) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U69 ( .A(add_x_735_n86), .B(add_x_735_n278), 
        .Y(add_x_735_n9) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U129 ( .A(add_x_735_n131), .B(add_x_735_n283), .Y(add_x_735_n14) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U235 ( .A(add_x_735_n210), .B(add_x_735_n292), .Y(add_x_735_n23) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U161 ( .A(add_x_735_n154), .B(
        add_x_735_n286), .Y(add_x_735_n17) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U183 ( .A1(
        DP_OP_1196_128_7433_n174), .A2(n23941), .B(DP_OP_1196_128_7433_n175), 
        .Y(DP_OP_1196_128_7433_n173) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U169 ( .A1(
        DP_OP_1196_128_7433_n163), .A2(n23941), .B(DP_OP_1196_128_7433_n164), 
        .Y(DP_OP_1196_128_7433_n162) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U135 ( .A1(
        DP_OP_1196_128_7433_n135), .A2(n23941), .B(DP_OP_1196_128_7433_n136), 
        .Y(DP_OP_1196_128_7433_n134) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U105 ( .A1(
        DP_OP_1196_128_7433_n111), .A2(n23941), .B(DP_OP_1196_128_7433_n112), 
        .Y(DP_OP_1196_128_7433_n110) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U291 ( .A(add_x_735_n248), .B(add_x_735_n298), .Y(add_x_735_n29) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U371 ( .A1(
        DP_OP_1196_128_7433_n329), .A2(n23941), .B(DP_OP_1196_128_7433_n330), 
        .Y(DP_OP_1196_128_7433_n328) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U274 ( .A(add_x_735_n237), .B(add_x_735_n296), .Y(add_x_735_n27) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U203 ( .A1(
        DP_OP_1196_128_7433_n191), .A2(n23941), .B(DP_OP_1196_128_7433_n192), 
        .Y(DP_OP_1196_128_7433_n190) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U303 ( .A1(
        DP_OP_1196_128_7433_n273), .A2(n23941), .B(DP_OP_1196_128_7433_n274), 
        .Y(DP_OP_1196_128_7433_n272) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U285 ( .A1(
        DP_OP_1196_128_7433_n258), .A2(n23941), .B(DP_OP_1196_128_7433_n259), 
        .Y(DP_OP_1196_128_7433_n257) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U235 ( .A1(
        DP_OP_1196_128_7433_n217), .A2(n23941), .B(DP_OP_1196_128_7433_n218), 
        .Y(DP_OP_1196_128_7433_n216) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U217 ( .A1(
        DP_OP_1196_128_7433_n202), .A2(n23941), .B(DP_OP_1196_128_7433_n203), 
        .Y(DP_OP_1196_128_7433_n201) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U241 ( .A(add_x_735_n213), .B(add_x_735_n293), .Y(add_x_735_n24) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U248 ( .A(add_x_735_n218), .B(add_x_735_n230), .Y(add_x_735_n216) );
  OAI21xp33_ASAP7_75t_SL add_x_735_U18 ( .A1(add_x_735_n57), .A2(add_x_735_n47), .B(add_x_735_n48), .Y(add_x_735_n46) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U211 ( .A(add_x_735_n192), .B(add_x_735_n290), .Y(add_x_735_n21) );
  OAI21xp33_ASAP7_75t_SL add_x_735_U259 ( .A1(add_x_735_n225), .A2(n18896), 
        .B(add_x_735_n228), .Y(add_x_735_n224) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U101 ( .A(add_x_735_n281), .B(
        add_x_735_n117), .Y(add_x_735_n108) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U1590 ( .A(mult_x_1196_n2689), .B(
        mult_x_1196_n2529), .Y(mult_x_1196_n1984) );
  AOI21xp33_ASAP7_75t_SL add_x_735_U52 ( .A1(add_x_735_n2), .A2(add_x_735_n72), 
        .B(add_x_735_n73), .Y(add_x_735_n71) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U55 ( .A(add_x_735_n75), .B(add_x_735_n72), 
        .Y(add_x_735_n8) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U19 ( .A(add_x_735_n48), .B(add_x_735_n274), 
        .Y(add_x_735_n5) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U371 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[0]), .B(u0_0_leon3x0_p0_div0_vaddsub), 
        .Y(DP_OP_5187J1_124_3275_n305) );
  NAND2xp33_ASAP7_75t_SL add_x_746_U44 ( .A(u0_0_leon3x0_p0_iu_fe_pc_25_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_24_), .Y(add_x_746_n37) );
  NAND2xp33_ASAP7_75t_SL add_x_746_U16 ( .A(u0_0_leon3x0_p0_iu_fe_pc_29_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_28_), .Y(add_x_746_n13) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U11 ( .A(n24315), .B(add_x_735_n3), .Y(
        add_x_735_n39) );
  OAI21xp33_ASAP7_75t_SL add_x_735_U28 ( .A1(add_x_735_n54), .A2(add_x_735_n64), .B(add_x_735_n57), .Y(add_x_735_n53) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U167 ( .A(add_x_735_n158), .B(
        add_x_735_n185), .Y(add_x_735_n156) );
  AOI21xp5_ASAP7_75t_SL add_x_735_U168 ( .A1(add_x_735_n186), .A2(
        add_x_735_n158), .B(add_x_735_n159), .Y(add_x_735_n157) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U162 ( .A(u0_0_leon3x0_p0_iu_fe_pc_7_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_6_), .Y(add_x_746_n135) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U139 ( .A(u0_0_leon3x0_p0_iu_fe_pc_11_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_10_), .Y(add_x_746_n116) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U58 ( .A(u0_0_leon3x0_p0_iu_fe_pc_22_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_23_), .Y(add_x_746_n47) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U111 ( .A(u0_0_leon3x0_p0_iu_fe_pc_14_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_15_), .Y(add_x_746_n92) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U86 ( .A(u0_0_leon3x0_p0_iu_fe_pc_19_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_18_), .Y(add_x_746_n71) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U173 ( .A(u0_0_leon3x0_p0_iu_fe_pc_5_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_4_), .Y(add_x_746_n146) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U150 ( .A(u0_0_leon3x0_p0_iu_fe_pc_8_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_9_), .Y(add_x_746_n127) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U228 ( .A(mult_x_1196_n839), .B(
        mult_x_1196_n837), .Y(mult_x_1196_n288) );
  FAx1_ASAP7_75t_SL mult_x_1196_U910 ( .A(mult_x_1196_n854), .B(
        mult_x_1196_n864), .CI(mult_x_1196_n862), .CON(mult_x_1196_n851), .SN(
        mult_x_1196_n852) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U271 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[11]), .B(u0_0_leon3x0_p0_div0_b[11]), .Y(
        DP_OP_5187J1_124_3275_n238) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U165 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[20]), .B(u0_0_leon3x0_p0_div0_b[20]), .Y(
        DP_OP_5187J1_124_3275_n159) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U247 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[13]), .B(u0_0_leon3x0_p0_div0_b[13]), .Y(
        DP_OP_5187J1_124_3275_n220) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U79 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[27]), .B(u0_0_leon3x0_p0_div0_b[27]), .Y(
        DP_OP_5187J1_124_3275_n94) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U221 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[15]), .B(u0_0_leon3x0_p0_div0_b[15]), .Y(
        DP_OP_5187J1_124_3275_n200) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U91 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[26]), .B(u0_0_leon3x0_p0_div0_b[26]), .Y(
        DP_OP_5187J1_124_3275_n103) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U334 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[5]), .B(u0_0_leon3x0_p0_div0_b[5]), .Y(
        DP_OP_5187J1_124_3275_n283) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U39 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[30]), .B(u0_0_leon3x0_p0_div0_b[30]), .Y(
        DP_OP_5187J1_124_3275_n63) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U351 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[3]), .B(u0_0_leon3x0_p0_div0_b[3]), .Y(
        DP_OP_5187J1_124_3275_n294) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U357 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[2]), .B(u0_0_leon3x0_p0_div0_b[2]), .Y(
        DP_OP_5187J1_124_3275_n297) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U364 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[1]), .B(u0_0_leon3x0_p0_div0_b[1]), .Y(
        DP_OP_5187J1_124_3275_n301) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U53 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[29]), .B(u0_0_leon3x0_p0_div0_b[29]), .Y(
        DP_OP_5187J1_124_3275_n74) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U225 ( .A(mult_x_1196_n288), .B(n24250), .Y(
        mult_x_1196_n224) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U25 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[31]), .B(u0_0_leon3x0_p0_div0_b[31]), .Y(
        DP_OP_5187J1_124_3275_n52) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U65 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[28]), .B(u0_0_leon3x0_p0_div0_b[28]), .Y(
        DP_OP_5187J1_124_3275_n83) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U141 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[22]), .B(u0_0_leon3x0_p0_div0_b[22]), .Y(
        DP_OP_5187J1_124_3275_n141) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U129 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[23]), .B(u0_0_leon3x0_p0_div0_b[23]), .Y(
        DP_OP_5187J1_124_3275_n132) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U155 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[21]), .B(u0_0_leon3x0_p0_div0_b[21]), .Y(
        DP_OP_5187J1_124_3275_n152) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U105 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[25]), .B(u0_0_leon3x0_p0_div0_b[25]), .Y(
        DP_OP_5187J1_124_3275_n114) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U115 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[24]), .B(u0_0_leon3x0_p0_div0_b[24]), .Y(
        DP_OP_5187J1_124_3275_n121) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U312 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[7]), .B(u0_0_leon3x0_p0_div0_b[7]), .Y(
        DP_OP_5187J1_124_3275_n267) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U49 ( .A1(
        DP_OP_5187J1_124_3275_n83), .A2(DP_OP_5187J1_124_3275_n73), .B(
        DP_OP_5187J1_124_3275_n74), .Y(DP_OP_5187J1_124_3275_n72) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U21 ( .A1(
        DP_OP_5187J1_124_3275_n63), .A2(DP_OP_5187J1_124_3275_n51), .B(
        DP_OP_5187J1_124_3275_n52), .Y(DP_OP_5187J1_124_3275_n50) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U75 ( .A1(
        DP_OP_5187J1_124_3275_n103), .A2(DP_OP_5187J1_124_3275_n93), .B(
        DP_OP_5187J1_124_3275_n94), .Y(DP_OP_5187J1_124_3275_n92) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U308 ( .A1(
        DP_OP_5187J1_124_3275_n274), .A2(DP_OP_5187J1_124_3275_n266), .B(
        DP_OP_5187J1_124_3275_n267), .Y(DP_OP_5187J1_124_3275_n265) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U125 ( .A1(
        DP_OP_5187J1_124_3275_n141), .A2(DP_OP_5187J1_124_3275_n131), .B(
        DP_OP_5187J1_124_3275_n132), .Y(DP_OP_5187J1_124_3275_n130) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U217 ( .A1(
        DP_OP_5187J1_124_3275_n209), .A2(DP_OP_5187J1_124_3275_n199), .B(
        DP_OP_5187J1_124_3275_n200), .Y(DP_OP_5187J1_124_3275_n198) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U175 ( .A1(
        DP_OP_5187J1_124_3275_n177), .A2(DP_OP_5187J1_124_3275_n169), .B(
        DP_OP_5187J1_124_3275_n170), .Y(DP_OP_5187J1_124_3275_n168) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U8 ( .A(
        DP_OP_5187J1_124_3275_n41), .B(n24316), .Y(DP_OP_5187J1_124_3275_n7)
         );
  OAI21xp5_ASAP7_75t_SL add_x_735_U216 ( .A1(add_x_735_n194), .A2(
        add_x_735_n214), .B(add_x_735_n195), .Y(add_x_735_n193) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U182 ( .A(
        DP_OP_5187J1_124_3275_n321), .B(DP_OP_5187J1_124_3275_n181), .Y(
        DP_OP_5187J1_124_3275_n172) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U102 ( .A(
        DP_OP_5187J1_124_3275_n114), .B(DP_OP_5187J1_124_3275_n314), .Y(
        DP_OP_5187J1_124_3275_n14) );
  AOI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U183 ( .A1(
        DP_OP_5187J1_124_3275_n182), .A2(DP_OP_5187J1_124_3275_n321), .B(
        DP_OP_5187J1_124_3275_n175), .Y(DP_OP_5187J1_124_3275_n173) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U62 ( .A(add_x_746_n53), .B(n18880), .Y(
        add_x_746_n52) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U48 ( .A(add_x_746_n41), .B(n18880), .Y(
        add_x_746_n40) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U135 ( .A(add_x_746_n115), .B(add_x_746_n124), .Y(add_x_746_n114) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U206 ( .A(
        DP_OP_5187J1_124_3275_n191), .B(DP_OP_5187J1_124_3275_n323), .Y(
        DP_OP_5187J1_124_3275_n23) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U305 ( .A(
        DP_OP_5187J1_124_3275_n264), .B(DP_OP_5187J1_124_3275_n276), .Y(
        DP_OP_5187J1_124_3275_n262) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U12 ( .A(n18880), .B(add_x_746_n10), .Y(
        add_x_746_n9) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U244 ( .A(
        DP_OP_5187J1_124_3275_n220), .B(DP_OP_5187J1_124_3275_n326), .Y(
        DP_OP_5187J1_124_3275_n26) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U107 ( .A(add_x_746_n124), .B(add_x_746_n91), 
        .Y(add_x_746_n90) );
  NAND2xp33_ASAP7_75t_SL mult_x_1196_U869 ( .A(mult_x_1196_n758), .B(n24261), 
        .Y(mult_x_1196_n282) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U331 ( .A(
        DP_OP_5187J1_124_3275_n283), .B(DP_OP_5187J1_124_3275_n334), .Y(
        DP_OP_5187J1_124_3275_n34) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U172 ( .A(
        DP_OP_5187J1_124_3275_n167), .B(DP_OP_5187J1_124_3275_n181), .Y(
        DP_OP_5187J1_124_3275_n161) );
  AOI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U215 ( .A1(
        DP_OP_5187J1_124_3275_n197), .A2(DP_OP_5187J1_124_3275_n214), .B(
        DP_OP_5187J1_124_3275_n198), .Y(DP_OP_5187J1_124_3275_n196) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U348 ( .A(
        DP_OP_5187J1_124_3275_n294), .B(DP_OP_5187J1_124_3275_n336), .Y(
        DP_OP_5187J1_124_3275_n36) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U214 ( .A(
        DP_OP_5187J1_124_3275_n197), .B(DP_OP_5187J1_124_3275_n213), .Y(
        DP_OP_5187J1_124_3275_n195) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U129 ( .A(add_x_746_n110), .B(add_x_746_n124), .Y(add_x_746_n109) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U88 ( .A(
        DP_OP_5187J1_124_3275_n103), .B(DP_OP_5187J1_124_3275_n313), .Y(
        DP_OP_5187J1_124_3275_n13) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U101 ( .A(add_x_746_n124), .B(add_x_746_n86), 
        .Y(add_x_746_n85) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U82 ( .A(add_x_746_n70), .B(n18880), .Y(
        add_x_746_n69) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U26 ( .A(n18880), .B(add_x_746_n22), .Y(
        add_x_746_n21) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U235 ( .A(mult_x_1196_n295), .B(
        mult_x_1196_n775), .Y(mult_x_1196_n225) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U309 ( .A(
        DP_OP_5187J1_124_3275_n267), .B(DP_OP_5187J1_124_3275_n332), .Y(
        DP_OP_5187J1_124_3275_n32) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U54 ( .A(add_x_746_n46), .B(n18880), .Y(
        add_x_746_n45) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U22 ( .A(
        DP_OP_5187J1_124_3275_n52), .B(DP_OP_5187J1_124_3275_n308), .Y(
        DP_OP_5187J1_124_3275_n8) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U32 ( .A(
        DP_OP_5187J1_124_3275_n60), .B(DP_OP_5187J1_124_3275_n71), .Y(
        DP_OP_5187J1_124_3275_n58) );
  AOI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U33 ( .A1(
        DP_OP_5187J1_124_3275_n72), .A2(DP_OP_5187J1_124_3275_n60), .B(
        DP_OP_5187J1_124_3275_n61), .Y(DP_OP_5187J1_124_3275_n59) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U18 ( .A(
        DP_OP_5187J1_124_3275_n49), .B(DP_OP_5187J1_124_3275_n71), .Y(
        DP_OP_5187J1_124_3275_n47) );
  NAND2xp33_ASAP7_75t_SL add_x_746_U143 ( .A(u0_0_leon3x0_p0_iu_fe_pc_10_), 
        .B(add_x_746_n124), .Y(add_x_746_n121) );
  NAND2xp33_ASAP7_75t_SL add_x_746_U121 ( .A(add_x_746_n103), .B(
        add_x_746_n124), .Y(add_x_746_n102) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U62 ( .A(
        DP_OP_5187J1_124_3275_n83), .B(DP_OP_5187J1_124_3275_n311), .Y(
        DP_OP_5187J1_124_3275_n11) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U115 ( .A(add_x_746_n124), .B(add_x_746_n98), 
        .Y(add_x_746_n97) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U31 ( .A1(
        DP_OP_5187J1_124_3275_n5), .A2(DP_OP_5187J1_124_3275_n58), .B(
        DP_OP_5187J1_124_3275_n59), .Y(DP_OP_5187J1_124_3275_n57) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U59 ( .A1(
        DP_OP_5187J1_124_3275_n80), .A2(DP_OP_5187J1_124_3275_n5), .B(
        DP_OP_5187J1_124_3275_n83), .Y(DP_OP_5187J1_124_3275_n79) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U135 ( .A1(
        DP_OP_5187J1_124_3275_n138), .A2(DP_OP_5187J1_124_3275_n148), .B(
        DP_OP_5187J1_124_3275_n141), .Y(DP_OP_5187J1_124_3275_n137) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U213 ( .A1(
        DP_OP_5187J1_124_3275_n230), .A2(DP_OP_5187J1_124_3275_n195), .B(
        DP_OP_5187J1_124_3275_n196), .Y(DP_OP_5187J1_124_3275_n194) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U85 ( .A1(
        DP_OP_5187J1_124_3275_n100), .A2(DP_OP_5187J1_124_3275_n110), .B(
        DP_OP_5187J1_124_3275_n103), .Y(DP_OP_5187J1_124_3275_n99) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U45 ( .A1(
        DP_OP_5187J1_124_3275_n69), .A2(DP_OP_5187J1_124_3275_n5), .B(
        DP_OP_5187J1_124_3275_n70), .Y(DP_OP_5187J1_124_3275_n68) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U316 ( .A1(
        DP_OP_5187J1_124_3275_n271), .A2(DP_OP_5187J1_124_3275_n279), .B(
        DP_OP_5187J1_124_3275_n274), .Y(DP_OP_5187J1_124_3275_n270) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U29 ( .A1(
        DP_OP_5187J1_124_3275_n56), .A2(DP_OP_5187J1_124_3275_n3), .B(
        DP_OP_5187J1_124_3275_n57), .Y(DP_OP_5187J1_124_3275_n55) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U94 ( .A(
        DP_OP_5187J1_124_3275_n107), .B(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n105) );
  AOI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U95 ( .A1(
        DP_OP_5187J1_124_3275_n3), .A2(DP_OP_5187J1_124_3275_n107), .B(
        DP_OP_5187J1_124_3275_n108), .Y(DP_OP_5187J1_124_3275_n106) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U56 ( .A(
        DP_OP_5187J1_124_3275_n78), .B(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n76) );
  AOI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U251 ( .A1(
        DP_OP_5187J1_124_3275_n232), .A2(DP_OP_5187J1_124_3275_n327), .B(
        DP_OP_5187J1_124_3275_n225), .Y(DP_OP_5187J1_124_3275_n223) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U28 ( .A(
        DP_OP_5187J1_124_3275_n56), .B(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n54) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U250 ( .A(
        DP_OP_5187J1_124_3275_n327), .B(DP_OP_5187J1_124_3275_n231), .Y(
        DP_OP_5187J1_124_3275_n222) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U144 ( .A(
        DP_OP_5187J1_124_3275_n145), .B(DP_OP_5187J1_124_3275_n163), .Y(
        DP_OP_5187J1_124_3275_n143) );
  AOI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U145 ( .A1(
        DP_OP_5187J1_124_3275_n164), .A2(DP_OP_5187J1_124_3275_n145), .B(
        DP_OP_5187J1_124_3275_n146), .Y(DP_OP_5187J1_124_3275_n144) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U108 ( .A(
        DP_OP_5187J1_124_3275_n315), .B(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n116) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U15 ( .A1(
        DP_OP_5187J1_124_3275_n45), .A2(DP_OP_5187J1_124_3275_n3), .B(
        DP_OP_5187J1_124_3275_n46), .Y(DP_OP_5187J1_124_3275_n44) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U69 ( .A1(
        DP_OP_5187J1_124_3275_n3), .A2(DP_OP_5187J1_124_3275_n87), .B(
        DP_OP_5187J1_124_3275_n88), .Y(DP_OP_5187J1_124_3275_n86) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U68 ( .A(
        DP_OP_5187J1_124_3275_n87), .B(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n85) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U42 ( .A(
        DP_OP_5187J1_124_3275_n67), .B(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n65) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U158 ( .A(
        DP_OP_5187J1_124_3275_n319), .B(DP_OP_5187J1_124_3275_n163), .Y(
        DP_OP_5187J1_124_3275_n154) );
  NAND2xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U82 ( .A(
        DP_OP_5187J1_124_3275_n98), .B(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n96) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U249 ( .A1(n23887), .A2(
        DP_OP_5187J1_124_3275_n222), .B(DP_OP_5187J1_124_3275_n223), .Y(
        DP_OP_5187J1_124_3275_n221) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U259 ( .A1(
        DP_OP_5187J1_124_3275_n229), .A2(n23887), .B(
        DP_OP_5187J1_124_3275_n230), .Y(DP_OP_5187J1_124_3275_n228) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U314 ( .A1(
        DP_OP_5187J1_124_3275_n269), .A2(DP_OP_5187J1_124_3275_n289), .B(
        DP_OP_5187J1_124_3275_n270), .Y(DP_OP_5187J1_124_3275_n268) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U117 ( .A1(
        DP_OP_5187J1_124_3275_n123), .A2(n22225), .B(
        DP_OP_5187J1_124_3275_n124), .Y(DP_OP_5187J1_124_3275_n122) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U181 ( .A1(
        DP_OP_5187J1_124_3275_n172), .A2(n22225), .B(
        DP_OP_5187J1_124_3275_n173), .Y(DP_OP_5187J1_124_3275_n171) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U143 ( .A1(
        DP_OP_5187J1_124_3275_n143), .A2(n22225), .B(
        DP_OP_5187J1_124_3275_n144), .Y(DP_OP_5187J1_124_3275_n142) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U167 ( .A1(
        DP_OP_5187J1_124_3275_n161), .A2(n22225), .B(
        DP_OP_5187J1_124_3275_n162), .Y(DP_OP_5187J1_124_3275_n160) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U107 ( .A1(n22225), .A2(
        DP_OP_5187J1_124_3275_n116), .B(DP_OP_5187J1_124_3275_n117), .Y(
        DP_OP_5187J1_124_3275_n115) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U131 ( .A1(
        DP_OP_5187J1_124_3275_n134), .A2(n22225), .B(
        DP_OP_5187J1_124_3275_n135), .Y(DP_OP_5187J1_124_3275_n133) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U93 ( .A1(n22225), .A2(
        DP_OP_5187J1_124_3275_n105), .B(DP_OP_5187J1_124_3275_n106), .Y(
        DP_OP_5187J1_124_3275_n104) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U27 ( .A1(n22225), .A2(
        DP_OP_5187J1_124_3275_n54), .B(DP_OP_5187J1_124_3275_n55), .Y(
        DP_OP_5187J1_124_3275_n53) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U55 ( .A1(n22225), .A2(
        DP_OP_5187J1_124_3275_n76), .B(DP_OP_5187J1_124_3275_n77), .Y(
        DP_OP_5187J1_124_3275_n75) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U41 ( .A1(n22225), .A2(
        DP_OP_5187J1_124_3275_n65), .B(DP_OP_5187J1_124_3275_n66), .Y(
        DP_OP_5187J1_124_3275_n64) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U157 ( .A1(
        DP_OP_5187J1_124_3275_n154), .A2(n22225), .B(
        DP_OP_5187J1_124_3275_n155), .Y(DP_OP_5187J1_124_3275_n153) );
  NAND2xp33_ASAP7_75t_SL mult_x_1196_U799 ( .A(mult_x_1196_n712), .B(
        mult_x_1196_n824), .Y(mult_x_1196_n274) );
  AOI21xp33_ASAP7_75t_SL mult_x_1196_U821 ( .A1(mult_x_1196_n729), .A2(n24276), 
        .B(mult_x_1196_n726), .Y(mult_x_1196_n724) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U700 ( .A(n22441), .B(mult_x_1196_n813), .Y(
        mult_x_1196_n263) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U624 ( .A(n22503), .B(mult_x_1196_n805), 
        .Y(mult_x_1196_n255) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U636 ( .A(mult_x_1196_n603), .B(
        mult_x_1196_n806), .Y(mult_x_1196_n256) );
  AOI21xp33_ASAP7_75t_SL mult_x_1196_U556 ( .A1(mult_x_1196_n552), .A2(
        mult_x_1196_n799), .B(mult_x_1196_n545), .Y(mult_x_1196_n543) );
  XNOR2xp5_ASAP7_75t_SL mult_x_1196_U449 ( .A(mult_x_1196_n241), .B(
        mult_x_1196_n476), .Y(u0_0_leon3x0_p0_mul0_m3232_dwm_N49) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77153 ( .A(uart1_uarto_SCALER__1_), .Y(
        n24608) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77146 ( .A(uart1_uarto_SCALER__8_), .Y(
        n24601) );
  INVx1_ASAP7_75t_SL sub_x_2325__cell_77147 ( .A(uart1_uarto_SCALER__7_), .Y(
        n24602) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U381 ( .A(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__5_), .B(u0_0_leon3x0_p0_ici[35]), 
        .Y(DP_OP_1196_128_7433_n336) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U366 ( .A(DP_OP_1196_128_7433_n327), .B(n23949), .Y(DP_OP_1196_128_7433_n32) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U378 ( .A(DP_OP_1196_128_7433_n336), .B(n23950), .Y(DP_OP_1196_128_7433_n33) );
  NOR2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U342 ( .A(DP_OP_1196_128_7433_n307), .B(DP_OP_1196_128_7433_n318), .Y(DP_OP_1196_128_7433_n305) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U331 ( .A1(n23948), .A2(
        DP_OP_1196_128_7433_n310), .B(DP_OP_1196_128_7433_n299), .Y(
        DP_OP_1196_128_7433_n297) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U312 ( .A(DP_OP_1196_128_7433_n278), .B(DP_OP_1196_128_7433_n378), .Y(DP_OP_1196_128_7433_n29) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U195 ( .A1(n23944), .A2(
        DP_OP_1196_128_7433_n198), .B(DP_OP_1196_128_7433_n187), .Y(
        DP_OP_1196_128_7433_n185) );
  INVxp67_ASAP7_75t_SL sub_x_2655__cell_77077 ( .A(timer0_N90), .Y(n24416) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77073 ( .A(timer0_N86), .Y(n24412) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77071 ( .A(timer0_N84), .Y(n24410) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U261 ( .A1(
        DP_OP_1196_128_7433_n267), .A2(DP_OP_1196_128_7433_n240), .B(
        DP_OP_1196_128_7433_n241), .Y(DP_OP_1196_128_7433_n239) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77074 ( .A(timer0_N87), .Y(n24413) );
  INVxp67_ASAP7_75t_SL sub_x_2655__cell_77056 ( .A(timer0_N69), .Y(n24395) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77070 ( .A(timer0_N83), .Y(n24409) );
  INVxp67_ASAP7_75t_SL sub_x_2655__cell_77059 ( .A(timer0_N72), .Y(n24398) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U75 ( .A1(DP_OP_1196_128_7433_n98), 
        .A2(DP_OP_1196_128_7433_n90), .B(DP_OP_1196_128_7433_n91), .Y(
        DP_OP_1196_128_7433_n85) );
  OAI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U408 ( .A1(
        DP_OP_1196_128_7433_n357), .A2(DP_OP_1196_128_7433_n354), .B(
        DP_OP_1196_128_7433_n355), .Y(DP_OP_1196_128_7433_n353) );
  OR2x2_ASAP7_75t_SL mult_x_1196_U1728 ( .A(n22227), .B(n23977), .Y(
        mult_x_1196_n2736) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U237 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n219), .B(DP_OP_1196_128_7433_n220), .Y(
        DP_OP_1196_128_7433_n218) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U287 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n260), .B(DP_OP_1196_128_7433_n261), .Y(
        DP_OP_1196_128_7433_n259) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U200 ( .A(n23964), .B(
        u0_0_leon3x0_p0_divi[14]), .Y(add_x_735_n181) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U176 ( .A(n23965), .B(
        u0_0_leon3x0_p0_divi[16]), .Y(add_x_735_n163) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U305 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n275), .B(DP_OP_1196_128_7433_n276), .Y(
        DP_OP_1196_128_7433_n274) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U273 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n249), .B(DP_OP_1196_128_7433_n250), .Y(
        DP_OP_1196_128_7433_n248) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U48 ( .A(add_x_735_A_29_), .B(
        u0_0_leon3x0_p0_divi[27]), .Y(add_x_735_n68) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U1875 ( .A1(mult_x_1196_n2807), .A2(n24034), .B1(n18402), .B2(mult_x_1196_n2806), .Y(mult_x_1196_n2241) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U185 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n176), .B(DP_OP_1196_128_7433_n177), .Y(
        DP_OP_1196_128_7433_n175) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U205 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n193), .B(DP_OP_1196_128_7433_n194), .Y(
        DP_OP_1196_128_7433_n192) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U219 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n204), .B(DP_OP_1196_128_7433_n205), .Y(
        DP_OP_1196_128_7433_n203) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U107 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n113), .B(DP_OP_1196_128_7433_n114), .Y(
        DP_OP_1196_128_7433_n112) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U123 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n126), .B(DP_OP_1196_128_7433_n127), .Y(
        DP_OP_1196_128_7433_n125) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U155 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n152), .B(DP_OP_1196_128_7433_n153), .Y(
        DP_OP_1196_128_7433_n151) );
  AOI21xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U171 ( .A1(DP_OP_1196_128_7433_n4), 
        .A2(DP_OP_1196_128_7433_n165), .B(DP_OP_1196_128_7433_n166), .Y(
        DP_OP_1196_128_7433_n164) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U81 ( .A(add_x_735_n95), .B(add_x_735_n279), 
        .Y(add_x_735_n10) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U173 ( .A(add_x_735_n163), .B(add_x_735_n287), .Y(add_x_735_n18) );
  OAI21xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U383 ( .A1(
        DP_OP_1196_128_7433_n338), .A2(n23941), .B(DP_OP_1196_128_7433_n339), 
        .Y(DP_OP_1196_128_7433_n337) );
  NAND2xp33_ASAP7_75t_SL add_x_735_U282 ( .A(n18895), .B(add_x_735_n297), .Y(
        add_x_735_n28) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U262 ( .A(add_x_735_n228), .B(add_x_735_n295), .Y(add_x_735_n26) );
  OAI21xp33_ASAP7_75t_SL add_x_735_U78 ( .A1(add_x_735_n92), .A2(
        add_x_735_n102), .B(add_x_735_n95), .Y(add_x_735_n91) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U45 ( .A(add_x_735_n68), .B(add_x_735_n276), 
        .Y(add_x_735_n7) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U30 ( .A(u0_0_leon3x0_p0_iu_fe_pc_27_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_26_), .Y(add_x_746_n23) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U317 ( .A1(add_x_735_n262), .A2(
        add_x_735_n264), .B(add_x_735_n263), .Y(add_x_735_n261) );
  AOI21xp33_ASAP7_75t_SL add_x_735_U88 ( .A1(add_x_735_n118), .A2(
        add_x_735_n99), .B(add_x_735_n100), .Y(add_x_735_n98) );
  AOI21xp5_ASAP7_75t_SL add_x_735_U102 ( .A1(add_x_735_n118), .A2(
        add_x_735_n281), .B(add_x_735_n111), .Y(add_x_735_n109) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U125 ( .A(u0_0_leon3x0_p0_iu_fe_pc_13_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_12_), .Y(add_x_746_n106) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U72 ( .A(u0_0_leon3x0_p0_iu_fe_pc_20_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_21_), .Y(add_x_746_n61) );
  AOI21xp5_ASAP7_75t_SL add_x_735_U12 ( .A1(n24315), .A2(add_x_735_n2), .B(
        n24314), .Y(add_x_735_n40) );
  AOI21xp5_ASAP7_75t_SL add_x_735_U194 ( .A1(add_x_735_n186), .A2(
        add_x_735_n289), .B(add_x_735_n179), .Y(add_x_735_n177) );
  AOI21xp33_ASAP7_75t_SL add_x_735_U26 ( .A1(add_x_735_n2), .A2(add_x_735_n52), 
        .B(add_x_735_n53), .Y(add_x_735_n51) );
  NOR2xp33_ASAP7_75t_SL mult_x_1196_U237 ( .A(mult_x_1196_n847), .B(
        mult_x_1196_n840), .Y(mult_x_1196_n294) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U238 ( .A(mult_x_1196_n847), .B(
        mult_x_1196_n840), .Y(mult_x_1196_n295) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U179 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[19]), .B(u0_0_leon3x0_p0_div0_b[19]), .Y(
        DP_OP_5187J1_124_3275_n170) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U189 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[18]), .B(u0_0_leon3x0_p0_div0_b[18]), .Y(
        DP_OP_5187J1_124_3275_n177) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U11 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[32]), .B(u0_0_leon3x0_p0_div0_b[32]), .Y(
        DP_OP_5187J1_124_3275_n41) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U203 ( .A(
        u0_0_leon3x0_p0_div0_vaddin1[17]), .B(u0_0_leon3x0_p0_div0_b[17]), .Y(
        DP_OP_5187J1_124_3275_n188) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U248 ( .A(mult_x_1196_n851), .B(
        mult_x_1196_n848), .Y(mult_x_1196_n302) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U60 ( .A1(add_x_735_n77), .A2(n22228), .B(
        add_x_735_n78), .Y(add_x_735_n76) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U134 ( .A1(add_x_735_n133), .A2(n22228), .B(
        add_x_735_n134), .Y(add_x_735_n132) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U36 ( .A1(n22228), .A2(add_x_735_n59), .B(
        add_x_735_n60), .Y(add_x_735_n58) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U6 ( .A(n18880), .B(add_x_746_n5), .Y(
        add_x_746_n4) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U192 ( .A1(add_x_735_n176), .A2(
        add_x_735_n214), .B(add_x_735_n177), .Y(add_x_735_n175) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U76 ( .A(add_x_746_n65), .B(n18880), .Y(
        add_x_746_n64) );
  OAI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U347 ( .A1(
        DP_OP_5187J1_124_3275_n297), .A2(DP_OP_5187J1_124_3275_n293), .B(
        DP_OP_5187J1_124_3275_n294), .Y(DP_OP_5187J1_124_3275_n292) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U20 ( .A(n18880), .B(add_x_746_n17), .Y(
        add_x_746_n16) );
  OAI21xp33_ASAP7_75t_SL add_x_735_U148 ( .A1(add_x_735_n144), .A2(n22228), 
        .B(n18889), .Y(add_x_735_n143) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U34 ( .A(n18880), .B(add_x_746_n29), .Y(
        add_x_746_n28) );
  AOI21xp33_ASAP7_75t_SL DP_OP_5187J1_124_3275_U19 ( .A1(
        DP_OP_5187J1_124_3275_n49), .A2(DP_OP_5187J1_124_3275_n72), .B(
        DP_OP_5187J1_124_3275_n50), .Y(DP_OP_5187J1_124_3275_n48) );
  AND2x2_ASAP7_75t_SL mult_x_1196_U245 ( .A(mult_x_1196_n302), .B(n22409), .Y(
        mult_x_1196_n226) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U276 ( .A(mult_x_1196_n869), .B(
        mult_x_1196_n860), .Y(mult_x_1196_n324) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U17 ( .A1(
        DP_OP_5187J1_124_3275_n5), .A2(DP_OP_5187J1_124_3275_n47), .B(
        DP_OP_5187J1_124_3275_n48), .Y(DP_OP_5187J1_124_3275_n46) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U57 ( .A1(
        DP_OP_5187J1_124_3275_n78), .A2(DP_OP_5187J1_124_3275_n3), .B(
        DP_OP_5187J1_124_3275_n79), .Y(DP_OP_5187J1_124_3275_n77) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U83 ( .A1(
        DP_OP_5187J1_124_3275_n3), .A2(DP_OP_5187J1_124_3275_n98), .B(
        DP_OP_5187J1_124_3275_n99), .Y(DP_OP_5187J1_124_3275_n97) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U133 ( .A1(
        DP_OP_5187J1_124_3275_n136), .A2(DP_OP_5187J1_124_3275_n164), .B(
        DP_OP_5187J1_124_3275_n137), .Y(DP_OP_5187J1_124_3275_n135) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U109 ( .A1(
        DP_OP_5187J1_124_3275_n3), .A2(DP_OP_5187J1_124_3275_n315), .B(
        DP_OP_5187J1_124_3275_n119), .Y(DP_OP_5187J1_124_3275_n117) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U43 ( .A1(
        DP_OP_5187J1_124_3275_n67), .A2(DP_OP_5187J1_124_3275_n3), .B(
        DP_OP_5187J1_124_3275_n68), .Y(DP_OP_5187J1_124_3275_n66) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U14 ( .A(
        DP_OP_5187J1_124_3275_n45), .B(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n43) );
  AOI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U159 ( .A1(
        DP_OP_5187J1_124_3275_n164), .A2(DP_OP_5187J1_124_3275_n319), .B(
        DP_OP_5187J1_124_3275_n157), .Y(DP_OP_5187J1_124_3275_n155) );
  OAI21xp33_ASAP7_75t_SL mult_x_1196_U262 ( .A1(mult_x_1196_n316), .A2(
        mult_x_1196_n324), .B(mult_x_1196_n317), .Y(mult_x_1196_n315) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U291 ( .A(mult_x_1196_n339), .B(n24252), 
        .Y(mult_x_1196_n229) );
  OAI21xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U81 ( .A1(n22225), .A2(
        DP_OP_5187J1_124_3275_n96), .B(DP_OP_5187J1_124_3275_n97), .Y(
        DP_OP_5187J1_124_3275_n95) );
  NAND2xp33_ASAP7_75t_SL mult_x_1196_U765 ( .A(mult_x_1196_n690), .B(
        mult_x_1196_n820), .Y(mult_x_1196_n270) );
  NOR2xp67_ASAP7_75t_SL mult_x_1196_U481 ( .A(mult_x_1196_n488), .B(
        mult_x_1196_n495), .Y(mult_x_1196_n486) );
  NAND2xp33_ASAP7_75t_SL mult_x_1196_U555 ( .A(mult_x_1196_n799), .B(n23914), 
        .Y(mult_x_1196_n542) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U469 ( .A(mult_x_1196_n792), .B(
        mult_x_1196_n486), .Y(mult_x_1196_n477) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U427 ( .A(n18533), .B(mult_x_1196_n455), 
        .Y(mult_x_1196_n444) );
  NAND2xp33_ASAP7_75t_SL DP_OP_1196_128_7433_U116 ( .A(
        DP_OP_1196_128_7433_n122), .B(n23942), .Y(DP_OP_1196_128_7433_n17) );
  INVxp67_ASAP7_75t_SL sub_x_2655__cell_77065 ( .A(timer0_N78), .Y(n24404) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U79 ( .A(u0_0_leon3x0_p0_ici[54]), 
        .B(DP_OP_1196_128_7433_n476), .Y(DP_OP_1196_128_7433_n91) );
  INVxp33_ASAP7_75t_SL sub_x_2655__cell_77051 ( .A(timer0_N64), .Y(n24391) );
  INVxp67_ASAP7_75t_SL sub_x_2655__cell_77058 ( .A(timer0_N71), .Y(n24397) );
  INVx1_ASAP7_75t_SL sub_x_2655__cell_77076 ( .A(timer0_N89), .Y(n24415) );
  INVxp67_ASAP7_75t_SL sub_x_2655__cell_77062 ( .A(timer0_N75), .Y(n24401) );
  NAND2xp5_ASAP7_75t_SL DP_OP_1196_128_7433_U417 ( .A(u0_0_leon3x0_p0_ici[30]), 
        .B(DP_OP_1196_128_7433_n452), .Y(DP_OP_1196_128_7433_n357) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U164 ( .A(add_x_735_A_19_), .B(
        u0_0_leon3x0_p0_divi[17]), .Y(add_x_735_n154) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U251 ( .A1(add_x_735_n228), .A2(
        add_x_735_n220), .B(add_x_735_n221), .Y(add_x_735_n219) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U160 ( .A1(add_x_735_n163), .A2(
        add_x_735_n153), .B(add_x_735_n154), .Y(add_x_735_n152) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U197 ( .A(add_x_735_n181), .B(add_x_735_n289), .Y(add_x_735_n20) );
  NAND2xp5_ASAP7_75t_SL add_x_735_U193 ( .A(add_x_735_n289), .B(add_x_735_n185), .Y(add_x_735_n176) );
  OAI21xp33_ASAP7_75t_SL add_x_735_U296 ( .A1(n18885), .A2(add_x_735_n252), 
        .B(add_x_735_n251), .Y(add_x_735_n249) );
  NAND2xp5_ASAP7_75t_SL add_x_746_U177 ( .A(u0_0_leon3x0_p0_iu_fe_pc_4_), .B(
        add_x_746_n152), .Y(add_x_746_n149) );
  OAI21xp5_ASAP7_75t_SL add_x_735_U74 ( .A1(add_x_735_n88), .A2(n22228), .B(
        add_x_735_n89), .Y(add_x_735_n87) );
  NAND2xp5_ASAP7_75t_SL DP_OP_5187J1_124_3275_U132 ( .A(
        DP_OP_5187J1_124_3275_n136), .B(DP_OP_5187J1_124_3275_n163), .Y(
        DP_OP_5187J1_124_3275_n134) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U389 ( .A(mult_x_1196_n416), .B(n18446), 
        .Y(mult_x_1196_n236) );
  NAND2xp33_ASAP7_75t_SL mult_x_1196_U583 ( .A(mult_x_1196_n565), .B(
        mult_x_1196_n801), .Y(mult_x_1196_n251) );
  NAND2xp33_ASAP7_75t_SL mult_x_1196_U692 ( .A(n18929), .B(mult_x_1196_n812), 
        .Y(mult_x_1196_n262) );
  AOI21xp5_ASAP7_75t_SL mult_x_1196_U428 ( .A1(mult_x_1196_n456), .A2(n18533), 
        .B(mult_x_1196_n449), .Y(mult_x_1196_n445) );
  DFFHQNx3_ASAP7_75t_SL uart1_r_reg_TXD_ ( .D(n22235), .CLK(clk), .QN(txd1) );
  SDFHx1_ASAP7_75t_SRAM u0_0_leon3x0_p0_iu_rp_reg_ERROR_ ( .D(
        u0_0_leon3x0_p0_iu_vp_ERROR_), .SI(n18295), .SE(n4818), .CLK(clk), 
        .QN(n4948) );
  DFFHQNx1_ASAP7_75t_SL ahb0_r_reg_HRDATAS__6_ ( .D(n22233), .CLK(clk), .QN(
        ahb0_r_HRDATAS__6_) );
  SDFHx4_ASAP7_75t_SL ahb0_r_reg_HRDATAS__11_ ( .D(n17271), .SI(n19002), .SE(
        n17270), .CLK(clk), .QN(ahb0_r_HRDATAS__11_) );
  DFFHQNx1_ASAP7_75t_SL apb0_r_reg_STATE__1_ ( .D(n22232), .CLK(clk), .QN(
        n4388) );
  SDFHx4_ASAP7_75t_SL ahb0_r_reg_HRDATAS__30_ ( .D(ahb0_r_HADDR__2_), .SI(
        n19002), .SE(n17273), .CLK(clk), .QN(ahb0_r_HRDATAS__30_) );
  SDFHx1_ASAP7_75t_SRAM u0_0_leon3x0_p0_iu_r_reg_W__S__S_ ( .D(n3366), .SI(
        n18295), .SE(n4818), .CLK(clk), .QN(u0_0_dbgo_SU_) );
  SDFHx1_ASAP7_75t_SRAM u0_0_leon3x0_p0_iu_r_reg_M__WERR_ ( .D(
        u0_0_leon3x0_p0_iu_v_M__WERR_), .SI(n18295), .SE(n22380), .CLK(clk), 
        .QN(n1769) );
  OAI22xp33_ASAP7_75t_SL apb0_r_reg_PRDATA__5__U3 ( .A1(n16599), .A2(
        apb0_r_CFGSEL_), .B1(n1637), .B2(n31954), .Y(n22231) );
  SDFHx4_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__INST__26_ ( .D(n3766), 
        .SI(n18295), .SE(n18295), .CLK(clk), .QN(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__26_) );
  DFFHQx4_ASAP7_75t_SL sr1_r_reg_READ_ ( .D(n22229), .CLK(clk), .Q(read) );
  SDFHx4_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_A__CTRL__CNT__1_ ( .D(n4165), 
        .SI(n18295), .SE(n18295), .CLK(clk), .QN(
        u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__1_) );
  DFFHQx4_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_icache0_r_reg_FLUSH2_ ( .D(n24555), .CLK(clk), .Q(n3065) );
  SDFHx4_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__LDBP1_ ( .D(n3314), .SI(
        n18295), .SE(n18295), .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__LDBP1_)
         );
  DFFHQNx2_ASAP7_75t_SL uart1_r_reg_TRADDR__0_ ( .D(n2238), .CLK(clk), .QN(
        uart1_r_TRADDR__0_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__CWP__0_ ( .D(n2788), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_A__CWP__0_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__CTRL__INST__19_ ( .D(n3604), .CLK(clk), .QN(u0_0_leon3x0_p0_muli[9]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP2__17_ ( .D(n2588), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP2__17_) );
  DFFHQNx2_ASAP7_75t_SL apb0_r_reg_PRDATA__5_ ( .D(n22230), .CLK(clk), .QN(
        ahbso_1__HRDATA__5_) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__55_ ( .D(
        n4199), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[54]) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__58_ ( .D(
        n4193), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[57]) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA2__9_ ( 
        .D(n4558), .CLK(clk), .QN(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__9_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__DATA1__1_ ( 
        .D(n4534), .CLK(clk), .QN(u0_0_leon3x0_p0_c0mmu_mcdi[5]) );
  SDFHx1_ASAP7_75t_SL u0_0_leon3x0_p0_c0mmu_dcache0_r_reg_WB__LOCK_ ( .D(n4074), .SI(n18295), .SE(n22380), .CLK(clk), .QN(n4076) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__ICC__2_ ( .D(n4579), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_de_icc_2_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__CNT__1_ ( .D(n4408), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_M__ICC__1_ ( .D(n4338), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_de_icc_1_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__19_ ( .D(n24446), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__31_ ( .D(n24442), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__31_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__22_ ( .D(n24450), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__22_) );
  DFFHQNx1_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_D__INST__0__21_ ( .D(n24447), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__21_) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__56_ ( .D(
        n4197), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[55]) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__61_ ( .D(
        n4187), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[60]) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__49_ ( .D(
        n4211), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[48]) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__60_ ( .D(
        n4189), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[59]) );
  NAND2x1_ASAP7_75t_SL mult_x_1196_U313 ( .A(mult_x_1196_n355), .B(
        mult_x_1196_n781), .Y(mult_x_1196_n231) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2289 ( .A(n24070), .B(n23965), .Y(
        mult_x_1196_n3001) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__63_ ( .D(
        n4183), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[62]) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__13_ ( .D(n4660), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__13_) );
  NAND2x1_ASAP7_75t_SL mult_x_1196_U778 ( .A(n24273), .B(n24310), .Y(
        mult_x_1196_n696) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U523 ( .A(mult_x_1196_n520), .B(
        mult_x_1196_n796), .Y(mult_x_1196_n246) );
  NOR2x1_ASAP7_75t_SL mult_x_1196_U797 ( .A(n22333), .B(mult_x_1196_n714), .Y(
        mult_x_1196_n709) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__51_ ( .D(
        n4207), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[50]) );
  OAI22x1_ASAP7_75t_SL mult_x_1196_U1890 ( .A1(mult_x_1196_n2822), .A2(n24034), 
        .B1(n22251), .B2(mult_x_1196_n2821), .Y(mult_x_1196_n2256) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U541 ( .A(n22264), .B(n23914), .Y(
        mult_x_1196_n531) );
  DFFHQNx3_ASAP7_75t_SL u0_0_leon3x0_p0_mul0_m3232_dwm_p_i_reg_1__41_ ( .D(
        n4227), .CLK(clk), .QN(u0_0_leon3x0_p0_mulo[40]) );
  OAI22x1_ASAP7_75t_SL mult_x_1196_U2305 ( .A1(mult_x_1196_n3015), .A2(n22563), 
        .B1(mult_x_1196_n3014), .B2(n22540), .Y(mult_x_1196_n2443) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2004 ( .A(n24069), .B(n23971), .Y(
        mult_x_1196_n2864) );
  NAND2x1p5_ASAP7_75t_SRAM mult_x_1196_U421 ( .A(mult_x_1196_n442), .B(
        mult_x_1196_n788), .Y(mult_x_1196_n238) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U1822 ( .A1(mult_x_1196_n2791), .A2(n24039), .B1(mult_x_1196_n2790), .B2(n22391), .Y(mult_x_1196_n2225) );
  NAND2xp33_ASAP7_75t_SL mult_x_1196_U433 ( .A(mult_x_1196_n451), .B(n23573), 
        .Y(mult_x_1196_n239) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__5_ ( .D(n4380), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__5_) );
  NAND2x1p5_ASAP7_75t_SRAM mult_x_1196_U403 ( .A(mult_x_1196_n423), .B(n18416), 
        .Y(mult_x_1196_n237) );
  AOI21xp5_ASAP7_75t_SRAM mult_x_1196_U470 ( .A1(mult_x_1196_n487), .A2(
        mult_x_1196_n792), .B(mult_x_1196_n480), .Y(mult_x_1196_n478) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2498 ( .A(n24066), .B(n23091), .Y(
        mult_x_1196_n3099) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2428 ( .A(n24067), .B(n24081), .Y(
        mult_x_1196_n3066) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__3_ ( .D(n3961), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__3_) );
  NAND2x1_ASAP7_75t_SRAM mult_x_1196_U445 ( .A(mult_x_1196_n460), .B(n23732), 
        .Y(mult_x_1196_n240) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__1_ ( .D(n4471), .CLK(
        clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__1_) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__11_ ( .D(n4461), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__11_) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U409 ( .A(n22676), .B(mult_x_1196_n464), 
        .Y(mult_x_1196_n429) );
  NAND2xp5_ASAP7_75t_SL mult_x_1196_U463 ( .A(mult_x_1196_n475), .B(
        mult_x_1196_n791), .Y(mult_x_1196_n241) );
  NAND2x2_ASAP7_75t_SRAM mult_x_1196_U341 ( .A(mult_x_1196_n377), .B(n24305), 
        .Y(mult_x_1196_n233) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__15_ ( .D(n4639), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__15_) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2620 ( .A(n24046), .B(n23960), .Y(
        mult_x_1196_n3147) );
  OAI22x1_ASAP7_75t_SL mult_x_1196_U2371 ( .A1(n18550), .A2(mult_x_1196_n3043), 
        .B1(mult_x_1196_n3044), .B2(n24007), .Y(mult_x_1196_n2472) );
  NOR2x1_ASAP7_75t_SL mult_x_1196_U531 ( .A(n22468), .B(mult_x_1196_n535), .Y(
        mult_x_1196_n524) );
  OAI22xp5_ASAP7_75t_SL mult_x_1196_U2184 ( .A1(mult_x_1196_n2968), .A2(n23141), .B1(n24017), .B2(mult_x_1196_n2967), .Y(mult_x_1196_n2396) );
  XNOR2x1_ASAP7_75t_SL mult_x_1196_U2072 ( .A(n24066), .B(n23089), .Y(
        mult_x_1196_n2895) );
  NAND2xp5_ASAP7_75t_SRAM mult_x_1196_U559 ( .A(mult_x_1196_n547), .B(
        mult_x_1196_n799), .Y(mult_x_1196_n249) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_E__OP1__24_ ( .D(n4509), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_E__OP1__24_) );
  XNOR2x1_ASAP7_75t_SL mult_x_1196_U2692 ( .A(n24047), .B(n23957), .Y(
        mult_x_1196_n3182) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2429 ( .A(n24068), .B(n24081), .Y(
        mult_x_1196_n3067) );
  XNOR2x2_ASAP7_75t_SL mult_x_1196_U2059 ( .A(n24053), .B(n23089), .Y(
        mult_x_1196_n2882) );
  DFFHQNx2_ASAP7_75t_SL u0_0_leon3x0_p0_iu_r_reg_X__DATA__0__26_ ( .D(n4611), 
        .CLK(clk), .QN(u0_0_leon3x0_p0_iu_r_X__DATA__0__26_) );
  XNOR2x1_ASAP7_75t_SL mult_x_1196_U2693 ( .A(n24048), .B(n23957), .Y(
        mult_x_1196_n3183) );
  TIELOx1_ASAP7_75t_SL U19751 ( .L(n18295) );
  TIEHIx1_ASAP7_75t_SL U19752 ( .H(n19002) );
  A2O1A1Ixp33_ASAP7_75t_SL U19753 ( .A1(n29517), .A2(n19002), .B(n22203), .C(
        n19002), .Y(n22204) );
  A2O1A1Ixp33_ASAP7_75t_SL U19754 ( .A1(n29516), .A2(n19002), .B(n30833), .C(
        n24694), .Y(n22205) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19755 ( .A1(n29521), .A2(n22202), .B(n22204), 
        .C(n19002), .D(n22205), .Y(n4780) );
  A2O1A1Ixp33_ASAP7_75t_SL U19756 ( .A1(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__3_), 
        .A2(n19002), .B(n29883), .C(n19002), .Y(n22191) );
  A2O1A1Ixp33_ASAP7_75t_SL U19757 ( .A1(n22191), .A2(n30677), .B(n22192), .C(
        n19002), .Y(n22193) );
  A2O1A1Ixp33_ASAP7_75t_SL U19758 ( .A1(n22191), .A2(n19002), .B(n29886), .C(
        n19002), .Y(n22194) );
  O2A1O1Ixp33_ASAP7_75t_SL U19759 ( .A1(n22193), .A2(n22194), .B(n19002), .C(
        n22197), .Y(n4762) );
  A2O1A1Ixp33_ASAP7_75t_SL U19760 ( .A1(n22427), .A2(n19002), .B(n32575), .C(
        n22190), .Y(n4760) );
  A2O1A1Ixp33_ASAP7_75t_SL U19761 ( .A1(n31940), .A2(n19002), .B(n31973), .C(
        n19002), .Y(n22188) );
  A2O1A1Ixp33_ASAP7_75t_SL U19762 ( .A1(n32004), .A2(n19002), .B(n31941), .C(
        n19002), .Y(n22189) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19763 ( .A1(n32008), .A2(n22187), .B(n22188), 
        .C(n19002), .D(n22189), .Y(n4740) );
  A2O1A1Ixp33_ASAP7_75t_SL U19764 ( .A1(uart1_r_TSHIFT__9_), .A2(n21967), .B(
        n29951), .C(n19002), .Y(n4709) );
  A2O1A1Ixp33_ASAP7_75t_SL U19765 ( .A1(n19002), .A2(uart1_r_LOOPB_), .B(
        n21727), .C(n21730), .Y(n4698) );
  A2O1A1Ixp33_ASAP7_75t_SL U19766 ( .A1(n31058), .A2(n19002), .B(n28224), .C(
        n19002), .Y(n22185) );
  A2O1A1Ixp33_ASAP7_75t_SL U19767 ( .A1(n31059), .A2(n19002), .B(n28225), .C(
        n19002), .Y(n22186) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19768 ( .A1(n31061), .A2(uart1_r_RHOLD__0__3_), 
        .B(n22185), .C(n19002), .D(n22186), .Y(n4695) );
  A2O1A1Ixp33_ASAP7_75t_SL U19769 ( .A1(n29744), .A2(n29745), .B(n22183), .C(
        n19002), .Y(n22184) );
  O2A1O1Ixp33_ASAP7_75t_SL U19770 ( .A1(n21962), .A2(n31047), .B(n19002), .C(
        n21965), .Y(n4660) );
  A2O1A1Ixp33_ASAP7_75t_SL U19771 ( .A1(n22422), .A2(n19002), .B(n27222), .C(
        n19002), .Y(n22181) );
  A2O1A1Ixp33_ASAP7_75t_SL U19772 ( .A1(n28330), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n22182) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19773 ( .A1(n31662), .A2(n23396), .B(n22181), 
        .C(n19002), .D(n22182), .Y(n4657) );
  A2O1A1Ixp33_ASAP7_75t_SL U19774 ( .A1(n28585), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n22172) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19775 ( .A1(n30644), .A2(n28586), .B(n22172), 
        .C(n19002), .D(n22175), .Y(n22176) );
  A2O1A1Ixp33_ASAP7_75t_SL U19776 ( .A1(n30645), .A2(n19002), .B(n30496), .C(
        n22176), .Y(n22177) );
  A2O1A1Ixp33_ASAP7_75t_SL U19777 ( .A1(n22432), .A2(n30495), .B(n22177), .C(
        n19002), .Y(n22178) );
  A2O1A1Ixp33_ASAP7_75t_SL U19778 ( .A1(n30595), .A2(n19002), .B(n22178), .C(
        n19002), .Y(n22179) );
  A2O1A1Ixp33_ASAP7_75t_SL U19779 ( .A1(n22178), .A2(n30593), .B(n22179), .C(
        n19002), .Y(n22180) );
  A2O1A1Ixp33_ASAP7_75t_SL U19780 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP2__14_), 
        .A2(n22171), .B(n22180), .C(n19002), .Y(n4654) );
  O2A1O1Ixp5_ASAP7_75t_SL U19781 ( .A1(n21955), .A2(n21956), .B(n19002), .C(
        n30580), .Y(n21957) );
  A2O1A1Ixp33_ASAP7_75t_SL U19782 ( .A1(n22422), .A2(n19002), .B(n29793), .C(
        n19002), .Y(n22161) );
  A2O1A1Ixp33_ASAP7_75t_SL U19783 ( .A1(n29794), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n22162) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19784 ( .A1(n31662), .A2(n18606), .B(n22161), 
        .C(n19002), .D(n22162), .Y(n4620) );
  A2O1A1Ixp33_ASAP7_75t_SL U19785 ( .A1(n19002), .A2(n24646), .B(n29787), .C(
        n20832), .Y(n4602) );
  A2O1A1Ixp33_ASAP7_75t_SL U19786 ( .A1(n24638), .A2(n19002), .B(n22154), .C(
        n19002), .Y(n22155) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19787 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__28_), .B(n24680), .C(n19002), .D(n22155), 
        .Y(n22156) );
  A2O1A1Ixp33_ASAP7_75t_SL U19788 ( .A1(n30394), .A2(n30236), .B(n22158), .C(
        n19002), .Y(n22159) );
  A2O1A1Ixp33_ASAP7_75t_SL U19789 ( .A1(n30426), .A2(n19002), .B(n30237), .C(
        n22159), .Y(n22160) );
  A2O1A1Ixp33_ASAP7_75t_SL U19790 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_divi[59]), .C(n22160), .Y(n4590) );
  A2O1A1Ixp33_ASAP7_75t_SL U19791 ( .A1(n24659), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__TT__5_), .B(n22153), .C(n19002), .Y(
        n4567) );
  A2O1A1Ixp33_ASAP7_75t_SL U19792 ( .A1(n22422), .A2(n19002), .B(n27176), .C(
        n19002), .Y(n22149) );
  A2O1A1Ixp33_ASAP7_75t_SL U19793 ( .A1(n27177), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n22150) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19794 ( .A1(n31662), .A2(n23658), .B(n22149), 
        .C(n19002), .D(n22150), .Y(n4554) );
  A2O1A1Ixp33_ASAP7_75t_SL U19795 ( .A1(n19002), .A2(n24646), .B(n31055), .C(
        n21441), .Y(n4549) );
  A2O1A1Ixp33_ASAP7_75t_SL U19796 ( .A1(u0_0_leon3x0_p0_div0_addout_31_), .A2(
        n24639), .B(n20674), .C(n19002), .Y(n4507) );
  A2O1A1Ixp33_ASAP7_75t_SL U19797 ( .A1(n22427), .A2(n19002), .B(rf_di_w[31]), 
        .C(n22148), .Y(n4490) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U19798 ( .A1(n30206), .A2(n22380), .B(n19002), 
        .C(u0_0_leon3x0_p0_c0mmu_dcache0_r_RBURST_), .Y(n21934) );
  A2O1A1Ixp33_ASAP7_75t_SL U19799 ( .A1(n19002), .A2(n30203), .B(n21934), .C(
        n21937), .Y(n4481) );
  A2O1A1Ixp33_ASAP7_75t_SL U19800 ( .A1(n22420), .A2(n19002), .B(n28353), .C(
        n31422), .Y(n22143) );
  A2O1A1Ixp33_ASAP7_75t_SL U19801 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[1]), 
        .B(n22143), .C(n19002), .Y(n22144) );
  A2O1A1Ixp33_ASAP7_75t_SL U19802 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_1_), .B(n22146), .C(n19002), .Y(n4473) );
  A2O1A1Ixp33_ASAP7_75t_SL U19803 ( .A1(n22420), .A2(n19002), .B(n29926), .C(
        n31422), .Y(n22139) );
  A2O1A1Ixp33_ASAP7_75t_SL U19804 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[8]), 
        .B(n22139), .C(n19002), .Y(n22140) );
  A2O1A1Ixp33_ASAP7_75t_SL U19805 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_8_), .B(n22142), .C(n19002), .Y(n4440) );
  A2O1A1Ixp33_ASAP7_75t_SL U19806 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[8]), .C(n22138), .Y(n4435) );
  A2O1A1Ixp33_ASAP7_75t_SL U19807 ( .A1(n24647), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), .B(n22136), .C(n19002), .Y(
        n4408) );
  A2O1A1Ixp33_ASAP7_75t_SL U19808 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__27_), .C(n22134), .Y(n4397) );
  A2O1A1Ixp33_ASAP7_75t_SL U19809 ( .A1(n22422), .A2(n19002), .B(n29692), .C(
        n19002), .Y(n22132) );
  A2O1A1Ixp33_ASAP7_75t_SL U19810 ( .A1(n29906), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n22133) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19811 ( .A1(n31662), .A2(n18325), .B(n22132), 
        .C(n19002), .D(n22133), .Y(n4379) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U19812 ( .A1(n31016), .A2(n31015), .B(n19002), 
        .C(n24677), .Y(n21695) );
  A2O1A1Ixp33_ASAP7_75t_SL U19813 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__21_), .C(n21924), .Y(n4341) );
  A2O1A1Ixp33_ASAP7_75t_SL U19814 ( .A1(n22379), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__30_), .C(n22131), .Y(n4322) );
  A2O1A1Ixp33_ASAP7_75t_SL U19815 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_), .B(n24650), .C(n21917), .Y(
        n4181) );
  A2O1A1Ixp33_ASAP7_75t_SL U19816 ( .A1(n19002), .A2(n18799), .B(n22377), .C(
        n21913), .Y(n4167) );
  A2O1A1Ixp33_ASAP7_75t_SL U19817 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .B(n24657), .C(n21001), .Y(
        n4157) );
  A2O1A1Ixp33_ASAP7_75t_SL U19818 ( .A1(n22427), .A2(n19002), .B(n27174), .C(
        n22127), .Y(n4145) );
  A2O1A1Ixp33_ASAP7_75t_SL U19819 ( .A1(n22427), .A2(n19002), .B(n30972), .C(
        n22126), .Y(n4143) );
  A2O1A1Ixp33_ASAP7_75t_SL U19820 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[12]), .B(n22379), .C(n21912), .Y(n4141)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U19821 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), .B(n24655), .C(n21410), .Y(
        n4099) );
  A2O1A1Ixp33_ASAP7_75t_SL U19822 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_), .B(n24654), .C(n21185), .Y(
        n4097) );
  A2O1A1Ixp33_ASAP7_75t_SL U19823 ( .A1(n19002), .A2(n22421), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__23_), .C(n21911), .Y(n4085) );
  A2O1A1Ixp33_ASAP7_75t_SL U19824 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__4_), .B(n24656), .C(n20640), .Y(
        n4057) );
  A2O1A1Ixp33_ASAP7_75t_SL U19825 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__19_), .C(n21910), .Y(n4042) );
  A2O1A1Ixp33_ASAP7_75t_SL U19826 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__17_), .A2(n19002), .B(n24649), .C(
        n22125), .Y(n4026) );
  A2O1A1Ixp33_ASAP7_75t_SL U19827 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[2]), .A2(
        n31429), .B(n21175), .C(n19002), .Y(n21176) );
  A2O1A1Ixp33_ASAP7_75t_SL U19828 ( .A1(n19002), .A2(n31428), .B(n21176), .C(
        n21179), .Y(n21180) );
  A2O1A1Ixp33_ASAP7_75t_SL U19829 ( .A1(u0_0_leon3x0_p0_iu_v_A__CWP__2_), .A2(
        n19002), .B(n22421), .C(n21180), .Y(n4018) );
  A2O1A1Ixp33_ASAP7_75t_SL U19830 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__18_), .C(n22124), .Y(n3998) );
  A2O1A1Ixp33_ASAP7_75t_SL U19831 ( .A1(n19002), .A2(n24646), .B(n29626), .C(
        n19880), .Y(n3963) );
  A2O1A1Ixp33_ASAP7_75t_SL U19832 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[34]), .C(n21904), .Y(n3942) );
  A2O1A1Ixp33_ASAP7_75t_SL U19833 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__5_), .C(n21170), .Y(n3917) );
  A2O1A1Ixp33_ASAP7_75t_SL U19834 ( .A1(n32564), .A2(n19002), .B(n32124), .C(
        n19002), .Y(n22122) );
  A2O1A1Ixp33_ASAP7_75t_SL U19835 ( .A1(n22405), .A2(n19002), .B(n22123), .C(
        n19002), .Y(n18248) );
  A2O1A1Ixp33_ASAP7_75t_SL U19836 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_), .A2(n19002), .B(n22377), .C(
        n22121), .Y(n3873) );
  A2O1A1Ixp33_ASAP7_75t_SL U19837 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__7_), .C(n21169), .Y(n3850) );
  A2O1A1Ixp33_ASAP7_75t_SL U19838 ( .A1(n19002), .A2(n22421), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__26_), .C(n20638), .Y(n3838) );
  A2O1A1Ixp33_ASAP7_75t_SL U19839 ( .A1(n19002), .A2(n24646), .B(n29866), .C(
        n21900), .Y(n3834) );
  A2O1A1Ixp33_ASAP7_75t_SL U19840 ( .A1(n19002), .A2(n24646), .B(n30609), .C(
        n21899), .Y(n3830) );
  A2O1A1Ixp33_ASAP7_75t_SL U19841 ( .A1(n19002), .A2(n24646), .B(n30452), .C(
        n21897), .Y(n3826) );
  A2O1A1Ixp33_ASAP7_75t_SL U19842 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_muli[6]), .C(n21398), .Y(n3822) );
  A2O1A1Ixp33_ASAP7_75t_SL U19843 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__9_), .C(n21653), .Y(n3816) );
  A2O1A1Ixp33_ASAP7_75t_SL U19844 ( .A1(n19002), .A2(n22378), .B(n30383), .C(
        n20986), .Y(n3812) );
  A2O1A1Ixp33_ASAP7_75t_SL U19845 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__12_), .C(n21896), .Y(n3810) );
  A2O1A1Ixp33_ASAP7_75t_SL U19846 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__13_), .C(n21895), .Y(n3808) );
  A2O1A1Ixp33_ASAP7_75t_SL U19847 ( .A1(n19002), .A2(n22378), .B(n30356), .C(
        n21652), .Y(n3806) );
  A2O1A1Ixp33_ASAP7_75t_SL U19848 ( .A1(n19002), .A2(n22378), .B(n30340), .C(
        n21396), .Y(n3804) );
  A2O1A1Ixp33_ASAP7_75t_SL U19849 ( .A1(n19002), .A2(n22428), .B(n30333), .C(
        n21651), .Y(n3802) );
  A2O1A1Ixp33_ASAP7_75t_SL U19850 ( .A1(n19002), .A2(n22428), .B(n30322), .C(
        n21894), .Y(n3800) );
  A2O1A1Ixp33_ASAP7_75t_SL U19851 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__20_), .C(n21893), .Y(n3794) );
  A2O1A1Ixp33_ASAP7_75t_SL U19852 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__5_), .C(n22120), .Y(n3691) );
  A2O1A1Ixp33_ASAP7_75t_SL U19853 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__6_), .B(n22377), .C(n21883), .Y(
        n3682) );
  A2O1A1Ixp33_ASAP7_75t_SL U19854 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__7_), .B(n22377), .C(n21881), .Y(
        n3673) );
  A2O1A1Ixp33_ASAP7_75t_SL U19855 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__9_), .B(n24652), .C(n21879), .Y(
        n3655) );
  A2O1A1Ixp33_ASAP7_75t_SL U19856 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__0_), 
        .A2(n19002), .B(n22377), .C(n22119), .Y(n3528) );
  A2O1A1Ixp33_ASAP7_75t_SL U19857 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__LD_), 
        .A2(n19002), .B(n22377), .C(n22118), .Y(n3512) );
  A2O1A1Ixp33_ASAP7_75t_SL U19858 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[32]), .C(n21381), .Y(n3468) );
  A2O1A1Ixp33_ASAP7_75t_SL U19859 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__7_), .B(n22428), .C(n19706), .Y(
        n3444) );
  A2O1A1Ixp33_ASAP7_75t_SL U19860 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[36]), .C(n20976), .Y(n3438) );
  A2O1A1Ixp33_ASAP7_75t_SL U19861 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[37]), .C(n21877), .Y(n3428) );
  A2O1A1Ixp33_ASAP7_75t_SL U19862 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[39]), .C(n21876), .Y(n3418) );
  A2O1A1Ixp33_ASAP7_75t_SL U19863 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[53]), .C(n21875), .Y(n3408) );
  A2O1A1Ixp33_ASAP7_75t_SL U19864 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[55]), .C(n21874), .Y(n3398) );
  A2O1A1Ixp33_ASAP7_75t_SL U19865 ( .A1(n19002), .A2(n24646), .B(rf_di_w[1]), 
        .C(n21873), .Y(n3387) );
  A2O1A1Ixp33_ASAP7_75t_SL U19866 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__ET_), .B(n22377), .C(n20971), .Y(n3372) );
  A2O1A1Ixp33_ASAP7_75t_SL U19867 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__TT__4_), .B(n22377), .C(n21641), .Y(
        n3348) );
  A2O1A1Ixp33_ASAP7_75t_SL U19868 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[57]), .C(n21374), .Y(n3290) );
  A2O1A1Ixp33_ASAP7_75t_SL U19869 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[56]), 
        .B(n24651), .C(n20074), .Y(n3276) );
  A2O1A1Ixp33_ASAP7_75t_SL U19870 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[51]), .C(n21871), .Y(n3250) );
  A2O1A1Ixp33_ASAP7_75t_SL U19871 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[49]), .C(n21870), .Y(n3238) );
  A2O1A1Ixp33_ASAP7_75t_SL U19872 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[43]), .C(n21869), .Y(n3226) );
  A2O1A1Ixp33_ASAP7_75t_SL U19873 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[42]), .C(n21868), .Y(n3214) );
  A2O1A1Ixp33_ASAP7_75t_SL U19874 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[30]), .C(n21867), .Y(n3200) );
  A2O1A1Ixp33_ASAP7_75t_SL U19875 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__3_), 
        .A2(n19002), .B(n24653), .C(n22117), .Y(n3184) );
  A2O1A1Ixp33_ASAP7_75t_SL U19876 ( .A1(n19002), .A2(n22428), .B(rf_di_w[10]), 
        .C(n21144), .Y(n3166) );
  A2O1A1Ixp33_ASAP7_75t_SL U19877 ( .A1(n19002), .A2(n30699), .B(n22414), .C(
        n20309), .Y(n20310) );
  A2O1A1Ixp33_ASAP7_75t_SL U19878 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__10_), .B(n20310), .C(n19002), .Y(n3145)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U19879 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[31]), .C(n22115), .Y(n3125) );
  A2O1A1Ixp33_ASAP7_75t_SL U19880 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[30]), .C(n22113), .Y(n3123) );
  A2O1A1Ixp33_ASAP7_75t_SL U19881 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[27]), .C(n22111), .Y(n3117) );
  A2O1A1Ixp33_ASAP7_75t_SL U19882 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[26]), .C(n22109), .Y(n3115) );
  A2O1A1Ixp33_ASAP7_75t_SL U19883 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[24]), .C(n22107), .Y(n3111) );
  A2O1A1Ixp33_ASAP7_75t_SL U19884 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[23]), .C(n21630), .Y(n3109) );
  A2O1A1Ixp33_ASAP7_75t_SL U19885 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[22]), .C(n21860), .Y(n3107) );
  A2O1A1Ixp33_ASAP7_75t_SL U19886 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[21]), .C(n22105), .Y(n3105) );
  A2O1A1Ixp33_ASAP7_75t_SL U19887 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[20]), .C(n21859), .Y(n3103) );
  A2O1A1Ixp33_ASAP7_75t_SL U19888 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[19]), .C(n22103), .Y(n3101) );
  A2O1A1Ixp33_ASAP7_75t_SL U19889 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[18]), .C(n22101), .Y(n3099) );
  A2O1A1Ixp33_ASAP7_75t_SL U19890 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[17]), .C(n22099), .Y(n3097) );
  A2O1A1Ixp33_ASAP7_75t_SL U19891 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[1]), .C(n21852), .Y(n3081) );
  A2O1A1Ixp33_ASAP7_75t_SL U19892 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[0]), .C(n21851), .Y(n3079) );
  A2O1A1Ixp33_ASAP7_75t_SL U19893 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_dci[37]), .C(n21359), .Y(n3077) );
  A2O1A1Ixp33_ASAP7_75t_SL U19894 ( .A1(n30186), .A2(n30165), .B(n30164), .C(
        n19002), .Y(n22096) );
  A2O1A1Ixp33_ASAP7_75t_SL U19895 ( .A1(n22422), .A2(n19002), .B(n30463), .C(
        n19002), .Y(n22092) );
  A2O1A1Ixp33_ASAP7_75t_SL U19896 ( .A1(n28357), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n22093) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19897 ( .A1(n31662), .A2(n22939), .B(n22092), 
        .C(n19002), .D(n22093), .Y(n3037) );
  A2O1A1Ixp33_ASAP7_75t_SL U19898 ( .A1(n31694), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n22090) );
  A2O1A1Ixp33_ASAP7_75t_SL U19899 ( .A1(n31703), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n22091) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19900 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__1_), .B(n22090), .C(n19002), .D(
        n22091), .Y(n2996) );
  A2O1A1Ixp33_ASAP7_75t_SL U19901 ( .A1(n31501), .A2(n19002), .B(apbi[27]), 
        .C(n22089), .Y(n2906) );
  A2O1A1Ixp33_ASAP7_75t_SL U19902 ( .A1(n28167), .A2(uart1_uarto_SCALER__7_), 
        .B(n22419), .C(n19002), .Y(n20780) );
  A2O1A1Ixp33_ASAP7_75t_SL U19903 ( .A1(n19002), .A2(uart1_r_RXCLK__0_), .B(
        uart1_r_TICK_), .C(n24694), .Y(n21616) );
  O2A1O1Ixp33_ASAP7_75t_SL U19904 ( .A1(n21616), .A2(n21617), .B(n19002), .C(
        n28186), .Y(n21618) );
  A2O1A1Ixp33_ASAP7_75t_SL U19905 ( .A1(n29383), .A2(n19002), .B(n30833), .C(
        n22085), .Y(n17785) );
  A2O1A1Ixp33_ASAP7_75t_SL U19906 ( .A1(n24646), .A2(n19002), .B(n32165), .C(
        n22083), .Y(n2782) );
  A2O1A1Ixp33_ASAP7_75t_SL U19907 ( .A1(n19002), .A2(n22421), .B(
        u0_0_leon3x0_p0_muli[3]), .C(n21831), .Y(n2745) );
  A2O1A1Ixp33_ASAP7_75t_SL U19908 ( .A1(n30428), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n22080) );
  A2O1A1Ixp33_ASAP7_75t_SL U19909 ( .A1(n30429), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n22081) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19910 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__4_), 
        .A2(n31403), .B(n22080), .C(n19002), .D(n22081), .Y(n2727) );
  A2O1A1Ixp33_ASAP7_75t_SL U19911 ( .A1(n22427), .A2(n19002), .B(rf_di_w[12]), 
        .C(n22079), .Y(n2665) );
  A2O1A1Ixp33_ASAP7_75t_SL U19912 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[41]), 
        .B(n22428), .C(n21826), .Y(n2649) );
  A2O1A1Ixp33_ASAP7_75t_SL U19913 ( .A1(n22422), .A2(n19002), .B(n27223), .C(
        n19002), .Y(n22076) );
  A2O1A1Ixp33_ASAP7_75t_SL U19914 ( .A1(n27264), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n22077) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19915 ( .A1(n31662), .A2(n23665), .B(n22076), 
        .C(n19002), .D(n22077), .Y(n2635) );
  A2O1A1Ixp33_ASAP7_75t_SL U19916 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[45]), .C(n21822), .Y(n2603) );
  A2O1A1Ixp33_ASAP7_75t_SL U19917 ( .A1(n22422), .A2(n19002), .B(n28320), .C(
        n19002), .Y(n22074) );
  A2O1A1Ixp33_ASAP7_75t_SL U19918 ( .A1(n27036), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n22075) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19919 ( .A1(n31662), .A2(n24231), .B(n22074), 
        .C(n19002), .D(n22075), .Y(n2564) );
  A2O1A1Ixp33_ASAP7_75t_SL U19920 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[47]), .C(n21818), .Y(n2554) );
  A2O1A1Ixp33_ASAP7_75t_SL U19921 ( .A1(n19002), .A2(n24646), .B(rf_di_w[20]), 
        .C(n21817), .Y(n2521) );
  A2O1A1Ixp33_ASAP7_75t_SL U19922 ( .A1(n19002), .A2(n24646), .B(n30272), .C(
        n21816), .Y(n2513) );
  A2O1A1Ixp33_ASAP7_75t_SL U19923 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[50]), 
        .B(n22428), .C(n21815), .Y(n2502) );
  A2O1A1Ixp33_ASAP7_75t_SL U19924 ( .A1(n22405), .A2(n19002), .B(n32538), .C(
        n19002), .Y(n22073) );
  A2O1A1Ixp33_ASAP7_75t_SL U19925 ( .A1(n32537), .A2(n19002), .B(n22073), .C(
        n19002), .Y(n2493) );
  A2O1A1Ixp33_ASAP7_75t_SL U19926 ( .A1(n19002), .A2(n22427), .B(n30257), .C(
        n21813), .Y(n2486) );
  A2O1A1Ixp33_ASAP7_75t_SL U19927 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[52]), 
        .B(n22428), .C(n21812), .Y(n2475) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19928 ( .A1(n25995), .A2(n2387), .B(n24695), .C(
        n19002), .D(n22072), .Y(n17457) );
  A2O1A1Ixp33_ASAP7_75t_SL U19929 ( .A1(n19002), .A2(n22427), .B(rf_di_w[30]), 
        .C(n21810), .Y(n2372) );
  A2O1A1Ixp33_ASAP7_75t_SL U19930 ( .A1(n19002), .A2(n27947), .B(
        uart1_r_THOLD__24__0_), .C(n21805), .Y(n2265) );
  A2O1A1Ixp33_ASAP7_75t_SL U19931 ( .A1(n29383), .A2(n19002), .B(n28116), .C(
        n22071), .Y(n17802) );
  A2O1A1Ixp33_ASAP7_75t_SL U19932 ( .A1(n19002), .A2(n22433), .B(n32922), .C(
        n21804), .Y(n1718) );
  A2O1A1Ixp33_ASAP7_75t_SL U19933 ( .A1(n19002), .A2(n22433), .B(n32911), .C(
        n21801), .Y(n1710) );
  A2O1A1Ixp33_ASAP7_75t_SL U19934 ( .A1(n32660), .A2(n19002), .B(n32654), .C(
        n22069), .Y(ic_data[28]) );
  A2O1A1Ixp33_ASAP7_75t_SL U19935 ( .A1(n32660), .A2(n19002), .B(n32630), .C(
        n22068), .Y(ic_data[16]) );
  A2O1A1Ixp33_ASAP7_75t_SL U19936 ( .A1(n32660), .A2(n19002), .B(n32624), .C(
        n22067), .Y(ic_data[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U19937 ( .A1(n19002), .A2(n32660), .B(n32604), .C(
        n21785), .Y(ic_data[3]) );
  A2O1A1Ixp33_ASAP7_75t_SL U19938 ( .A1(n32628), .A2(n19002), .B(n32543), .C(
        n22066), .Y(it_data[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL U19939 ( .A1(n32162), .A2(n19002), .B(n32158), .C(
        n22060), .Y(rf_addr_w[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U19940 ( .A1(n32162), .A2(n19002), .B(n32157), .C(
        n22059), .Y(rf_addr_w[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U19941 ( .A1(irqctrl0_r_ILEVEL__2_), .A2(n19002), 
        .B(n29400), .C(n19002), .Y(n22057) );
  O2A1O1Ixp5_ASAP7_75t_SL U19942 ( .A1(timer0_N63), .A2(timer0_N64), .B(n19002), .C(n21770), .Y(n24367) );
  A2O1A1Ixp33_ASAP7_75t_SL U19943 ( .A1(n22373), .A2(n19002), .B(n25314), .C(
        n22055), .Y(n30249) );
  A2O1A1Ixp33_ASAP7_75t_SL U19944 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__19_), 
        .A2(n31824), .B(n24680), .C(n19002), .Y(n20550) );
  A2O1A1Ixp33_ASAP7_75t_SL U19945 ( .A1(n19002), .A2(n24585), .B(n31687), .C(
        n20550), .Y(n31682) );
  A2O1A1Ixp33_ASAP7_75t_SL U19946 ( .A1(n19002), .A2(n22214), .B(n23213), .C(
        n21560), .Y(n23211) );
  A2O1A1Ixp33_ASAP7_75t_SL U19947 ( .A1(n22373), .A2(n19002), .B(n25302), .C(
        n19002), .Y(n22053) );
  A2O1A1Ixp33_ASAP7_75t_SL U19948 ( .A1(u0_0_leon3x0_p0_divi[49]), .A2(n22373), 
        .B(n22053), .C(n19002), .Y(n30312) );
  A2O1A1Ixp33_ASAP7_75t_SL U19949 ( .A1(n31266), .A2(n19002), .B(n22051), .C(
        n19002), .Y(n30562) );
  A2O1A1Ixp33_ASAP7_75t_SL U19950 ( .A1(n27501), .A2(n19002), .B(n22050), .C(
        n19002), .Y(n27508) );
  A2O1A1Ixp33_ASAP7_75t_SL U19951 ( .A1(mult_x_1196_n323), .A2(n19002), .B(
        n22049), .C(n19002), .Y(mult_x_1196_n228) );
  A2O1A1Ixp33_ASAP7_75t_SL U19952 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[5]), .B(n32353), .C(n20176), .Y(n32408)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U19953 ( .A1(n32290), .A2(n19002), .B(n32150), .C(
        n19002), .Y(n22048) );
  A2O1A1Ixp33_ASAP7_75t_SL U19954 ( .A1(n32427), .A2(n19002), .B(n22048), .C(
        n19002), .Y(n32388) );
  A2O1A1Ixp33_ASAP7_75t_SL U19955 ( .A1(uart1_r_TRADDR__4_), .A2(n19002), .B(
        uart1_r_TRADDR__2_), .C(n19002), .Y(n22047) );
  A2O1A1Ixp33_ASAP7_75t_SL U19956 ( .A1(u0_0_leon3x0_p0_divi[26]), .A2(n19002), 
        .B(n24630), .C(n19002), .Y(n22046) );
  A2O1A1Ixp33_ASAP7_75t_SL U19957 ( .A1(u0_0_leon3x0_p0_divi[20]), .A2(n19002), 
        .B(n24630), .C(n19002), .Y(n22045) );
  A2O1A1Ixp33_ASAP7_75t_SL U19958 ( .A1(n22481), .A2(n22412), .B(
        mult_x_1196_n2771), .C(n19002), .Y(n22042) );
  A2O1A1Ixp33_ASAP7_75t_SL U19959 ( .A1(n24043), .A2(n19002), .B(n22041), .C(
        n19002), .Y(mult_x_1196_n2153) );
  A2O1A1Ixp33_ASAP7_75t_SL U19960 ( .A1(n4824), .A2(n19002), .B(n4821), .C(
        n19002), .Y(n22040) );
  A2O1A1Ixp33_ASAP7_75t_SL U19961 ( .A1(timer0_r_SCALER__7_), .A2(n31245), .B(
        n21982), .C(n19002), .Y(n21983) );
  A2O1A1Ixp33_ASAP7_75t_SL U19962 ( .A1(n4775), .A2(n19002), .B(n21984), .C(
        n19002), .Y(n21985) );
  A2O1A1Ixp33_ASAP7_75t_SL U19963 ( .A1(irqctrl0_r_IFORCE__0__7_), .A2(n31251), 
        .B(n21985), .C(n19002), .Y(n21986) );
  A2O1A1Ixp33_ASAP7_75t_SL U19964 ( .A1(n2851), .A2(n19002), .B(n30983), .C(
        n21986), .Y(n21987) );
  A2O1A1Ixp33_ASAP7_75t_SL U19965 ( .A1(n31237), .A2(timer0_r_RELOAD__7_), .B(
        n21987), .C(n19002), .Y(n21988) );
  A2O1A1Ixp33_ASAP7_75t_SL U19966 ( .A1(n31216), .A2(uart1_r_RHOLD__3__7_), 
        .B(n21992), .C(n19002), .Y(n21993) );
  A2O1A1Ixp33_ASAP7_75t_SL U19967 ( .A1(uart1_r_RHOLD__31__7_), .A2(n31221), 
        .B(n21997), .C(n19002), .Y(n21998) );
  A2O1A1Ixp33_ASAP7_75t_SL U19968 ( .A1(n31213), .A2(uart1_r_RHOLD__15__7_), 
        .B(n22002), .C(n19002), .Y(n22003) );
  A2O1A1Ixp33_ASAP7_75t_SL U19969 ( .A1(n31208), .A2(uart1_r_RHOLD__19__7_), 
        .B(n22007), .C(n19002), .Y(n22008) );
  A2O1A1Ixp33_ASAP7_75t_SL U19970 ( .A1(uart1_r_RHOLD__6__7_), .A2(n31226), 
        .B(n22014), .C(n19002), .Y(n22015) );
  A2O1A1Ixp33_ASAP7_75t_SL U19971 ( .A1(n31230), .A2(uart1_r_RHOLD__27__7_), 
        .B(n22019), .C(n19002), .Y(n22020) );
  A2O1A1Ixp33_ASAP7_75t_SL U19972 ( .A1(n31200), .A2(uart1_r_RHOLD__5__7_), 
        .B(n22024), .C(n19002), .Y(n22025) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19973 ( .A1(uart1_r_RHOLD__14__7_), .A2(n31203), 
        .B(n22010), .C(n19002), .D(n22026), .Y(n22027) );
  A2O1A1Ixp33_ASAP7_75t_SL U19974 ( .A1(n30872), .A2(n19002), .B(n30871), .C(
        n19002), .Y(n22029) );
  A2O1A1Ixp33_ASAP7_75t_SL U19975 ( .A1(n1626), .A2(n19002), .B(n31953), .C(
        n19002), .Y(n22030) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19976 ( .A1(n30870), .A2(n22028), .B(n22029), 
        .C(n19002), .D(n22030), .Y(n22031) );
  A2O1A1Ixp33_ASAP7_75t_SL U19977 ( .A1(n31241), .A2(uart1_r_RHOLD__24__7_), 
        .B(n22033), .C(n19002), .Y(n22034) );
  A2O1A1Ixp33_ASAP7_75t_SL U19978 ( .A1(n32004), .A2(n19002), .B(n30874), .C(
        n19002), .Y(n22037) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19979 ( .A1(n32003), .A2(sr1_r_MCFG1__ROMWWS__3_), .B(n31849), .C(n19002), .D(n22037), .Y(n22038) );
  A2O1A1Ixp33_ASAP7_75t_SL U19980 ( .A1(n31973), .A2(n19002), .B(n22036), .C(
        n22038), .Y(n22039) );
  A2O1A1Ixp33_ASAP7_75t_SL U19981 ( .A1(n31954), .A2(n22035), .B(n22039), .C(
        n19002), .Y(n4779) );
  A2O1A1Ixp33_ASAP7_75t_SL U19982 ( .A1(n30738), .A2(apbi[4]), .B(n24695), .C(
        n19002), .Y(n21978) );
  A2O1A1Ixp33_ASAP7_75t_SL U19983 ( .A1(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__1_), 
        .A2(n19002), .B(n29883), .C(n19002), .Y(n21974) );
  A2O1A1Ixp33_ASAP7_75t_SL U19984 ( .A1(n30211), .A2(n21974), .B(n30706), .C(
        n19002), .Y(n21975) );
  A2O1A1Ixp33_ASAP7_75t_SL U19985 ( .A1(n4752), .A2(n19002), .B(n21976), .C(
        n19002), .Y(n21977) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U19986 ( .A1(n24649), .A2(
        u0_0_leon3x0_p0_iu_r_X__CTRL__TT__1_), .B(n21975), .C(n19002), .D(
        n21977), .Y(n4751) );
  A2O1A1Ixp33_ASAP7_75t_SL U19987 ( .A1(n22393), .A2(n19002), .B(n32992), .C(
        n19002), .Y(n21972) );
  A2O1A1Ixp33_ASAP7_75t_SL U19988 ( .A1(n32705), .A2(n19002), .B(n31949), .C(
        n19002), .Y(n21973) );
  A2O1A1Ixp33_ASAP7_75t_SL U19989 ( .A1(n21972), .A2(n19002), .B(n21973), .C(
        n19002), .Y(n4747) );
  A2O1A1Ixp33_ASAP7_75t_SL U19990 ( .A1(n30026), .A2(n19002), .B(n31045), .C(
        n19002), .Y(n21962) );
  A2O1A1Ixp33_ASAP7_75t_SL U19991 ( .A1(n22420), .A2(n19002), .B(n28330), .C(
        n31422), .Y(n21958) );
  A2O1A1Ixp33_ASAP7_75t_SL U19992 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[14]), 
        .B(n21958), .C(n19002), .Y(n21959) );
  A2O1A1Ixp33_ASAP7_75t_SL U19993 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_14_), .B(n21961), .C(n19002), .Y(n4656) );
  A2O1A1Ixp33_ASAP7_75t_SL U19994 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__15_), .A2(n19002), .B(n24495), .C(
        n19002), .Y(n21955) );
  A2O1A1Ixp33_ASAP7_75t_SL U19995 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_A__IMM__25_), .C(n19002), .Y(n21956) );
  A2O1A1Ixp33_ASAP7_75t_SL U19996 ( .A1(n29805), .A2(n24647), .B(n21953), .C(
        n19002), .Y(n21954) );
  A2O1A1Ixp33_ASAP7_75t_SL U19997 ( .A1(n31343), .A2(n19002), .B(n29806), .C(
        n21954), .Y(n4627) );
  O2A1O1Ixp5_ASAP7_75t_SL U19998 ( .A1(n29803), .A2(n32110), .B(n19002), .C(
        n21952), .Y(n21953) );
  A2O1A1Ixp33_ASAP7_75t_SL U19999 ( .A1(n22420), .A2(n19002), .B(n28282), .C(
        n31422), .Y(n21948) );
  A2O1A1Ixp33_ASAP7_75t_SL U20000 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[28]), 
        .B(n21948), .C(n19002), .Y(n21949) );
  A2O1A1Ixp33_ASAP7_75t_SL U20001 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_28_), .B(n21951), .C(n19002), .Y(n4589) );
  A2O1A1Ixp33_ASAP7_75t_SL U20002 ( .A1(n24646), .A2(n19002), .B(n18844), .C(
        n19002), .Y(n21947) );
  A2O1A1Ixp33_ASAP7_75t_SL U20003 ( .A1(n28713), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n21938) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20004 ( .A1(n30644), .A2(n28714), .B(n21938), 
        .C(n19002), .D(n21941), .Y(n21942) );
  A2O1A1Ixp33_ASAP7_75t_SL U20005 ( .A1(n30645), .A2(n19002), .B(n30385), .C(
        n21942), .Y(n21943) );
  A2O1A1Ixp33_ASAP7_75t_SL U20006 ( .A1(n31055), .A2(n22432), .B(n21943), .C(
        n19002), .Y(n21944) );
  A2O1A1Ixp33_ASAP7_75t_SL U20007 ( .A1(n28715), .A2(n19002), .B(n22379), .C(
        n19002), .Y(n21946) );
  A2O1A1Ixp33_ASAP7_75t_SL U20008 ( .A1(u0_0_leon3x0_p0_c0mmu_dcache0_r_MEXC_), 
        .A2(n19002), .B(n21935), .C(n19002), .Y(n21936) );
  A2O1A1Ixp33_ASAP7_75t_SL U20009 ( .A1(n28353), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21932) );
  A2O1A1Ixp33_ASAP7_75t_SL U20010 ( .A1(n23980), .A2(n19002), .B(n31677), .C(
        n19002), .Y(n21933) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20011 ( .A1(n29114), .A2(n24517), .B(n21932), 
        .C(n19002), .D(n21933), .Y(n4474) );
  A2O1A1Ixp33_ASAP7_75t_SL U20012 ( .A1(n22422), .A2(n19002), .B(n27177), .C(
        n19002), .Y(n21930) );
  A2O1A1Ixp33_ASAP7_75t_SL U20013 ( .A1(n28337), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21931) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20014 ( .A1(n31662), .A2(n22837), .B(n21930), 
        .C(n19002), .D(n21931), .Y(n4452) );
  A2O1A1Ixp33_ASAP7_75t_SL U20015 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__9_), .A2(
        n22429), .B(n19749), .C(n19002), .Y(n19750) );
  A2O1A1Ixp33_ASAP7_75t_SL U20016 ( .A1(n19002), .A2(n30446), .B(n30391), .C(
        n19753), .Y(n19754) );
  A2O1A1Ixp33_ASAP7_75t_SL U20017 ( .A1(n22427), .A2(n19002), .B(n30736), .C(
        n21929), .Y(n4436) );
  A2O1A1Ixp33_ASAP7_75t_SL U20018 ( .A1(n22420), .A2(n19002), .B(n29906), .C(
        n31422), .Y(n21925) );
  A2O1A1Ixp33_ASAP7_75t_SL U20019 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[6]), 
        .B(n21925), .C(n19002), .Y(n21926) );
  A2O1A1Ixp33_ASAP7_75t_SL U20020 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_6_), .B(n21928), .C(n19002), .Y(n4378) );
  A2O1A1Ixp33_ASAP7_75t_SL U20021 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[6]), .C(n21421), .Y(n4373) );
  A2O1A1Ixp33_ASAP7_75t_SL U20022 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[59]), .C(n21694), .Y(n4332) );
  A2O1A1Ixp33_ASAP7_75t_SL U20023 ( .A1(n32125), .A2(n19002), .B(n21922), .C(
        n32129), .Y(u0_0_leon3x0_p0_c0mmu_icache0_v_HOLDN_) );
  A2O1A1Ixp33_ASAP7_75t_SL U20024 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_div0_v_ZERO2_), .B(n24657), .C(n21680), .Y(n4311) );
  A2O1A1Ixp33_ASAP7_75t_SL U20025 ( .A1(n19002), .A2(n22427), .B(n21417), .C(
        n21418), .Y(n4303) );
  A2O1A1Ixp33_ASAP7_75t_SL U20026 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), .B(n24654), .C(n21674), .Y(
        n4175) );
  A2O1A1Ixp33_ASAP7_75t_SL U20027 ( .A1(n19002), .A2(n22378), .B(n31947), .C(
        n21411), .Y(n4147) );
  A2O1A1Ixp33_ASAP7_75t_SL U20028 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__20_), .B(n22377), .C(n21671), .Y(
        n4101) );
  A2O1A1Ixp33_ASAP7_75t_SL U20029 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__RD__4_), .B(n22377), .C(n21409), .Y(
        n4055) );
  A2O1A1Ixp33_ASAP7_75t_SL U20030 ( .A1(n30306), .A2(n19002), .B(n22414), .C(
        n21908), .Y(n21909) );
  A2O1A1Ixp33_ASAP7_75t_SL U20031 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__18_), .B(n21909), .C(n19002), .Y(n3997)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20032 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__16_), .C(n21906), .Y(n3988) );
  A2O1A1Ixp33_ASAP7_75t_SL U20033 ( .A1(n22427), .A2(n19002), .B(n30799), .C(
        n21905), .Y(n3967) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20034 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TT__6_), 
        .A2(u0_0_leon3x0_p0_iu_r_W__S__TT__7_), .B(n19002), .C(n21901), .Y(
        n21902) );
  A2O1A1Ixp33_ASAP7_75t_SL U20035 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_A__CTRL__RETT_), .C(n21660), .Y(n3883) );
  A2O1A1Ixp33_ASAP7_75t_SL U20036 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__11_), .C(n21659), .Y(n3844) );
  A2O1A1Ixp33_ASAP7_75t_SL U20037 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__15_), .C(n21658), .Y(n3840) );
  A2O1A1Ixp33_ASAP7_75t_SL U20038 ( .A1(n22427), .A2(n19002), .B(n30613), .C(
        n21898), .Y(n3828) );
  A2O1A1Ixp33_ASAP7_75t_SL U20039 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_muli[7]), .C(n21656), .Y(n3820) );
  A2O1A1Ixp33_ASAP7_75t_SL U20040 ( .A1(n19002), .A2(n24646), .B(n30244), .C(
        n21390), .Y(n3786) );
  A2O1A1Ixp33_ASAP7_75t_SL U20041 ( .A1(n19002), .A2(n24646), .B(n30240), .C(
        n21650), .Y(n3784) );
  A2O1A1Ixp33_ASAP7_75t_SL U20042 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__1_), .B(n22377), .C(n21166), .Y(
        n3754) );
  A2O1A1Ixp33_ASAP7_75t_SL U20043 ( .A1(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__29_), .A2(n19002), .B(n24655), .C(
        n21889), .Y(n3741) );
  A2O1A1Ixp33_ASAP7_75t_SL U20044 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_r_A__DIVSTART_), .B(n23229), .C(n21647), .Y(n3717)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20045 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__5_), .B(n22428), .C(n21646), .Y(
        n3689) );
  A2O1A1Ixp33_ASAP7_75t_SL U20046 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[35]), .C(n21642), .Y(n3448) );
  A2O1A1Ixp33_ASAP7_75t_SL U20047 ( .A1(n22427), .A2(n19002), .B(rf_di_w[5]), 
        .C(n21872), .Y(n3381) );
  A2O1A1Ixp33_ASAP7_75t_SL U20048 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_dci[1]), .C(n20967), .Y(n3320) );
  A2O1A1Ixp33_ASAP7_75t_SL U20049 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[57]), 
        .B(n22428), .C(n21639), .Y(n3288) );
  A2O1A1Ixp33_ASAP7_75t_SL U20050 ( .A1(n19002), .A2(n22427), .B(rf_di_w[28]), 
        .C(n20620), .Y(n3268) );
  A2O1A1Ixp33_ASAP7_75t_SL U20051 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[38]), 
        .B(n24653), .C(n19309), .Y(n3174) );
  A2O1A1Ixp33_ASAP7_75t_SL U20052 ( .A1(n30417), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21865) );
  A2O1A1Ixp33_ASAP7_75t_SL U20053 ( .A1(n30418), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21866) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20054 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__5_), 
        .A2(n31403), .B(n21865), .C(n19002), .D(n21866), .Y(n3149) );
  A2O1A1Ixp33_ASAP7_75t_SL U20055 ( .A1(n30247), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21863) );
  A2O1A1Ixp33_ASAP7_75t_SL U20056 ( .A1(n30248), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21864) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20057 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__25_), 
        .A2(n31403), .B(n21863), .C(n19002), .D(n21864), .Y(n3139) );
  A2O1A1Ixp33_ASAP7_75t_SL U20058 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_dci[5]), .C(n20785), .Y(n3129) );
  A2O1A1Ixp33_ASAP7_75t_SL U20059 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[28]), .C(n21862), .Y(n3119) );
  A2O1A1Ixp33_ASAP7_75t_SL U20060 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[16]), .C(n21858), .Y(n3095) );
  A2O1A1Ixp33_ASAP7_75t_SL U20061 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[15]), .C(n21856), .Y(n3093) );
  A2O1A1Ixp33_ASAP7_75t_SL U20062 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[14]), .C(n21854), .Y(n3091) );
  A2O1A1Ixp33_ASAP7_75t_SL U20063 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[11]), .C(n21625), .Y(n3072) );
  A2O1A1Ixp33_ASAP7_75t_SL U20064 ( .A1(n22422), .A2(n19002), .B(n28357), .C(
        n19002), .Y(n21849) );
  A2O1A1Ixp33_ASAP7_75t_SL U20065 ( .A1(n29691), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21850) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20066 ( .A1(n31662), .A2(n22449), .B(n21849), 
        .C(n19002), .D(n21850), .Y(n3035) );
  A2O1A1Ixp33_ASAP7_75t_SL U20067 ( .A1(n19002), .A2(n22427), .B(rf_di_w[8]), 
        .C(n21624), .Y(n3028) );
  A2O1A1Ixp33_ASAP7_75t_SL U20068 ( .A1(n22422), .A2(n19002), .B(n28328), .C(
        n19002), .Y(n21847) );
  A2O1A1Ixp33_ASAP7_75t_SL U20069 ( .A1(n27223), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21848) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20070 ( .A1(n31662), .A2(n23964), .B(n21847), 
        .C(n19002), .D(n21848), .Y(n3019) );
  A2O1A1Ixp33_ASAP7_75t_SL U20071 ( .A1(n22422), .A2(n19002), .B(n29022), .C(
        n19002), .Y(n21845) );
  A2O1A1Ixp33_ASAP7_75t_SL U20072 ( .A1(n28298), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21846) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20073 ( .A1(n31662), .A2(n22968), .B(n21845), 
        .C(n19002), .D(n21846), .Y(n3001) );
  A2O1A1Ixp33_ASAP7_75t_SL U20074 ( .A1(n32730), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n21843) );
  A2O1A1Ixp33_ASAP7_75t_SL U20075 ( .A1(n32733), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n21844) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20076 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__0_), .B(n21843), .C(n19002), .D(
        n21844), .Y(n2997) );
  A2O1A1Ixp33_ASAP7_75t_SL U20077 ( .A1(n32616), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n21841) );
  A2O1A1Ixp33_ASAP7_75t_SL U20078 ( .A1(n31971), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n21842) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20079 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__9_), .B(n21841), .C(n19002), .D(
        n21842), .Y(n2991) );
  A2O1A1Ixp33_ASAP7_75t_SL U20080 ( .A1(n22405), .A2(n19002), .B(n21839), .C(
        n32550), .Y(n21840) );
  A2O1A1Ixp33_ASAP7_75t_SL U20081 ( .A1(n19002), .A2(n31198), .B(
        sr1_r_MCFG2__RMW_), .C(n21128), .Y(n2915) );
  A2O1A1Ixp33_ASAP7_75t_SL U20082 ( .A1(n28167), .A2(uart1_uarto_SCALER__8_), 
        .B(n22419), .C(n19002), .Y(n21124) );
  A2O1A1Ixp33_ASAP7_75t_SL U20083 ( .A1(n19002), .A2(n24633), .B(
        uart1_r_RFIFOIRQEN_), .C(n21345), .Y(n2871) );
  A2O1A1Ixp33_ASAP7_75t_SL U20084 ( .A1(n19002), .A2(n24633), .B(
        uart1_r_PAREN_), .C(n21344), .Y(n2868) );
  A2O1A1Ixp33_ASAP7_75t_SL U20085 ( .A1(n29383), .A2(n19002), .B(apbi[12]), 
        .C(n21838), .Y(n2849) );
  A2O1A1Ixp33_ASAP7_75t_SL U20086 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__31_), .C(n21836), .Y(n2813) );
  A2O1A1Ixp33_ASAP7_75t_SL U20087 ( .A1(n24646), .A2(n19002), .B(n32185), .C(
        n19002), .Y(n21832) );
  A2O1A1Ixp33_ASAP7_75t_SL U20088 ( .A1(n24660), .A2(
        u0_0_leon3x0_p0_iu_r_A__RFA1__6_), .B(n21832), .C(n19002), .Y(n2774)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20089 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__30_), .C(n21343), .Y(n2758) );
  A2O1A1Ixp33_ASAP7_75t_SL U20090 ( .A1(n19002), .A2(n22428), .B(n30435), .C(
        n21605), .Y(n2749) );
  A2O1A1Ixp33_ASAP7_75t_SL U20091 ( .A1(n22428), .A2(n19002), .B(rf_di_w[3]), 
        .C(n21830), .Y(n2740) );
  A2O1A1Ixp33_ASAP7_75t_SL U20092 ( .A1(n19002), .A2(n24646), .B(rf_di_w[4]), 
        .C(n21600), .Y(n2728) );
  A2O1A1Ixp33_ASAP7_75t_SL U20093 ( .A1(n22422), .A2(n19002), .B(n29924), .C(
        n19002), .Y(n21827) );
  A2O1A1Ixp33_ASAP7_75t_SL U20094 ( .A1(n29926), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21828) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20095 ( .A1(n31662), .A2(n23960), .B(n21827), 
        .C(n19002), .D(n21828), .Y(n2683) );
  A2O1A1Ixp33_ASAP7_75t_SL U20096 ( .A1(n22422), .A2(n19002), .B(n28322), .C(
        n19002), .Y(n21823) );
  A2O1A1Ixp33_ASAP7_75t_SL U20097 ( .A1(n28320), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21824) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20098 ( .A1(n31662), .A2(n24571), .B(n21823), 
        .C(n19002), .D(n21824), .Y(n2633) );
  A2O1A1Ixp33_ASAP7_75t_SL U20099 ( .A1(n22427), .A2(n19002), .B(rf_di_w[18]), 
        .C(n21821), .Y(n2572) );
  A2O1A1Ixp33_ASAP7_75t_SL U20100 ( .A1(n22422), .A2(n19002), .B(n28306), .C(
        n19002), .Y(n21819) );
  A2O1A1Ixp33_ASAP7_75t_SL U20101 ( .A1(n28312), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21820) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20102 ( .A1(n31662), .A2(n23969), .B(n21819), 
        .C(n19002), .D(n21820), .Y(n2562) );
  A2O1A1Ixp33_ASAP7_75t_SL U20103 ( .A1(n19002), .A2(n27513), .B(n29987), .C(
        n21585), .Y(n2461) );
  A2O1A1Ixp33_ASAP7_75t_SL U20104 ( .A1(n22405), .A2(n19002), .B(n21808), .C(
        n32556), .Y(n21809) );
  A2O1A1Ixp33_ASAP7_75t_SL U20105 ( .A1(n19002), .A2(n27018), .B(n30654), .C(
        n20286), .Y(n20287) );
  A2O1A1Ixp33_ASAP7_75t_SL U20106 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__20_), 
        .A2(n30655), .B(n20287), .C(n19002), .Y(n2278) );
  A2O1A1Ixp33_ASAP7_75t_SL U20107 ( .A1(n22422), .A2(n19002), .B(n29792), .C(
        n19002), .Y(n21806) );
  A2O1A1Ixp33_ASAP7_75t_SL U20108 ( .A1(n29793), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21807) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20109 ( .A1(n31662), .A2(n23002), .B(n21806), 
        .C(n19002), .D(n21807), .Y(n2275) );
  A2O1A1Ixp33_ASAP7_75t_SL U20110 ( .A1(dataout[0]), .A2(n19002), .B(n21802), 
        .C(n19002), .Y(n21803) );
  A2O1A1Ixp33_ASAP7_75t_SL U20111 ( .A1(dataout[8]), .A2(n19002), .B(n21799), 
        .C(n19002), .Y(n21800) );
  A2O1A1Ixp33_ASAP7_75t_SL U20112 ( .A1(n32586), .A2(n19002), .B(n32585), .C(
        n19002), .Y(n21792) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20113 ( .A1(n32590), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__10_), .B(n21792), .C(n19002), 
        .D(n21795), .Y(n21796) );
  A2O1A1Ixp33_ASAP7_75t_SL U20114 ( .A1(n32660), .A2(n19002), .B(n32661), .C(
        n21791), .Y(ic_data[31]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20115 ( .A1(n32660), .A2(n19002), .B(n32652), .C(
        n21790), .Y(ic_data[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20116 ( .A1(n32660), .A2(n19002), .B(n32650), .C(
        n21789), .Y(ic_data[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20117 ( .A1(n32660), .A2(n19002), .B(n32648), .C(
        n21788), .Y(ic_data[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20118 ( .A1(n32660), .A2(n19002), .B(n32646), .C(
        n21787), .Y(ic_data[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20119 ( .A1(n32660), .A2(n19002), .B(n32632), .C(
        n21786), .Y(ic_data[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20120 ( .A1(n19002), .A2(n32660), .B(n32606), .C(
        n20428), .Y(ic_data[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20121 ( .A1(n19002), .A2(n32660), .B(n32602), .C(
        n21575), .Y(ic_data[2]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20122 ( .A1(n32348), .A2(n19002), .B(n32426), .C(
        n19002), .Y(n21779) );
  A2O1A1Ixp33_ASAP7_75t_SL U20123 ( .A1(n21779), .A2(n19002), .B(n21782), .C(
        n19002), .Y(n21783) );
  A2O1A1Ixp33_ASAP7_75t_SL U20124 ( .A1(n32418), .A2(n19002), .B(n32232), .C(
        n19002), .Y(n21776) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20125 ( .A1(n32239), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__30_), .B(n33067), .C(n19002), .D(
        n21776), .Y(n21777) );
  A2O1A1Ixp33_ASAP7_75t_SL U20126 ( .A1(n22377), .A2(n19002), .B(n21774), .C(
        n21775), .Y(rf_addr_b[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20127 ( .A1(n19002), .A2(n32166), .B(n22377), .C(
        n21568), .Y(rf_addr_b[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20128 ( .A1(n32162), .A2(n19002), .B(n32159), .C(
        n21773), .Y(rf_addr_w[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20129 ( .A1(n28829), .A2(n19002), .B(n29909), .C(
        n25871), .Y(n21772) );
  A2O1A1Ixp33_ASAP7_75t_SL U20130 ( .A1(n25874), .A2(n19002), .B(n21772), .C(
        n19002), .Y(n32307) );
  A2O1A1Ixp33_ASAP7_75t_SL U20131 ( .A1(n19002), .A2(n29468), .B(n19820), .C(
        n29727), .Y(n30704) );
  A2O1A1Ixp33_ASAP7_75t_SL U20132 ( .A1(n22373), .A2(n19002), .B(n25307), .C(
        n19002), .Y(n21769) );
  A2O1A1Ixp33_ASAP7_75t_SL U20133 ( .A1(u0_0_leon3x0_p0_divi[52]), .A2(n22373), 
        .B(n21769), .C(n19002), .Y(n30282) );
  A2O1A1Ixp33_ASAP7_75t_SL U20134 ( .A1(n31263), .A2(n19002), .B(n31573), .C(
        n19002), .Y(n21768) );
  A2O1A1Ixp33_ASAP7_75t_SL U20135 ( .A1(n22373), .A2(n19002), .B(n25304), .C(
        n21767), .Y(n30302) );
  A2O1A1Ixp33_ASAP7_75t_SL U20136 ( .A1(n32503), .A2(n19002), .B(n21762), .C(
        n19002), .Y(n21763) );
  A2O1A1Ixp33_ASAP7_75t_SL U20137 ( .A1(n32491), .A2(n19002), .B(n32490), .C(
        n19002), .Y(n21764) );
  A2O1A1Ixp33_ASAP7_75t_SL U20138 ( .A1(n21763), .A2(n19002), .B(n21764), .C(
        n19002), .Y(n21765) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20139 ( .A1(n1724), .A2(sr1_r_BUSW__1_), .B(
        n19002), .C(sr1_r_BUSW__0_), .Y(n21761) );
  A2O1A1Ixp33_ASAP7_75t_SL U20140 ( .A1(n21761), .A2(n19002), .B(n22433), .C(
        n19002), .Y(n32906) );
  A2O1A1Ixp33_ASAP7_75t_SL U20141 ( .A1(n24642), .A2(n19002), .B(n32329), .C(
        n21760), .Y(n32400) );
  A2O1A1Ixp33_ASAP7_75t_SL U20142 ( .A1(n22373), .A2(n19002), .B(n25321), .C(
        n19002), .Y(n21759) );
  A2O1A1Ixp33_ASAP7_75t_SL U20143 ( .A1(u0_0_leon3x0_p0_divi[60]), .A2(n22373), 
        .B(n21759), .C(n19002), .Y(n25897) );
  A2O1A1Ixp33_ASAP7_75t_SL U20144 ( .A1(n22468), .A2(n19002), .B(n21758), .C(
        n18988), .Y(mult_x_1196_n525) );
  A2O1A1Ixp33_ASAP7_75t_SL U20145 ( .A1(mult_x_1196_n387), .A2(n19002), .B(
        mult_x_1196_n361), .C(n19002), .Y(n21757) );
  A2O1A1Ixp33_ASAP7_75t_SL U20146 ( .A1(n22376), .A2(n19002), .B(n31423), .C(
        n21756), .Y(n29012) );
  A2O1A1Ixp33_ASAP7_75t_SL U20147 ( .A1(u0_0_leon3x0_p0_divi[28]), .A2(n19002), 
        .B(n24630), .C(n19002), .Y(n21754) );
  A2O1A1Ixp33_ASAP7_75t_SL U20148 ( .A1(n18364), .A2(n24040), .B(
        mult_x_1196_n2737), .C(n19002), .Y(n21749) );
  A2O1A1Ixp33_ASAP7_75t_SL U20149 ( .A1(mult_x_1196_n2813), .A2(n19002), .B(
        n22251), .C(n19002), .Y(n21748) );
  A2O1A1Ixp33_ASAP7_75t_SL U20150 ( .A1(n19002), .A2(n21747), .B(n21748), .C(
        n19002), .Y(n23301) );
  A2O1A1Ixp33_ASAP7_75t_SL U20151 ( .A1(mult_x_1196_n2814), .A2(n19002), .B(
        n24034), .C(n19002), .Y(n21747) );
  A2O1A1Ixp33_ASAP7_75t_SL U20152 ( .A1(uart1_r_RHOLD__19__4_), .A2(n31208), 
        .B(n21490), .C(n19002), .Y(n21491) );
  A2O1A1Ixp33_ASAP7_75t_SL U20153 ( .A1(uart1_r_RHOLD__15__4_), .A2(n31213), 
        .B(n21495), .C(n19002), .Y(n21496) );
  A2O1A1Ixp33_ASAP7_75t_SL U20154 ( .A1(n31205), .A2(uart1_r_RHOLD__16__4_), 
        .B(n21500), .C(n19002), .Y(n21501) );
  O2A1O1Ixp5_ASAP7_75t_SL U20155 ( .A1(n21485), .A2(n21486), .B(n19002), .C(
        n21517), .Y(n21518) );
  A2O1A1Ixp33_ASAP7_75t_SL U20156 ( .A1(irqctrl0_r_IFORCE__0__4_), .A2(n31251), 
        .B(n21529), .C(n19002), .Y(n21530) );
  A2O1A1Ixp33_ASAP7_75t_SL U20157 ( .A1(timer0_vtimers_1__RELOAD__4_), .A2(
        n31956), .B(n21532), .C(n19002), .Y(n21533) );
  A2O1A1Ixp33_ASAP7_75t_SL U20158 ( .A1(uart1_r_RHOLD__0__4_), .A2(n31242), 
        .B(n21537), .C(n19002), .Y(n21538) );
  A2O1A1Ixp33_ASAP7_75t_SL U20159 ( .A1(n31954), .A2(n21539), .B(n31849), .C(
        n19002), .Y(n4768) );
  A2O1A1Ixp33_ASAP7_75t_SL U20160 ( .A1(n29663), .A2(n21740), .B(n29662), .C(
        n19002), .Y(n21741) );
  A2O1A1Ixp33_ASAP7_75t_SL U20161 ( .A1(n21741), .A2(n19002), .B(n29661), .C(
        n19002), .Y(n21742) );
  A2O1A1Ixp33_ASAP7_75t_SL U20162 ( .A1(n29662), .A2(n19002), .B(n29658), .C(
        n19002), .Y(n21743) );
  A2O1A1Ixp33_ASAP7_75t_SL U20163 ( .A1(n32669), .A2(n19002), .B(n32677), .C(
        n19002), .Y(n21734) );
  A2O1A1Ixp33_ASAP7_75t_SL U20164 ( .A1(n19002), .A2(n21243), .B(n21245), .C(
        n31756), .Y(n4726) );
  A2O1A1Ixp33_ASAP7_75t_SL U20165 ( .A1(uart1_r_RXF__4_), .A2(n19002), .B(
        uart1_r_RXF__3_), .C(n19002), .Y(n21725) );
  A2O1A1Ixp33_ASAP7_75t_SL U20166 ( .A1(uart1_r_RXF__3_), .A2(uart1_r_RXF__4_), 
        .B(uart1_r_RXF__2_), .C(n19002), .Y(n21726) );
  A2O1A1Ixp33_ASAP7_75t_SL U20167 ( .A1(n21725), .A2(n19002), .B(n21726), .C(
        n19002), .Y(n21727) );
  A2O1A1Ixp33_ASAP7_75t_SL U20168 ( .A1(uart1_r_TSHIFT__0_), .A2(n19002), .B(
        n21728), .C(n19002), .Y(n21729) );
  A2O1A1Ixp33_ASAP7_75t_SL U20169 ( .A1(n24681), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_E__OP1__13_), .C(n19002), .Y(n21722) );
  A2O1A1Ixp33_ASAP7_75t_SL U20170 ( .A1(n31054), .A2(n30490), .B(n21722), .C(
        n19002), .Y(n21723) );
  A2O1A1Ixp33_ASAP7_75t_SL U20171 ( .A1(n31802), .A2(n19002), .B(n21720), .C(
        n19002), .Y(n21721) );
  O2A1O1Ixp33_ASAP7_75t_SL U20172 ( .A1(n21460), .A2(n21461), .B(n19002), .C(
        n30578), .Y(n4641) );
  A2O1A1Ixp33_ASAP7_75t_SL U20173 ( .A1(n29787), .A2(n31868), .B(n21455), .C(
        n19002), .Y(n21456) );
  A2O1A1Ixp33_ASAP7_75t_SL U20174 ( .A1(n19002), .A2(n24541), .B(n29789), .C(
        n21456), .Y(n21457) );
  A2O1A1Ixp33_ASAP7_75t_SL U20175 ( .A1(n22420), .A2(n19002), .B(n29794), .C(
        n31422), .Y(n21716) );
  A2O1A1Ixp33_ASAP7_75t_SL U20176 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[26]), 
        .B(n21716), .C(n19002), .Y(n21717) );
  A2O1A1Ixp33_ASAP7_75t_SL U20177 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_26_), .B(n21719), .C(n19002), .Y(n4619) );
  A2O1A1Ixp33_ASAP7_75t_SL U20178 ( .A1(n22422), .A2(n19002), .B(n28282), .C(
        n19002), .Y(n21714) );
  A2O1A1Ixp33_ASAP7_75t_SL U20179 ( .A1(n29022), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21715) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20180 ( .A1(n31662), .A2(n22906), .B(n21714), 
        .C(n19002), .D(n21715), .Y(n4586) );
  A2O1A1Ixp33_ASAP7_75t_SL U20181 ( .A1(n31641), .A2(n19002), .B(n22397), .C(
        n19002), .Y(n21713) );
  A2O1A1Ixp33_ASAP7_75t_SL U20182 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__5_), 
        .A2(n19002), .B(n22428), .C(n21712), .Y(n4565) );
  A2O1A1Ixp33_ASAP7_75t_SL U20183 ( .A1(n22420), .A2(n19002), .B(n27177), .C(
        n31422), .Y(n21707) );
  A2O1A1Ixp33_ASAP7_75t_SL U20184 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[10]), 
        .B(n21707), .C(n19002), .Y(n21708) );
  A2O1A1Ixp33_ASAP7_75t_SL U20185 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_10_), .B(n21710), .C(n19002), .Y(n4553) );
  A2O1A1Ixp33_ASAP7_75t_SL U20186 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[10]), .C(n21706), .Y(n4548) );
  A2O1A1Ixp33_ASAP7_75t_SL U20187 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_de_icc_0_), .B(n22379), .C(n21437), .Y(n4503) );
  A2O1A1Ixp33_ASAP7_75t_SL U20188 ( .A1(u0_0_leon3x0_p0_iu_r_X__NPC__0_), .A2(
        n25725), .B(n21704), .C(n19002), .Y(n4492) );
  A2O1A1Ixp33_ASAP7_75t_SL U20189 ( .A1(n31404), .A2(n19002), .B(n30459), .C(
        n22379), .Y(n21429) );
  A2O1A1Ixp33_ASAP7_75t_SL U20190 ( .A1(n30613), .A2(n30394), .B(n21429), .C(
        n19002), .Y(n21430) );
  A2O1A1Ixp33_ASAP7_75t_SL U20191 ( .A1(n19002), .A2(n24514), .B(n26369), .C(
        n21430), .Y(n21431) );
  A2O1A1Ixp33_ASAP7_75t_SL U20192 ( .A1(n24428), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__1_), .B(n21431), .C(n19002), .Y(n21432)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20193 ( .A1(n32614), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n21702) );
  A2O1A1Ixp33_ASAP7_75t_SL U20194 ( .A1(n30737), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n21703) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20195 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__8_), .B(n21702), .C(n19002), .D(
        n21703), .Y(n4434) );
  A2O1A1Ixp33_ASAP7_75t_SL U20196 ( .A1(n22422), .A2(n19002), .B(n28330), .C(
        n19002), .Y(n21700) );
  A2O1A1Ixp33_ASAP7_75t_SL U20197 ( .A1(n28328), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21701) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20198 ( .A1(n31662), .A2(n18610), .B(n21700), 
        .C(n19002), .D(n21701), .Y(n4428) );
  A2O1A1Ixp33_ASAP7_75t_SL U20199 ( .A1(n32443), .A2(n19002), .B(n31446), .C(
        n19002), .Y(n21681) );
  A2O1A1Ixp33_ASAP7_75t_SL U20200 ( .A1(n31447), .A2(n19002), .B(n32200), .C(
        n19002), .Y(n21682) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20201 ( .A1(n21681), .A2(n21682), .B(n19002), 
        .C(n31464), .Y(n21683) );
  A2O1A1Ixp33_ASAP7_75t_SL U20202 ( .A1(n31583), .A2(n31455), .B(n21683), .C(
        n19002), .Y(n21684) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20203 ( .A1(n31585), .A2(n32729), .B(n19002), 
        .C(u0_0_leon3x0_p0_dci[2]), .Y(n21687) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20204 ( .A1(n31462), .A2(n31461), .B(n31460), 
        .C(n19002), .D(n21689), .Y(n21690) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20205 ( .A1(n31601), .A2(n21684), .B(n19002), 
        .C(n21691), .Y(n21692) );
  A2O1A1Ixp33_ASAP7_75t_SL U20206 ( .A1(n19002), .A2(n24646), .B(n31545), .C(
        n19737), .Y(n4131) );
  A2O1A1Ixp33_ASAP7_75t_SL U20207 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__0_), 
        .A2(n19002), .B(n24656), .C(n21673), .Y(n4111) );
  A2O1A1Ixp33_ASAP7_75t_SL U20208 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__4_), 
        .A2(n19002), .B(n24655), .C(n21670), .Y(n4053) );
  A2O1A1Ixp33_ASAP7_75t_SL U20209 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_), .B(n24650), .C(n21408), .Y(
        n4028) );
  A2O1A1Ixp33_ASAP7_75t_SL U20210 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_A__CWP__2_), .B(n24651), .C(n21406), .Y(n4016) );
  A2O1A1Ixp33_ASAP7_75t_SL U20211 ( .A1(n19002), .A2(n24646), .B(n29846), .C(
        n21404), .Y(n3971) );
  A2O1A1Ixp33_ASAP7_75t_SL U20212 ( .A1(n22427), .A2(n19002), .B(rf_di_w[6]), 
        .C(n21668), .Y(n3932) );
  A2O1A1Ixp33_ASAP7_75t_SL U20213 ( .A1(n22422), .A2(n19002), .B(n29906), .C(
        n19002), .Y(n21665) );
  A2O1A1Ixp33_ASAP7_75t_SL U20214 ( .A1(n29924), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21666) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20215 ( .A1(n31662), .A2(n23375), .B(n21665), 
        .C(n19002), .D(n21666), .Y(n3929) );
  A2O1A1Ixp33_ASAP7_75t_SL U20216 ( .A1(n22420), .A2(n19002), .B(n29692), .C(
        n31422), .Y(n21661) );
  A2O1A1Ixp33_ASAP7_75t_SL U20217 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[5]), 
        .B(n21661), .C(n19002), .Y(n21662) );
  A2O1A1Ixp33_ASAP7_75t_SL U20218 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_5_), .B(n21664), .C(n19002), .Y(n3919) );
  A2O1A1Ixp33_ASAP7_75t_SL U20219 ( .A1(n22379), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__28_), .C(n21657), .Y(n3836) );
  A2O1A1Ixp33_ASAP7_75t_SL U20220 ( .A1(n19002), .A2(n24646), .B(n31681), .C(
        n21399), .Y(n3832) );
  A2O1A1Ixp33_ASAP7_75t_SL U20221 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__8_), .C(n21655), .Y(n3818) );
  A2O1A1Ixp33_ASAP7_75t_SL U20222 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__18_), .C(n21395), .Y(n3798) );
  A2O1A1Ixp33_ASAP7_75t_SL U20223 ( .A1(n19002), .A2(n24646), .B(n30302), .C(
        n21394), .Y(n3796) );
  A2O1A1Ixp33_ASAP7_75t_SL U20224 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__21_), .C(n21393), .Y(n3792) );
  A2O1A1Ixp33_ASAP7_75t_SL U20225 ( .A1(n19002), .A2(n22427), .B(n30264), .C(
        n21392), .Y(n3790) );
  A2O1A1Ixp33_ASAP7_75t_SL U20226 ( .A1(n19002), .A2(n22427), .B(n30249), .C(
        n21391), .Y(n3788) );
  A2O1A1Ixp33_ASAP7_75t_SL U20227 ( .A1(n19002), .A2(n24909), .B(
        u0_0_leon3x0_p0_div0_r_CNT__0_), .C(n20088), .Y(n3724) );
  O2A1O1Ixp5_ASAP7_75t_SL U20228 ( .A1(n21386), .A2(n21387), .B(n19002), .C(
        n30580), .Y(n21388) );
  A2O1A1Ixp33_ASAP7_75t_SL U20229 ( .A1(n31873), .A2(n19002), .B(n31013), .C(
        n19002), .Y(n21643) );
  A2O1A1Ixp33_ASAP7_75t_SL U20230 ( .A1(n31012), .A2(n19002), .B(n31872), .C(
        n21644), .Y(n21645) );
  A2O1A1Ixp33_ASAP7_75t_SL U20231 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_E__SHCNT__2_), .C(n21645), .Y(n3564) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20232 ( .A1(n32103), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_), .B(n19002), .C(n26826), .Y(
        n19713) );
  A2O1A1Ixp33_ASAP7_75t_SL U20233 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__5_), .B(n24652), .C(n20625), .Y(
        n3454) );
  A2O1A1Ixp33_ASAP7_75t_SL U20234 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[39]), 
        .B(n24653), .C(n21378), .Y(n3416) );
  A2O1A1Ixp33_ASAP7_75t_SL U20235 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[56]), .C(n21373), .Y(n3278) );
  A2O1A1Ixp33_ASAP7_75t_SL U20236 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[54]), .C(n21372), .Y(n3264) );
  A2O1A1Ixp33_ASAP7_75t_SL U20237 ( .A1(u0_0_leon3x0_p0_ici[43]), .A2(n19002), 
        .B(n22428), .C(n21637), .Y(n3224) );
  A2O1A1Ixp33_ASAP7_75t_SL U20238 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[38]), .C(n21369), .Y(n3176) );
  A2O1A1Ixp33_ASAP7_75t_SL U20239 ( .A1(n30407), .A2(n19002), .B(n22414), .C(
        n21634), .Y(n21635) );
  A2O1A1Ixp33_ASAP7_75t_SL U20240 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__6_), .B(n21635), .C(n19002), .Y(n3148)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20241 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[29]), .C(n21632), .Y(n3121) );
  A2O1A1Ixp33_ASAP7_75t_SL U20242 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[7]), .C(n21629), .Y(n3074) );
  A2O1A1Ixp33_ASAP7_75t_SL U20243 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[9]), .C(n21627), .Y(n3073) );
  A2O1A1Ixp33_ASAP7_75t_SL U20244 ( .A1(n22422), .A2(n19002), .B(n28337), .C(
        n19002), .Y(n21622) );
  A2O1A1Ixp33_ASAP7_75t_SL U20245 ( .A1(n28335), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21623) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20246 ( .A1(n31662), .A2(n22394), .B(n21622), 
        .C(n19002), .D(n21623), .Y(n3024) );
  A2O1A1Ixp33_ASAP7_75t_SL U20247 ( .A1(n22427), .A2(n19002), .B(rf_di_w[21]), 
        .C(n21621), .Y(n3013) );
  A2O1A1Ixp33_ASAP7_75t_SL U20248 ( .A1(n19002), .A2(n24646), .B(rf_di_w[23]), 
        .C(n21353), .Y(n3009) );
  A2O1A1Ixp33_ASAP7_75t_SL U20249 ( .A1(n19002), .A2(n24646), .B(rf_di_w[27]), 
        .C(n21136), .Y(n3006) );
  A2O1A1Ixp33_ASAP7_75t_SL U20250 ( .A1(n32608), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n21619) );
  A2O1A1Ixp33_ASAP7_75t_SL U20251 ( .A1(n31948), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n21620) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20252 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__5_), .B(n21619), .C(n19002), .D(
        n21620), .Y(n2995) );
  A2O1A1Ixp33_ASAP7_75t_SL U20253 ( .A1(n19002), .A2(uart1_uarto_SCALER__6_), 
        .B(n21120), .C(n19002), .Y(n21121) );
  A2O1A1Ixp33_ASAP7_75t_SL U20254 ( .A1(n19002), .A2(n29383), .B(apbi[10]), 
        .C(n20295), .Y(n2850) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20255 ( .A1(n32181), .A2(n32180), .B(n19002), 
        .C(n22378), .Y(n21614) );
  A2O1A1Ixp33_ASAP7_75t_SL U20256 ( .A1(n21614), .A2(n19002), .B(n32182), .C(
        n19002), .Y(n21615) );
  A2O1A1Ixp33_ASAP7_75t_SL U20257 ( .A1(n22428), .A2(n19002), .B(rf_di_w[0]), 
        .C(n21610), .Y(n2770) );
  A2O1A1Ixp33_ASAP7_75t_SL U20258 ( .A1(n30213), .A2(n19002), .B(n22414), .C(
        n21607), .Y(n21608) );
  A2O1A1Ixp33_ASAP7_75t_SL U20259 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__30_), .B(n21608), .C(n19002), .Y(n2757)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20260 ( .A1(n22420), .A2(n19002), .B(n28357), .C(
        n31422), .Y(n21601) );
  A2O1A1Ixp33_ASAP7_75t_SL U20261 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[3]), 
        .B(n21601), .C(n19002), .Y(n21602) );
  A2O1A1Ixp33_ASAP7_75t_SL U20262 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_3_), .B(n21604), .C(n19002), .Y(n2744) );
  A2O1A1Ixp33_ASAP7_75t_SL U20263 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[40]), .C(n21335), .Y(n2675) );
  A2O1A1Ixp33_ASAP7_75t_SL U20264 ( .A1(n30361), .A2(n19002), .B(n22414), .C(
        n21597), .Y(n21598) );
  A2O1A1Ixp33_ASAP7_75t_SL U20265 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__13_), .B(n21598), .C(n19002), .Y(n2656)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20266 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[41]), .C(n21334), .Y(n2651) );
  A2O1A1Ixp33_ASAP7_75t_SL U20267 ( .A1(n22422), .A2(n19002), .B(n27264), .C(
        n19002), .Y(n21594) );
  A2O1A1Ixp33_ASAP7_75t_SL U20268 ( .A1(n28322), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21595) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20269 ( .A1(n31662), .A2(n23965), .B(n21594), 
        .C(n19002), .D(n21595), .Y(n2634) );
  A2O1A1Ixp33_ASAP7_75t_SL U20270 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[44]), .C(n21331), .Y(n2627) );
  A2O1A1Ixp33_ASAP7_75t_SL U20271 ( .A1(n19002), .A2(n22421), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__17_), .C(n21330), .Y(n2609) );
  A2O1A1Ixp33_ASAP7_75t_SL U20272 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[46]), .C(n21329), .Y(n2582) );
  A2O1A1Ixp33_ASAP7_75t_SL U20273 ( .A1(n22422), .A2(n19002), .B(n27036), .C(
        n19002), .Y(n21592) );
  A2O1A1Ixp33_ASAP7_75t_SL U20274 ( .A1(n28306), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21593) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20275 ( .A1(n31662), .A2(n23161), .B(n21592), 
        .C(n19002), .D(n21593), .Y(n2563) );
  A2O1A1Ixp33_ASAP7_75t_SL U20276 ( .A1(n22422), .A2(n19002), .B(n28309), .C(
        n19002), .Y(n21590) );
  A2O1A1Ixp33_ASAP7_75t_SL U20277 ( .A1(n29792), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21591) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20278 ( .A1(n31662), .A2(n18296), .B(n21590), 
        .C(n19002), .D(n21591), .Y(n2560) );
  A2O1A1Ixp33_ASAP7_75t_SL U20279 ( .A1(n22427), .A2(n19002), .B(rf_di_w[19]), 
        .C(n21589), .Y(n2544) );
  A2O1A1Ixp33_ASAP7_75t_SL U20280 ( .A1(n30285), .A2(n19002), .B(n22414), .C(
        n21587), .Y(n21588) );
  A2O1A1Ixp33_ASAP7_75t_SL U20281 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__20_), .B(n21588), .C(n19002), .Y(n2536)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20282 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[48]), .C(n21328), .Y(n2531) );
  A2O1A1Ixp33_ASAP7_75t_SL U20283 ( .A1(n19002), .A2(n22421), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__22_), .C(n21327), .Y(n2510) );
  A2O1A1Ixp33_ASAP7_75t_SL U20284 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[50]), .C(n21326), .Y(n2504) );
  A2O1A1Ixp33_ASAP7_75t_SL U20285 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__24_), .C(n21325), .Y(n2483) );
  A2O1A1Ixp33_ASAP7_75t_SL U20286 ( .A1(n19002), .A2(n18830), .B(
        u0_0_leon3x0_p0_ici[52]), .C(n21324), .Y(n2477) );
  A2O1A1Ixp33_ASAP7_75t_SL U20287 ( .A1(n31019), .A2(n19002), .B(n21584), .C(
        n19002), .Y(n33062) );
  A2O1A1Ixp33_ASAP7_75t_SL U20288 ( .A1(n19002), .A2(n24646), .B(rf_di_w[9]), 
        .C(n20931), .Y(n2314) );
  A2O1A1Ixp33_ASAP7_75t_SL U20289 ( .A1(n19002), .A2(n27952), .B(
        uart1_r_THOLD__22__0_), .C(n21315), .Y(n2264) );
  A2O1A1Ixp33_ASAP7_75t_SL U20290 ( .A1(n30224), .A2(n19002), .B(n22414), .C(
        n21582), .Y(n21583) );
  A2O1A1Ixp33_ASAP7_75t_SL U20291 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__29_), .B(n21583), .C(n19002), .Y(n1783)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20292 ( .A1(n29334), .A2(n29335), .B(n29338), .C(
        n19002), .Y(n19685) );
  A2O1A1Ixp33_ASAP7_75t_SL U20293 ( .A1(n19002), .A2(n22433), .B(n32930), .C(
        n21314), .Y(n1717) );
  A2O1A1Ixp33_ASAP7_75t_SL U20294 ( .A1(n19002), .A2(n22433), .B(n32923), .C(
        n21311), .Y(n1709) );
  A2O1A1Ixp33_ASAP7_75t_SL U20295 ( .A1(n32660), .A2(n19002), .B(n32658), .C(
        n21580), .Y(ic_data[30]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20296 ( .A1(n32660), .A2(n19002), .B(n32638), .C(
        n21579), .Y(ic_data[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20297 ( .A1(n32660), .A2(n19002), .B(n32636), .C(
        n21578), .Y(ic_data[19]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20298 ( .A1(n32660), .A2(n19002), .B(n32634), .C(
        n21577), .Y(ic_data[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20299 ( .A1(n32660), .A2(n19002), .B(n32626), .C(
        n21576), .Y(ic_data[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20300 ( .A1(n19002), .A2(n32660), .B(n32713), .C(
        n21297), .Y(ic_data[0]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20301 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__28_), .A2(n19002), .B(n32565), .C(n19002), .Y(n21573) );
  A2O1A1Ixp33_ASAP7_75t_SL U20302 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[28]), 
        .A2(n19002), .B(n32593), .C(n19002), .Y(n21574) );
  O2A1O1Ixp33_ASAP7_75t_SL U20303 ( .A1(n32559), .A2(n21573), .B(n19002), .C(
        n21574), .Y(it_data[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20304 ( .A1(n29939), .A2(n19002), .B(n21567), .C(
        n19002), .Y(n32317) );
  A2O1A1Ixp33_ASAP7_75t_SL U20305 ( .A1(timer0_N68), .A2(n19002), .B(n21564), 
        .C(n19002), .Y(n24361) );
  A2O1A1Ixp33_ASAP7_75t_SL U20306 ( .A1(n22373), .A2(n19002), .B(n25319), .C(
        n21563), .Y(n30236) );
  A2O1A1Ixp33_ASAP7_75t_SL U20307 ( .A1(n31654), .A2(n19002), .B(
        u0_0_leon3x0_p0_muli[10]), .C(n19002), .Y(n21561) );
  A2O1A1Ixp33_ASAP7_75t_SL U20308 ( .A1(n22380), .A2(n19002), .B(n4325), .C(
        n19002), .Y(n21562) );
  A2O1A1Ixp33_ASAP7_75t_SL U20309 ( .A1(n22373), .A2(n19002), .B(n25300), .C(
        n21559), .Y(n30322) );
  A2O1A1Ixp33_ASAP7_75t_SL U20310 ( .A1(n22373), .A2(n19002), .B(n25296), .C(
        n21558), .Y(n30340) );
  A2O1A1Ixp33_ASAP7_75t_SL U20311 ( .A1(n22373), .A2(n19002), .B(n25290), .C(
        n19002), .Y(n21557) );
  A2O1A1Ixp33_ASAP7_75t_SL U20312 ( .A1(u0_0_leon3x0_p0_divi[43]), .A2(n22373), 
        .B(n21557), .C(n19002), .Y(n30376) );
  O2A1O1Ixp5_ASAP7_75t_SL U20313 ( .A1(n31559), .A2(n21555), .B(n19002), .C(
        n21556), .Y(n31562) );
  A2O1A1Ixp33_ASAP7_75t_SL U20314 ( .A1(n22373), .A2(n19002), .B(n25309), .C(
        n21554), .Y(n30272) );
  A2O1A1Ixp33_ASAP7_75t_SL U20315 ( .A1(n22373), .A2(n19002), .B(n25313), .C(
        n21553), .Y(n30257) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20316 ( .A1(n22433), .A2(n32918), .B(n19002), 
        .C(n32908), .Y(n32983) );
  A2O1A1Ixp33_ASAP7_75t_SL U20317 ( .A1(n32353), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[4]), .C(n19002), .Y(n21552) );
  A2O1A1Ixp33_ASAP7_75t_SL U20318 ( .A1(n32307), .A2(n32353), .B(n21552), .C(
        n19002), .Y(n32406) );
  A2O1A1Ixp33_ASAP7_75t_SL U20319 ( .A1(n22376), .A2(n19002), .B(n30439), .C(
        n21551), .Y(n29490) );
  A2O1A1Ixp33_ASAP7_75t_SL U20320 ( .A1(n24630), .A2(n19002), .B(n21549), .C(
        n19002), .Y(n21550) );
  A2O1A1Ixp33_ASAP7_75t_SL U20321 ( .A1(n19002), .A2(n22373), .B(n26371), .C(
        n21261), .Y(n31401) );
  A2O1A1Ixp33_ASAP7_75t_SL U20322 ( .A1(add_x_735_n54), .A2(n19002), .B(n21548), .C(n19002), .Y(add_x_735_n52) );
  A2O1A1Ixp33_ASAP7_75t_SL U20323 ( .A1(n24630), .A2(n19002), .B(
        u0_0_leon3x0_p0_divi[29]), .C(n19002), .Y(n21547) );
  O2A1O1Ixp33_ASAP7_75t_SL U20324 ( .A1(n22367), .A2(n22427), .B(n19002), .C(
        n23225), .Y(n20875) );
  A2O1A1Ixp33_ASAP7_75t_SL U20325 ( .A1(n24041), .A2(n19002), .B(
        mult_x_1196_n2750), .C(n19002), .Y(n21546) );
  A2O1A1Ixp33_ASAP7_75t_SL U20326 ( .A1(n18339), .A2(n21545), .B(n21546), .C(
        n19002), .Y(n23172) );
  A2O1A1Ixp33_ASAP7_75t_SL U20327 ( .A1(mult_x_1196_n2535), .A2(n19002), .B(
        n21543), .C(n19002), .Y(n21544) );
  A2O1A1Ixp33_ASAP7_75t_SL U20328 ( .A1(mult_x_1196_n1248), .A2(n21542), .B(
        n21544), .C(n19002), .Y(mult_x_1196_n1214) );
  A2O1A1Ixp33_ASAP7_75t_SL U20329 ( .A1(uart1_r_PARSEL_), .A2(n31950), .B(
        n21481), .C(n19002), .Y(n21482) );
  A2O1A1Ixp33_ASAP7_75t_SL U20330 ( .A1(uart1_r_RHOLD__9__4_), .A2(n31204), 
        .B(n21503), .C(n19002), .Y(n21504) );
  A2O1A1Ixp33_ASAP7_75t_SL U20331 ( .A1(n21509), .A2(n19002), .B(n21512), .C(
        n19002), .Y(n21513) );
  A2O1A1Ixp33_ASAP7_75t_SL U20332 ( .A1(n21505), .A2(n19002), .B(n21515), .C(
        n19002), .Y(n21516) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20333 ( .A1(n30789), .A2(n21484), .B(n21520), 
        .C(n19002), .D(n21523), .Y(n21524) );
  A2O1A1Ixp33_ASAP7_75t_SL U20334 ( .A1(n21483), .A2(n19002), .B(n21534), .C(
        n19002), .Y(n21535) );
  A2O1A1Ixp33_ASAP7_75t_SL U20335 ( .A1(n29406), .A2(n29405), .B(n29422), .C(
        n19002), .Y(n20860) );
  A2O1A1Ixp33_ASAP7_75t_SL U20336 ( .A1(n19002), .A2(n29429), .B(n29413), .C(
        n29433), .Y(n20862) );
  A2O1A1Ixp33_ASAP7_75t_SL U20337 ( .A1(n19002), .A2(n20863), .B(n29630), .C(
        n29629), .Y(n20864) );
  A2O1A1Ixp33_ASAP7_75t_SL U20338 ( .A1(n32786), .A2(n19002), .B(n21474), .C(
        n21475), .Y(n4729) );
  A2O1A1Ixp33_ASAP7_75t_SL U20339 ( .A1(n31722), .A2(n19002), .B(n31717), .C(
        n31740), .Y(n21467) );
  A2O1A1Ixp33_ASAP7_75t_SL U20340 ( .A1(n29949), .A2(n19002), .B(n30871), .C(
        n19002), .Y(n21463) );
  A2O1A1Ixp33_ASAP7_75t_SL U20341 ( .A1(n21463), .A2(n19002), .B(n21466), .C(
        n19002), .Y(n24528) );
  A2O1A1Ixp33_ASAP7_75t_SL U20342 ( .A1(n22427), .A2(n19002), .B(n30495), .C(
        n21462), .Y(n4652) );
  A2O1A1Ixp33_ASAP7_75t_SL U20343 ( .A1(n19002), .A2(n24646), .B(n32578), .C(
        n21235), .Y(n4646) );
  A2O1A1Ixp33_ASAP7_75t_SL U20344 ( .A1(n30577), .A2(n19002), .B(n30477), .C(
        n19002), .Y(n21460) );
  A2O1A1Ixp33_ASAP7_75t_SL U20345 ( .A1(n26680), .A2(n19002), .B(n30575), .C(
        n19002), .Y(n21461) );
  A2O1A1Ixp33_ASAP7_75t_SL U20346 ( .A1(n30644), .A2(n29783), .B(n21452), .C(
        n19002), .Y(n21453) );
  A2O1A1Ixp33_ASAP7_75t_SL U20347 ( .A1(n28808), .A2(n19002), .B(n21457), .C(
        n19002), .Y(n21458) );
  A2O1A1Ixp33_ASAP7_75t_SL U20348 ( .A1(n29801), .A2(n19002), .B(n22421), .C(
        n19002), .Y(n21448) );
  A2O1A1Ixp33_ASAP7_75t_SL U20349 ( .A1(n32110), .A2(n19002), .B(n29802), .C(
        n19002), .Y(n21449) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20350 ( .A1(n31542), .A2(n21447), .B(n21448), 
        .C(n19002), .D(n21449), .Y(n4617) );
  A2O1A1Ixp33_ASAP7_75t_SL U20351 ( .A1(n22420), .A2(n19002), .B(n29022), .C(
        n31422), .Y(n21442) );
  A2O1A1Ixp33_ASAP7_75t_SL U20352 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[29]), 
        .B(n21442), .C(n19002), .Y(n21443) );
  A2O1A1Ixp33_ASAP7_75t_SL U20353 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_29_), .B(n21445), .C(n19002), .Y(n4585) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20354 ( .A1(n26092), .A2(n26095), .B(n19002), 
        .C(n29337), .Y(n21438) );
  A2O1A1Ixp33_ASAP7_75t_SL U20355 ( .A1(n29955), .A2(n19002), .B(n30865), .C(
        n19002), .Y(n21439) );
  O2A1O1Ixp5_ASAP7_75t_SL U20356 ( .A1(n21438), .A2(n21439), .B(n19002), .C(
        n21440), .Y(n4544) );
  A2O1A1Ixp33_ASAP7_75t_SL U20357 ( .A1(n30679), .A2(n27019), .B(n21435), .C(
        n19002), .Y(n21436) );
  A2O1A1Ixp33_ASAP7_75t_SL U20358 ( .A1(n22420), .A2(n19002), .B(n28337), .C(
        n31422), .Y(n21422) );
  A2O1A1Ixp33_ASAP7_75t_SL U20359 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[11]), 
        .B(n21422), .C(n19002), .Y(n21423) );
  A2O1A1Ixp33_ASAP7_75t_SL U20360 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_11_), .B(n21425), .C(n19002), .Y(n4451) );
  A2O1A1Ixp33_ASAP7_75t_SL U20361 ( .A1(u0_0_leon3x0_p0_ici[59]), .A2(n19002), 
        .B(n24657), .C(n21420), .Y(n4330) );
  A2O1A1Ixp33_ASAP7_75t_SL U20362 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__1_), 
        .A2(n19002), .B(n24654), .C(n21412), .Y(n4161) );
  A2O1A1Ixp33_ASAP7_75t_SL U20363 ( .A1(n22420), .A2(n19002), .B(n29924), .C(
        n31422), .Y(n21400) );
  A2O1A1Ixp33_ASAP7_75t_SL U20364 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[7]), 
        .B(n21400), .C(n19002), .Y(n21401) );
  A2O1A1Ixp33_ASAP7_75t_SL U20365 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_7_), .B(n21403), .C(n19002), .Y(n3928) );
  A2O1A1Ixp33_ASAP7_75t_SL U20366 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__8_), .C(n21168), .Y(n3848) );
  A2O1A1Ixp33_ASAP7_75t_SL U20367 ( .A1(n19002), .A2(n22428), .B(n30423), .C(
        n20987), .Y(n3824) );
  A2O1A1Ixp33_ASAP7_75t_SL U20368 ( .A1(n22379), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__Y__10_), .C(n21397), .Y(n3814) );
  A2O1A1Ixp33_ASAP7_75t_SL U20369 ( .A1(n19002), .A2(n24646), .B(n30236), .C(
        n21167), .Y(n3782) );
  O2A1O1Ixp33_ASAP7_75t_SL U20370 ( .A1(n31443), .A2(n31442), .B(n19002), .C(
        n24510), .Y(n20090) );
  A2O1A1Ixp33_ASAP7_75t_SL U20371 ( .A1(n19002), .A2(n20458), .B(n22380), .C(
        n31663), .Y(n18175) );
  A2O1A1Ixp33_ASAP7_75t_SL U20372 ( .A1(u0_0_leon3x0_p0_div0_r_CNT__2_), .A2(
        n19002), .B(n24905), .C(n21389), .Y(n3722) );
  A2O1A1Ixp33_ASAP7_75t_SL U20373 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__6_), .A2(n19002), .B(n24495), .C(n19002), .Y(n21386) );
  A2O1A1Ixp33_ASAP7_75t_SL U20374 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_A__IMM__16_), .C(n19002), .Y(n21387) );
  A2O1A1Ixp33_ASAP7_75t_SL U20375 ( .A1(n22379), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__19_), .C(n21385), .Y(n3602) );
  A2O1A1Ixp33_ASAP7_75t_SL U20376 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[33]), 
        .B(n24652), .C(n20798), .Y(n3456) );
  A2O1A1Ixp33_ASAP7_75t_SL U20377 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__7_), 
        .A2(n19002), .B(n22428), .C(n21380), .Y(n3442) );
  A2O1A1Ixp33_ASAP7_75t_SL U20378 ( .A1(n19002), .A2(n29737), .B(
        u0_0_leon3x0_p0_iu_r_W__S__TT__7_), .C(n20794), .Y(n3323) );
  A2O1A1Ixp33_ASAP7_75t_SL U20379 ( .A1(n22422), .A2(n19002), .B(n29794), .C(
        n19002), .Y(n21375) );
  A2O1A1Ixp33_ASAP7_75t_SL U20380 ( .A1(n28276), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21376) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20381 ( .A1(n31662), .A2(n22556), .B(n21375), 
        .C(n19002), .D(n21376), .Y(n3313) );
  A2O1A1Ixp33_ASAP7_75t_SL U20382 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__15_), 
        .A2(n19002), .B(n22428), .C(n21371), .Y(n3222) );
  A2O1A1Ixp33_ASAP7_75t_SL U20383 ( .A1(n19002), .A2(n24646), .B(rf_di_w[14]), 
        .C(n20619), .Y(n3204) );
  A2O1A1Ixp33_ASAP7_75t_SL U20384 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[31]), .C(n21145), .Y(n3188) );
  A2O1A1Ixp33_ASAP7_75t_SL U20385 ( .A1(n30350), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21367) );
  A2O1A1Ixp33_ASAP7_75t_SL U20386 ( .A1(n30351), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21368) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20387 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__14_), 
        .A2(n31403), .B(n21367), .C(n19002), .D(n21368), .Y(n3143) );
  A2O1A1Ixp33_ASAP7_75t_SL U20388 ( .A1(n30238), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21365) );
  A2O1A1Ixp33_ASAP7_75t_SL U20389 ( .A1(n30239), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21366) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20390 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__27_), 
        .A2(n31403), .B(n21365), .C(n19002), .D(n21366), .Y(n3137) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20391 ( .A1(n32729), .A2(u0_0_leon3x0_p0_dci[2]), 
        .B(n19002), .C(n31585), .Y(n21362) );
  A2O1A1Ixp33_ASAP7_75t_SL U20392 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[13]), .C(n21361), .Y(n3089) );
  A2O1A1Ixp33_ASAP7_75t_SL U20393 ( .A1(n30181), .A2(n3054), .B(n30183), .C(
        n19002), .Y(n21356) );
  A2O1A1Ixp33_ASAP7_75t_SL U20394 ( .A1(n19002), .A2(n22428), .B(rf_di_w[2]), 
        .C(n21137), .Y(n3038) );
  A2O1A1Ixp33_ASAP7_75t_SL U20395 ( .A1(n32612), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n21351) );
  A2O1A1Ixp33_ASAP7_75t_SL U20396 ( .A1(n30800), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n21352) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20397 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__7_), .B(n21351), .C(n19002), .D(
        n21352), .Y(n2993) );
  A2O1A1Ixp33_ASAP7_75t_SL U20398 ( .A1(n22405), .A2(n19002), .B(n21349), .C(
        n32547), .Y(n21350) );
  A2O1A1Ixp33_ASAP7_75t_SL U20399 ( .A1(n19002), .A2(n31840), .B(apbi[15]), 
        .C(n20776), .Y(n2836) );
  A2O1A1Ixp33_ASAP7_75t_SL U20400 ( .A1(n30439), .A2(n19002), .B(n22414), .C(
        n21341), .Y(n21342) );
  A2O1A1Ixp33_ASAP7_75t_SL U20401 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__3_), .B(n21342), .C(n19002), .Y(n2739)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20402 ( .A1(n19002), .A2(n24646), .B(n29623), .C(
        n20771), .Y(n2733) );
  A2O1A1Ixp33_ASAP7_75t_SL U20403 ( .A1(n22422), .A2(n19002), .B(n29691), .C(
        n19002), .Y(n21338) );
  A2O1A1Ixp33_ASAP7_75t_SL U20404 ( .A1(n29692), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21339) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20405 ( .A1(n31662), .A2(
        u0_0_leon3x0_p0_muli[41]), .B(n21338), .C(n19002), .D(n21339), .Y(
        n2730) );
  A2O1A1Ixp33_ASAP7_75t_SL U20406 ( .A1(n22422), .A2(n19002), .B(n28335), .C(
        n19002), .Y(n21336) );
  A2O1A1Ixp33_ASAP7_75t_SL U20407 ( .A1(n27222), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21337) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20408 ( .A1(n31662), .A2(n22721), .B(n21336), 
        .C(n19002), .D(n21337), .Y(n2681) );
  A2O1A1Ixp33_ASAP7_75t_SL U20409 ( .A1(n30327), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21332) );
  A2O1A1Ixp33_ASAP7_75t_SL U20410 ( .A1(n30328), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21333) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20411 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__16_), 
        .A2(n31403), .B(n21332), .C(n19002), .D(n21333), .Y(n2632) );
  A2O1A1Ixp33_ASAP7_75t_SL U20412 ( .A1(n27524), .A2(n19002), .B(n27502), .C(
        n27500), .Y(n21321) );
  A2O1A1Ixp33_ASAP7_75t_SL U20413 ( .A1(n27517), .A2(n19002), .B(n21322), .C(
        n19002), .Y(n21323) );
  A2O1A1Ixp33_ASAP7_75t_SL U20414 ( .A1(n21320), .A2(n19002), .B(n21321), .C(
        n21323), .Y(n2460) );
  A2O1A1Ixp33_ASAP7_75t_SL U20415 ( .A1(n17270), .A2(n19002), .B(n30802), .C(
        n19002), .Y(n21319) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20416 ( .A1(n31019), .A2(n30801), .B(n19002), 
        .C(n21319), .Y(n2330) );
  A2O1A1Ixp33_ASAP7_75t_SL U20417 ( .A1(n19002), .A2(n22421), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__9_), .C(n21095), .Y(n2316) );
  A2O1A1Ixp33_ASAP7_75t_SL U20418 ( .A1(n22422), .A2(n19002), .B(n28298), .C(
        n19002), .Y(n21317) );
  A2O1A1Ixp33_ASAP7_75t_SL U20419 ( .A1(n28283), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21318) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20420 ( .A1(n31662), .A2(n23365), .B(n21317), 
        .C(n19002), .D(n21318), .Y(n2309) );
  A2O1A1Ixp33_ASAP7_75t_SL U20421 ( .A1(n32831), .A2(n19002), .B(datadir[0]), 
        .C(n21316), .Y(n2299) );
  A2O1A1Ixp33_ASAP7_75t_SL U20422 ( .A1(dataout[1]), .A2(n19002), .B(n21312), 
        .C(n19002), .Y(n21313) );
  A2O1A1Ixp33_ASAP7_75t_SL U20423 ( .A1(dataout[9]), .A2(n19002), .B(n21309), 
        .C(n19002), .Y(n21310) );
  A2O1A1Ixp33_ASAP7_75t_SL U20424 ( .A1(n12995), .A2(n19002), .B(n21308), .C(
        n19002), .Y(n22232) );
  A2O1A1Ixp33_ASAP7_75t_SL U20425 ( .A1(n32580), .A2(n19002), .B(n32585), .C(
        n19002), .Y(n21302) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20426 ( .A1(n32590), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__9_), .B(n21302), .C(n19002), 
        .D(n21305), .Y(n21306) );
  A2O1A1Ixp33_ASAP7_75t_SL U20427 ( .A1(n32660), .A2(n19002), .B(n32656), .C(
        n21301), .Y(ic_data[29]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20428 ( .A1(n32660), .A2(n19002), .B(n32644), .C(
        n21300), .Y(ic_data[23]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20429 ( .A1(n32660), .A2(n19002), .B(n32640), .C(
        n21299), .Y(ic_data[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20430 ( .A1(n32660), .A2(n19002), .B(n32628), .C(
        n21298), .Y(ic_data[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20431 ( .A1(n19002), .A2(n32660), .B(n32620), .C(
        n20921), .Y(ic_data[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20432 ( .A1(n19002), .A2(n32660), .B(n32734), .C(
        n20046), .Y(ic_data[1]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20433 ( .A1(n32654), .A2(n19002), .B(n32429), .C(
        n21292), .Y(n21293) );
  A2O1A1Ixp33_ASAP7_75t_SL U20434 ( .A1(n32434), .A2(n32406), .B(n21293), .C(
        n19002), .Y(n21294) );
  A2O1A1Ixp33_ASAP7_75t_SL U20435 ( .A1(n32405), .A2(n19002), .B(n32431), .C(
        n21294), .Y(n21295) );
  A2O1A1Ixp33_ASAP7_75t_SL U20436 ( .A1(n33069), .A2(dc_q[28]), .B(n21295), 
        .C(n19002), .Y(n21296) );
  A2O1A1Ixp33_ASAP7_75t_SL U20437 ( .A1(n32425), .A2(n19002), .B(n32407), .C(
        n21296), .Y(dc_data[28]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20438 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__6_), 
        .A2(n30725), .B(n20567), .C(n19002), .Y(n20568) );
  A2O1A1Ixp33_ASAP7_75t_SL U20439 ( .A1(n24641), .A2(n19002), .B(n21291), .C(
        n19002), .Y(rf_di_w[1]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20440 ( .A1(n22902), .A2(n19002), .B(n29909), .C(
        n25857), .Y(n21290) );
  A2O1A1Ixp33_ASAP7_75t_SL U20441 ( .A1(n25860), .A2(n19002), .B(n21290), .C(
        n19002), .Y(n32314) );
  A2O1A1Ixp33_ASAP7_75t_SL U20442 ( .A1(n31340), .A2(n19002), .B(n30592), .C(
        n19002), .Y(n21286) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20443 ( .A1(n31342), .A2(n30597), .B(n21286), 
        .C(n19002), .D(n21289), .Y(n30600) );
  A2O1A1Ixp33_ASAP7_75t_SL U20444 ( .A1(timer0_N66), .A2(n19002), .B(n21285), 
        .C(n19002), .Y(n24366) );
  A2O1A1Ixp33_ASAP7_75t_SL U20445 ( .A1(n18890), .A2(n28830), .B(n22578), .C(
        n19002), .Y(n21279) );
  A2O1A1Ixp33_ASAP7_75t_SL U20446 ( .A1(n18890), .A2(n19002), .B(n29150), .C(
        n21279), .Y(n21280) );
  A2O1A1Ixp33_ASAP7_75t_SL U20447 ( .A1(n18890), .A2(n19002), .B(n29148), .C(
        n19002), .Y(n21281) );
  A2O1A1Ixp33_ASAP7_75t_SL U20448 ( .A1(n18890), .A2(n19002), .B(n24631), .C(
        n19002), .Y(n21283) );
  A2O1A1Ixp33_ASAP7_75t_SL U20449 ( .A1(n28680), .A2(n18890), .B(n21283), .C(
        n19002), .Y(n21284) );
  A2O1A1Ixp33_ASAP7_75t_SL U20450 ( .A1(n21280), .A2(n21282), .B(n21284), .C(
        n19002), .Y(n30389) );
  A2O1A1Ixp33_ASAP7_75t_SL U20451 ( .A1(n22374), .A2(n19002), .B(n28321), .C(
        n19002), .Y(n21274) );
  A2O1A1Ixp33_ASAP7_75t_SL U20452 ( .A1(n18805), .A2(n19002), .B(n32638), .C(
        n19002), .Y(n21275) );
  A2O1A1Ixp33_ASAP7_75t_SL U20453 ( .A1(n22373), .A2(n19002), .B(n27025), .C(
        n19002), .Y(n21276) );
  O2A1O1Ixp5_ASAP7_75t_SL U20454 ( .A1(n21274), .A2(n21275), .B(n19002), .C(
        n21276), .Y(n27030) );
  A2O1A1Ixp33_ASAP7_75t_SL U20455 ( .A1(n22374), .A2(n19002), .B(n28324), .C(
        n19002), .Y(n21271) );
  A2O1A1Ixp33_ASAP7_75t_SL U20456 ( .A1(n18806), .A2(n19002), .B(n32634), .C(
        n19002), .Y(n21272) );
  A2O1A1Ixp33_ASAP7_75t_SL U20457 ( .A1(n22373), .A2(n19002), .B(n29094), .C(
        n19002), .Y(n21273) );
  O2A1O1Ixp5_ASAP7_75t_SL U20458 ( .A1(n21271), .A2(n21272), .B(n19002), .C(
        n21273), .Y(n31823) );
  A2O1A1Ixp33_ASAP7_75t_SL U20459 ( .A1(n19002), .A2(uart1_uarto_SCALER__10_), 
        .B(n19235), .C(uart1_uarto_SCALER__11_), .Y(n19236) );
  A2O1A1Ixp33_ASAP7_75t_SL U20460 ( .A1(n22373), .A2(n19002), .B(n25279), .C(
        n21267), .Y(n30435) );
  A2O1A1Ixp33_ASAP7_75t_SL U20461 ( .A1(n32722), .A2(n19002), .B(n21266), .C(
        n19002), .Y(n32698) );
  A2O1A1Ixp33_ASAP7_75t_SL U20462 ( .A1(n22433), .A2(n19002), .B(n32918), .C(
        n19002), .Y(n21265) );
  A2O1A1Ixp33_ASAP7_75t_SL U20463 ( .A1(n32353), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[3]), .C(n19002), .Y(n21264) );
  A2O1A1Ixp33_ASAP7_75t_SL U20464 ( .A1(n32305), .A2(n32353), .B(n21264), .C(
        n19002), .Y(n32403) );
  A2O1A1Ixp33_ASAP7_75t_SL U20465 ( .A1(n32325), .A2(n19002), .B(n24642), .C(
        n19002), .Y(n21263) );
  A2O1A1Ixp33_ASAP7_75t_SL U20466 ( .A1(n24642), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[9]), .B(n21263), .C(n19002), .Y(n32397)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20467 ( .A1(n23387), .A2(n19002), .B(n21262), .C(
        n19002), .Y(n23674) );
  A2O1A1Ixp33_ASAP7_75t_SL U20468 ( .A1(mult_x_1196_n881), .A2(n19002), .B(
        n21257), .C(mult_x_1196_n872), .Y(n21258) );
  A2O1A1Ixp33_ASAP7_75t_SL U20469 ( .A1(mult_x_1196_n874), .A2(n19002), .B(
        n21256), .C(n21258), .Y(mult_x_1196_n869) );
  A2O1A1Ixp33_ASAP7_75t_SL U20470 ( .A1(n21252), .A2(n19002), .B(n21253), .C(
        n21251), .Y(n21254) );
  A2O1A1Ixp33_ASAP7_75t_SL U20471 ( .A1(n29384), .A2(n19002), .B(n30780), .C(
        n19002), .Y(n21249) );
  A2O1A1Ixp33_ASAP7_75t_SL U20472 ( .A1(n29402), .A2(n19002), .B(n29385), .C(
        n19002), .Y(n21250) );
  A2O1A1Ixp33_ASAP7_75t_SL U20473 ( .A1(n21249), .A2(n19002), .B(n21250), .C(
        n19002), .Y(n4764) );
  A2O1A1Ixp33_ASAP7_75t_SL U20474 ( .A1(apbi[14]), .A2(n19002), .B(n29745), 
        .C(n19002), .Y(n21246) );
  A2O1A1Ixp33_ASAP7_75t_SL U20475 ( .A1(n29745), .A2(n19002), .B(
        irqctrl0_r_IPEND__14_), .C(n19002), .Y(n21247) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20476 ( .A1(n29655), .A2(n29656), .B(n21247), 
        .C(n19002), .D(n24695), .Y(n21248) );
  A2O1A1Ixp33_ASAP7_75t_SL U20477 ( .A1(n31754), .A2(n31755), .B(n31753), .C(
        n19002), .Y(n21243) );
  A2O1A1Ixp33_ASAP7_75t_SL U20478 ( .A1(n32790), .A2(n31752), .B(n31757), .C(
        n19002), .Y(n21244) );
  A2O1A1Ixp33_ASAP7_75t_SL U20479 ( .A1(n22408), .A2(n19002), .B(apbi[45]), 
        .C(n21242), .Y(n4719) );
  A2O1A1Ixp33_ASAP7_75t_SL U20480 ( .A1(n31058), .A2(n19002), .B(n29555), .C(
        n19002), .Y(n21239) );
  A2O1A1Ixp33_ASAP7_75t_SL U20481 ( .A1(n31059), .A2(n19002), .B(n29556), .C(
        n19002), .Y(n21240) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20482 ( .A1(n31061), .A2(uart1_r_RHOLD__0__2_), 
        .B(n21239), .C(n19002), .D(n21240), .Y(n4675) );
  A2O1A1Ixp33_ASAP7_75t_SL U20483 ( .A1(n31602), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mcdi[0]), .C(n19002), .Y(n21236) );
  A2O1A1Ixp33_ASAP7_75t_SL U20484 ( .A1(n21236), .A2(n19002), .B(n25597), .C(
        n19002), .Y(n21237) );
  A2O1A1Ixp33_ASAP7_75t_SL U20485 ( .A1(n18800), .A2(n19002), .B(n21237), .C(
        n19002), .Y(n21238) );
  A2O1A1Ixp33_ASAP7_75t_SL U20486 ( .A1(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__4_), 
        .A2(n30707), .B(n30706), .C(n19002), .Y(n20685) );
  A2O1A1Ixp33_ASAP7_75t_SL U20487 ( .A1(n28425), .A2(n19002), .B(n30575), .C(
        n19002), .Y(n21234) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20488 ( .A1(n28411), .A2(n31357), .B(n21234), 
        .C(n19002), .D(n30578), .Y(n4621) );
  A2O1A1Ixp33_ASAP7_75t_SL U20489 ( .A1(n28400), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n21225) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20490 ( .A1(n30644), .A2(n29796), .B(n21225), 
        .C(n19002), .D(n21228), .Y(n21229) );
  A2O1A1Ixp33_ASAP7_75t_SL U20491 ( .A1(n30645), .A2(n19002), .B(n29795), .C(
        n21229), .Y(n21230) );
  A2O1A1Ixp33_ASAP7_75t_SL U20492 ( .A1(n22432), .A2(n29800), .B(n21230), .C(
        n19002), .Y(n21231) );
  A2O1A1Ixp33_ASAP7_75t_SL U20493 ( .A1(n28799), .A2(n19002), .B(n21231), .C(
        n21232), .Y(n21233) );
  A2O1A1Ixp33_ASAP7_75t_SL U20494 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP2__26_), 
        .A2(n19002), .B(n21224), .C(n21233), .Y(n4609) );
  A2O1A1Ixp33_ASAP7_75t_SL U20495 ( .A1(n22420), .A2(n19002), .B(n29793), .C(
        n31422), .Y(n21220) );
  A2O1A1Ixp33_ASAP7_75t_SL U20496 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[25]), 
        .B(n21220), .C(n19002), .Y(n21221) );
  A2O1A1Ixp33_ASAP7_75t_SL U20497 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_25_), .B(n21223), .C(n19002), .Y(n4604) );
  A2O1A1Ixp33_ASAP7_75t_SL U20498 ( .A1(n24681), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_E__OP1__28_), .C(n19002), .Y(n21217) );
  A2O1A1Ixp33_ASAP7_75t_SL U20499 ( .A1(n32618), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n21215) );
  A2O1A1Ixp33_ASAP7_75t_SL U20500 ( .A1(n31056), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n21216) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20501 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__10_), .B(n21215), .C(n19002), .D(
        n21216), .Y(n4547) );
  A2O1A1Ixp33_ASAP7_75t_SL U20502 ( .A1(n31182), .A2(n19002), .B(n29955), .C(
        n19002), .Y(n21214) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20503 ( .A1(n29959), .A2(uart1_r_RSHIFT__7_), 
        .B(n21214), .C(n19002), .D(n29958), .Y(n4543) );
  A2O1A1Ixp33_ASAP7_75t_SL U20504 ( .A1(n25217), .A2(n25216), .B(n25215), .C(
        n19002), .Y(n21209) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20505 ( .A1(n30909), .A2(
        u0_0_leon3x0_p0_iu_r_D__ANNUL_), .B(n19002), .C(n21209), .Y(n21210) );
  A2O1A1Ixp33_ASAP7_75t_SL U20506 ( .A1(n25218), .A2(n19002), .B(n21210), .C(
        n32091), .Y(n21211) );
  A2O1A1Ixp33_ASAP7_75t_SL U20507 ( .A1(n30681), .A2(n19002), .B(n22379), .C(
        n19002), .Y(n21212) );
  A2O1A1Ixp33_ASAP7_75t_SL U20508 ( .A1(n30382), .A2(n19002), .B(n24514), .C(
        n19002), .Y(n21203) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20509 ( .A1(n24428), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__11_), .B(n24679), .C(n19002), .D(n21203), 
        .Y(n21204) );
  A2O1A1Ixp33_ASAP7_75t_SL U20510 ( .A1(n30453), .A2(n30383), .B(n21206), .C(
        n19002), .Y(n21207) );
  A2O1A1Ixp33_ASAP7_75t_SL U20511 ( .A1(n30426), .A2(n19002), .B(n30384), .C(
        n21207), .Y(n21208) );
  A2O1A1Ixp33_ASAP7_75t_SL U20512 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_divi[42]), .C(n21208), .Y(n4447) );
  A2O1A1Ixp33_ASAP7_75t_SL U20513 ( .A1(n22420), .A2(n19002), .B(n28328), .C(
        n31422), .Y(n21199) );
  A2O1A1Ixp33_ASAP7_75t_SL U20514 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[15]), 
        .B(n21199), .C(n19002), .Y(n21200) );
  A2O1A1Ixp33_ASAP7_75t_SL U20515 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_15_), .B(n21202), .C(n19002), .Y(n4427) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20516 ( .A1(n32705), .A2(n24695), .B(n19002), 
        .C(n4391), .Y(n21005) );
  A2O1A1Ixp33_ASAP7_75t_SL U20517 ( .A1(n19002), .A2(n32040), .B(n32002), .C(
        n21006), .Y(ahb0_v_HSLAVE__0_) );
  A2O1A1Ixp33_ASAP7_75t_SL U20518 ( .A1(n32610), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n21197) );
  A2O1A1Ixp33_ASAP7_75t_SL U20519 ( .A1(n31017), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n21198) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20520 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__6_), .B(n21197), .C(n19002), .D(
        n21198), .Y(n4372) );
  A2O1A1Ixp33_ASAP7_75t_SL U20521 ( .A1(n4354), .A2(n19002), .B(n21195), .C(
        n19002), .Y(n21196) );
  A2O1A1Ixp33_ASAP7_75t_SL U20522 ( .A1(timer0_vtimers_1__RELOAD__18_), .A2(
        n30993), .B(n21196), .C(n19002), .Y(n4353) );
  A2O1A1Ixp33_ASAP7_75t_SL U20523 ( .A1(n30669), .A2(n19002), .B(n30654), .C(
        n19002), .Y(n21192) );
  A2O1A1Ixp33_ASAP7_75t_SL U20524 ( .A1(n30653), .A2(n19002), .B(n21193), .C(
        n19002), .Y(n21194) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20525 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__21_), 
        .A2(n30655), .B(n21192), .C(n19002), .D(n21194), .Y(n4340) );
  A2O1A1Ixp33_ASAP7_75t_SL U20526 ( .A1(mult_x_1196_n2703), .A2(n19002), .B(
        mult_x_1196_n2143), .C(n19002), .Y(n21189) );
  A2O1A1Ixp33_ASAP7_75t_SL U20527 ( .A1(n18384), .A2(n19002), .B(n21189), .C(
        n19002), .Y(n21190) );
  A2O1A1Ixp33_ASAP7_75t_SL U20528 ( .A1(n21190), .A2(n19002), .B(n22427), .C(
        n21191), .Y(n4307) );
  A2O1A1Ixp33_ASAP7_75t_SL U20529 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__18_), .A2(n19002), .B(n24649), .C(
        n21187), .Y(n4159) );
  A2O1A1Ixp33_ASAP7_75t_SL U20530 ( .A1(n19002), .A2(n24646), .B(n28608), .C(
        n21000), .Y(n4139) );
  A2O1A1Ixp33_ASAP7_75t_SL U20531 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[1]), .B(n24657), .C(n20472), .Y(n4087) );
  A2O1A1Ixp33_ASAP7_75t_SL U20532 ( .A1(n21182), .A2(n19002), .B(n30190), .C(
        n19002), .Y(n21183) );
  A2O1A1Ixp33_ASAP7_75t_SL U20533 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[3]), .A2(
        n32120), .B(n21183), .C(n19002), .Y(n4084) );
  A2O1A1Ixp33_ASAP7_75t_SL U20534 ( .A1(n26807), .A2(n19002), .B(n26808), .C(
        n19002), .Y(n21175) );
  A2O1A1Ixp33_ASAP7_75t_SL U20535 ( .A1(n32169), .A2(n19002), .B(n31435), .C(
        n19002), .Y(n21177) );
  A2O1A1Ixp33_ASAP7_75t_SL U20536 ( .A1(n31427), .A2(n19002), .B(n26802), .C(
        n19002), .Y(n21178) );
  A2O1A1Ixp33_ASAP7_75t_SL U20537 ( .A1(n21177), .A2(n19002), .B(n21178), .C(
        n19002), .Y(n21179) );
  A2O1A1Ixp33_ASAP7_75t_SL U20538 ( .A1(n22420), .A2(n19002), .B(n30463), .C(
        n31422), .Y(n21171) );
  A2O1A1Ixp33_ASAP7_75t_SL U20539 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[2]), 
        .B(n21171), .C(n19002), .Y(n21172) );
  A2O1A1Ixp33_ASAP7_75t_SL U20540 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_2_), .B(n21174), .C(n19002), .Y(n3948) );
  A2O1A1Ixp33_ASAP7_75t_SL U20541 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[0]), .B(n24656), .C(n20811), .Y(n3908) );
  A2O1A1Ixp33_ASAP7_75t_SL U20542 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__14_), .C(n20988), .Y(n3842) );
  A2O1A1Ixp33_ASAP7_75t_SL U20543 ( .A1(n22378), .A2(n31441), .B(n31440), .C(
        n19002), .Y(n20092) );
  A2O1A1Ixp33_ASAP7_75t_SL U20544 ( .A1(n24646), .A2(n19002), .B(n21160), .C(
        n19002), .Y(n21161) );
  A2O1A1Ixp33_ASAP7_75t_SL U20545 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_), .B(n24655), .C(n19518), .Y(
        n3505) );
  A2O1A1Ixp33_ASAP7_75t_SL U20546 ( .A1(u0_0_leon3x0_p0_ici[32]), .A2(n19002), 
        .B(n24651), .C(n21153), .Y(n3466) );
  A2O1A1Ixp33_ASAP7_75t_SL U20547 ( .A1(n19002), .A2(n18829), .B(
        u0_0_leon3x0_p0_ici[33]), .C(n20979), .Y(n3458) );
  A2O1A1Ixp33_ASAP7_75t_SL U20548 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[35]), 
        .B(n24652), .C(n19872), .Y(n3446) );
  A2O1A1Ixp33_ASAP7_75t_SL U20549 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__11_), 
        .A2(n19002), .B(n24653), .C(n21151), .Y(n3412) );
  A2O1A1Ixp33_ASAP7_75t_SL U20550 ( .A1(n22427), .A2(n19002), .B(n31014), .C(
        n21149), .Y(n3332) );
  A2O1A1Ixp33_ASAP7_75t_SL U20551 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__15_), 
        .A2(n19002), .B(n22428), .C(n21147), .Y(n3220) );
  A2O1A1Ixp33_ASAP7_75t_SL U20552 ( .A1(n26369), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21142) );
  A2O1A1Ixp33_ASAP7_75t_SL U20553 ( .A1(n29180), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21143) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20554 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__1_), 
        .A2(n31403), .B(n21142), .C(n19002), .D(n21143), .Y(n3151) );
  A2O1A1Ixp33_ASAP7_75t_SL U20555 ( .A1(n30262), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21140) );
  A2O1A1Ixp33_ASAP7_75t_SL U20556 ( .A1(n30263), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21141) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20557 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__23_), 
        .A2(n31403), .B(n21140), .C(n19002), .D(n21141), .Y(n3140) );
  A2O1A1Ixp33_ASAP7_75t_SL U20558 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[12]), .C(n21139), .Y(n3087) );
  A2O1A1Ixp33_ASAP7_75t_SL U20559 ( .A1(n22422), .A2(n19002), .B(n28276), .C(
        n19002), .Y(n21134) );
  A2O1A1Ixp33_ASAP7_75t_SL U20560 ( .A1(n28282), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21135) );
  A2O1A1Ixp33_ASAP7_75t_SL U20561 ( .A1(n18491), .A2(n31662), .B(n21134), .C(
        n19002), .Y(n18495) );
  A2O1A1Ixp33_ASAP7_75t_SL U20562 ( .A1(n32620), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n21132) );
  A2O1A1Ixp33_ASAP7_75t_SL U20563 ( .A1(n30973), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n21133) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20564 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__11_), .B(n21132), .C(n19002), .D(
        n21133), .Y(n2990) );
  A2O1A1Ixp33_ASAP7_75t_SL U20565 ( .A1(n19002), .A2(n24633), .B(
        uart1_r_PARSEL_), .C(n20941), .Y(n2860) );
  A2O1A1Ixp33_ASAP7_75t_SL U20566 ( .A1(n29383), .A2(n19002), .B(apbi[1]), .C(
        n21119), .Y(n2856) );
  A2O1A1Ixp33_ASAP7_75t_SL U20567 ( .A1(n31680), .A2(n19002), .B(n22414), .C(
        n21116), .Y(n21117) );
  A2O1A1Ixp33_ASAP7_75t_SL U20568 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__31_), .B(n21117), .C(n19002), .Y(n2812)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20569 ( .A1(n20056), .A2(
        u0_0_leon3x0_p0_div0_addout_0_), .B(n20060), .C(n19002), .Y(n2810) );
  A2O1A1Ixp33_ASAP7_75t_SL U20570 ( .A1(n22420), .A2(n19002), .B(n29691), .C(
        n31422), .Y(n21111) );
  A2O1A1Ixp33_ASAP7_75t_SL U20571 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[4]), 
        .B(n21111), .C(n19002), .Y(n21112) );
  A2O1A1Ixp33_ASAP7_75t_SL U20572 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_4_), .B(n21114), .C(n19002), .Y(n2735) );
  A2O1A1Ixp33_ASAP7_75t_SL U20573 ( .A1(n22422), .A2(n19002), .B(n29926), .C(
        n19002), .Y(n21109) );
  A2O1A1Ixp33_ASAP7_75t_SL U20574 ( .A1(n27176), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n21110) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20575 ( .A1(n31662), .A2(add_x_735_A_9_), .B(
        n21109), .C(n19002), .D(n21110), .Y(n2682) );
  A2O1A1Ixp33_ASAP7_75t_SL U20576 ( .A1(n22427), .A2(n19002), .B(rf_di_w[13]), 
        .C(n21108), .Y(n2641) );
  A2O1A1Ixp33_ASAP7_75t_SL U20577 ( .A1(n19002), .A2(n24646), .B(rf_di_w[16]), 
        .C(n20937), .Y(n2617) );
  A2O1A1Ixp33_ASAP7_75t_SL U20578 ( .A1(n30320), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21105) );
  A2O1A1Ixp33_ASAP7_75t_SL U20579 ( .A1(n30317), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21106) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20580 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__17_), .B(n21105), .C(n19002), .D(n21106), 
        .Y(n2608) );
  A2O1A1Ixp33_ASAP7_75t_SL U20581 ( .A1(n19002), .A2(n24646), .B(rf_di_w[17]), 
        .C(n20936), .Y(n2593) );
  A2O1A1Ixp33_ASAP7_75t_SL U20582 ( .A1(n30296), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21103) );
  A2O1A1Ixp33_ASAP7_75t_SL U20583 ( .A1(n30297), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21104) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20584 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__19_), 
        .A2(n31403), .B(n21103), .C(n19002), .D(n21104), .Y(n2559) );
  A2O1A1Ixp33_ASAP7_75t_SL U20585 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__20_), .C(n20935), .Y(n2537) );
  A2O1A1Ixp33_ASAP7_75t_SL U20586 ( .A1(n30270), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21101) );
  A2O1A1Ixp33_ASAP7_75t_SL U20587 ( .A1(n30267), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21102) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20588 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__22_), 
        .A2(n31403), .B(n21101), .C(n19002), .D(n21102), .Y(n2509) );
  A2O1A1Ixp33_ASAP7_75t_SL U20589 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__22_), 
        .A2(n19002), .B(n22428), .C(n21100), .Y(n2500) );
  A2O1A1Ixp33_ASAP7_75t_SL U20590 ( .A1(n30251), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n21097) );
  A2O1A1Ixp33_ASAP7_75t_SL U20591 ( .A1(n30252), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n21098) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20592 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__24_), 
        .A2(n31403), .B(n21097), .C(n19002), .D(n21098), .Y(n2482) );
  A2O1A1Ixp33_ASAP7_75t_SL U20593 ( .A1(n19002), .A2(n24646), .B(rf_di_w[24]), 
        .C(n20932), .Y(n2467) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20594 ( .A1(n25412), .A2(n31949), .B(n19002), 
        .C(n2926), .Y(n20598) );
  A2O1A1Ixp33_ASAP7_75t_SL U20595 ( .A1(n20597), .A2(n20598), .B(n22234), .C(
        n19002), .Y(n33063) );
  A2O1A1Ixp33_ASAP7_75t_SL U20596 ( .A1(n30801), .A2(n19002), .B(n21096), .C(
        n19002), .Y(n2329) );
  A2O1A1Ixp33_ASAP7_75t_SL U20597 ( .A1(n19002), .A2(n27926), .B(
        uart1_r_THOLD__21__0_), .C(n19849), .Y(n2263) );
  A2O1A1Ixp33_ASAP7_75t_SL U20598 ( .A1(n19002), .A2(n27948), .B(
        uart1_r_THOLD__10__0_), .C(n19848), .Y(n2256) );
  A2O1A1Ixp33_ASAP7_75t_SL U20599 ( .A1(n29341), .A2(n29340), .B(n29344), .C(
        n19002), .Y(n21094) );
  A2O1A1Ixp33_ASAP7_75t_SL U20600 ( .A1(n19002), .A2(n22433), .B(n32938), .C(
        n20925), .Y(n1716) );
  A2O1A1Ixp33_ASAP7_75t_SL U20601 ( .A1(n19002), .A2(n22433), .B(n32939), .C(
        n20759), .Y(n1707) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20602 ( .A1(uart1_r_LOOPB_), .A2(n33068), .B(
        n19002), .C(uart1_r_TSHIFT__0_), .Y(n22235) );
  A2O1A1Ixp33_ASAP7_75t_SL U20603 ( .A1(timer0_N61), .A2(n19002), .B(n21092), 
        .C(timer0_N60), .Y(n21093) );
  A2O1A1Ixp33_ASAP7_75t_SL U20604 ( .A1(timer0_N61), .A2(n19002), .B(n21091), 
        .C(n21093), .Y(timer0_res_31_) );
  A2O1A1Ixp33_ASAP7_75t_SL U20605 ( .A1(n32574), .A2(n19002), .B(n32585), .C(
        n19002), .Y(n21084) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20606 ( .A1(n32590), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__7_), .B(n21084), .C(n19002), 
        .D(n21087), .Y(n21088) );
  A2O1A1Ixp33_ASAP7_75t_SL U20607 ( .A1(n32660), .A2(n19002), .B(n32642), .C(
        n21083), .Y(ic_data[22]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20608 ( .A1(n32444), .A2(u0_0_leon3x0_p0_dci[14]), 
        .B(n19478), .C(n19002), .Y(n19479) );
  A2O1A1Ixp33_ASAP7_75t_SL U20609 ( .A1(n19002), .A2(n33067), .B(n19479), .C(
        n19480), .Y(dc_address[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20610 ( .A1(n32432), .A2(n19002), .B(n32431), .C(
        n20579), .Y(n20580) );
  A2O1A1Ixp33_ASAP7_75t_SL U20611 ( .A1(n32217), .A2(n19002), .B(n32640), .C(
        n20744), .Y(dt_data[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20612 ( .A1(timer0_r_SCALER__7_), .A2(n19002), .B(
        n21082), .C(n19002), .Y(timer0_v_TICK_) );
  A2O1A1Ixp33_ASAP7_75t_SL U20613 ( .A1(n23954), .A2(n19002), .B(n30008), .C(
        n19002), .Y(n21079) );
  A2O1A1Ixp33_ASAP7_75t_SL U20614 ( .A1(n21079), .A2(n19002), .B(n21080), .C(
        n19002), .Y(n32305) );
  A2O1A1Ixp33_ASAP7_75t_SL U20615 ( .A1(n31340), .A2(n19002), .B(n29808), .C(
        n19002), .Y(n21075) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20616 ( .A1(n31342), .A2(n29807), .B(n21075), 
        .C(n19002), .D(n21078), .Y(n29073) );
  A2O1A1Ixp33_ASAP7_75t_SL U20617 ( .A1(u0_0_leon3x0_p0_iu_r_E__CTRL__WICC_), 
        .A2(n19002), .B(n21074), .C(n19002), .Y(n30946) );
  A2O1A1Ixp33_ASAP7_75t_SL U20618 ( .A1(n31579), .A2(n19002), .B(n21073), .C(
        n19002), .Y(n31456) );
  A2O1A1Ixp33_ASAP7_75t_SL U20619 ( .A1(n22374), .A2(n19002), .B(n28301), .C(
        n19002), .Y(n21070) );
  A2O1A1Ixp33_ASAP7_75t_SL U20620 ( .A1(n18806), .A2(n19002), .B(n32658), .C(
        n19002), .Y(n21071) );
  A2O1A1Ixp33_ASAP7_75t_SL U20621 ( .A1(n22373), .A2(n19002), .B(n29084), .C(
        n19002), .Y(n21072) );
  O2A1O1Ixp5_ASAP7_75t_SL U20622 ( .A1(n21070), .A2(n21071), .B(n19002), .C(
        n21072), .Y(n30592) );
  A2O1A1Ixp33_ASAP7_75t_SL U20623 ( .A1(timer0_N70), .A2(n19002), .B(n21069), 
        .C(n19002), .Y(n24356) );
  A2O1A1Ixp33_ASAP7_75t_SL U20624 ( .A1(n22373), .A2(n19002), .B(n25317), .C(
        n21068), .Y(n30240) );
  A2O1A1Ixp33_ASAP7_75t_SL U20625 ( .A1(n31340), .A2(n19002), .B(n31823), .C(
        n19002), .Y(n21064) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20626 ( .A1(n31342), .A2(n28546), .B(n21064), 
        .C(n19002), .D(n21067), .Y(n27282) );
  A2O1A1Ixp33_ASAP7_75t_SL U20627 ( .A1(add_x_746_n2), .A2(n19002), .B(n21063), 
        .C(n19002), .Y(add_x_746_n5) );
  A2O1A1Ixp33_ASAP7_75t_SL U20628 ( .A1(n22373), .A2(n19002), .B(n25306), .C(
        n19002), .Y(n21059) );
  A2O1A1Ixp33_ASAP7_75t_SL U20629 ( .A1(u0_0_leon3x0_p0_divi[51]), .A2(n22373), 
        .B(n21059), .C(n19002), .Y(n30291) );
  A2O1A1Ixp33_ASAP7_75t_SL U20630 ( .A1(n22373), .A2(n19002), .B(n25298), .C(
        n21058), .Y(n30333) );
  A2O1A1Ixp33_ASAP7_75t_SL U20631 ( .A1(n22373), .A2(n19002), .B(n25294), .C(
        n21057), .Y(n30356) );
  A2O1A1Ixp33_ASAP7_75t_SL U20632 ( .A1(n22373), .A2(n19002), .B(n25283), .C(
        n19002), .Y(n21056) );
  A2O1A1Ixp33_ASAP7_75t_SL U20633 ( .A1(u0_0_leon3x0_p0_divi[38]), .A2(n22373), 
        .B(n21056), .C(n19002), .Y(n30402) );
  A2O1A1Ixp33_ASAP7_75t_SL U20634 ( .A1(n22373), .A2(n19002), .B(n25280), .C(
        n21055), .Y(n30423) );
  A2O1A1Ixp33_ASAP7_75t_SL U20635 ( .A1(n22373), .A2(n19002), .B(n25322), .C(
        n19002), .Y(n21054) );
  A2O1A1Ixp33_ASAP7_75t_SL U20636 ( .A1(u0_0_leon3x0_p0_divi[61]), .A2(n22373), 
        .B(n21054), .C(n19002), .Y(n30219) );
  A2O1A1Ixp33_ASAP7_75t_SL U20637 ( .A1(n32320), .A2(n19002), .B(n24642), .C(
        n19002), .Y(n21053) );
  A2O1A1Ixp33_ASAP7_75t_SL U20638 ( .A1(n24642), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[8]), .B(n21053), .C(n19002), .Y(n32394)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20639 ( .A1(n32580), .A2(n19002), .B(n18876), .C(
        n20526), .Y(u0_0_leon3x0_p0_iu_fe_pc_9_) );
  A2O1A1Ixp33_ASAP7_75t_SL U20640 ( .A1(sr1_r_BUSW__1_), .A2(n19002), .B(n1723), .C(n19002), .Y(n21052) );
  A2O1A1Ixp33_ASAP7_75t_SL U20641 ( .A1(n2357), .A2(n19002), .B(n32884), .C(
        n21052), .Y(n32885) );
  A2O1A1Ixp33_ASAP7_75t_SL U20642 ( .A1(u0_0_leon3x0_p0_divi[30]), .A2(n19002), 
        .B(n24630), .C(n19002), .Y(n21051) );
  A2O1A1Ixp33_ASAP7_75t_SL U20643 ( .A1(n29384), .A2(n19002), .B(n29851), .C(
        n19002), .Y(n21048) );
  A2O1A1Ixp33_ASAP7_75t_SL U20644 ( .A1(n29399), .A2(n19002), .B(n29385), .C(
        n19002), .Y(n21049) );
  A2O1A1Ixp33_ASAP7_75t_SL U20645 ( .A1(n21048), .A2(n19002), .B(n21049), .C(
        n19002), .Y(n4753) );
  A2O1A1Ixp33_ASAP7_75t_SL U20646 ( .A1(n29883), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_M__CTRL__TT__0_), .C(n19002), .Y(n21042) );
  A2O1A1Ixp33_ASAP7_75t_SL U20647 ( .A1(n29639), .A2(n18845), .B(n29726), .C(
        n19002), .Y(n21043) );
  A2O1A1Ixp33_ASAP7_75t_SL U20648 ( .A1(n21042), .A2(n19002), .B(n21043), .C(
        n19002), .Y(n21044) );
  A2O1A1Ixp33_ASAP7_75t_SL U20649 ( .A1(n21044), .A2(n19002), .B(n21047), .C(
        n19002), .Y(n4733) );
  A2O1A1Ixp33_ASAP7_75t_SL U20650 ( .A1(sr1_r_MCFG1__ROMWWS__1_), .A2(n31725), 
        .B(n20854), .C(n19002), .Y(n20855) );
  A2O1A1Ixp33_ASAP7_75t_SL U20651 ( .A1(n29949), .A2(n19002), .B(n30077), .C(
        n19002), .Y(n21037) );
  A2O1A1Ixp33_ASAP7_75t_SL U20652 ( .A1(n21037), .A2(n19002), .B(n21040), .C(
        n19002), .Y(n24525) );
  A2O1A1Ixp33_ASAP7_75t_SL U20653 ( .A1(n22393), .A2(n19002), .B(n32996), .C(
        n19002), .Y(n21036) );
  A2O1A1Ixp33_ASAP7_75t_SL U20654 ( .A1(ahb0_r_HADDR__8_), .A2(n21035), .B(
        n21036), .C(n19002), .Y(n4644) );
  A2O1A1Ixp33_ASAP7_75t_SL U20655 ( .A1(n26236), .A2(n19002), .B(n30575), .C(
        n19002), .Y(n21034) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20656 ( .A1(n28411), .A2(n31044), .B(n21034), 
        .C(n19002), .D(n30578), .Y(n4611) );
  A2O1A1Ixp33_ASAP7_75t_SL U20657 ( .A1(n24638), .A2(n19002), .B(n21027), .C(
        n19002), .Y(n21028) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20658 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__25_), .B(n24680), .C(n19002), .D(n21028), 
        .Y(n21029) );
  A2O1A1Ixp33_ASAP7_75t_SL U20659 ( .A1(n30453), .A2(n30249), .B(n21031), .C(
        n19002), .Y(n21032) );
  A2O1A1Ixp33_ASAP7_75t_SL U20660 ( .A1(n30426), .A2(n19002), .B(n30250), .C(
        n21032), .Y(n21033) );
  A2O1A1Ixp33_ASAP7_75t_SL U20661 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_divi[56]), .C(n21033), .Y(n4605) );
  A2O1A1Ixp33_ASAP7_75t_SL U20662 ( .A1(n28271), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n21018) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20663 ( .A1(n28272), .A2(n30644), .B(n21018), 
        .C(n19002), .D(n21021), .Y(n21022) );
  A2O1A1Ixp33_ASAP7_75t_SL U20664 ( .A1(n30645), .A2(n19002), .B(n28273), .C(
        n21022), .Y(n21023) );
  A2O1A1Ixp33_ASAP7_75t_SL U20665 ( .A1(n28275), .A2(n22432), .B(n21023), .C(
        n19002), .Y(n21024) );
  A2O1A1Ixp33_ASAP7_75t_SL U20666 ( .A1(n28799), .A2(n19002), .B(n21024), .C(
        n19002), .Y(n21025) );
  A2O1A1Ixp33_ASAP7_75t_SL U20667 ( .A1(n24681), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_E__OP1__29_), .C(n19002), .Y(n21015) );
  A2O1A1Ixp33_ASAP7_75t_SL U20668 ( .A1(n22427), .A2(n19002), .B(n32581), .C(
        n21014), .Y(n4562) );
  A2O1A1Ixp33_ASAP7_75t_SL U20669 ( .A1(n30062), .A2(n19002), .B(n29955), .C(
        n19002), .Y(n21013) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20670 ( .A1(n29959), .A2(uart1_r_RSHIFT__6_), 
        .B(n21013), .C(n19002), .D(n29958), .Y(n4542) );
  A2O1A1Ixp33_ASAP7_75t_SL U20671 ( .A1(n31058), .A2(n19002), .B(n26126), .C(
        n19002), .Y(n21011) );
  A2O1A1Ixp33_ASAP7_75t_SL U20672 ( .A1(n31059), .A2(n19002), .B(n26127), .C(
        n19002), .Y(n21012) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20673 ( .A1(n31061), .A2(uart1_r_RHOLD__0__1_), 
        .B(n21011), .C(n19002), .D(n21012), .Y(n4537) );
  A2O1A1Ixp33_ASAP7_75t_SL U20674 ( .A1(n22420), .A2(n19002), .B(n28309), .C(
        n31422), .Y(n21007) );
  A2O1A1Ixp33_ASAP7_75t_SL U20675 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[23]), 
        .B(n21007), .C(n19002), .Y(n21008) );
  A2O1A1Ixp33_ASAP7_75t_SL U20676 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_23_), .B(n21010), .C(n19002), .Y(n4420) );
  A2O1A1Ixp33_ASAP7_75t_SL U20677 ( .A1(n22431), .A2(n19002), .B(n31659), .C(
        n19002), .Y(n21003) );
  A2O1A1Ixp33_ASAP7_75t_SL U20678 ( .A1(n22427), .A2(n19002), .B(n20654), .C(
        n20655), .Y(n4305) );
  A2O1A1Ixp33_ASAP7_75t_SL U20679 ( .A1(n4032), .A2(n19002), .B(n20998), .C(
        n19002), .Y(n20999) );
  A2O1A1Ixp33_ASAP7_75t_SL U20680 ( .A1(timer0_vtimers_1__RELOAD__17_), .A2(
        n30993), .B(n20999), .C(n19002), .Y(n4031) );
  A2O1A1Ixp33_ASAP7_75t_SL U20681 ( .A1(u0_0_leon3x0_p0_iu_v_E__CWP__2_), .A2(
        n19002), .B(n24651), .C(n20997), .Y(n4014) );
  A2O1A1Ixp33_ASAP7_75t_SL U20682 ( .A1(n22420), .A2(n19002), .B(n28335), .C(
        n31422), .Y(n20992) );
  A2O1A1Ixp33_ASAP7_75t_SL U20683 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[12]), 
        .B(n20992), .C(n19002), .Y(n20993) );
  A2O1A1Ixp33_ASAP7_75t_SL U20684 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_12_), .B(n20995), .C(n19002), .Y(n3973) );
  A2O1A1Ixp33_ASAP7_75t_SL U20685 ( .A1(n32121), .A2(n20989), .B(n20991), .C(
        n19002), .Y(n3913) );
  A2O1A1Ixp33_ASAP7_75t_SL U20686 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__21_), .B(n24655), .C(n20803), .Y(
        n3869) );
  A2O1A1Ixp33_ASAP7_75t_SL U20687 ( .A1(n19002), .A2(n24646), .B(n28806), .C(
        n20800), .Y(n3852) );
  A2O1A1Ixp33_ASAP7_75t_SL U20688 ( .A1(n19002), .A2(n22421), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__10_), .C(n20799), .Y(n3846) );
  A2O1A1Ixp33_ASAP7_75t_SL U20689 ( .A1(u0_0_leon3x0_p0_iu_v_M__MUL_), .A2(
        n19002), .B(n24656), .C(n20985), .Y(n3778) );
  A2O1A1Ixp33_ASAP7_75t_SL U20690 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__9_), .B(n24652), .C(n20454), .Y(
        n3657) );
  A2O1A1Ixp33_ASAP7_75t_SL U20691 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__1_), .A2(
        n19002), .B(n30813), .C(n19002), .Y(n20982) );
  A2O1A1Ixp33_ASAP7_75t_SL U20692 ( .A1(n20982), .A2(n19002), .B(n30814), .C(
        n19002), .Y(n20983) );
  A2O1A1Ixp33_ASAP7_75t_SL U20693 ( .A1(n24646), .A2(n19002), .B(
        DP_OP_1196_128_7433_n453), .C(n20983), .Y(n3546) );
  A2O1A1Ixp33_ASAP7_75t_SL U20694 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__4_), 
        .A2(n19002), .B(n24650), .C(n20981), .Y(n3460) );
  A2O1A1Ixp33_ASAP7_75t_SL U20695 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__7_), 
        .A2(n19002), .B(n22428), .C(n20978), .Y(n3440) );
  A2O1A1Ixp33_ASAP7_75t_SL U20696 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__11_), 
        .A2(n19002), .B(n24653), .C(n20975), .Y(n3414) );
  A2O1A1Ixp33_ASAP7_75t_SL U20697 ( .A1(n24646), .A2(n19002), .B(rf_di_w[25]), 
        .C(n20973), .Y(n3379) );
  A2O1A1Ixp33_ASAP7_75t_SL U20698 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__3_), 
        .A2(n19002), .B(n22428), .C(n20969), .Y(n3344) );
  A2O1A1Ixp33_ASAP7_75t_SL U20699 ( .A1(n22422), .A2(n19002), .B(n28353), .C(
        n19002), .Y(n20962) );
  A2O1A1Ixp33_ASAP7_75t_SL U20700 ( .A1(n30463), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n20963) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20701 ( .A1(n31662), .A2(add_x_735_A_2_), .B(
        n20962), .C(n19002), .D(n20963), .Y(n3312) );
  A2O1A1Ixp33_ASAP7_75t_SL U20702 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_), .C(n20961), .Y(n3310) );
  A2O1A1Ixp33_ASAP7_75t_SL U20703 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__15_), 
        .A2(n19002), .B(n22428), .C(n20959), .Y(n3218) );
  A2O1A1Ixp33_ASAP7_75t_SL U20704 ( .A1(n30458), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n20956) );
  A2O1A1Ixp33_ASAP7_75t_SL U20705 ( .A1(n30450), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n20957) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20706 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__2_), 
        .A2(n31403), .B(n20956), .C(n19002), .D(n20957), .Y(n3150) );
  A2O1A1Ixp33_ASAP7_75t_SL U20707 ( .A1(n19002), .A2(n30397), .B(n22414), .C(
        n20616), .Y(n20617) );
  A2O1A1Ixp33_ASAP7_75t_SL U20708 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__7_), .B(n20617), .C(n19002), .Y(n3147)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20709 ( .A1(n30392), .A2(n19002), .B(n22414), .C(
        n20954), .Y(n20955) );
  A2O1A1Ixp33_ASAP7_75t_SL U20710 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__8_), .B(n20955), .C(n19002), .Y(n3146)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20711 ( .A1(n30338), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n20951) );
  A2O1A1Ixp33_ASAP7_75t_SL U20712 ( .A1(n30339), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n20952) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20713 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__15_), 
        .A2(n31403), .B(n20951), .C(n19002), .D(n20952), .Y(n3142) );
  A2O1A1Ixp33_ASAP7_75t_SL U20714 ( .A1(n30277), .A2(n19002), .B(n22414), .C(
        n20949), .Y(n20950) );
  A2O1A1Ixp33_ASAP7_75t_SL U20715 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__21_), .B(n20950), .C(n19002), .Y(n3141)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20716 ( .A1(n30234), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n20946) );
  A2O1A1Ixp33_ASAP7_75t_SL U20717 ( .A1(n30235), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n20947) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20718 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__28_), 
        .A2(n31403), .B(n20946), .C(n19002), .D(n20947), .Y(n3136) );
  A2O1A1Ixp33_ASAP7_75t_SL U20719 ( .A1(n32622), .A2(n19002), .B(n32729), .C(
        n19002), .Y(n20944) );
  A2O1A1Ixp33_ASAP7_75t_SL U20720 ( .A1(n31790), .A2(n19002), .B(n24645), .C(
        n19002), .Y(n20945) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20721 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__12_), .B(n20944), .C(n19002), .D(
        n20945), .Y(n2988) );
  A2O1A1Ixp33_ASAP7_75t_SL U20722 ( .A1(n31198), .A2(n19002), .B(
        sr1_r_MCFG2__RAMBANKSZ__1_), .C(n20064), .Y(n2914) );
  A2O1A1Ixp33_ASAP7_75t_SL U20723 ( .A1(n28056), .A2(n19002), .B(apbi[11]), 
        .C(n20943), .Y(n2884) );
  A2O1A1Ixp33_ASAP7_75t_SL U20724 ( .A1(n19002), .A2(n24633), .B(
        uart1_r_TIRQEN_), .C(n20777), .Y(n2858) );
  A2O1A1Ixp33_ASAP7_75t_SL U20725 ( .A1(n30610), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n20939) );
  A2O1A1Ixp33_ASAP7_75t_SL U20726 ( .A1(n31423), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n20940) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20727 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__0_), 
        .A2(n31403), .B(n20939), .C(n19002), .D(n20940), .Y(n2769) );
  A2O1A1Ixp33_ASAP7_75t_SL U20728 ( .A1(n22427), .A2(n19002), .B(n29887), .C(
        n20938), .Y(n2742) );
  A2O1A1Ixp33_ASAP7_75t_SL U20729 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__22_), 
        .A2(n19002), .B(n22428), .C(n20934), .Y(n2498) );
  A2O1A1Ixp33_ASAP7_75t_SL U20730 ( .A1(n19002), .A2(n29812), .B(n30654), .C(
        n20602), .Y(n20603) );
  A2O1A1Ixp33_ASAP7_75t_SL U20731 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__23_), 
        .A2(n30655), .B(n20603), .C(n19002), .Y(n2366) );
  A2O1A1Ixp33_ASAP7_75t_SL U20732 ( .A1(n30388), .A2(n19002), .B(n22414), .C(
        n20929), .Y(n20930) );
  A2O1A1Ixp33_ASAP7_75t_SL U20733 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__9_), .B(n20930), .C(n19002), .Y(n2313)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20734 ( .A1(n22422), .A2(n19002), .B(n28283), .C(
        n19002), .Y(n20926) );
  A2O1A1Ixp33_ASAP7_75t_SL U20735 ( .A1(n28295), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n20927) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20736 ( .A1(n31662), .A2(n18530), .B(n20926), 
        .C(n19002), .D(n20927), .Y(n2308) );
  A2O1A1Ixp33_ASAP7_75t_SL U20737 ( .A1(dataout[2]), .A2(n19002), .B(n20923), 
        .C(n19002), .Y(n20924) );
  A2O1A1Ixp33_ASAP7_75t_SL U20738 ( .A1(n19002), .A2(n22433), .B(n32947), .C(
        n20588), .Y(n1706) );
  A2O1A1Ixp33_ASAP7_75t_SL U20739 ( .A1(n30555), .A2(n19002), .B(n20922), .C(
        n19002), .Y(n4431) );
  A2O1A1Ixp33_ASAP7_75t_SL U20740 ( .A1(n19002), .A2(n32660), .B(n32614), .C(
        n20584), .Y(ic_data[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20741 ( .A1(n32660), .A2(n19002), .B(n32612), .C(
        n20920), .Y(ic_data[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20742 ( .A1(n19002), .A2(n32660), .B(n32608), .C(
        n20754), .Y(ic_data[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20743 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__31_), .A2(n19002), .B(n32565), .C(n19002), .Y(n20918) );
  A2O1A1Ixp33_ASAP7_75t_SL U20744 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[31]), 
        .A2(n19002), .B(n32593), .C(n19002), .Y(n20919) );
  O2A1O1Ixp33_ASAP7_75t_SL U20745 ( .A1(n32559), .A2(n20918), .B(n19002), .C(
        n20919), .Y(it_data[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20746 ( .A1(n32640), .A2(n19002), .B(n32543), .C(
        n20917), .Y(it_data[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20747 ( .A1(n32648), .A2(n19002), .B(n32429), .C(
        n20911), .Y(n20912) );
  A2O1A1Ixp33_ASAP7_75t_SL U20748 ( .A1(n32434), .A2(n32396), .B(n20912), .C(
        n19002), .Y(n20913) );
  A2O1A1Ixp33_ASAP7_75t_SL U20749 ( .A1(n32395), .A2(n19002), .B(n32431), .C(
        n20913), .Y(n20914) );
  A2O1A1Ixp33_ASAP7_75t_SL U20750 ( .A1(n33069), .A2(dc_q[25]), .B(n20914), 
        .C(n19002), .Y(n20915) );
  A2O1A1Ixp33_ASAP7_75t_SL U20751 ( .A1(n32425), .A2(n19002), .B(n32397), .C(
        n20915), .Y(dc_data[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20752 ( .A1(n32636), .A2(n19002), .B(n32217), .C(
        n20263), .Y(dt_data[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20753 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__27_), 
        .A2(n30725), .B(n20738), .C(n19002), .Y(n20739) );
  O2A1O1Ixp5_ASAP7_75t_SL U20754 ( .A1(timer0_N60), .A2(n20909), .B(n19002), 
        .C(n20910), .Y(n30739) );
  A2O1A1Ixp33_ASAP7_75t_SL U20755 ( .A1(n30009), .A2(n19002), .B(n30010), .C(
        n19002), .Y(n20906) );
  A2O1A1Ixp33_ASAP7_75t_SL U20756 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__5_), .A2(
        n22375), .B(n30006), .C(n19002), .Y(n20907) );
  A2O1A1Ixp33_ASAP7_75t_SL U20757 ( .A1(n18314), .A2(n19002), .B(n30008), .C(
        n20907), .Y(n20908) );
  A2O1A1Ixp33_ASAP7_75t_SL U20758 ( .A1(n20906), .A2(n19002), .B(n20908), .C(
        n19002), .Y(n32310) );
  A2O1A1Ixp33_ASAP7_75t_SL U20759 ( .A1(apb0_r_STATE__0_), .A2(n19002), .B(
        n20904), .C(n20905), .Y(n31838) );
  A2O1A1Ixp33_ASAP7_75t_SL U20760 ( .A1(n22374), .A2(n19002), .B(n28305), .C(
        n19002), .Y(n20901) );
  A2O1A1Ixp33_ASAP7_75t_SL U20761 ( .A1(n18806), .A2(n19002), .B(n32650), .C(
        n19002), .Y(n20902) );
  A2O1A1Ixp33_ASAP7_75t_SL U20762 ( .A1(n22373), .A2(n19002), .B(n29086), .C(
        n19002), .Y(n20903) );
  O2A1O1Ixp5_ASAP7_75t_SL U20763 ( .A1(n20901), .A2(n20902), .B(n19002), .C(
        n20903), .Y(n29795) );
  A2O1A1Ixp33_ASAP7_75t_SL U20764 ( .A1(u0_0_leon3x0_p0_iu_r_A__WUNF_), .A2(
        n19002), .B(n20900), .C(n19002), .Y(n29698) );
  A2O1A1Ixp33_ASAP7_75t_SL U20765 ( .A1(n30195), .A2(n19002), .B(n20899), .C(
        n19002), .Y(n32280) );
  O2A1O1Ixp33_ASAP7_75t_SL U20766 ( .A1(n22374), .A2(n31673), .B(n19002), .C(
        n31982), .Y(n19456) );
  A2O1A1Ixp33_ASAP7_75t_SL U20767 ( .A1(add_x_746_n2), .A2(n19002), .B(n20898), 
        .C(n19002), .Y(add_x_746_n10) );
  A2O1A1Ixp33_ASAP7_75t_SL U20768 ( .A1(n22752), .A2(n19002), .B(
        mult_x_1196_n580), .C(n20897), .Y(mult_x_1196_n548) );
  A2O1A1Ixp33_ASAP7_75t_SL U20769 ( .A1(n23213), .A2(n19002), .B(n20896), .C(
        n19002), .Y(n23212) );
  A2O1A1Ixp33_ASAP7_75t_SL U20770 ( .A1(n23941), .A2(n19002), .B(n20889), .C(
        n19002), .Y(n20890) );
  A2O1A1Ixp33_ASAP7_75t_SL U20771 ( .A1(n20890), .A2(n19002), .B(n20892), .C(
        n19002), .Y(n20893) );
  A2O1A1Ixp33_ASAP7_75t_SL U20772 ( .A1(n30517), .A2(n19002), .B(n18876), .C(
        n20004), .Y(u0_0_leon3x0_p0_iu_fe_pc_15_) );
  A2O1A1Ixp33_ASAP7_75t_SL U20773 ( .A1(n22373), .A2(n19002), .B(n25278), .C(
        n19002), .Y(n20887) );
  A2O1A1Ixp33_ASAP7_75t_SL U20774 ( .A1(u0_0_leon3x0_p0_divi[34]), .A2(n22373), 
        .B(n20887), .C(n19002), .Y(n30445) );
  A2O1A1Ixp33_ASAP7_75t_SL U20775 ( .A1(n22374), .A2(n19002), .B(n28507), .C(
        n19002), .Y(n20882) );
  A2O1A1Ixp33_ASAP7_75t_SL U20776 ( .A1(n18805), .A2(n19002), .B(n32642), .C(
        n19002), .Y(n20883) );
  A2O1A1Ixp33_ASAP7_75t_SL U20777 ( .A1(n22373), .A2(n19002), .B(n29079), .C(
        n19002), .Y(n20884) );
  O2A1O1Ixp5_ASAP7_75t_SL U20778 ( .A1(n20882), .A2(n20883), .B(n19002), .C(
        n20884), .Y(n29081) );
  A2O1A1Ixp33_ASAP7_75t_SL U20779 ( .A1(n32353), .A2(n32343), .B(n19631), .C(
        n19002), .Y(n32436) );
  A2O1A1Ixp33_ASAP7_75t_SL U20780 ( .A1(n27109), .A2(n19002), .B(n27108), .C(
        n19002), .Y(n20878) );
  A2O1A1Ixp33_ASAP7_75t_SL U20781 ( .A1(n28986), .A2(n19002), .B(n27106), .C(
        n19002), .Y(n20879) );
  A2O1A1Ixp33_ASAP7_75t_SL U20782 ( .A1(n28850), .A2(n19002), .B(n27107), .C(
        n19002), .Y(n20880) );
  O2A1O1Ixp5_ASAP7_75t_SL U20783 ( .A1(n20878), .A2(n20879), .B(n19002), .C(
        n20880), .Y(n20881) );
  A2O1A1Ixp33_ASAP7_75t_SL U20784 ( .A1(n28869), .A2(n19002), .B(n28916), .C(
        n20881), .Y(n28761) );
  A2O1A1Ixp33_ASAP7_75t_SL U20785 ( .A1(n19002), .A2(n28301), .B(n31660), .C(
        n20367), .Y(n20368) );
  A2O1A1Ixp33_ASAP7_75t_SL U20786 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[29]), 
        .B(n20368), .C(n19002), .Y(n20369) );
  A2O1A1Ixp33_ASAP7_75t_SL U20787 ( .A1(n19002), .A2(n28324), .B(n31660), .C(
        n20510), .Y(n20511) );
  A2O1A1Ixp33_ASAP7_75t_SL U20788 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[17]), 
        .B(n20511), .C(n19002), .Y(n20512) );
  A2O1A1Ixp33_ASAP7_75t_SL U20789 ( .A1(n18364), .A2(n19002), .B(
        mult_x_1196_n2738), .C(n19002), .Y(n20870) );
  A2O1A1Ixp33_ASAP7_75t_SL U20790 ( .A1(n24040), .A2(n19002), .B(
        mult_x_1196_n2737), .C(n19002), .Y(n20871) );
  A2O1A1Ixp33_ASAP7_75t_SL U20791 ( .A1(n20870), .A2(n19002), .B(n20871), .C(
        n19002), .Y(n20872) );
  A2O1A1Ixp33_ASAP7_75t_SL U20792 ( .A1(n20872), .A2(n19002), .B(
        mult_x_1196_n844), .C(mult_x_1196_n849), .Y(n20873) );
  A2O1A1Ixp33_ASAP7_75t_SL U20793 ( .A1(n24043), .A2(n19002), .B(n20869), .C(
        n19002), .Y(mult_x_1196_n2151) );
  A2O1A1Ixp33_ASAP7_75t_SL U20794 ( .A1(n19002), .A2(mult_x_1196_n2914), .B(
        n18471), .C(n20868), .Y(mult_x_1196_n2343) );
  OAI21xp5_ASAP7_75t_SL U20795 ( .A1(n22781), .A2(mult_x_1196_n2915), .B(
        n19002), .Y(n20867) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20796 ( .A1(n30107), .A2(n30073), .B(n19002), 
        .C(n30134), .Y(n20695) );
  A2O1A1Ixp33_ASAP7_75t_SL U20797 ( .A1(n29632), .A2(n20865), .B(n29627), .C(
        n19002), .Y(n20866) );
  A2O1A1Ixp33_ASAP7_75t_SL U20798 ( .A1(n29628), .A2(n19002), .B(n20866), .C(
        n19002), .Y(n4734) );
  A2O1A1Ixp33_ASAP7_75t_SL U20799 ( .A1(n31727), .A2(n19002), .B(n20846), .C(
        n19002), .Y(n20847) );
  A2O1A1Ixp33_ASAP7_75t_SL U20800 ( .A1(n31728), .A2(n19002), .B(n20848), .C(
        n19002), .Y(n20849) );
  A2O1A1Ixp33_ASAP7_75t_SL U20801 ( .A1(n31721), .A2(n19002), .B(n20850), .C(
        n19002), .Y(n20851) );
  A2O1A1Ixp33_ASAP7_75t_SL U20802 ( .A1(n4724), .A2(n19002), .B(n31740), .C(
        n19002), .Y(n20852) );
  A2O1A1Ixp33_ASAP7_75t_SL U20803 ( .A1(n20858), .A2(n19002), .B(n24695), .C(
        n19002), .Y(n17422) );
  A2O1A1Ixp33_ASAP7_75t_SL U20804 ( .A1(n20843), .A2(n19002), .B(n20844), .C(
        n19002), .Y(n20845) );
  A2O1A1Ixp33_ASAP7_75t_SL U20805 ( .A1(n29949), .A2(n19002), .B(n28249), .C(
        n19002), .Y(n20839) );
  A2O1A1Ixp33_ASAP7_75t_SL U20806 ( .A1(n20839), .A2(n19002), .B(n20842), .C(
        n19002), .Y(n24521) );
  A2O1A1Ixp33_ASAP7_75t_SL U20807 ( .A1(n24428), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__26_), .B(n24680), .C(n19002), .Y(n20833)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20808 ( .A1(n24514), .A2(n19002), .B(n30243), .C(
        n20833), .Y(n20834) );
  A2O1A1Ixp33_ASAP7_75t_SL U20809 ( .A1(u0_0_leon3x0_p0_divi[58]), .A2(n30430), 
        .B(n20834), .C(n19002), .Y(n20835) );
  A2O1A1Ixp33_ASAP7_75t_SL U20810 ( .A1(n26916), .A2(n19002), .B(n30575), .C(
        n19002), .Y(n20831) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20811 ( .A1(n28411), .A2(n31477), .B(n20831), 
        .C(n19002), .D(n30578), .Y(n4594) );
  A2O1A1Ixp33_ASAP7_75t_SL U20812 ( .A1(n29865), .A2(n19002), .B(n29864), .C(
        n19002), .Y(n20821) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20813 ( .A1(u0_0_leon3x0_p0_iu_r_W__RESULT__29_), 
        .A2(n29863), .B(n20821), .C(n19002), .D(n20824), .Y(n20825) );
  A2O1A1Ixp33_ASAP7_75t_SL U20814 ( .A1(n22432), .A2(n29867), .B(n20827), .C(
        n19002), .Y(n20828) );
  A2O1A1Ixp33_ASAP7_75t_SL U20815 ( .A1(n30595), .A2(n19002), .B(n20828), .C(
        n19002), .Y(n20829) );
  A2O1A1Ixp33_ASAP7_75t_SL U20816 ( .A1(n20828), .A2(n30593), .B(n20829), .C(
        n19002), .Y(n20830) );
  A2O1A1Ixp33_ASAP7_75t_SL U20817 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP2__29_), 
        .A2(n20820), .B(n20830), .C(n19002), .Y(n4581) );
  A2O1A1Ixp33_ASAP7_75t_SL U20818 ( .A1(n19002), .A2(n22408), .B(apbi[36]), 
        .C(n20501), .Y(n4546) );
  A2O1A1Ixp33_ASAP7_75t_SL U20819 ( .A1(n30771), .A2(n19002), .B(n29955), .C(
        n19002), .Y(n20819) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20820 ( .A1(n29959), .A2(uart1_r_RSHIFT__5_), 
        .B(n20819), .C(n19002), .D(n29958), .Y(n4541) );
  A2O1A1Ixp33_ASAP7_75t_SL U20821 ( .A1(n31678), .A2(n19002), .B(n31677), .C(
        n19002), .Y(n20672) );
  A2O1A1Ixp33_ASAP7_75t_SL U20822 ( .A1(n31526), .A2(n19002), .B(n22397), .C(
        n19002), .Y(n20818) );
  A2O1A1Ixp33_ASAP7_75t_SL U20823 ( .A1(n24646), .A2(n19002), .B(n31350), .C(
        n20817), .Y(n4149) );
  A2O1A1Ixp33_ASAP7_75t_SL U20824 ( .A1(n19002), .A2(n24646), .B(n31875), .C(
        n20649), .Y(n4137) );
  A2O1A1Ixp33_ASAP7_75t_SL U20825 ( .A1(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__31_), .A2(n19002), .B(n24657), .C(
        n20816), .Y(n4063) );
  A2O1A1Ixp33_ASAP7_75t_SL U20826 ( .A1(n25004), .A2(n19002), .B(n25003), .C(
        n26810), .Y(n20812) );
  A2O1A1Ixp33_ASAP7_75t_SL U20827 ( .A1(n20812), .A2(n19002), .B(n20813), .C(
        n19002), .Y(n20814) );
  A2O1A1Ixp33_ASAP7_75t_SL U20828 ( .A1(n24649), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__4_), .B(n20814), .C(n19002), .Y(
        n4059) );
  A2O1A1Ixp33_ASAP7_75t_SL U20829 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__4_), .B(n24651), .C(n20627), .Y(
        n3464) );
  A2O1A1Ixp33_ASAP7_75t_SL U20830 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__11_), 
        .A2(n19002), .B(n24653), .C(n20796), .Y(n3410) );
  A2O1A1Ixp33_ASAP7_75t_SL U20831 ( .A1(n19002), .A2(n24646), .B(rf_di_w[26]), 
        .C(n20450), .Y(n3254) );
  A2O1A1Ixp33_ASAP7_75t_SL U20832 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__14_), 
        .A2(n19002), .B(n24650), .C(n20793), .Y(n3210) );
  A2O1A1Ixp33_ASAP7_75t_SL U20833 ( .A1(n24646), .A2(n19002), .B(n32679), .C(
        n20791), .Y(n3190) );
  A2O1A1Ixp33_ASAP7_75t_SL U20834 ( .A1(n30382), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n20789) );
  A2O1A1Ixp33_ASAP7_75t_SL U20835 ( .A1(n30696), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n20790) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20836 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__11_), 
        .A2(n31403), .B(n20789), .C(n19002), .D(n20790), .Y(n3144) );
  A2O1A1Ixp33_ASAP7_75t_SL U20837 ( .A1(n22427), .A2(n19002), .B(rf_di_w[7]), 
        .C(n20784), .Y(n3031) );
  A2O1A1Ixp33_ASAP7_75t_SL U20838 ( .A1(n19002), .A2(n22427), .B(rf_di_w[15]), 
        .C(n20612), .Y(n3020) );
  A2O1A1Ixp33_ASAP7_75t_SL U20839 ( .A1(n19002), .A2(n31198), .B(
        sr1_r_MCFG2__RAMBANKSZ__3_), .C(n20610), .Y(n2913) );
  A2O1A1Ixp33_ASAP7_75t_SL U20840 ( .A1(n32169), .A2(n19002), .B(n32168), .C(
        n19002), .Y(n20772) );
  A2O1A1Ixp33_ASAP7_75t_SL U20841 ( .A1(n20772), .A2(n19002), .B(n20773), .C(
        n19002), .Y(n20774) );
  A2O1A1Ixp33_ASAP7_75t_SL U20842 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_A__RFA2__6_), .C(n20775), .Y(n2780) );
  A2O1A1Ixp33_ASAP7_75t_SL U20843 ( .A1(n19002), .A2(n30370), .B(n22414), .C(
        n20607), .Y(n20608) );
  A2O1A1Ixp33_ASAP7_75t_SL U20844 ( .A1(n31403), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__12_), .B(n20608), .C(n19002), .Y(n2680)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U20845 ( .A1(n22420), .A2(n19002), .B(n27222), .C(
        n31422), .Y(n20765) );
  A2O1A1Ixp33_ASAP7_75t_SL U20846 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[13]), 
        .B(n20765), .C(n19002), .Y(n20766) );
  A2O1A1Ixp33_ASAP7_75t_SL U20847 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_13_), .B(n20768), .C(n19002), .Y(n2659) );
  A2O1A1Ixp33_ASAP7_75t_SL U20848 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__13_), .B(n22428), .C(n20604), .Y(
        n2647) );
  A2O1A1Ixp33_ASAP7_75t_SL U20849 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__22_), 
        .A2(n19002), .B(n22428), .C(n20761), .Y(n2496) );
  A2O1A1Ixp33_ASAP7_75t_SL U20850 ( .A1(n27508), .A2(n19853), .B(n19858), .C(
        n19002), .Y(n2459) );
  A2O1A1Ixp33_ASAP7_75t_SL U20851 ( .A1(n19002), .A2(n22433), .B(n32946), .C(
        n20591), .Y(n1715) );
  A2O1A1Ixp33_ASAP7_75t_SL U20852 ( .A1(dataout[11]), .A2(n19002), .B(n20757), 
        .C(n19002), .Y(n20758) );
  A2O1A1Ixp33_ASAP7_75t_SL U20853 ( .A1(n32660), .A2(n19002), .B(n32622), .C(
        n20755), .Y(ic_data[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20854 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__30_), .A2(n19002), .B(n32565), .C(n19002), .Y(n20752) );
  A2O1A1Ixp33_ASAP7_75t_SL U20855 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[30]), 
        .A2(n19002), .B(n32593), .C(n19002), .Y(n20753) );
  O2A1O1Ixp33_ASAP7_75t_SL U20856 ( .A1(n32559), .A2(n20752), .B(n19002), .C(
        n20753), .Y(it_data[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20857 ( .A1(n32636), .A2(n19002), .B(n32543), .C(
        n20751), .Y(it_data[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20858 ( .A1(n32652), .A2(n19002), .B(n32429), .C(
        n20745), .Y(n20746) );
  A2O1A1Ixp33_ASAP7_75t_SL U20859 ( .A1(n32434), .A2(n32403), .B(n20746), .C(
        n19002), .Y(n20747) );
  A2O1A1Ixp33_ASAP7_75t_SL U20860 ( .A1(n32402), .A2(n19002), .B(n32431), .C(
        n20747), .Y(n20748) );
  A2O1A1Ixp33_ASAP7_75t_SL U20861 ( .A1(n33069), .A2(dc_q[27]), .B(n20748), 
        .C(n19002), .Y(n20749) );
  A2O1A1Ixp33_ASAP7_75t_SL U20862 ( .A1(n32425), .A2(n19002), .B(n32404), .C(
        n20749), .Y(dc_data[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20863 ( .A1(n30725), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__PC__9_), .B(n20730), .C(n19002), .Y(
        n20731) );
  A2O1A1Ixp33_ASAP7_75t_SL U20864 ( .A1(n27472), .A2(n19002), .B(n27471), .C(
        n19002), .Y(n20726) );
  A2O1A1Ixp33_ASAP7_75t_SL U20865 ( .A1(n22374), .A2(n19002), .B(n28334), .C(
        n19002), .Y(n20723) );
  A2O1A1Ixp33_ASAP7_75t_SL U20866 ( .A1(n18806), .A2(n19002), .B(n32626), .C(
        n19002), .Y(n20724) );
  A2O1A1Ixp33_ASAP7_75t_SL U20867 ( .A1(n22373), .A2(n19002), .B(n29096), .C(
        n19002), .Y(n20725) );
  O2A1O1Ixp5_ASAP7_75t_SL U20868 ( .A1(n20723), .A2(n20724), .B(n19002), .C(
        n20725), .Y(n30496) );
  A2O1A1Ixp33_ASAP7_75t_SL U20869 ( .A1(add_x_746_n92), .A2(n19002), .B(n20720), .C(n19002), .Y(n20721) );
  A2O1A1Ixp33_ASAP7_75t_SL U20870 ( .A1(add_x_746_n125), .A2(n19002), .B(
        n20722), .C(n19002), .Y(add_x_746_n1) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20871 ( .A1(n28405), .A2(n28736), .B(n26509), 
        .C(n19002), .D(n20719), .Y(n32392) );
  A2O1A1Ixp33_ASAP7_75t_SL U20872 ( .A1(n22373), .A2(n19002), .B(n25285), .C(
        n19002), .Y(n20715) );
  A2O1A1Ixp33_ASAP7_75t_SL U20873 ( .A1(u0_0_leon3x0_p0_divi[40]), .A2(n22373), 
        .B(n20715), .C(n19002), .Y(n30391) );
  A2O1A1Ixp33_ASAP7_75t_SL U20874 ( .A1(u0_0_leon3x0_p0_dci[38]), .A2(n19002), 
        .B(n20713), .C(n19002), .Y(n20714) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20875 ( .A1(n25585), .A2(n20714), .B(n25584), 
        .C(n19002), .D(n32280), .Y(n31457) );
  A2O1A1Ixp33_ASAP7_75t_SL U20876 ( .A1(n22373), .A2(n19002), .B(n25273), .C(
        n20712), .Y(n30452) );
  A2O1A1Ixp33_ASAP7_75t_SL U20877 ( .A1(n22373), .A2(n19002), .B(n25281), .C(
        n19002), .Y(n20711) );
  A2O1A1Ixp33_ASAP7_75t_SL U20878 ( .A1(u0_0_leon3x0_p0_divi[37]), .A2(n22373), 
        .B(n20711), .C(n19002), .Y(n30412) );
  A2O1A1Ixp33_ASAP7_75t_SL U20879 ( .A1(n22374), .A2(n19002), .B(n28749), .C(
        n19002), .Y(n20708) );
  A2O1A1Ixp33_ASAP7_75t_SL U20880 ( .A1(n18805), .A2(n19002), .B(n32614), .C(
        n19002), .Y(n20709) );
  A2O1A1Ixp33_ASAP7_75t_SL U20881 ( .A1(n22373), .A2(n19002), .B(n29100), .C(
        n19002), .Y(n20710) );
  O2A1O1Ixp5_ASAP7_75t_SL U20882 ( .A1(n20708), .A2(n20709), .B(n19002), .C(
        n20710), .Y(n29932) );
  A2O1A1Ixp33_ASAP7_75t_SL U20883 ( .A1(n22374), .A2(n19002), .B(n28327), .C(
        n19002), .Y(n20705) );
  A2O1A1Ixp33_ASAP7_75t_SL U20884 ( .A1(n18805), .A2(n19002), .B(n32632), .C(
        n19002), .Y(n20706) );
  A2O1A1Ixp33_ASAP7_75t_SL U20885 ( .A1(n22373), .A2(n19002), .B(n27265), .C(
        n19002), .Y(n20707) );
  O2A1O1Ixp5_ASAP7_75t_SL U20886 ( .A1(n20705), .A2(n20706), .B(n19002), .C(
        n20707), .Y(n27267) );
  A2O1A1Ixp33_ASAP7_75t_SL U20887 ( .A1(n32353), .A2(n19002), .B(n32624), .C(
        n20703), .Y(n32413) );
  A2O1A1Ixp33_ASAP7_75t_SL U20888 ( .A1(n32353), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[2]), .C(n20702), .Y(n32398) );
  A2O1A1Ixp33_ASAP7_75t_SL U20889 ( .A1(n22373), .A2(n19002), .B(n25286), .C(
        n20701), .Y(n27147) );
  A2O1A1Ixp33_ASAP7_75t_SL U20890 ( .A1(n18891), .A2(n19002), .B(n28720), .C(
        n19002), .Y(n20699) );
  A2O1A1Ixp33_ASAP7_75t_SL U20891 ( .A1(n28769), .A2(n19002), .B(
        u0_0_leon3x0_p0_muli[18]), .C(n19002), .Y(n20700) );
  A2O1A1Ixp33_ASAP7_75t_SL U20892 ( .A1(n20699), .A2(n19002), .B(n20700), .C(
        n19002), .Y(u0_0_leon3x0_p0_divi[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20893 ( .A1(n26009), .A2(n19002), .B(n20698), .C(
        n19002), .Y(n26045) );
  A2O1A1Ixp33_ASAP7_75t_SL U20894 ( .A1(n19002), .A2(n28310), .B(n31660), .C(
        n19986), .Y(n19987) );
  A2O1A1Ixp33_ASAP7_75t_SL U20895 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[23]), 
        .B(n19987), .C(n19002), .Y(n19988) );
  A2O1A1Ixp33_ASAP7_75t_SL U20896 ( .A1(n19002), .A2(n28323), .B(n31660), .C(
        n20158), .Y(n20159) );
  A2O1A1Ixp33_ASAP7_75t_SL U20897 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[18]), 
        .B(n20159), .C(n19002), .Y(n20160) );
  O2A1O1Ixp33_ASAP7_75t_SL U20898 ( .A1(n20870), .A2(mult_x_1196_n844), .B(
        n19002), .C(n20871), .Y(n20505) );
  A2O1A1Ixp33_ASAP7_75t_SL U20899 ( .A1(n19002), .A2(n20871), .B(n20870), .C(
        mult_x_1196_n844), .Y(n20507) );
  A2O1A1Ixp33_ASAP7_75t_SL U20900 ( .A1(n31718), .A2(n20141), .B(sr1_r_WS__0_), 
        .C(n19002), .Y(n20142) );
  A2O1A1Ixp33_ASAP7_75t_SL U20901 ( .A1(sr1_r_MCFG1__ROMRWS__0_), .A2(n31726), 
        .B(n20148), .C(n19002), .Y(n20149) );
  A2O1A1Ixp33_ASAP7_75t_SL U20902 ( .A1(n28030), .A2(n27915), .B(n20362), .C(
        n19002), .Y(n4702) );
  A2O1A1Ixp33_ASAP7_75t_SL U20903 ( .A1(apbi[13]), .A2(n19002), .B(n29745), 
        .C(n19002), .Y(n20689) );
  A2O1A1Ixp33_ASAP7_75t_SL U20904 ( .A1(n29745), .A2(n19002), .B(
        irqctrl0_r_IPEND__13_), .C(n19002), .Y(n20691) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20905 ( .A1(n29238), .A2(n20690), .B(n20691), 
        .C(n19002), .D(n24695), .Y(n20692) );
  A2O1A1Ixp33_ASAP7_75t_SL U20906 ( .A1(n30705), .A2(n24662), .B(n20685), .C(
        n19002), .Y(n20686) );
  A2O1A1Ixp33_ASAP7_75t_SL U20907 ( .A1(n30704), .A2(n19002), .B(n30703), .C(
        n19002), .Y(n20687) );
  A2O1A1Ixp33_ASAP7_75t_SL U20908 ( .A1(n22408), .A2(n19002), .B(apbi[44]), 
        .C(n20684), .Y(n4597) );
  A2O1A1Ixp33_ASAP7_75t_SL U20909 ( .A1(n24681), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_E__OP1__22_), .C(n19002), .Y(n20680) );
  A2O1A1Ixp33_ASAP7_75t_SL U20910 ( .A1(n31540), .A2(n31542), .B(n20680), .C(
        n19002), .Y(n20681) );
  A2O1A1Ixp33_ASAP7_75t_SL U20911 ( .A1(n31359), .A2(n19002), .B(n31045), .C(
        n19002), .Y(n20676) );
  O2A1O1Ixp33_ASAP7_75t_SL U20912 ( .A1(n20676), .A2(n31047), .B(n19002), .C(
        n20679), .Y(n4557) );
  A2O1A1Ixp33_ASAP7_75t_SL U20913 ( .A1(n28224), .A2(n19002), .B(n29955), .C(
        n19002), .Y(n20675) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20914 ( .A1(n29959), .A2(uart1_r_RSHIFT__4_), 
        .B(n20675), .C(n19002), .D(n29958), .Y(n4540) );
  A2O1A1Ixp33_ASAP7_75t_SL U20915 ( .A1(n31676), .A2(n19002), .B(n31675), .C(
        n20668), .Y(n20669) );
  A2O1A1Ixp33_ASAP7_75t_SL U20916 ( .A1(n19002), .A2(n20671), .B(n20672), .C(
        n19002), .Y(n20673) );
  A2O1A1Ixp33_ASAP7_75t_SL U20917 ( .A1(n30590), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n20656) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20918 ( .A1(n30591), .A2(n30644), .B(n20656), 
        .C(n19002), .D(n20659), .Y(n20660) );
  A2O1A1Ixp33_ASAP7_75t_SL U20919 ( .A1(n30645), .A2(n19002), .B(n30592), .C(
        n20660), .Y(n20661) );
  A2O1A1Ixp33_ASAP7_75t_SL U20920 ( .A1(n30597), .A2(n22432), .B(n20661), .C(
        n19002), .Y(n20662) );
  A2O1A1Ixp33_ASAP7_75t_SL U20921 ( .A1(n30594), .A2(n19002), .B(n23229), .C(
        n19002), .Y(n20664) );
  A2O1A1Ixp33_ASAP7_75t_SL U20922 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__10_), .B(n19354), .C(n19002), .Y(n19355) );
  A2O1A1Ixp33_ASAP7_75t_SL U20923 ( .A1(n19002), .A2(n31412), .B(n30387), .C(
        n19355), .Y(n19356) );
  A2O1A1Ixp33_ASAP7_75t_SL U20924 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_), .B(n24654), .C(n20474), .Y(
        n4153) );
  A2O1A1Ixp33_ASAP7_75t_SL U20925 ( .A1(n27522), .A2(n19002), .B(n20643), .C(
        n20644), .Y(n20645) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20926 ( .A1(n31940), .A2(n27521), .B(n30980), 
        .C(n19002), .D(n27522), .Y(n20646) );
  A2O1A1Ixp33_ASAP7_75t_SL U20927 ( .A1(n29978), .A2(n20647), .B(n27524), .C(
        n19002), .Y(n20648) );
  A2O1A1Ixp33_ASAP7_75t_SL U20928 ( .A1(n29985), .A2(n20645), .B(n20648), .C(
        n19002), .Y(n4071) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20929 ( .A1(n30680), .A2(n30682), .B(n19002), 
        .C(n30681), .Y(n19730) );
  A2O1A1Ixp33_ASAP7_75t_SL U20930 ( .A1(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__30_), .A2(n19002), .B(n24657), .C(
        n20639), .Y(n3887) );
  A2O1A1Ixp33_ASAP7_75t_SL U20931 ( .A1(n19002), .A2(n22379), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__1_), .C(n20462), .Y(n3854) );
  A2O1A1Ixp33_ASAP7_75t_SL U20932 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_), .A2(n19002), .B(n24655), .C(
        n20637), .Y(n3775) );
  A2O1A1Ixp33_ASAP7_75t_SL U20933 ( .A1(n26195), .A2(n19002), .B(n24981), .C(
        n19002), .Y(n20635) );
  A2O1A1Ixp33_ASAP7_75t_SL U20934 ( .A1(n22379), .A2(n19002), .B(n25050), .C(
        n19002), .Y(n20636) );
  A2O1A1Ixp33_ASAP7_75t_SL U20935 ( .A1(n20635), .A2(n19002), .B(n20636), .C(
        n19002), .Y(n3580) );
  A2O1A1Ixp33_ASAP7_75t_SL U20936 ( .A1(n31873), .A2(n19002), .B(n31874), .C(
        n19002), .Y(n20631) );
  A2O1A1Ixp33_ASAP7_75t_SL U20937 ( .A1(n31872), .A2(n19002), .B(n20632), .C(
        n19002), .Y(n20633) );
  A2O1A1Ixp33_ASAP7_75t_SL U20938 ( .A1(n20631), .A2(n19002), .B(n20633), .C(
        n20634), .Y(n3566) );
  A2O1A1Ixp33_ASAP7_75t_SL U20939 ( .A1(n19002), .A2(n32057), .B(n29177), .C(
        n23229), .Y(n19875) );
  A2O1A1Ixp33_ASAP7_75t_SL U20940 ( .A1(n19002), .A2(n23229), .B(
        u0_0_leon3x0_p0_iu_r_A__TICC_), .C(n19875), .Y(n3556) );
  A2O1A1Ixp33_ASAP7_75t_SL U20941 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_W__S__WIM__2_), .C(n20623), .Y(n3336) );
  A2O1A1Ixp33_ASAP7_75t_SL U20942 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__29_), 
        .A2(n19002), .B(n24650), .C(n20622), .Y(n3286) );
  A2O1A1Ixp33_ASAP7_75t_SL U20943 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[30]), 
        .B(n24653), .C(n20449), .Y(n3198) );
  A2O1A1Ixp33_ASAP7_75t_SL U20944 ( .A1(n22427), .A2(n19002), .B(n32587), .C(
        n20618), .Y(n3178) );
  A2O1A1Ixp33_ASAP7_75t_SL U20945 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[25]), .C(n20614), .Y(n3113) );
  A2O1A1Ixp33_ASAP7_75t_SL U20946 ( .A1(n19002), .A2(n22427), .B(rf_di_w[11]), 
        .C(n20438), .Y(n3025) );
  A2O1A1Ixp33_ASAP7_75t_SL U20947 ( .A1(n32673), .A2(n19002), .B(n32674), .C(
        n32682), .Y(n20611) );
  A2O1A1Ixp33_ASAP7_75t_SL U20948 ( .A1(n22405), .A2(n19002), .B(n20611), .C(
        n32675), .Y(u0_0_leon3x0_p0_c0mmu_icache0_v_VADDRESS__3_) );
  A2O1A1Ixp33_ASAP7_75t_SL U20949 ( .A1(n28167), .A2(uart1_uarto_SCALER__6_), 
        .B(n22419), .C(n19002), .Y(n20299) );
  A2O1A1Ixp33_ASAP7_75t_SL U20950 ( .A1(n19002), .A2(n24633), .B(
        uart1_r_RIRQEN_), .C(n20061), .Y(n2857) );
  A2O1A1Ixp33_ASAP7_75t_SL U20951 ( .A1(n19002), .A2(n24646), .B(n31424), .C(
        n20437), .Y(n2808) );
  A2O1A1Ixp33_ASAP7_75t_SL U20952 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_W__S__CWP__2_), .C(n20609), .Y(n2684) );
  A2O1A1Ixp33_ASAP7_75t_SL U20953 ( .A1(n22427), .A2(n19002), .B(n28601), .C(
        n20605), .Y(n2657) );
  A2O1A1Ixp33_ASAP7_75t_SL U20954 ( .A1(n32733), .A2(n19002), .B(n32732), .C(
        n19002), .Y(n20599) );
  A2O1A1Ixp33_ASAP7_75t_SL U20955 ( .A1(n20595), .A2(n19002), .B(n20596), .C(
        n19002), .Y(n20597) );
  A2O1A1Ixp33_ASAP7_75t_SL U20956 ( .A1(dataout[3]), .A2(n19002), .B(n20589), 
        .C(n19002), .Y(n20590) );
  A2O1A1Ixp33_ASAP7_75t_SL U20957 ( .A1(dataout[12]), .A2(n19002), .B(n20586), 
        .C(n19002), .Y(n20587) );
  A2O1A1Ixp33_ASAP7_75t_SL U20958 ( .A1(n31452), .A2(n19002), .B(n32443), .C(
        n19002), .Y(n20585) );
  A2O1A1Ixp33_ASAP7_75t_SL U20959 ( .A1(n25513), .A2(n19002), .B(n20585), .C(
        n19002), .Y(n31570) );
  A2O1A1Ixp33_ASAP7_75t_SL U20960 ( .A1(n19002), .A2(n32660), .B(n32618), .C(
        n20430), .Y(ic_data[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20961 ( .A1(n19002), .A2(n32660), .B(n32610), .C(
        n20429), .Y(ic_data[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20962 ( .A1(n32634), .A2(n19002), .B(n32543), .C(
        n20583), .Y(it_data[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U20963 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__0_), .A2(n19002), .B(n32427), 
        .C(n19002), .Y(n20570) );
  A2O1A1Ixp33_ASAP7_75t_SL U20964 ( .A1(n32436), .A2(n19002), .B(n20570), .C(
        n19002), .Y(n20571) );
  A2O1A1Ixp33_ASAP7_75t_SL U20965 ( .A1(n32428), .A2(n19002), .B(
        u0_0_leon3x0_p0_dci[4]), .C(n19002), .Y(n20573) );
  O2A1O1Ixp33_ASAP7_75t_SL U20966 ( .A1(n32435), .A2(n20572), .B(n19002), .C(
        n20573), .Y(n20574) );
  A2O1A1Ixp33_ASAP7_75t_SL U20967 ( .A1(n32430), .A2(n19002), .B(n24543), .C(
        n19002), .Y(n20578) );
  A2O1A1Ixp33_ASAP7_75t_SL U20968 ( .A1(n20577), .A2(n19002), .B(n20578), .C(
        n19002), .Y(n20579) );
  A2O1A1Ixp33_ASAP7_75t_SL U20969 ( .A1(n32434), .A2(n32433), .B(n20580), .C(
        n19002), .Y(n20581) );
  A2O1A1Ixp33_ASAP7_75t_SL U20970 ( .A1(n28725), .A2(n19002), .B(n29909), .C(
        n28748), .Y(n20562) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20971 ( .A1(n28736), .A2(n28132), .B(n26509), 
        .C(n19002), .D(n20562), .Y(n32320) );
  A2O1A1Ixp33_ASAP7_75t_SL U20972 ( .A1(n23887), .A2(n19002), .B(n20557), .C(
        n19002), .Y(n20558) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U20973 ( .A1(DP_OP_5187J1_124_3275_n213), .A2(
        DP_OP_5187J1_124_3275_n232), .B(n20558), .C(n19002), .D(
        DP_OP_5187J1_124_3275_n214), .Y(n20559) );
  A2O1A1Ixp33_ASAP7_75t_SL U20974 ( .A1(n22373), .A2(n19002), .B(n25315), .C(
        n20556), .Y(n30244) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20975 ( .A1(add_x_746_n47), .A2(add_x_746_n59), 
        .B(n19002), .C(n20555), .Y(add_x_746_n41) );
  A2O1A1Ixp33_ASAP7_75t_SL U20976 ( .A1(n22374), .A2(n19002), .B(n28304), .C(
        n19002), .Y(n20552) );
  A2O1A1Ixp33_ASAP7_75t_SL U20977 ( .A1(n18806), .A2(n19002), .B(n32652), .C(
        n19002), .Y(n20553) );
  A2O1A1Ixp33_ASAP7_75t_SL U20978 ( .A1(n22373), .A2(n19002), .B(n26912), .C(
        n19002), .Y(n20554) );
  O2A1O1Ixp5_ASAP7_75t_SL U20979 ( .A1(n20552), .A2(n20553), .B(n19002), .C(
        n20554), .Y(n26953) );
  A2O1A1Ixp33_ASAP7_75t_SL U20980 ( .A1(n19002), .A2(n31786), .B(n18876), .C(
        n20190), .Y(u0_0_leon3x0_p0_iu_fe_pc_27_) );
  A2O1A1Ixp33_ASAP7_75t_SL U20981 ( .A1(n22376), .A2(n19002), .B(n30277), .C(
        n20551), .Y(n28521) );
  A2O1A1Ixp33_ASAP7_75t_SL U20982 ( .A1(n31895), .A2(n31896), .B(n20549), .C(
        n19002), .Y(n32128) );
  A2O1A1Ixp33_ASAP7_75t_SL U20983 ( .A1(mult_x_1196_n524), .A2(
        mult_x_1196_n552), .B(mult_x_1196_n525), .C(n19002), .Y(n20548) );
  A2O1A1Ixp33_ASAP7_75t_SL U20984 ( .A1(n19002), .A2(mult_x_1196_n580), .B(
        n20547), .C(n20548), .Y(n18448) );
  A2O1A1Ixp33_ASAP7_75t_SL U20985 ( .A1(n22374), .A2(n19002), .B(n28323), .C(
        n19002), .Y(n20544) );
  A2O1A1Ixp33_ASAP7_75t_SL U20986 ( .A1(n18806), .A2(n19002), .B(n32636), .C(
        n19002), .Y(n20545) );
  A2O1A1Ixp33_ASAP7_75t_SL U20987 ( .A1(n22373), .A2(n19002), .B(n29092), .C(
        n19002), .Y(n20546) );
  O2A1O1Ixp5_ASAP7_75t_SL U20988 ( .A1(n20544), .A2(n20545), .B(n19002), .C(
        n20546), .Y(n30821) );
  A2O1A1Ixp33_ASAP7_75t_SL U20989 ( .A1(n29887), .A2(n31868), .B(n19647), .C(
        n19002), .Y(n19648) );
  A2O1A1Ixp33_ASAP7_75t_SL U20990 ( .A1(n22374), .A2(n19002), .B(n28356), .C(
        n19002), .Y(n20541) );
  A2O1A1Ixp33_ASAP7_75t_SL U20991 ( .A1(n18806), .A2(n19002), .B(n32608), .C(
        n19002), .Y(n20542) );
  A2O1A1Ixp33_ASAP7_75t_SL U20992 ( .A1(n22373), .A2(n19002), .B(n29102), .C(
        n19002), .Y(n20543) );
  O2A1O1Ixp5_ASAP7_75t_SL U20993 ( .A1(n20541), .A2(n20542), .B(n19002), .C(
        n20543), .Y(n29693) );
  A2O1A1Ixp33_ASAP7_75t_SL U20994 ( .A1(u0_0_leon3x0_p0_iu_r_M__CTRL__RETT_), 
        .A2(n19002), .B(u0_0_leon3x0_p0_iu_r_E__CTRL__RETT_), .C(n19002), .Y(
        n20537) );
  A2O1A1Ixp33_ASAP7_75t_SL U20995 ( .A1(u0_0_leon3x0_p0_iu_r_A__CTRL__RETT_), 
        .A2(n19002), .B(u0_0_leon3x0_p0_iu_r_X__CTRL__RETT_), .C(n19002), .Y(
        n20538) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U20996 ( .A1(add_x_746_n92), .A2(add_x_746_n104), 
        .B(n19002), .C(n20535), .Y(add_x_746_n86) );
  A2O1A1Ixp33_ASAP7_75t_SL U20997 ( .A1(n22374), .A2(n19002), .B(n28310), .C(
        n19002), .Y(n20532) );
  A2O1A1Ixp33_ASAP7_75t_SL U20998 ( .A1(n18805), .A2(n19002), .B(n32646), .C(
        n19002), .Y(n20533) );
  A2O1A1Ixp33_ASAP7_75t_SL U20999 ( .A1(n22373), .A2(n19002), .B(n29088), .C(
        n19002), .Y(n20534) );
  O2A1O1Ixp5_ASAP7_75t_SL U21000 ( .A1(n20532), .A2(n20533), .B(n19002), .C(
        n20534), .Y(n29768) );
  O2A1O1Ixp33_ASAP7_75t_SL U21001 ( .A1(n32255), .A2(n20529), .B(n19002), .C(
        n20530), .Y(n32444) );
  A2O1A1Ixp33_ASAP7_75t_SL U21002 ( .A1(n32353), .A2(n32342), .B(n20177), .C(
        n19002), .Y(n32426) );
  A2O1A1Ixp33_ASAP7_75t_SL U21003 ( .A1(n32353), .A2(n32336), .B(n20175), .C(
        n19002), .Y(n32407) );
  A2O1A1Ixp33_ASAP7_75t_SL U21004 ( .A1(n32332), .A2(n19002), .B(n24642), .C(
        n19002), .Y(n20528) );
  A2O1A1Ixp33_ASAP7_75t_SL U21005 ( .A1(n24642), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[11]), .B(n20528), .C(n19002), .Y(n32404)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21006 ( .A1(n32353), .A2(n32300), .B(n19630), .C(
        n19002), .Y(n32396) );
  A2O1A1Ixp33_ASAP7_75t_SL U21007 ( .A1(n28967), .A2(n26258), .B(n20520), .C(
        n19002), .Y(n20521) );
  A2O1A1Ixp33_ASAP7_75t_SL U21008 ( .A1(n19002), .A2(n28507), .B(n31660), .C(
        n19784), .Y(n19785) );
  A2O1A1Ixp33_ASAP7_75t_SL U21009 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[21]), 
        .B(n19785), .C(n19002), .Y(n19786) );
  A2O1A1Ixp33_ASAP7_75t_SL U21010 ( .A1(n20502), .A2(n19002), .B(n20503), .C(
        n20504), .Y(n4736) );
  O2A1O1Ixp5_ASAP7_75t_SL U21011 ( .A1(n20132), .A2(n20133), .B(n19002), .C(
        n20135), .Y(n4668) );
  A2O1A1Ixp33_ASAP7_75t_SL U21012 ( .A1(n19002), .A2(n22421), .B(n29728), .C(
        n29885), .Y(n20357) );
  O2A1O1Ixp5_ASAP7_75t_SL U21013 ( .A1(n31050), .A2(n31048), .B(n19002), .C(
        n32110), .Y(n20124) );
  A2O1A1Ixp33_ASAP7_75t_SL U21014 ( .A1(n29555), .A2(n19002), .B(n29955), .C(
        n19002), .Y(n20500) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21015 ( .A1(n29959), .A2(uart1_r_RSHIFT__3_), 
        .B(n20500), .C(n19002), .D(n29958), .Y(n4539) );
  A2O1A1Ixp33_ASAP7_75t_SL U21016 ( .A1(n26514), .A2(n19002), .B(n30575), .C(
        n19002), .Y(n20499) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21017 ( .A1(n28411), .A2(n30479), .B(n20499), 
        .C(n19002), .D(n30578), .Y(n4511) );
  A2O1A1Ixp33_ASAP7_75t_SL U21018 ( .A1(n29865), .A2(n19002), .B(n26734), .C(
        n19002), .Y(n20489) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21019 ( .A1(u0_0_leon3x0_p0_iu_r_W__RESULT__31_), 
        .A2(n29863), .B(n20489), .C(n19002), .D(n20492), .Y(n20493) );
  A2O1A1Ixp33_ASAP7_75t_SL U21020 ( .A1(n22432), .A2(n26735), .B(n20495), .C(
        n19002), .Y(n20496) );
  A2O1A1Ixp33_ASAP7_75t_SL U21021 ( .A1(n30595), .A2(n19002), .B(n20496), .C(
        n19002), .Y(n20497) );
  A2O1A1Ixp33_ASAP7_75t_SL U21022 ( .A1(n20496), .A2(n30593), .B(n20497), .C(
        n19002), .Y(n20498) );
  A2O1A1Ixp33_ASAP7_75t_SL U21023 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP2__31_), 
        .A2(n20488), .B(n20498), .C(n19002), .Y(n4505) );
  A2O1A1Ixp33_ASAP7_75t_SL U21024 ( .A1(n24638), .A2(n19002), .B(n20481), .C(
        n19002), .Y(n20482) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21025 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__8_), .B(n24679), .C(n19002), .D(n20482), 
        .Y(n20483) );
  A2O1A1Ixp33_ASAP7_75t_SL U21026 ( .A1(n30426), .A2(n19002), .B(n30396), .C(
        n20486), .Y(n20487) );
  A2O1A1Ixp33_ASAP7_75t_SL U21027 ( .A1(u0_0_leon3x0_p0_divi[39]), .A2(n19002), 
        .B(n23229), .C(n20487), .Y(n4441) );
  A2O1A1Ixp33_ASAP7_75t_SL U21028 ( .A1(n26530), .A2(n19002), .B(n22397), .C(
        n19002), .Y(n20479) );
  A2O1A1Ixp33_ASAP7_75t_SL U21029 ( .A1(n22420), .A2(n19002), .B(n28276), .C(
        n31422), .Y(n20475) );
  A2O1A1Ixp33_ASAP7_75t_SL U21030 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[27]), 
        .B(n20475), .C(n19002), .Y(n20476) );
  A2O1A1Ixp33_ASAP7_75t_SL U21031 ( .A1(n31679), .A2(
        u0_0_leon3x0_p0_div0_addout_27_), .B(n20478), .C(n19002), .Y(n4399) );
  A2O1A1Ixp33_ASAP7_75t_SL U21032 ( .A1(n19002), .A2(n22427), .B(n20334), .C(
        n20335), .Y(n4301) );
  A2O1A1Ixp33_ASAP7_75t_SL U21033 ( .A1(n22427), .A2(n19002), .B(n30820), .C(
        n20473), .Y(n4135) );
  A2O1A1Ixp33_ASAP7_75t_SL U21034 ( .A1(n22379), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__2_), .C(n19725), .Y(n3946) );
  A2O1A1Ixp33_ASAP7_75t_SL U21035 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_), .A2(n19002), .B(n32123), 
        .C(n20464), .Y(n3879) );
  A2O1A1Ixp33_ASAP7_75t_SL U21036 ( .A1(n18842), .A2(n19002), .B(n24658), .C(
        n20463), .Y(n3875) );
  A2O1A1Ixp33_ASAP7_75t_SL U21037 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__26_), .B(n24655), .C(n19135), .Y(
        n3764) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21038 ( .A1(n24646), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__ET_), .B(n19002), .C(n32077), .Y(n20459) );
  A2O1A1Ixp33_ASAP7_75t_SL U21039 ( .A1(n20459), .A2(n19002), .B(n20460), .C(
        n19002), .Y(n20461) );
  A2O1A1Ixp33_ASAP7_75t_SL U21040 ( .A1(n32076), .A2(n19002), .B(n20461), .C(
        n19002), .Y(n18277) );
  A2O1A1Ixp33_ASAP7_75t_SL U21041 ( .A1(n3727), .A2(n19002), .B(n22379), .C(
        n19002), .Y(n20457) );
  A2O1A1Ixp33_ASAP7_75t_SL U21042 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__8_), .B(n24656), .C(n19316), .Y(
        n3664) );
  A2O1A1Ixp33_ASAP7_75t_SL U21043 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__14_), .B(n24649), .C(n19716), .Y(
        n3616) );
  A2O1A1Ixp33_ASAP7_75t_SL U21044 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__4_), .B(n24650), .C(n19708), .Y(
        n3462) );
  A2O1A1Ixp33_ASAP7_75t_SL U21045 ( .A1(n30243), .A2(n19002), .B(n22390), .C(
        n19002), .Y(n20446) );
  A2O1A1Ixp33_ASAP7_75t_SL U21046 ( .A1(n30242), .A2(n19002), .B(n22414), .C(
        n19002), .Y(n20447) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21047 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__26_), 
        .A2(n31403), .B(n20446), .C(n19002), .D(n20447), .Y(n3138) );
  A2O1A1Ixp33_ASAP7_75t_SL U21048 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_dci[4]), .C(n20305), .Y(n3127) );
  A2O1A1Ixp33_ASAP7_75t_SL U21049 ( .A1(n22396), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[5]), .C(n20445), .Y(n3075) );
  A2O1A1Ixp33_ASAP7_75t_SL U21050 ( .A1(n32446), .A2(n19002), .B(n31568), .C(
        n24684), .Y(n20439) );
  A2O1A1Ixp33_ASAP7_75t_SL U21051 ( .A1(n24684), .A2(n31617), .B(n20440), .C(
        n19002), .Y(n20441) );
  A2O1A1Ixp33_ASAP7_75t_SL U21052 ( .A1(n31298), .A2(n19002), .B(n20440), .C(
        n19002), .Y(n20442) );
  A2O1A1Ixp33_ASAP7_75t_SL U21053 ( .A1(n3068), .A2(n19002), .B(n20441), .C(
        n20443), .Y(n18047) );
  A2O1A1Ixp33_ASAP7_75t_SL U21054 ( .A1(n19002), .A2(n24646), .B(rf_di_w[29]), 
        .C(n20304), .Y(n3002) );
  A2O1A1Ixp33_ASAP7_75t_SL U21055 ( .A1(n19002), .A2(n24633), .B(
        uart1_r_BREAKIRQEN_), .C(n20296), .Y(n2870) );
  A2O1A1Ixp33_ASAP7_75t_SL U21056 ( .A1(n19002), .A2(n31662), .B(
        u0_0_leon3x0_p0_div0_r_NEG_), .C(n19504), .Y(n2815) );
  A2O1A1Ixp33_ASAP7_75t_SL U21057 ( .A1(n22422), .A2(n19002), .B(n28312), .C(
        n19002), .Y(n20435) );
  A2O1A1Ixp33_ASAP7_75t_SL U21058 ( .A1(n28309), .A2(n19002), .B(n29925), .C(
        n19002), .Y(n20436) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21059 ( .A1(n31662), .A2(n22436), .B(n20435), 
        .C(n19002), .D(n20436), .Y(n2561) );
  A2O1A1Ixp33_ASAP7_75t_SL U21060 ( .A1(n19002), .A2(n24646), .B(rf_di_w[22]), 
        .C(n20290), .Y(n2494) );
  A2O1A1Ixp33_ASAP7_75t_SL U21061 ( .A1(n29956), .A2(n19002), .B(n31114), .C(
        n19002), .Y(n20433) );
  A2O1A1Ixp33_ASAP7_75t_SL U21062 ( .A1(n31115), .A2(n19002), .B(n26069), .C(
        n19002), .Y(n20434) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21063 ( .A1(n31117), .A2(uart1_r_RHOLD__15__0_), 
        .B(n20433), .C(n19002), .D(n20434), .Y(n2452) );
  A2O1A1Ixp33_ASAP7_75t_SL U21064 ( .A1(n32463), .A2(n19002), .B(n32513), .C(
        n19002), .Y(n20431) );
  A2O1A1Ixp33_ASAP7_75t_SL U21065 ( .A1(n32465), .A2(n19002), .B(n32512), .C(
        n19002), .Y(n20432) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21066 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__0_), .A2(n32517), .B(n20431), 
        .C(n19002), .D(n20432), .Y(n2287) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21067 ( .A1(n27305), .A2(n27320), .B(n19002), 
        .C(n24695), .Y(n20053) );
  A2O1A1Ixp33_ASAP7_75t_SL U21068 ( .A1(n19002), .A2(n22433), .B(n32954), .C(
        n20281), .Y(n1714) );
  A2O1A1Ixp33_ASAP7_75t_SL U21069 ( .A1(n19002), .A2(n22433), .B(n32955), .C(
        n20278), .Y(n1705) );
  A2O1A1Ixp33_ASAP7_75t_SL U21070 ( .A1(n32632), .A2(n19002), .B(n32543), .C(
        n20427), .Y(it_data[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21071 ( .A1(n32401), .A2(n19002), .B(n32431), .C(
        n19002), .Y(n20419) );
  A2O1A1Ixp33_ASAP7_75t_SL U21072 ( .A1(n32399), .A2(n19002), .B(n24543), .C(
        n19002), .Y(n20420) );
  A2O1A1Ixp33_ASAP7_75t_SL U21073 ( .A1(n32398), .A2(n19002), .B(n32409), .C(
        n19002), .Y(n20421) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21074 ( .A1(dc_q[26]), .A2(n33069), .B(n20420), 
        .C(n19002), .D(n20421), .Y(n20422) );
  A2O1A1Ixp33_ASAP7_75t_SL U21075 ( .A1(n32650), .A2(n19002), .B(n32429), .C(
        n20422), .Y(n20423) );
  A2O1A1Ixp33_ASAP7_75t_SL U21076 ( .A1(n20419), .A2(n19002), .B(n20423), .C(
        n19002), .Y(n20424) );
  A2O1A1Ixp33_ASAP7_75t_SL U21077 ( .A1(n32634), .A2(n19002), .B(n32217), .C(
        n19663), .Y(dt_data[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21078 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__15_), 
        .A2(n30725), .B(n20257), .C(n19002), .Y(n20258) );
  A2O1A1Ixp33_ASAP7_75t_SL U21079 ( .A1(n22376), .A2(n19002), .B(n30351), .C(
        n20414), .Y(n28586) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21080 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__25_), 
        .A2(n22375), .B(n28406), .C(n19002), .D(n20413), .Y(n32395) );
  A2O1A1Ixp33_ASAP7_75t_SL U21081 ( .A1(DP_OP_1196_128_7433_n8), .A2(n20200), 
        .B(DP_OP_1196_128_7433_n7), .C(n19002), .Y(n20201) );
  A2O1A1Ixp33_ASAP7_75t_SL U21082 ( .A1(n22374), .A2(n19002), .B(n28303), .C(
        n19002), .Y(n20408) );
  A2O1A1Ixp33_ASAP7_75t_SL U21083 ( .A1(n18806), .A2(n19002), .B(n32654), .C(
        n19002), .Y(n20409) );
  A2O1A1Ixp33_ASAP7_75t_SL U21084 ( .A1(n22373), .A2(n19002), .B(n28277), .C(
        n19002), .Y(n20410) );
  O2A1O1Ixp5_ASAP7_75t_SL U21085 ( .A1(n20408), .A2(n20409), .B(n19002), .C(
        n20410), .Y(n28273) );
  A2O1A1Ixp33_ASAP7_75t_SL U21086 ( .A1(n31340), .A2(n19002), .B(n28522), .C(
        n19002), .Y(n20402) );
  A2O1A1Ixp33_ASAP7_75t_SL U21087 ( .A1(n20402), .A2(n19002), .B(n20405), .C(
        n19002), .Y(n20406) );
  A2O1A1Ixp33_ASAP7_75t_SL U21088 ( .A1(n22373), .A2(n19002), .B(n25288), .C(
        n20401), .Y(n30383) );
  A2O1A1Ixp33_ASAP7_75t_SL U21089 ( .A1(DP_OP_5187J1_124_3275_n206), .A2(
        n19002), .B(n20391), .C(n19002), .Y(n20392) );
  A2O1A1Ixp33_ASAP7_75t_SL U21090 ( .A1(n23887), .A2(n19002), .B(n20393), .C(
        n19002), .Y(n20394) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21091 ( .A1(n20392), .A2(
        DP_OP_5187J1_124_3275_n232), .B(n20394), .C(n19002), .D(n20397), .Y(
        n20398) );
  A2O1A1Ixp33_ASAP7_75t_SL U21092 ( .A1(n22373), .A2(n19002), .B(n25311), .C(
        n20390), .Y(n30264) );
  A2O1A1Ixp33_ASAP7_75t_SL U21093 ( .A1(n22376), .A2(n19002), .B(n30407), .C(
        n20389), .Y(n28805) );
  A2O1A1Ixp33_ASAP7_75t_SL U21094 ( .A1(n22374), .A2(n19002), .B(n28329), .C(
        n19002), .Y(n20381) );
  A2O1A1Ixp33_ASAP7_75t_SL U21095 ( .A1(n18806), .A2(n19002), .B(n32630), .C(
        n19002), .Y(n20382) );
  A2O1A1Ixp33_ASAP7_75t_SL U21096 ( .A1(n22373), .A2(n19002), .B(n27224), .C(
        n19002), .Y(n20383) );
  O2A1O1Ixp5_ASAP7_75t_SL U21097 ( .A1(n20381), .A2(n20382), .B(n19002), .C(
        n20383), .Y(n28556) );
  A2O1A1Ixp33_ASAP7_75t_SL U21098 ( .A1(n22373), .A2(n19002), .B(n25292), .C(
        n19002), .Y(n20380) );
  A2O1A1Ixp33_ASAP7_75t_SL U21099 ( .A1(u0_0_leon3x0_p0_divi[44]), .A2(n22373), 
        .B(n20380), .C(n19002), .Y(n30366) );
  A2O1A1Ixp33_ASAP7_75t_SL U21100 ( .A1(n22374), .A2(n19002), .B(n28794), .C(
        n19002), .Y(n20377) );
  A2O1A1Ixp33_ASAP7_75t_SL U21101 ( .A1(n18806), .A2(n19002), .B(n32612), .C(
        n19002), .Y(n20378) );
  A2O1A1Ixp33_ASAP7_75t_SL U21102 ( .A1(n22373), .A2(n19002), .B(n29101), .C(
        n19002), .Y(n20379) );
  O2A1O1Ixp5_ASAP7_75t_SL U21103 ( .A1(n20377), .A2(n20378), .B(n19002), .C(
        n20379), .Y(n29907) );
  A2O1A1Ixp33_ASAP7_75t_SL U21104 ( .A1(n22376), .A2(n19002), .B(n30370), .C(
        n19002), .Y(n20374) );
  A2O1A1Ixp33_ASAP7_75t_SL U21105 ( .A1(n28623), .A2(n19002), .B(n24425), .C(
        n19002), .Y(n20375) );
  A2O1A1Ixp33_ASAP7_75t_SL U21106 ( .A1(n20374), .A2(n19002), .B(n20375), .C(
        n19002), .Y(n29831) );
  A2O1A1Ixp33_ASAP7_75t_SL U21107 ( .A1(n30526), .A2(n19002), .B(n18876), .C(
        n20183), .Y(u0_0_leon3x0_p0_iu_fe_pc_13_) );
  A2O1A1Ixp33_ASAP7_75t_SL U21108 ( .A1(uart1_r_RWADDR__1_), .A2(n19002), .B(
        n20371), .C(n19002), .Y(n26049) );
  A2O1A1Ixp33_ASAP7_75t_SL U21109 ( .A1(n19002), .A2(n28321), .B(n31660), .C(
        n19620), .Y(n19621) );
  A2O1A1Ixp33_ASAP7_75t_SL U21110 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[19]), 
        .B(n19621), .C(n19002), .Y(n19622) );
  A2O1A1Ixp33_ASAP7_75t_SL U21111 ( .A1(n24043), .A2(n19002), .B(n20365), .C(
        n19002), .Y(mult_x_1196_n855) );
  A2O1A1Ixp33_ASAP7_75t_SL U21112 ( .A1(n24043), .A2(n19002), .B(n20364), .C(
        n19002), .Y(mult_x_1196_n2157) );
  A2O1A1Ixp33_ASAP7_75t_SL U21113 ( .A1(n24043), .A2(n19002), .B(n20363), .C(
        n19002), .Y(mult_x_1196_n2152) );
  A2O1A1Ixp33_ASAP7_75t_SL U21114 ( .A1(n29510), .A2(n19002), .B(n30030), .C(
        n19002), .Y(n20358) );
  A2O1A1Ixp33_ASAP7_75t_SL U21115 ( .A1(n22408), .A2(n19002), .B(apbi[35]), 
        .C(n20353), .Y(n4560) );
  A2O1A1Ixp33_ASAP7_75t_SL U21116 ( .A1(n26126), .A2(n19002), .B(n29955), .C(
        n19002), .Y(n20352) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21117 ( .A1(n29959), .A2(uart1_r_RSHIFT__2_), 
        .B(n20352), .C(n19002), .D(n29958), .Y(n4538) );
  A2O1A1Ixp33_ASAP7_75t_SL U21118 ( .A1(n25237), .A2(n19002), .B(n30575), .C(
        n19002), .Y(n20351) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21119 ( .A1(n28411), .A2(n31035), .B(n20351), 
        .C(n19002), .D(n30578), .Y(n4475) );
  A2O1A1Ixp33_ASAP7_75t_SL U21120 ( .A1(n28699), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n20342) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21121 ( .A1(n30644), .A2(n29837), .B(n20342), 
        .C(n19002), .D(n20345), .Y(n20346) );
  A2O1A1Ixp33_ASAP7_75t_SL U21122 ( .A1(n30645), .A2(n19002), .B(n30381), .C(
        n20346), .Y(n20347) );
  A2O1A1Ixp33_ASAP7_75t_SL U21123 ( .A1(n22432), .A2(n30972), .B(n20347), .C(
        n19002), .Y(n20348) );
  A2O1A1Ixp33_ASAP7_75t_SL U21124 ( .A1(n30595), .A2(n19002), .B(n20348), .C(
        n19002), .Y(n20349) );
  A2O1A1Ixp33_ASAP7_75t_SL U21125 ( .A1(n20348), .A2(n30593), .B(n20349), .C(
        n19002), .Y(n20350) );
  A2O1A1Ixp33_ASAP7_75t_SL U21126 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP2__11_), 
        .A2(n20341), .B(n20350), .C(n19002), .Y(n4449) );
  A2O1A1Ixp33_ASAP7_75t_SL U21127 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__23_), .B(n24680), .C(n19002), .Y(n19158) );
  A2O1A1Ixp33_ASAP7_75t_SL U21128 ( .A1(n31842), .A2(n19002), .B(n22397), .C(
        n19002), .Y(n20340) );
  A2O1A1Ixp33_ASAP7_75t_SL U21129 ( .A1(n22420), .A2(n19002), .B(n28306), .C(
        n31422), .Y(n20336) );
  A2O1A1Ixp33_ASAP7_75t_SL U21130 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[21]), 
        .B(n20336), .C(n19002), .Y(n20337) );
  A2O1A1Ixp33_ASAP7_75t_SL U21131 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_21_), .B(n20339), .C(n19002), .Y(n4343) );
  A2O1A1Ixp33_ASAP7_75t_SL U21132 ( .A1(n19002), .A2(n24646), .B(n27032), .C(
        n20097), .Y(n4133) );
  A2O1A1Ixp33_ASAP7_75t_SL U21133 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_), .B(n24654), .C(n19532), .Y(
        n4065) );
  A2O1A1Ixp33_ASAP7_75t_SL U21134 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__RD__6_), .B(n24658), .C(n19137), .Y(
        n4008) );
  A2O1A1Ixp33_ASAP7_75t_SL U21135 ( .A1(n32039), .A2(n19002), .B(n32040), .C(
        n20331), .Y(ahb0_v_CFGSEL_) );
  A2O1A1Ixp33_ASAP7_75t_SL U21136 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__30_), .B(n24655), .C(n19879), .Y(
        n3885) );
  A2O1A1Ixp33_ASAP7_75t_SL U21137 ( .A1(n19002), .A2(n31809), .B(n19317), .C(
        n31815), .Y(n19318) );
  A2O1A1Ixp33_ASAP7_75t_SL U21138 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_r_A__CTRL__ANNUL_), .B(n31810), .C(n19318), .Y(
        n19319) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21139 ( .A1(n31814), .A2(n31813), .B(n19002), 
        .C(n19323), .Y(n19324) );
  A2O1A1Ixp33_ASAP7_75t_SL U21140 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_D__INULL_), .C(n19326), .Y(n3881) );
  A2O1A1Ixp33_ASAP7_75t_SL U21141 ( .A1(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__26_), .A2(n19002), .B(n24656), .C(
        n20329), .Y(n3760) );
  A2O1A1Ixp33_ASAP7_75t_SL U21142 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__11_), .C(n20325), .Y(n3645) );
  A2O1A1Ixp33_ASAP7_75t_SL U21143 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_A__IMM__30_), .C(n19002), .Y(n20321) );
  A2O1A1Ixp33_ASAP7_75t_SL U21144 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), .A2(n19002), .B(n24495), .C(
        n19002), .Y(n20322) );
  A2O1A1Ixp33_ASAP7_75t_SL U21145 ( .A1(n20321), .A2(n19002), .B(n20322), .C(
        n19002), .Y(n20323) );
  A2O1A1Ixp33_ASAP7_75t_SL U21146 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__14_), .A2(n19002), .B(n24650), .C(
        n20320), .Y(n3614) );
  A2O1A1Ixp33_ASAP7_75t_SL U21147 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__5_), 
        .A2(n19002), .B(n24652), .C(n20319), .Y(n3452) );
  A2O1A1Ixp33_ASAP7_75t_SL U21148 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__1_), 
        .A2(n19002), .B(n24651), .C(n20317), .Y(n3356) );
  A2O1A1Ixp33_ASAP7_75t_SL U21149 ( .A1(n22427), .A2(n19002), .B(n30796), .C(
        n20315), .Y(n3330) );
  A2O1A1Ixp33_ASAP7_75t_SL U21150 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__2_), .B(n24653), .C(n20072), .Y(
        n3196) );
  A2O1A1Ixp33_ASAP7_75t_SL U21151 ( .A1(n31257), .A2(n19002), .B(n20306), .C(
        n19002), .Y(n20307) );
  A2O1A1Ixp33_ASAP7_75t_SL U21152 ( .A1(n19002), .A2(n20069), .B(n22405), .C(
        n32675), .Y(n20070) );
  A2O1A1Ixp33_ASAP7_75t_SL U21153 ( .A1(n27493), .A2(n19002), .B(n29376), .C(
        n19002), .Y(n20291) );
  A2O1A1Ixp33_ASAP7_75t_SL U21154 ( .A1(irqctrl0_r_IPEND__1_), .A2(n19002), 
        .B(n29745), .C(n19002), .Y(n20292) );
  A2O1A1Ixp33_ASAP7_75t_SL U21155 ( .A1(irqctrl0_r_IFORCE__0__1_), .A2(n19002), 
        .B(n27297), .C(n24694), .Y(n20293) );
  A2O1A1Ixp33_ASAP7_75t_SL U21156 ( .A1(n20292), .A2(n19002), .B(n20293), .C(
        n19002), .Y(n20294) );
  A2O1A1Ixp33_ASAP7_75t_SL U21157 ( .A1(n29982), .A2(n19002), .B(n29983), .C(
        n20288), .Y(n20289) );
  A2O1A1Ixp33_ASAP7_75t_SL U21158 ( .A1(dataout[4]), .A2(n19002), .B(n20279), 
        .C(n19002), .Y(n20280) );
  A2O1A1Ixp33_ASAP7_75t_SL U21159 ( .A1(dataout[13]), .A2(n19002), .B(n20276), 
        .C(n19002), .Y(n20277) );
  A2O1A1Ixp33_ASAP7_75t_SL U21160 ( .A1(n32592), .A2(n19002), .B(n32593), .C(
        n19002), .Y(n20272) );
  A2O1A1Ixp33_ASAP7_75t_SL U21161 ( .A1(n32590), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__11_), .B(n20272), .C(n19002), 
        .Y(n20273) );
  A2O1A1Ixp33_ASAP7_75t_SL U21162 ( .A1(u0_0_leon3x0_p0_ici[69]), .A2(n32594), 
        .B(n20274), .C(n19002), .Y(n20275) );
  A2O1A1Ixp33_ASAP7_75t_SL U21163 ( .A1(n32596), .A2(n19002), .B(n32595), .C(
        n20275), .Y(ic_address[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21164 ( .A1(n32444), .A2(u0_0_leon3x0_p0_dci[15]), 
        .B(n19675), .C(n19002), .Y(n19676) );
  A2O1A1Ixp33_ASAP7_75t_SL U21165 ( .A1(n19002), .A2(n33067), .B(n19676), .C(
        n19677), .Y(dc_address[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21166 ( .A1(n32383), .A2(n19002), .B(n32431), .C(
        n19002), .Y(n20264) );
  A2O1A1Ixp33_ASAP7_75t_SL U21167 ( .A1(n32642), .A2(n19002), .B(n32429), .C(
        n19002), .Y(n20265) );
  A2O1A1Ixp33_ASAP7_75t_SL U21168 ( .A1(n32382), .A2(n19002), .B(n24543), .C(
        n19002), .Y(n20266) );
  A2O1A1Ixp33_ASAP7_75t_SL U21169 ( .A1(n20265), .A2(n19002), .B(n20266), .C(
        n19002), .Y(n20267) );
  A2O1A1Ixp33_ASAP7_75t_SL U21170 ( .A1(n20264), .A2(n19002), .B(n20269), .C(
        n19002), .Y(n20270) );
  A2O1A1Ixp33_ASAP7_75t_SL U21171 ( .A1(n28000), .A2(uart1_r_THOLD__9__7_), 
        .B(n20210), .C(n19002), .Y(n20211) );
  A2O1A1Ixp33_ASAP7_75t_SL U21172 ( .A1(n28002), .A2(uart1_r_THOLD__5__7_), 
        .B(n20215), .C(n19002), .Y(n20216) );
  A2O1A1Ixp33_ASAP7_75t_SL U21173 ( .A1(n28010), .A2(uart1_r_THOLD__16__7_), 
        .B(uart1_r_TRADDR__1_), .C(n19002), .Y(n20218) );
  A2O1A1Ixp33_ASAP7_75t_SL U21174 ( .A1(n28017), .A2(uart1_r_THOLD__24__7_), 
        .B(n20222), .C(n19002), .Y(n20223) );
  A2O1A1Ixp33_ASAP7_75t_SL U21175 ( .A1(n28018), .A2(uart1_r_THOLD__28__7_), 
        .B(n20227), .C(n19002), .Y(n20228) );
  A2O1A1Ixp33_ASAP7_75t_SL U21176 ( .A1(n27998), .A2(uart1_r_THOLD__27__7_), 
        .B(n20233), .C(n19002), .Y(n20234) );
  A2O1A1Ixp33_ASAP7_75t_SL U21177 ( .A1(n28002), .A2(uart1_r_THOLD__7__7_), 
        .B(n20238), .C(n19002), .Y(n20239) );
  A2O1A1Ixp33_ASAP7_75t_SL U21178 ( .A1(n28018), .A2(uart1_r_THOLD__30__7_), 
        .B(n28016), .C(n19002), .Y(n20241) );
  A2O1A1Ixp33_ASAP7_75t_SL U21179 ( .A1(n28017), .A2(uart1_r_THOLD__26__7_), 
        .B(n20244), .C(n19002), .Y(n20245) );
  A2O1A1Ixp33_ASAP7_75t_SL U21180 ( .A1(uart1_r_TRADDR__0_), .A2(n20240), .B(
        n20248), .C(n19002), .Y(n20249) );
  A2O1A1Ixp33_ASAP7_75t_SL U21181 ( .A1(n31340), .A2(n19002), .B(n28556), .C(
        n19002), .Y(n20203) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21182 ( .A1(n31342), .A2(n31875), .B(n20203), 
        .C(n19002), .D(n20206), .Y(n27240) );
  A2O1A1Ixp33_ASAP7_75t_SL U21183 ( .A1(DP_OP_5187J1_124_3275_n249), .A2(
        n20197), .B(n18833), .C(n19002), .Y(n20198) );
  A2O1A1Ixp33_ASAP7_75t_SL U21184 ( .A1(n30619), .A2(n29563), .B(n20196), .C(
        n19002), .Y(n32300) );
  O2A1O1Ixp33_ASAP7_75t_SL U21185 ( .A1(n18610), .A2(add_x_735_A_19_), .B(
        n19002), .C(n20194), .Y(n31665) );
  A2O1A1Ixp33_ASAP7_75t_SL U21186 ( .A1(n22373), .A2(n19002), .B(n26350), .C(
        n20191), .Y(n30613) );
  A2O1A1Ixp33_ASAP7_75t_SL U21187 ( .A1(n22373), .A2(n19002), .B(n30607), .C(
        n20186), .Y(n30609) );
  A2O1A1Ixp33_ASAP7_75t_SL U21188 ( .A1(n30205), .A2(n19002), .B(n20185), .C(
        n19002), .Y(n31549) );
  A2O1A1Ixp33_ASAP7_75t_SL U21189 ( .A1(n31945), .A2(n19002), .B(n20184), .C(
        n19002), .Y(n30488) );
  A2O1A1Ixp33_ASAP7_75t_SL U21190 ( .A1(n22376), .A2(n19002), .B(n30361), .C(
        n20179), .Y(n28602) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21191 ( .A1(n32786), .A2(n32802), .B(n19002), 
        .C(n32801), .Y(n20178) );
  A2O1A1Ixp33_ASAP7_75t_SL U21192 ( .A1(n19002), .A2(n28334), .B(n31660), .C(
        n19794), .Y(n19795) );
  A2O1A1Ixp33_ASAP7_75t_SL U21193 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[13]), 
        .B(n19795), .C(n19002), .Y(n19796) );
  A2O1A1Ixp33_ASAP7_75t_SL U21194 ( .A1(n32353), .A2(n19002), .B(n32626), .C(
        n19002), .Y(n20177) );
  A2O1A1Ixp33_ASAP7_75t_SL U21195 ( .A1(n32353), .A2(n19002), .B(n32622), .C(
        n19002), .Y(n20175) );
  A2O1A1Ixp33_ASAP7_75t_SL U21196 ( .A1(n32353), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[0]), .C(n19002), .Y(n20174) );
  A2O1A1Ixp33_ASAP7_75t_SL U21197 ( .A1(n32293), .A2(n32353), .B(n20174), .C(
        n19002), .Y(n32393) );
  A2O1A1Ixp33_ASAP7_75t_SL U21198 ( .A1(n22376), .A2(n19002), .B(n30429), .C(
        n19002), .Y(n20172) );
  A2O1A1Ixp33_ASAP7_75t_SL U21199 ( .A1(n31475), .A2(n19002), .B(n24425), .C(
        n19002), .Y(n20173) );
  A2O1A1Ixp33_ASAP7_75t_SL U21200 ( .A1(n20172), .A2(n19002), .B(n20173), .C(
        n19002), .Y(n29499) );
  O2A1O1Ixp33_ASAP7_75t_SL U21201 ( .A1(n26009), .A2(uart1_r_RWADDR__0_), .B(
        n19002), .C(uart1_r_RWADDR__2_), .Y(n26055) );
  A2O1A1Ixp33_ASAP7_75t_SL U21202 ( .A1(n28305), .A2(n19002), .B(n31660), .C(
        n20167), .Y(n20168) );
  A2O1A1Ixp33_ASAP7_75t_SL U21203 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[25]), 
        .B(n20168), .C(n19002), .Y(n20169) );
  A2O1A1Ixp33_ASAP7_75t_SL U21204 ( .A1(n28302), .A2(n19002), .B(n31660), .C(
        n20162), .Y(n20163) );
  A2O1A1Ixp33_ASAP7_75t_SL U21205 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[28]), 
        .B(n20163), .C(n19002), .Y(n20164) );
  A2O1A1Ixp33_ASAP7_75t_SL U21206 ( .A1(n24046), .A2(n19002), .B(n22642), .C(
        n19002), .Y(n20153) );
  A2O1A1Ixp33_ASAP7_75t_SL U21207 ( .A1(n24043), .A2(n19002), .B(n20153), .C(
        n19002), .Y(n20154) );
  A2O1A1Ixp33_ASAP7_75t_SL U21208 ( .A1(n24043), .A2(n19002), .B(n20152), .C(
        n19002), .Y(mult_x_1196_n2149) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21209 ( .A1(n4701), .A2(n29945), .B(n19002), .C(
        n4519), .Y(n20136) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21210 ( .A1(n4701), .A2(n29947), .B(n29953), .C(
        n19002), .D(n29946), .Y(n20137) );
  A2O1A1Ixp33_ASAP7_75t_SL U21211 ( .A1(n29950), .A2(n19002), .B(n29949), .C(
        n19002), .Y(n20139) );
  A2O1A1Ixp33_ASAP7_75t_SL U21212 ( .A1(n31973), .A2(n19002), .B(n20131), .C(
        n19002), .Y(n20132) );
  A2O1A1Ixp33_ASAP7_75t_SL U21213 ( .A1(n32004), .A2(n19002), .B(n29988), .C(
        n19002), .Y(n20133) );
  A2O1A1Ixp33_ASAP7_75t_SL U21214 ( .A1(n4669), .A2(n19002), .B(n20134), .C(
        n19002), .Y(n20135) );
  A2O1A1Ixp33_ASAP7_75t_SL U21215 ( .A1(apbi[29]), .A2(n19002), .B(n29650), 
        .C(n29649), .Y(n20128) );
  A2O1A1Ixp33_ASAP7_75t_SL U21216 ( .A1(n32280), .A2(n33067), .B(n31456), .C(
        n19002), .Y(n20119) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21217 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_MEXC_), .A2(n30207), .B(n30208), .C(
        n19002), .D(n32199), .Y(n20121) );
  A2O1A1Ixp33_ASAP7_75t_SL U21218 ( .A1(n29071), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n20110) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21219 ( .A1(n29067), .A2(n30644), .B(n20110), 
        .C(n19002), .D(n20113), .Y(n20114) );
  A2O1A1Ixp33_ASAP7_75t_SL U21220 ( .A1(n30645), .A2(n19002), .B(n29808), .C(
        n20114), .Y(n20115) );
  A2O1A1Ixp33_ASAP7_75t_SL U21221 ( .A1(n29807), .A2(n22432), .B(n20115), .C(
        n19002), .Y(n20116) );
  A2O1A1Ixp33_ASAP7_75t_SL U21222 ( .A1(n28472), .A2(n19002), .B(n22379), .C(
        n19002), .Y(n20118) );
  A2O1A1Ixp33_ASAP7_75t_SL U21223 ( .A1(n24638), .A2(n19002), .B(n20103), .C(
        n19002), .Y(n20104) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21224 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__27_), .B(n24680), .C(n19002), .D(n20104), 
        .Y(n20105) );
  A2O1A1Ixp33_ASAP7_75t_SL U21225 ( .A1(n30453), .A2(n30240), .B(n20107), .C(
        n19002), .Y(n20108) );
  A2O1A1Ixp33_ASAP7_75t_SL U21226 ( .A1(n30426), .A2(n19002), .B(n30241), .C(
        n20108), .Y(n20109) );
  A2O1A1Ixp33_ASAP7_75t_SL U21227 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_divi[58]), .C(n20109), .Y(n4400) );
  A2O1A1Ixp33_ASAP7_75t_SL U21228 ( .A1(n22420), .A2(n19002), .B(n28298), .C(
        n31422), .Y(n20098) );
  A2O1A1Ixp33_ASAP7_75t_SL U21229 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[30]), 
        .B(n20098), .C(n19002), .Y(n20099) );
  A2O1A1Ixp33_ASAP7_75t_SL U21230 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_30_), .B(n20101), .C(n19002), .Y(n4324) );
  A2O1A1Ixp33_ASAP7_75t_SL U21231 ( .A1(n24646), .A2(n19002), .B(n19742), .C(
        n19743), .Y(n4297) );
  A2O1A1Ixp33_ASAP7_75t_SL U21232 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__1_), .B(n24650), .C(n19890), .Y(
        n4109) );
  A2O1A1Ixp33_ASAP7_75t_SL U21233 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PV_), .B(n24649), .C(n19531), .Y(n4022)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21234 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__6_), 
        .A2(n19002), .B(n24658), .C(n20094), .Y(n4010) );
  A2O1A1Ixp33_ASAP7_75t_SL U21235 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__26_), .B(n24656), .C(n19723), .Y(
        n3762) );
  A2O1A1Ixp33_ASAP7_75t_SL U21236 ( .A1(n33055), .A2(n19002), .B(n23229), .C(
        n19002), .Y(n20089) );
  A2O1A1Ixp33_ASAP7_75t_SL U21237 ( .A1(u0_0_leon3x0_p0_iu_v_X__DCI__SIGNED_), 
        .A2(n19002), .B(n24657), .C(n20079), .Y(n3578) );
  A2O1A1Ixp33_ASAP7_75t_SL U21238 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__5_), 
        .A2(n19002), .B(n22428), .C(n20077), .Y(n3450) );
  A2O1A1Ixp33_ASAP7_75t_SL U21239 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_W__S__WIM__1_), .C(n20075), .Y(n3338) );
  A2O1A1Ixp33_ASAP7_75t_SL U21240 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[4]), .C(n19702), .Y(n3085) );
  A2O1A1Ixp33_ASAP7_75t_SL U21241 ( .A1(n31318), .A2(n19002), .B(n20065), .C(
        n19002), .Y(n20066) );
  A2O1A1Ixp33_ASAP7_75t_SL U21242 ( .A1(n32467), .A2(n31892), .B(
        u0_0_leon3x0_p0_c0mmu_mcii[1]), .C(n19002), .Y(n20067) );
  A2O1A1Ixp33_ASAP7_75t_SL U21243 ( .A1(n20066), .A2(n19002), .B(n20067), .C(
        n19002), .Y(n20068) );
  A2O1A1Ixp33_ASAP7_75t_SL U21244 ( .A1(n28167), .A2(uart1_uarto_SCALER__5_), 
        .B(n22419), .C(n19002), .Y(n19867) );
  A2O1A1Ixp33_ASAP7_75t_SL U21245 ( .A1(uart1_r_RXSTATE__0_), .A2(n19002), .B(
        n29972), .C(n20062), .Y(n20063) );
  A2O1A1Ixp33_ASAP7_75t_SL U21246 ( .A1(n29974), .A2(n19002), .B(n20063), .C(
        n29973), .Y(n17450) );
  A2O1A1Ixp33_ASAP7_75t_SL U21247 ( .A1(u0_0_leon3x0_p0_divo[0]), .A2(n31421), 
        .B(n20057), .C(n19002), .Y(n20058) );
  A2O1A1Ixp33_ASAP7_75t_SL U21248 ( .A1(n19002), .A2(n22433), .B(n32962), .C(
        n19684), .Y(n1713) );
  A2O1A1Ixp33_ASAP7_75t_SL U21249 ( .A1(n19002), .A2(n22433), .B(n32963), .C(
        n19845), .Y(n1704) );
  A2O1A1Ixp33_ASAP7_75t_SL U21250 ( .A1(n32577), .A2(n19002), .B(n32585), .C(
        n19002), .Y(n20047) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21251 ( .A1(n32590), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__8_), .B(n20047), .C(n19002), 
        .D(n20050), .Y(n20051) );
  A2O1A1Ixp33_ASAP7_75t_SL U21252 ( .A1(n19002), .A2(n32660), .B(n32616), .C(
        n19831), .Y(ic_data[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21253 ( .A1(n32646), .A2(n19002), .B(n32429), .C(
        n19002), .Y(n20041) );
  A2O1A1Ixp33_ASAP7_75t_SL U21254 ( .A1(n32391), .A2(n19002), .B(n24543), .C(
        n19002), .Y(n20042) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21255 ( .A1(dc_q[24]), .A2(n33069), .B(n20041), 
        .C(n19002), .D(n20042), .Y(n20043) );
  A2O1A1Ixp33_ASAP7_75t_SL U21256 ( .A1(n32392), .A2(n19002), .B(n32431), .C(
        n20043), .Y(n20044) );
  A2O1A1Ixp33_ASAP7_75t_SL U21257 ( .A1(n32434), .A2(n32393), .B(n20044), .C(
        n19002), .Y(n20045) );
  A2O1A1Ixp33_ASAP7_75t_SL U21258 ( .A1(n32425), .A2(n19002), .B(n32394), .C(
        n20045), .Y(dc_data[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21259 ( .A1(n32405), .A2(n19002), .B(n32232), .C(
        n19002), .Y(n20038) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21260 ( .A1(n32239), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__28_), .B(n33067), .C(n19002), .D(
        n20038), .Y(n20039) );
  A2O1A1Ixp33_ASAP7_75t_SL U21261 ( .A1(n30725), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__PC__22_), .B(n20034), .C(n19002), .Y(
        n20035) );
  A2O1A1Ixp33_ASAP7_75t_SL U21262 ( .A1(n22375), .A2(n30598), .B(n19063), .C(
        n19002), .Y(n19064) );
  O2A1O1Ixp5_ASAP7_75t_SL U21263 ( .A1(n19061), .A2(n19062), .B(n19002), .C(
        n19064), .Y(n32418) );
  A2O1A1Ixp33_ASAP7_75t_SL U21264 ( .A1(n31340), .A2(n19002), .B(n28576), .C(
        n19002), .Y(n20027) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21265 ( .A1(n31342), .A2(n28578), .B(n20027), 
        .C(n19002), .D(n20030), .Y(n30492) );
  A2O1A1Ixp33_ASAP7_75t_SL U21266 ( .A1(n22376), .A2(n19002), .B(n30248), .C(
        n20026), .Y(n29783) );
  A2O1A1Ixp33_ASAP7_75t_SL U21267 ( .A1(n23887), .A2(n19002), .B(n20019), .C(
        n19002), .Y(n20020) );
  A2O1A1Ixp33_ASAP7_75t_SL U21268 ( .A1(n20020), .A2(n19002), .B(n20022), .C(
        n19002), .Y(n20023) );
  A2O1A1Ixp33_ASAP7_75t_SL U21269 ( .A1(n22376), .A2(n19002), .B(n30696), .C(
        n20018), .Y(n29837) );
  A2O1A1Ixp33_ASAP7_75t_SL U21270 ( .A1(n23941), .A2(n19002), .B(n20014), .C(
        n19002), .Y(n20015) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21271 ( .A1(DP_OP_1196_128_7433_n84), .A2(
        DP_OP_1196_128_7433_n7), .B(n20015), .C(n19002), .D(
        DP_OP_1196_128_7433_n85), .Y(n20016) );
  A2O1A1Ixp33_ASAP7_75t_SL U21272 ( .A1(n22374), .A2(n19002), .B(n28319), .C(
        n19002), .Y(n20010) );
  A2O1A1Ixp33_ASAP7_75t_SL U21273 ( .A1(n18805), .A2(n19002), .B(n32640), .C(
        n19002), .Y(n20011) );
  A2O1A1Ixp33_ASAP7_75t_SL U21274 ( .A1(n22373), .A2(n19002), .B(n27037), .C(
        n19002), .Y(n20012) );
  O2A1O1Ixp5_ASAP7_75t_SL U21275 ( .A1(n20010), .A2(n20011), .B(n19002), .C(
        n20012), .Y(n28522) );
  A2O1A1Ixp33_ASAP7_75t_SL U21276 ( .A1(n22374), .A2(n19002), .B(n28364), .C(
        n19002), .Y(n20005) );
  A2O1A1Ixp33_ASAP7_75t_SL U21277 ( .A1(n18805), .A2(n19002), .B(n32602), .C(
        n19002), .Y(n20006) );
  A2O1A1Ixp33_ASAP7_75t_SL U21278 ( .A1(n22373), .A2(n19002), .B(n29106), .C(
        n19002), .Y(n20007) );
  O2A1O1Ixp5_ASAP7_75t_SL U21279 ( .A1(n20005), .A2(n20006), .B(n19002), .C(
        n20007), .Y(n30464) );
  A2O1A1Ixp33_ASAP7_75t_SL U21280 ( .A1(n31690), .A2(n19002), .B(n18876), .C(
        n19036), .Y(u0_0_leon3x0_p0_iu_fe_pc_29_) );
  A2O1A1Ixp33_ASAP7_75t_SL U21281 ( .A1(n19002), .A2(n29773), .B(n18876), .C(
        n19441), .Y(u0_0_leon3x0_p0_iu_fe_pc_24_) );
  A2O1A1Ixp33_ASAP7_75t_SL U21282 ( .A1(n27503), .A2(n19002), .B(n20000), .C(
        n19002), .Y(n27501) );
  A2O1A1Ixp33_ASAP7_75t_SL U21283 ( .A1(n22906), .A2(n22416), .B(n18813), .C(
        n19002), .Y(n19993) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21284 ( .A1(n28847), .A2(n26424), .B(n19994), 
        .C(n19002), .D(n19997), .Y(n19998) );
  A2O1A1Ixp33_ASAP7_75t_SL U21285 ( .A1(n22374), .A2(n19002), .B(n31675), .C(
        n19002), .Y(n19991) );
  A2O1A1Ixp33_ASAP7_75t_SL U21286 ( .A1(n29082), .A2(n19002), .B(n22373), .C(
        n19002), .Y(n19992) );
  A2O1A1Ixp33_ASAP7_75t_SL U21287 ( .A1(n19991), .A2(n19002), .B(n19992), .C(
        n19002), .Y(n29810) );
  A2O1A1Ixp33_ASAP7_75t_SL U21288 ( .A1(uart1_r_RWADDR__1_), .A2(n19002), .B(
        n19990), .C(n19002), .Y(n26062) );
  A2O1A1Ixp33_ASAP7_75t_SL U21289 ( .A1(n28329), .A2(n19002), .B(n31660), .C(
        n19980), .Y(n19981) );
  A2O1A1Ixp33_ASAP7_75t_SL U21290 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[15]), 
        .B(n19981), .C(n19002), .Y(n19982) );
  A2O1A1Ixp33_ASAP7_75t_SL U21291 ( .A1(n24047), .A2(n19002), .B(n24043), .C(
        n22642), .Y(n19979) );
  A2O1A1Ixp33_ASAP7_75t_SL U21292 ( .A1(n24043), .A2(n19002), .B(n19977), .C(
        n19002), .Y(mult_x_1196_n2158) );
  A2O1A1Ixp33_ASAP7_75t_SL U21293 ( .A1(n1728), .A2(n19002), .B(n31953), .C(
        n19002), .Y(n19918) );
  A2O1A1Ixp33_ASAP7_75t_SL U21294 ( .A1(n31243), .A2(n19002), .B(n31244), .C(
        n19002), .Y(n19919) );
  A2O1A1Ixp33_ASAP7_75t_SL U21295 ( .A1(n31248), .A2(irqctrl0_r_ILEVEL__6_), 
        .B(apb0_r_CFGSEL_), .C(n19002), .Y(n19920) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21296 ( .A1(uart1_r_FLOW_), .A2(n31950), .B(
        n19923), .C(n19002), .D(n19927), .Y(n19928) );
  O2A1O1Ixp33_ASAP7_75t_SL U21297 ( .A1(n19918), .A2(n19919), .B(n19002), .C(
        n19931), .Y(n19932) );
  A2O1A1Ixp33_ASAP7_75t_SL U21298 ( .A1(n31208), .A2(uart1_r_RHOLD__19__6_), 
        .B(n19938), .C(n19002), .Y(n19939) );
  A2O1A1Ixp33_ASAP7_75t_SL U21299 ( .A1(n31212), .A2(uart1_r_RHOLD__26__6_), 
        .B(n19943), .C(n19002), .Y(n19944) );
  A2O1A1Ixp33_ASAP7_75t_SL U21300 ( .A1(n31204), .A2(uart1_r_RHOLD__9__6_), 
        .B(n19947), .C(n19002), .Y(n19948) );
  A2O1A1Ixp33_ASAP7_75t_SL U21301 ( .A1(n19954), .A2(n19002), .B(n19957), .C(
        n19002), .Y(n19958) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21302 ( .A1(n31205), .A2(uart1_r_RHOLD__16__6_), 
        .B(n19951), .C(n19002), .D(n19961), .Y(n19962) );
  O2A1O1Ixp5_ASAP7_75t_SL U21303 ( .A1(n19933), .A2(n19934), .B(n19002), .C(
        n19963), .Y(n19964) );
  A2O1A1Ixp33_ASAP7_75t_SL U21304 ( .A1(n31237), .A2(timer0_r_RELOAD__6_), .B(
        n19966), .C(n19002), .Y(n19967) );
  A2O1A1Ixp33_ASAP7_75t_SL U21305 ( .A1(n31238), .A2(n19002), .B(n19964), .C(
        n19967), .Y(n19968) );
  A2O1A1Ixp33_ASAP7_75t_SL U21306 ( .A1(n31239), .A2(n31240), .B(n19968), .C(
        n19002), .Y(n19969) );
  A2O1A1Ixp33_ASAP7_75t_SL U21307 ( .A1(n31241), .A2(uart1_r_RHOLD__24__6_), 
        .B(n19971), .C(n19002), .Y(n19972) );
  A2O1A1Ixp33_ASAP7_75t_SL U21308 ( .A1(n31252), .A2(n19002), .B(n19917), .C(
        n19973), .Y(n4714) );
  A2O1A1Ixp33_ASAP7_75t_SL U21309 ( .A1(n29951), .A2(n28031), .B(n24695), .C(
        n19002), .Y(n19915) );
  A2O1A1Ixp33_ASAP7_75t_SL U21310 ( .A1(uart1_r_TSHIFT__0_), .A2(n29954), .B(
        n19916), .C(n19002), .Y(n4699) );
  O2A1O1Ixp33_ASAP7_75t_SL U21311 ( .A1(n29790), .A2(n29791), .B(n19002), .C(
        n31343), .Y(n19550) );
  O2A1O1Ixp33_ASAP7_75t_SL U21312 ( .A1(n19762), .A2(n19765), .B(n19002), .C(
        n19769), .Y(n19770) );
  A2O1A1Ixp33_ASAP7_75t_SL U21313 ( .A1(n32311), .A2(n19002), .B(n31470), .C(
        n19002), .Y(n19901) );
  A2O1A1Ixp33_ASAP7_75t_SL U21314 ( .A1(n30012), .A2(n19002), .B(n31466), .C(
        n31465), .Y(n19902) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21315 ( .A1(n22387), .A2(ic_q[5]), .B(n19901), 
        .C(n19002), .D(n19902), .Y(n19903) );
  A2O1A1Ixp33_ASAP7_75t_SL U21316 ( .A1(n32497), .A2(n19002), .B(n24426), .C(
        n19903), .Y(n19904) );
  A2O1A1Ixp33_ASAP7_75t_SL U21317 ( .A1(dc_q[5]), .A2(n31473), .B(n19904), .C(
        n19002), .Y(n19905) );
  A2O1A1Ixp33_ASAP7_75t_SL U21318 ( .A1(n30026), .A2(n19002), .B(n31483), .C(
        n19002), .Y(n19906) );
  A2O1A1Ixp33_ASAP7_75t_SL U21319 ( .A1(n19906), .A2(n19002), .B(n19909), .C(
        n19002), .Y(n19910) );
  A2O1A1Ixp33_ASAP7_75t_SL U21320 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__5_), .A2(n31486), .B(n19912), .C(n19002), .Y(n19913) );
  A2O1A1Ixp33_ASAP7_75t_SL U21321 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__5_), 
        .A2(n19002), .B(n31491), .C(n19914), .Y(n4382) );
  A2O1A1Ixp33_ASAP7_75t_SL U21322 ( .A1(n29570), .A2(n19002), .B(n22397), .C(
        n19002), .Y(n19900) );
  A2O1A1Ixp33_ASAP7_75t_SL U21323 ( .A1(n28520), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n19891) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21324 ( .A1(n30644), .A2(n28521), .B(n19891), 
        .C(n19002), .D(n19894), .Y(n19895) );
  A2O1A1Ixp33_ASAP7_75t_SL U21325 ( .A1(n30645), .A2(n19002), .B(n28522), .C(
        n19895), .Y(n19896) );
  A2O1A1Ixp33_ASAP7_75t_SL U21326 ( .A1(n31545), .A2(n22432), .B(n19896), .C(
        n19002), .Y(n19897) );
  A2O1A1Ixp33_ASAP7_75t_SL U21327 ( .A1(n28523), .A2(n19002), .B(n22379), .C(
        n19002), .Y(n19899) );
  A2O1A1Ixp33_ASAP7_75t_SL U21328 ( .A1(n19002), .A2(n24646), .B(n29078), .C(
        n19533), .Y(n4129) );
  A2O1A1Ixp33_ASAP7_75t_SL U21329 ( .A1(n22420), .A2(n19002), .B(n28320), .C(
        n31422), .Y(n19885) );
  A2O1A1Ixp33_ASAP7_75t_SL U21330 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[19]), 
        .B(n19885), .C(n19002), .Y(n19886) );
  A2O1A1Ixp33_ASAP7_75t_SL U21331 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_19_), .B(n19888), .C(n19002), .Y(n4044) );
  A2O1A1Ixp33_ASAP7_75t_SL U21332 ( .A1(n26872), .A2(n19002), .B(n23229), .C(
        n19002), .Y(n19881) );
  A2O1A1Ixp33_ASAP7_75t_SL U21333 ( .A1(n30810), .A2(n19882), .B(n30811), .C(
        n19002), .Y(n19883) );
  A2O1A1Ixp33_ASAP7_75t_SL U21334 ( .A1(n19883), .A2(n19002), .B(n30812), .C(
        n19002), .Y(n19884) );
  A2O1A1Ixp33_ASAP7_75t_SL U21335 ( .A1(n19881), .A2(n19002), .B(n19884), .C(
        n19002), .Y(n4004) );
  A2O1A1Ixp33_ASAP7_75t_SL U21336 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__TRAP_), .B(n24656), .C(n19528), .Y(n3735) );
  A2O1A1Ixp33_ASAP7_75t_SL U21337 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__10_), .A2(n19002), .B(n24649), .C(
        n19877), .Y(n3648) );
  A2O1A1Ixp33_ASAP7_75t_SL U21338 ( .A1(n24495), .A2(n19002), .B(
        DP_OP_1196_128_7433_n453), .C(n19874), .Y(n3538) );
  A2O1A1Ixp33_ASAP7_75t_SL U21339 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__23_), 
        .A2(n19002), .B(n24651), .C(n19870), .Y(n3246) );
  A2O1A1Ixp33_ASAP7_75t_SL U21340 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__2_), .B(n24653), .C(n19704), .Y(
        n3194) );
  A2O1A1Ixp33_ASAP7_75t_SL U21341 ( .A1(uart1_uarto_SCALER__3_), .A2(n19002), 
        .B(n19861), .C(n19002), .Y(n19862) );
  A2O1A1Ixp33_ASAP7_75t_SL U21342 ( .A1(n28182), .A2(n28181), .B(n28185), .C(
        n19002), .Y(n19860) );
  A2O1A1Ixp33_ASAP7_75t_SL U21343 ( .A1(n19002), .A2(n29383), .B(apbi[15]), 
        .C(n19693), .Y(n2848) );
  A2O1A1Ixp33_ASAP7_75t_SL U21344 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_W__S__WIM__0_), .C(n19859), .Y(n2767) );
  A2O1A1Ixp33_ASAP7_75t_SL U21345 ( .A1(n27524), .A2(n19002), .B(n27515), .C(
        n19002), .Y(n19853) );
  A2O1A1Ixp33_ASAP7_75t_SL U21346 ( .A1(n19002), .A2(n24633), .B(
        uart1_r_TSEMPTYIRQEN_), .C(n19688), .Y(n2325) );
  A2O1A1Ixp33_ASAP7_75t_SL U21347 ( .A1(n32454), .A2(n3135), .B(n32660), .C(
        n19002), .Y(n19850) );
  A2O1A1Ixp33_ASAP7_75t_SL U21348 ( .A1(n32564), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_icache0_r_HIT_), .C(n19002), .Y(n19851) );
  A2O1A1Ixp33_ASAP7_75t_SL U21349 ( .A1(n19850), .A2(n19002), .B(n19851), .C(
        n19002), .Y(n19852) );
  A2O1A1Ixp33_ASAP7_75t_SL U21350 ( .A1(n19852), .A2(n19002), .B(n32458), .C(
        n19002), .Y(n2289) );
  A2O1A1Ixp33_ASAP7_75t_SL U21351 ( .A1(n22393), .A2(n19002), .B(n33000), .C(
        n19002), .Y(n19847) );
  A2O1A1Ixp33_ASAP7_75t_SL U21352 ( .A1(ahb0_r_HADDR__10_), .A2(n19846), .B(
        n19847), .C(n19002), .Y(n1806) );
  A2O1A1Ixp33_ASAP7_75t_SL U21353 ( .A1(n19002), .A2(n22433), .B(n32970), .C(
        n19488), .Y(n1712) );
  A2O1A1Ixp33_ASAP7_75t_SL U21354 ( .A1(dataout[14]), .A2(n19002), .B(n19843), 
        .C(n19002), .Y(n19844) );
  A2O1A1Ixp33_ASAP7_75t_SL U21355 ( .A1(n22379), .A2(n19002), .B(
        u0_0_leon3x0_p0_dci[2]), .C(n19842), .Y(n3302) );
  A2O1A1Ixp33_ASAP7_75t_SL U21356 ( .A1(n32572), .A2(n19002), .B(n32595), .C(
        n19002), .Y(n19832) );
  A2O1A1Ixp33_ASAP7_75t_SL U21357 ( .A1(n32570), .A2(n19002), .B(n32593), .C(
        n19002), .Y(n19833) );
  A2O1A1Ixp33_ASAP7_75t_SL U21358 ( .A1(n3065), .A2(n19002), .B(n32571), .C(
        n19002), .Y(n19834) );
  A2O1A1Ixp33_ASAP7_75t_SL U21359 ( .A1(n19833), .A2(n19002), .B(n19834), .C(
        n19002), .Y(n19835) );
  A2O1A1Ixp33_ASAP7_75t_SL U21360 ( .A1(n19832), .A2(n19002), .B(n19837), .C(
        n19002), .Y(n19838) );
  A2O1A1Ixp33_ASAP7_75t_SL U21361 ( .A1(n32408), .A2(n19002), .B(n32341), .C(
        n19002), .Y(n19825) );
  A2O1A1Ixp33_ASAP7_75t_SL U21362 ( .A1(n19825), .A2(n19002), .B(n19828), .C(
        n19002), .Y(n19829) );
  A2O1A1Ixp33_ASAP7_75t_SL U21363 ( .A1(n32661), .A2(n19002), .B(n32235), .C(
        n19002), .Y(n19822) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21364 ( .A1(n32239), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__31_), .B(n33067), .C(n19002), .D(
        n19822), .Y(n19823) );
  A2O1A1Ixp33_ASAP7_75t_SL U21365 ( .A1(n29413), .A2(n19002), .B(n19821), .C(
        n19002), .Y(n29663) );
  A2O1A1Ixp33_ASAP7_75t_SL U21366 ( .A1(n22376), .A2(n19002), .B(n30242), .C(
        n19819), .Y(n29796) );
  A2O1A1Ixp33_ASAP7_75t_SL U21367 ( .A1(n22374), .A2(n19002), .B(n28344), .C(
        n19002), .Y(n19816) );
  A2O1A1Ixp33_ASAP7_75t_SL U21368 ( .A1(n18805), .A2(n19002), .B(n32618), .C(
        n19002), .Y(n19817) );
  A2O1A1Ixp33_ASAP7_75t_SL U21369 ( .A1(n22373), .A2(n19002), .B(n27168), .C(
        n19002), .Y(n19818) );
  O2A1O1Ixp5_ASAP7_75t_SL U21370 ( .A1(n19816), .A2(n19817), .B(n19002), .C(
        n19818), .Y(n30385) );
  A2O1A1Ixp33_ASAP7_75t_SL U21371 ( .A1(n22374), .A2(n19002), .B(n28316), .C(
        n19002), .Y(n19813) );
  A2O1A1Ixp33_ASAP7_75t_SL U21372 ( .A1(n18805), .A2(n19002), .B(n32644), .C(
        n19002), .Y(n19814) );
  A2O1A1Ixp33_ASAP7_75t_SL U21373 ( .A1(n22373), .A2(n19002), .B(n29090), .C(
        n19002), .Y(n19815) );
  O2A1O1Ixp5_ASAP7_75t_SL U21374 ( .A1(n19813), .A2(n19814), .B(n19002), .C(
        n19815), .Y(n29808) );
  A2O1A1Ixp33_ASAP7_75t_SL U21375 ( .A1(DP_OP_5187J1_124_3275_n276), .A2(
        DP_OP_5187J1_124_3275_n289), .B(n18835), .C(n19002), .Y(n19651) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21376 ( .A1(DP_OP_1196_128_7433_n57), .A2(
        DP_OP_1196_128_7433_n50), .B(n19002), .C(DP_OP_1196_128_7433_n66), .Y(
        n19242) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21377 ( .A1(DP_OP_1196_128_7433_n57), .A2(
        DP_OP_1196_128_7433_n50), .B(n19002), .C(DP_OP_1196_128_7433_n67), .Y(
        n19245) );
  A2O1A1Ixp33_ASAP7_75t_SL U21378 ( .A1(n19002), .A2(DP_OP_1196_128_7433_n50), 
        .B(DP_OP_1196_128_7433_n60), .C(DP_OP_1196_128_7433_n51), .Y(n19246)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21379 ( .A1(u0_0_leon3x0_p0_ici[59]), .A2(n19252), 
        .B(n19253), .C(n19002), .Y(n19254) );
  A2O1A1Ixp33_ASAP7_75t_SL U21380 ( .A1(n23965), .A2(n19002), .B(n28821), .C(
        n19807), .Y(n19808) );
  A2O1A1Ixp33_ASAP7_75t_SL U21381 ( .A1(n22216), .A2(n19002), .B(n28928), .C(
        n19002), .Y(n19809) );
  A2O1A1Ixp33_ASAP7_75t_SL U21382 ( .A1(n23965), .A2(n19002), .B(n29148), .C(
        n19002), .Y(n19810) );
  A2O1A1Ixp33_ASAP7_75t_SL U21383 ( .A1(n19809), .A2(n19002), .B(n19810), .C(
        n19002), .Y(n19811) );
  O2A1O1Ixp33_ASAP7_75t_SL U21384 ( .A1(u0_0_leon3x0_p0_divi[16]), .A2(n19811), 
        .B(n19002), .C(n24631), .Y(n19812) );
  A2O1A1Ixp33_ASAP7_75t_SL U21385 ( .A1(n22374), .A2(n19002), .B(n28333), .C(
        n19002), .Y(n19804) );
  A2O1A1Ixp33_ASAP7_75t_SL U21386 ( .A1(n18805), .A2(n19002), .B(n32628), .C(
        n19002), .Y(n19805) );
  A2O1A1Ixp33_ASAP7_75t_SL U21387 ( .A1(n22373), .A2(n19002), .B(n28563), .C(
        n19002), .Y(n19806) );
  O2A1O1Ixp5_ASAP7_75t_SL U21388 ( .A1(n19804), .A2(n19805), .B(n19002), .C(
        n19806), .Y(n28576) );
  A2O1A1Ixp33_ASAP7_75t_SL U21389 ( .A1(n22374), .A2(n19002), .B(n28370), .C(
        n19002), .Y(n19801) );
  A2O1A1Ixp33_ASAP7_75t_SL U21390 ( .A1(n18806), .A2(n19002), .B(n32734), .C(
        n19002), .Y(n19802) );
  A2O1A1Ixp33_ASAP7_75t_SL U21391 ( .A1(n22373), .A2(n19002), .B(n26752), .C(
        n19002), .Y(n19803) );
  O2A1O1Ixp5_ASAP7_75t_SL U21392 ( .A1(n19801), .A2(n19802), .B(n19002), .C(
        n19803), .Y(n31339) );
  O2A1O1Ixp33_ASAP7_75t_SL U21393 ( .A1(add_x_746_n23), .A2(add_x_746_n2), .B(
        n19002), .C(n19800), .Y(add_x_746_n17) );
  A2O1A1Ixp33_ASAP7_75t_SL U21394 ( .A1(uart1_r_RXSTATE__1_), .A2(n19002), .B(
        n19799), .C(n19002), .Y(n29966) );
  A2O1A1Ixp33_ASAP7_75t_SL U21395 ( .A1(n22376), .A2(n19002), .B(n30388), .C(
        n19798), .Y(n27169) );
  INVx1_ASAP7_75t_SL U21396 ( .A(n22392), .Y(n18661) );
  A2O1A1Ixp33_ASAP7_75t_SL U21397 ( .A1(n19002), .A2(n24796), .B(n30906), .C(
        n19427), .Y(n30938) );
  O2A1O1Ixp33_ASAP7_75t_SL U21398 ( .A1(n28833), .A2(n29307), .B(n19002), .C(
        n19791), .Y(n29279) );
  A2O1A1Ixp33_ASAP7_75t_SL U21399 ( .A1(n19002), .A2(n28452), .B(n31660), .C(
        n19625), .Y(n19626) );
  A2O1A1Ixp33_ASAP7_75t_SL U21400 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[24]), 
        .B(n19626), .C(n19002), .Y(n19627) );
  A2O1A1Ixp33_ASAP7_75t_SL U21401 ( .A1(n18364), .A2(n19002), .B(
        mult_x_1196_n2739), .C(n19002), .Y(n19781) );
  A2O1A1Ixp33_ASAP7_75t_SL U21402 ( .A1(n24040), .A2(n19002), .B(
        mult_x_1196_n2738), .C(n19002), .Y(n19782) );
  A2O1A1Ixp33_ASAP7_75t_SL U21403 ( .A1(n19781), .A2(n19002), .B(n19782), .C(
        n19002), .Y(n21251) );
  A2O1A1Ixp33_ASAP7_75t_SL U21404 ( .A1(n24043), .A2(n19002), .B(n19780), .C(
        n19002), .Y(mult_x_1196_n2150) );
  A2O1A1Ixp33_ASAP7_75t_SL U21405 ( .A1(uart1_r_RSEMPTY_), .A2(n19184), .B(
        n19191), .C(n19002), .Y(n4696) );
  A2O1A1Ixp33_ASAP7_75t_SL U21406 ( .A1(uart1_r_RHOLD__15__3_), .A2(n31213), 
        .B(n19565), .C(n19002), .Y(n19566) );
  A2O1A1Ixp33_ASAP7_75t_SL U21407 ( .A1(uart1_r_RHOLD__19__3_), .A2(n31208), 
        .B(n19570), .C(n19002), .Y(n19571) );
  A2O1A1Ixp33_ASAP7_75t_SL U21408 ( .A1(uart1_r_RHOLD__6__3_), .A2(n31226), 
        .B(n19576), .C(n19002), .Y(n19577) );
  A2O1A1Ixp33_ASAP7_75t_SL U21409 ( .A1(uart1_r_RHOLD__16__3_), .A2(n31205), 
        .B(n19581), .C(n19002), .Y(n19582) );
  A2O1A1Ixp33_ASAP7_75t_SL U21410 ( .A1(uart1_r_RHOLD__9__3_), .A2(n31204), 
        .B(n19584), .C(n19002), .Y(n19585) );
  A2O1A1Ixp33_ASAP7_75t_SL U21411 ( .A1(uart1_r_RHOLD__27__3_), .A2(n31230), 
        .B(n19589), .C(n19002), .Y(n19590) );
  O2A1O1Ixp33_ASAP7_75t_SL U21412 ( .A1(n19555), .A2(n19604), .B(n19002), .C(
        n19605), .Y(n19606) );
  A2O1A1Ixp33_ASAP7_75t_SL U21413 ( .A1(uart1_r_RHOLD__0__3_), .A2(n31242), 
        .B(n19615), .C(n19002), .Y(n19616) );
  A2O1A1Ixp33_ASAP7_75t_SL U21414 ( .A1(n19002), .A2(n32004), .B(n28254), .C(
        n28253), .Y(n19618) );
  A2O1A1Ixp33_ASAP7_75t_SL U21415 ( .A1(n31954), .A2(n19617), .B(n19618), .C(
        n19002), .Y(n4694) );
  A2O1A1Ixp33_ASAP7_75t_SL U21416 ( .A1(n4519), .A2(n19002), .B(n4518), .C(
        n19002), .Y(n19779) );
  A2O1A1Ixp33_ASAP7_75t_SL U21417 ( .A1(n19002), .A2(n19549), .B(n19550), .C(
        n19002), .Y(n19551) );
  A2O1A1Ixp33_ASAP7_75t_SL U21418 ( .A1(u0_0_leon3x0_p0_div0_addout_32_), .A2(
        n19757), .B(n31677), .C(n19002), .Y(n19758) );
  A2O1A1Ixp33_ASAP7_75t_SL U21419 ( .A1(u0_0_leon3x0_p0_div0_addout_32_), .A2(
        n19002), .B(n19757), .C(n19758), .Y(n19759) );
  A2O1A1Ixp33_ASAP7_75t_SL U21420 ( .A1(n23375), .A2(n19002), .B(
        add_x_735_A_2_), .C(n19002), .Y(n19760) );
  A2O1A1Ixp33_ASAP7_75t_SL U21421 ( .A1(u0_0_leon3x0_p0_muli[41]), .A2(n19002), 
        .B(n22837), .C(n19002), .Y(n19761) );
  A2O1A1Ixp33_ASAP7_75t_SL U21422 ( .A1(n23964), .A2(n19002), .B(n18296), .C(
        n19002), .Y(n19763) );
  A2O1A1Ixp33_ASAP7_75t_SL U21423 ( .A1(n23960), .A2(n19002), .B(n22939), .C(
        n19002), .Y(n19764) );
  A2O1A1Ixp33_ASAP7_75t_SL U21424 ( .A1(n19766), .A2(n19002), .B(n19767), .C(
        n19002), .Y(n19768) );
  A2O1A1Ixp33_ASAP7_75t_SL U21425 ( .A1(n24231), .A2(n19002), .B(n18606), .C(
        n19002), .Y(n19771) );
  A2O1A1Ixp33_ASAP7_75t_SL U21426 ( .A1(n22968), .A2(n19002), .B(n23665), .C(
        n19002), .Y(n19772) );
  A2O1A1Ixp33_ASAP7_75t_SL U21427 ( .A1(n23091), .A2(n19002), .B(n23965), .C(
        n19002), .Y(n19775) );
  A2O1A1Ixp33_ASAP7_75t_SL U21428 ( .A1(n19773), .A2(n19002), .B(n19776), .C(
        n19002), .Y(n19777) );
  OAI21xp5_ASAP7_75t_SL U21429 ( .A1(n18491), .A2(n23396), .B(n19002), .Y(
        n19774) );
  A2O1A1Ixp33_ASAP7_75t_SL U21430 ( .A1(n30390), .A2(n19002), .B(n31404), .C(
        n19002), .Y(n19749) );
  A2O1A1Ixp33_ASAP7_75t_SL U21431 ( .A1(n19751), .A2(n19002), .B(n19754), .C(
        n19002), .Y(n19755) );
  A2O1A1Ixp33_ASAP7_75t_SL U21432 ( .A1(n25768), .A2(n19002), .B(n30575), .C(
        n19002), .Y(n19744) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21433 ( .A1(n28411), .A2(n30885), .B(n19744), 
        .C(n19002), .D(n30578), .Y(n4360) );
  A2O1A1Ixp33_ASAP7_75t_SL U21434 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_M__NALIGN_), .C(n19736), .Y(n4091) );
  A2O1A1Ixp33_ASAP7_75t_SL U21435 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__31_), .B(n24654), .C(n19327), .Y(
        n4067) );
  A2O1A1Ixp33_ASAP7_75t_SL U21436 ( .A1(n22420), .A2(n19002), .B(n27223), .C(
        n31422), .Y(n19726) );
  A2O1A1Ixp33_ASAP7_75t_SL U21437 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[16]), 
        .B(n19726), .C(n19002), .Y(n19727) );
  A2O1A1Ixp33_ASAP7_75t_SL U21438 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_16_), .B(n19729), .C(n19002), .Y(n3990) );
  A2O1A1Ixp33_ASAP7_75t_SL U21439 ( .A1(n22393), .A2(n19002), .B(n3905), .C(
        n19002), .Y(n19724) );
  A2O1A1Ixp33_ASAP7_75t_SL U21440 ( .A1(n32042), .A2(
        u0_0_leon3x0_p0_c0mmu_a0_r_BO__0_), .B(n19724), .C(n19002), .Y(n3904)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21441 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__TRAP_), 
        .A2(n19002), .B(n23229), .C(n19721), .Y(n3733) );
  O2A1O1Ixp5_ASAP7_75t_SL U21442 ( .A1(n31263), .A2(n30210), .B(n19002), .C(
        n19696), .Y(n19697) );
  A2O1A1Ixp33_ASAP7_75t_SL U21443 ( .A1(n24549), .A2(n19002), .B(n19699), .C(
        n19002), .Y(n19700) );
  A2O1A1Ixp33_ASAP7_75t_SL U21444 ( .A1(n19700), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_RBURST_), .C(n19701), .Y(n2971) );
  A2O1A1Ixp33_ASAP7_75t_SL U21445 ( .A1(n29383), .A2(n19002), .B(apbi[2]), .C(
        n19695), .Y(n2855) );
  A2O1A1Ixp33_ASAP7_75t_SL U21446 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_A__CWP__1_), .B(n24657), .C(n19303), .Y(n2800) );
  A2O1A1Ixp33_ASAP7_75t_SL U21447 ( .A1(n29956), .A2(n19002), .B(n31098), .C(
        n19002), .Y(n19691) );
  A2O1A1Ixp33_ASAP7_75t_SL U21448 ( .A1(n31099), .A2(n19002), .B(n26069), .C(
        n19002), .Y(n19692) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21449 ( .A1(n31101), .A2(uart1_r_RHOLD__29__0_), 
        .B(n19691), .C(n19002), .D(n19692), .Y(n2443) );
  A2O1A1Ixp33_ASAP7_75t_SL U21450 ( .A1(n32875), .A2(n19002), .B(n2357), .C(
        n19690), .Y(n17778) );
  A2O1A1Ixp33_ASAP7_75t_SL U21451 ( .A1(n19002), .A2(n27968), .B(
        uart1_r_THOLD__19__0_), .C(n19490), .Y(n2262) );
  A2O1A1Ixp33_ASAP7_75t_SL U21452 ( .A1(n19002), .A2(n27929), .B(
        uart1_r_THOLD__9__0_), .C(n19489), .Y(n2255) );
  A2O1A1Ixp33_ASAP7_75t_SL U21453 ( .A1(dataout[5]), .A2(n19002), .B(n19682), 
        .C(n19002), .Y(n19683) );
  A2O1A1Ixp33_ASAP7_75t_SL U21454 ( .A1(n32567), .A2(n19002), .B(n32585), .C(
        n19002), .Y(n19678) );
  A2O1A1Ixp33_ASAP7_75t_SL U21455 ( .A1(n32584), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__5_), .B(n19678), .C(n19002), .Y(
        n19679) );
  A2O1A1Ixp33_ASAP7_75t_SL U21456 ( .A1(n32590), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__5_), .B(n19680), .C(n19002), 
        .Y(n19681) );
  A2O1A1Ixp33_ASAP7_75t_SL U21457 ( .A1(n32568), .A2(n19002), .B(n32595), .C(
        n19681), .Y(ic_address[3]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21458 ( .A1(n32387), .A2(n19002), .B(n32431), .C(
        n19002), .Y(n19664) );
  A2O1A1Ixp33_ASAP7_75t_SL U21459 ( .A1(n32644), .A2(n19002), .B(n32429), .C(
        n19002), .Y(n19665) );
  A2O1A1Ixp33_ASAP7_75t_SL U21460 ( .A1(n32384), .A2(n19002), .B(n24543), .C(
        n19002), .Y(n19666) );
  A2O1A1Ixp33_ASAP7_75t_SL U21461 ( .A1(n19665), .A2(n19002), .B(n19666), .C(
        n19002), .Y(n19667) );
  A2O1A1Ixp33_ASAP7_75t_SL U21462 ( .A1(n19664), .A2(n19002), .B(n19669), .C(
        n19002), .Y(n19670) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21463 ( .A1(n29721), .A2(n29719), .B(n19002), 
        .C(n30704), .Y(n19659) );
  A2O1A1Ixp33_ASAP7_75t_SL U21464 ( .A1(n29999), .A2(ahbso_0__HRDATA__13_), 
        .B(n19658), .C(n19002), .Y(n30808) );
  A2O1A1Ixp33_ASAP7_75t_SL U21465 ( .A1(n22376), .A2(n19002), .B(n30699), .C(
        n19654), .Y(n28714) );
  A2O1A1Ixp33_ASAP7_75t_SL U21466 ( .A1(n22375), .A2(n19002), .B(n29815), .C(
        n19653), .Y(n26735) );
  O2A1O1Ixp5_ASAP7_75t_SL U21467 ( .A1(n19459), .A2(n19460), .B(n19002), .C(
        n19461), .Y(n30381) );
  A2O1A1Ixp33_ASAP7_75t_SL U21468 ( .A1(DP_OP_5187J1_124_3275_n271), .A2(
        n19002), .B(n19649), .C(n19002), .Y(n19650) );
  A2O1A1Ixp33_ASAP7_75t_SL U21469 ( .A1(n19650), .A2(n19002), .B(n19651), .C(
        n19652), .Y(u0_0_leon3x0_p0_div0_addout_6_) );
  A2O1A1Ixp33_ASAP7_75t_SL U21470 ( .A1(n19002), .A2(DP_OP_1196_128_7433_n57), 
        .B(DP_OP_1196_128_7433_n67), .C(DP_OP_1196_128_7433_n60), .Y(n19450)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21471 ( .A1(n29865), .A2(n19002), .B(n29495), .C(
        n19002), .Y(n19641) );
  A2O1A1Ixp33_ASAP7_75t_SL U21472 ( .A1(n19641), .A2(n19002), .B(n19644), .C(
        n19002), .Y(n19645) );
  A2O1A1Ixp33_ASAP7_75t_SL U21473 ( .A1(n29728), .A2(n19002), .B(n29733), .C(
        n19640), .Y(n29729) );
  A2O1A1Ixp33_ASAP7_75t_SL U21474 ( .A1(n22968), .A2(n19002), .B(n29148), .C(
        n19002), .Y(n19633) );
  A2O1A1Ixp33_ASAP7_75t_SL U21475 ( .A1(n29150), .A2(n22968), .B(n19633), .C(
        n19002), .Y(n19634) );
  O2A1O1Ixp33_ASAP7_75t_SL U21476 ( .A1(u0_0_leon3x0_p0_divi[28]), .A2(n19634), 
        .B(n19002), .C(n24631), .Y(n19635) );
  A2O1A1Ixp33_ASAP7_75t_SL U21477 ( .A1(n24690), .A2(n19002), .B(n29146), .C(
        n24579), .Y(n19637) );
  A2O1A1Ixp33_ASAP7_75t_SL U21478 ( .A1(n19636), .A2(n19002), .B(n19637), .C(
        n19002), .Y(n19638) );
  A2O1A1Ixp33_ASAP7_75t_SL U21479 ( .A1(n19635), .A2(n19002), .B(n19638), .C(
        n19002), .Y(n19639) );
  A2O1A1Ixp33_ASAP7_75t_SL U21480 ( .A1(n24690), .A2(n25900), .B(n19639), .C(
        n19002), .Y(n30225) );
  A2O1A1Ixp33_ASAP7_75t_SL U21481 ( .A1(n32459), .A2(n19002), .B(n19632), .C(
        n19002), .Y(n32518) );
  A2O1A1Ixp33_ASAP7_75t_SL U21482 ( .A1(n32353), .A2(n19002), .B(n32628), .C(
        n19002), .Y(n19631) );
  A2O1A1Ixp33_ASAP7_75t_SL U21483 ( .A1(n32353), .A2(n19002), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[1]), .C(n19002), .Y(n19630) );
  A2O1A1Ixp33_ASAP7_75t_SL U21484 ( .A1(n29307), .A2(n19002), .B(irqo[0]), .C(
        n19002), .Y(n19629) );
  A2O1A1Ixp33_ASAP7_75t_SL U21485 ( .A1(n19186), .A2(n19187), .B(n19190), .C(
        n19002), .Y(n19191) );
  A2O1A1Ixp33_ASAP7_75t_SL U21486 ( .A1(n2840), .A2(n19002), .B(n19554), .C(
        n19002), .Y(n19555) );
  A2O1A1Ixp33_ASAP7_75t_SL U21487 ( .A1(n19556), .A2(n19002), .B(n19559), .C(
        n19002), .Y(n19560) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21488 ( .A1(n19002), .A2(n19561), .B(n19572), 
        .C(n19002), .D(n19591), .Y(n19592) );
  A2O1A1Ixp33_ASAP7_75t_SL U21489 ( .A1(n31238), .A2(n19002), .B(n19592), .C(
        n19593), .Y(n19594) );
  A2O1A1Ixp33_ASAP7_75t_SL U21490 ( .A1(sr1_r_MCFG2__RAMWWS__1_), .A2(n31250), 
        .B(n19597), .C(n19002), .Y(n19598) );
  A2O1A1Ixp33_ASAP7_75t_SL U21491 ( .A1(n19002), .A2(n19594), .B(n19600), .C(
        n19002), .Y(n19601) );
  A2O1A1Ixp33_ASAP7_75t_SL U21492 ( .A1(n19002), .A2(n30872), .B(n28249), .C(
        n19002), .Y(n19605) );
  A2O1A1Ixp33_ASAP7_75t_SL U21493 ( .A1(irqctrl0_r_ILEVEL__3_), .A2(n31248), 
        .B(n19612), .C(n19002), .Y(n19613) );
  A2O1A1Ixp33_ASAP7_75t_SL U21494 ( .A1(n29806), .A2(n19002), .B(n32110), .C(
        n19002), .Y(n19549) );
  A2O1A1Ixp33_ASAP7_75t_SL U21495 ( .A1(n31046), .A2(n19002), .B(n31045), .C(
        n19002), .Y(n19543) );
  O2A1O1Ixp33_ASAP7_75t_SL U21496 ( .A1(n19543), .A2(n31047), .B(n19002), .C(
        n19546), .Y(n4453) );
  A2O1A1Ixp33_ASAP7_75t_SL U21497 ( .A1(u0_0_leon3x0_p0_divi[55]), .A2(n30430), 
        .B(n19161), .C(n19002), .Y(n19162) );
  A2O1A1Ixp33_ASAP7_75t_SL U21498 ( .A1(n26910), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n19534) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21499 ( .A1(n30644), .A2(n26950), .B(n19534), 
        .C(n19002), .D(n19537), .Y(n19538) );
  A2O1A1Ixp33_ASAP7_75t_SL U21500 ( .A1(n30645), .A2(n19002), .B(n26953), .C(
        n19538), .Y(n19539) );
  A2O1A1Ixp33_ASAP7_75t_SL U21501 ( .A1(n26955), .A2(n22432), .B(n19539), .C(
        n19002), .Y(n19540) );
  A2O1A1Ixp33_ASAP7_75t_SL U21502 ( .A1(n28799), .A2(n19002), .B(n19540), .C(
        n19002), .Y(n19541) );
  A2O1A1Ixp33_ASAP7_75t_SL U21503 ( .A1(n32043), .A2(n19002), .B(n10988), .C(
        n19530), .Y(u0_0_leon3x0_p0_c0mmu_a0_v_BO__1_) );
  A2O1A1Ixp33_ASAP7_75t_SL U21504 ( .A1(n19002), .A2(n19320), .B(n19321), .C(
        n19002), .Y(n19322) );
  A2O1A1Ixp33_ASAP7_75t_SL U21505 ( .A1(n22427), .A2(n19002), .B(n31657), .C(
        n19527), .Y(n3719) );
  A2O1A1Ixp33_ASAP7_75t_SL U21506 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__12_), .A2(n19002), .B(n22428), .C(
        n19525), .Y(n3642) );
  A2O1A1Ixp33_ASAP7_75t_SL U21507 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_), .A2(n19002), .B(n24657), .C(
        n19523), .Y(n3621) );
  A2O1A1Ixp33_ASAP7_75t_SL U21508 ( .A1(n19002), .A2(u0_0_leon3x0_p0_ici[36]), 
        .B(n24652), .C(n19313), .Y(n3436) );
  A2O1A1Ixp33_ASAP7_75t_SL U21509 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_W__S__WIM__5_), .C(n19516), .Y(n3334) );
  A2O1A1Ixp33_ASAP7_75t_SL U21510 ( .A1(n30701), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__8_), .C(n19515), .Y(n3329) );
  A2O1A1Ixp33_ASAP7_75t_SL U21511 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__29_), 
        .A2(n19002), .B(n24650), .C(n19514), .Y(n3284) );
  A2O1A1Ixp33_ASAP7_75t_SL U21512 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__23_), 
        .A2(n19002), .B(n24651), .C(n19512), .Y(n3244) );
  A2O1A1Ixp33_ASAP7_75t_SL U21513 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__2_), 
        .A2(n19002), .B(n24653), .C(n19510), .Y(n3192) );
  A2O1A1Ixp33_ASAP7_75t_SL U21514 ( .A1(n19002), .A2(n19508), .B(n22380), .C(
        n19002), .Y(n18096) );
  A2O1A1Ixp33_ASAP7_75t_SL U21515 ( .A1(n29383), .A2(n19002), .B(apbi[4]), .C(
        n19506), .Y(n2853) );
  A2O1A1Ixp33_ASAP7_75t_SL U21516 ( .A1(n19002), .A2(n31840), .B(apbi[10]), 
        .C(n19307), .Y(n2837) );
  A2O1A1Ixp33_ASAP7_75t_SL U21517 ( .A1(n31664), .A2(n19002), .B(n31418), .C(
        n19002), .Y(n19503) );
  A2O1A1Ixp33_ASAP7_75t_SL U21518 ( .A1(n22421), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_W__S__CWP__1_), .C(n19501), .Y(n2804) );
  A2O1A1Ixp33_ASAP7_75t_SL U21519 ( .A1(n22420), .A2(n19002), .B(n27264), .C(
        n31422), .Y(n19497) );
  A2O1A1Ixp33_ASAP7_75t_SL U21520 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[17]), 
        .B(n19497), .C(n19002), .Y(n19498) );
  A2O1A1Ixp33_ASAP7_75t_SL U21521 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_17_), .B(n19500), .C(n19002), .Y(n2611) );
  A2O1A1Ixp33_ASAP7_75t_SL U21522 ( .A1(n31098), .A2(n19002), .B(n26126), .C(
        n19002), .Y(n19495) );
  A2O1A1Ixp33_ASAP7_75t_SL U21523 ( .A1(n31099), .A2(n19002), .B(n26127), .C(
        n19002), .Y(n19496) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21524 ( .A1(n31101), .A2(uart1_r_RHOLD__29__1_), 
        .B(n19495), .C(n19002), .D(n19496), .Y(n2442) );
  A2O1A1Ixp33_ASAP7_75t_SL U21525 ( .A1(n22420), .A2(n19002), .B(n27176), .C(
        n31422), .Y(n19491) );
  A2O1A1Ixp33_ASAP7_75t_SL U21526 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[9]), 
        .B(n19491), .C(n19002), .Y(n19492) );
  A2O1A1Ixp33_ASAP7_75t_SL U21527 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_9_), .B(n19494), .C(n19002), .Y(n2318) );
  A2O1A1Ixp33_ASAP7_75t_SL U21528 ( .A1(n5014), .A2(n26086), .B(n26087), .C(
        n19002), .Y(n19293) );
  A2O1A1Ixp33_ASAP7_75t_SL U21529 ( .A1(n19002), .A2(n24633), .B(
        uart1_r_TFIFOIRQEN_), .C(n19292), .Y(n1801) );
  A2O1A1Ixp33_ASAP7_75t_SL U21530 ( .A1(dataout[6]), .A2(n19002), .B(n19486), 
        .C(n19002), .Y(n19487) );
  A2O1A1Ixp33_ASAP7_75t_SL U21531 ( .A1(n19002), .A2(n22433), .B(n32971), .C(
        n19289), .Y(n1703) );
  A2O1A1Ixp33_ASAP7_75t_SL U21532 ( .A1(n22386), .A2(n19002), .B(n33008), .C(
        n19485), .Y(n1677) );
  A2O1A1Ixp33_ASAP7_75t_SL U21533 ( .A1(n19002), .A2(n22421), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[0]), .C(n19286), .Y(n3910) );
  A2O1A1Ixp33_ASAP7_75t_SL U21534 ( .A1(n32630), .A2(n19002), .B(n32543), .C(
        n19482), .Y(it_data[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21535 ( .A1(n32638), .A2(n19002), .B(n32429), .C(
        n19002), .Y(n19470) );
  A2O1A1Ixp33_ASAP7_75t_SL U21536 ( .A1(n32376), .A2(n19002), .B(n32431), .C(
        n19002), .Y(n19471) );
  A2O1A1Ixp33_ASAP7_75t_SL U21537 ( .A1(dc_q[20]), .A2(n32385), .B(n19471), 
        .C(n19002), .Y(n19472) );
  A2O1A1Ixp33_ASAP7_75t_SL U21538 ( .A1(n32377), .A2(n19002), .B(n24543), .C(
        n19472), .Y(n19473) );
  A2O1A1Ixp33_ASAP7_75t_SL U21539 ( .A1(n19470), .A2(n19002), .B(n19473), .C(
        n19002), .Y(n19474) );
  A2O1A1Ixp33_ASAP7_75t_SL U21540 ( .A1(n32381), .A2(n19002), .B(n32378), .C(
        n19474), .Y(dc_data[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21541 ( .A1(n31680), .A2(n19002), .B(n22376), .C(
        n19002), .Y(n19468) );
  A2O1A1Ixp33_ASAP7_75t_SL U21542 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__31_), .B(n19468), .C(n19002), .Y(
        n26734) );
  A2O1A1Ixp33_ASAP7_75t_SL U21543 ( .A1(n30643), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n19462) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21544 ( .A1(n30644), .A2(n31335), .B(n19462), 
        .C(n19002), .D(n19465), .Y(n19466) );
  A2O1A1Ixp33_ASAP7_75t_SL U21545 ( .A1(n30645), .A2(n19002), .B(n31339), .C(
        n19466), .Y(n19467) );
  A2O1A1Ixp33_ASAP7_75t_SL U21546 ( .A1(n22432), .A2(n31350), .B(n19467), .C(
        n19002), .Y(n30646) );
  A2O1A1Ixp33_ASAP7_75t_SL U21547 ( .A1(n18805), .A2(n19002), .B(n32620), .C(
        n19002), .Y(n19459) );
  A2O1A1Ixp33_ASAP7_75t_SL U21548 ( .A1(n22374), .A2(n19002), .B(n28697), .C(
        n19002), .Y(n19460) );
  A2O1A1Ixp33_ASAP7_75t_SL U21549 ( .A1(n22373), .A2(n19002), .B(n28698), .C(
        n19002), .Y(n19461) );
  A2O1A1Ixp33_ASAP7_75t_SL U21550 ( .A1(u0_0_leon3x0_p0_iu_de_icc_1_), .A2(
        n30652), .B(n24680), .C(n19002), .Y(n19458) );
  A2O1A1Ixp33_ASAP7_75t_SL U21551 ( .A1(DP_OP_1196_128_7433_n57), .A2(n19002), 
        .B(DP_OP_1196_128_7433_n66), .C(n19002), .Y(n19446) );
  A2O1A1Ixp33_ASAP7_75t_SL U21552 ( .A1(n19449), .A2(n19002), .B(n19450), .C(
        n19002), .Y(n19451) );
  A2O1A1Ixp33_ASAP7_75t_SL U21553 ( .A1(n19449), .A2(n19002), .B(n19450), .C(
        n19454), .Y(n19455) );
  A2O1A1Ixp33_ASAP7_75t_SL U21554 ( .A1(DP_OP_1196_128_7433_n50), .A2(n19002), 
        .B(n19452), .C(n19455), .Y(u0_0_leon3x0_p0_iu_N5494) );
  A2O1A1Ixp33_ASAP7_75t_SL U21555 ( .A1(n29733), .A2(n19002), .B(n29640), .C(
        n19443), .Y(n29648) );
  A2O1A1Ixp33_ASAP7_75t_SL U21556 ( .A1(n29195), .A2(n19002), .B(n29206), .C(
        n19002), .Y(n19442) );
  A2O1A1Ixp33_ASAP7_75t_SL U21557 ( .A1(n29206), .A2(
        u0_0_leon3x0_p0_iu_v_A__CWP__1_), .B(n19442), .C(n19002), .Y(n26813)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21558 ( .A1(n28352), .A2(n19002), .B(n31660), .C(
        n19432), .Y(n19433) );
  A2O1A1Ixp33_ASAP7_75t_SL U21559 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[5]), 
        .B(n19433), .C(n19002), .Y(n19434) );
  A2O1A1Ixp33_ASAP7_75t_SL U21560 ( .A1(n32200), .A2(n19002), .B(n32455), .C(
        n19002), .Y(n19428) );
  A2O1A1Ixp33_ASAP7_75t_SL U21561 ( .A1(n19002), .A2(n22392), .B(n23164), .C(
        n19011), .Y(n26597) );
  A2O1A1Ixp33_ASAP7_75t_SL U21562 ( .A1(n19002), .A2(n28336), .B(n31660), .C(
        n19213), .Y(n19214) );
  A2O1A1Ixp33_ASAP7_75t_SL U21563 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[12]), 
        .B(n19214), .C(n19002), .Y(n19215) );
  A2O1A1Ixp33_ASAP7_75t_SL U21564 ( .A1(n28303), .A2(n19002), .B(n31660), .C(
        n19422), .Y(n19423) );
  A2O1A1Ixp33_ASAP7_75t_SL U21565 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[27]), 
        .B(n19423), .C(n19002), .Y(n19424) );
  A2O1A1Ixp33_ASAP7_75t_SL U21566 ( .A1(n31250), .A2(sr1_r_MCFG2__RAMWWS__0_), 
        .B(n19362), .C(n19002), .Y(n19363) );
  A2O1A1Ixp33_ASAP7_75t_SL U21567 ( .A1(uart1_r_RHOLD__0__2_), .A2(n31242), 
        .B(n19365), .C(n19002), .Y(n19366) );
  A2O1A1Ixp33_ASAP7_75t_SL U21568 ( .A1(n2842), .A2(n19002), .B(n31953), .C(
        n19366), .Y(n19367) );
  A2O1A1Ixp33_ASAP7_75t_SL U21569 ( .A1(n31225), .A2(uart1_r_RHOLD__10__2_), 
        .B(n19371), .C(n19002), .Y(n19372) );
  A2O1A1Ixp33_ASAP7_75t_SL U21570 ( .A1(n31229), .A2(uart1_r_RHOLD__22__2_), 
        .B(n19376), .C(n19002), .Y(n19377) );
  A2O1A1Ixp33_ASAP7_75t_SL U21571 ( .A1(n31212), .A2(uart1_r_RHOLD__26__2_), 
        .B(n19381), .C(n19002), .Y(n19382) );
  A2O1A1Ixp33_ASAP7_75t_SL U21572 ( .A1(n31208), .A2(uart1_r_RHOLD__19__2_), 
        .B(n19386), .C(n19002), .Y(n19387) );
  A2O1A1Ixp33_ASAP7_75t_SL U21573 ( .A1(n31200), .A2(uart1_r_RHOLD__5__2_), 
        .B(n19393), .C(n19002), .Y(n19394) );
  A2O1A1Ixp33_ASAP7_75t_SL U21574 ( .A1(n31216), .A2(uart1_r_RHOLD__3__2_), 
        .B(n19398), .C(n19002), .Y(n19399) );
  A2O1A1Ixp33_ASAP7_75t_SL U21575 ( .A1(n31220), .A2(uart1_r_RHOLD__13__2_), 
        .B(n19403), .C(n19002), .Y(n19404) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21576 ( .A1(n31202), .A2(uart1_r_RHOLD__12__2_), 
        .B(n19389), .C(n19002), .D(n19405), .Y(n19406) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21577 ( .A1(n30870), .A2(n19407), .B(n19410), 
        .C(n19002), .D(n19413), .Y(n19414) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21578 ( .A1(n31241), .A2(uart1_r_RHOLD__24__2_), 
        .B(n19367), .C(n19002), .D(n19417), .Y(n19418) );
  A2O1A1Ixp33_ASAP7_75t_SL U21579 ( .A1(n29559), .A2(n31240), .B(n19421), .C(
        n19002), .Y(n16838) );
  O2A1O1Ixp33_ASAP7_75t_SL U21580 ( .A1(n31543), .A2(n31544), .B(n19002), .C(
        n32110), .Y(n19166) );
  A2O1A1Ixp33_ASAP7_75t_SL U21581 ( .A1(n31759), .A2(n19002), .B(n31758), .C(
        n19002), .Y(n19358) );
  A2O1A1Ixp33_ASAP7_75t_SL U21582 ( .A1(n31760), .A2(n19002), .B(n19358), .C(
        n19002), .Y(n33061) );
  A2O1A1Ixp33_ASAP7_75t_SL U21583 ( .A1(n30566), .A2(n19002), .B(n31045), .C(
        n19002), .Y(n19345) );
  O2A1O1Ixp33_ASAP7_75t_SL U21584 ( .A1(n19345), .A2(n31047), .B(n19002), .C(
        n19348), .Y(n4429) );
  A2O1A1Ixp33_ASAP7_75t_SL U21585 ( .A1(n28805), .A2(n30644), .B(n19337), .C(
        n19002), .Y(n19338) );
  A2O1A1Ixp33_ASAP7_75t_SL U21586 ( .A1(n31868), .A2(n28806), .B(n19340), .C(
        n19002), .Y(n19341) );
  A2O1A1Ixp33_ASAP7_75t_SL U21587 ( .A1(n24541), .A2(n19002), .B(n28807), .C(
        n19341), .Y(n19342) );
  A2O1A1Ixp33_ASAP7_75t_SL U21588 ( .A1(n28808), .A2(n19002), .B(n19342), .C(
        n19002), .Y(n19343) );
  A2O1A1Ixp33_ASAP7_75t_SL U21589 ( .A1(mult_x_1196_n744), .A2(n19002), .B(
        mult_x_1196_n747), .C(n19002), .Y(n19332) );
  A2O1A1Ixp33_ASAP7_75t_SL U21590 ( .A1(n24646), .A2(n19002), .B(n29807), .C(
        n19328), .Y(n4127) );
  A2O1A1Ixp33_ASAP7_75t_SL U21591 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PV_), .B(n24650), .C(n19138), .Y(n4020)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21592 ( .A1(u0_0_leon3x0_p0_iu_r_E__CTRL__ANNUL_), 
        .A2(n19002), .B(n31812), .C(n19002), .Y(n19320) );
  A2O1A1Ixp33_ASAP7_75t_SL U21593 ( .A1(u0_0_leon3x0_p0_iu_r_A__JMPL_), .A2(
        n19002), .B(u0_0_leon3x0_p0_iu_r_A__CTRL__RETT_), .C(n19002), .Y(
        n19321) );
  A2O1A1Ixp33_ASAP7_75t_SL U21594 ( .A1(n19324), .A2(n19002), .B(n24646), .C(
        n19002), .Y(n19325) );
  O2A1O1Ixp5_ASAP7_75t_SL U21595 ( .A1(n19130), .A2(n19131), .B(n19002), .C(
        n30580), .Y(n19132) );
  A2O1A1Ixp33_ASAP7_75t_SL U21596 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__0_), 
        .A2(n19002), .B(n24655), .C(n19314), .Y(n3526) );
  A2O1A1Ixp33_ASAP7_75t_SL U21597 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__23_), 
        .A2(n19002), .B(n24651), .C(n19311), .Y(n3242) );
  A2O1A1Ixp33_ASAP7_75t_SL U21598 ( .A1(n19002), .A2(n22396), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[3]), .C(n19115), .Y(n3083) );
  A2O1A1Ixp33_ASAP7_75t_SL U21599 ( .A1(n19002), .A2(n29383), .B(apbi[3]), .C(
        n19113), .Y(n2854) );
  A2O1A1Ixp33_ASAP7_75t_SL U21600 ( .A1(n22422), .A2(n19002), .B(n4325), .C(
        n19002), .Y(n19304) );
  A2O1A1Ixp33_ASAP7_75t_SL U21601 ( .A1(n22422), .A2(n19002), .B(n4325), .C(
        n28379), .Y(n19305) );
  A2O1A1Ixp33_ASAP7_75t_SL U21602 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_W__S__WIM__3_), .C(n19301), .Y(n2737) );
  A2O1A1Ixp33_ASAP7_75t_SL U21603 ( .A1(n22420), .A2(n19002), .B(n28322), .C(
        n31422), .Y(n19297) );
  A2O1A1Ixp33_ASAP7_75t_SL U21604 ( .A1(n31421), .A2(u0_0_leon3x0_p0_divo[18]), 
        .B(n19297), .C(n19002), .Y(n19298) );
  A2O1A1Ixp33_ASAP7_75t_SL U21605 ( .A1(n24639), .A2(
        u0_0_leon3x0_p0_div0_addout_18_), .B(n19300), .C(n19002), .Y(n2587) );
  A2O1A1Ixp33_ASAP7_75t_SL U21606 ( .A1(n32786), .A2(n19002), .B(n32728), .C(
        n19296), .Y(n2361) );
  A2O1A1Ixp33_ASAP7_75t_SL U21607 ( .A1(n32749), .A2(writen), .B(n19295), .C(
        n19002), .Y(n2301) );
  A2O1A1Ixp33_ASAP7_75t_SL U21608 ( .A1(n19002), .A2(n27946), .B(
        uart1_r_THOLD__16__0_), .C(n19105), .Y(n2261) );
  A2O1A1Ixp33_ASAP7_75t_SL U21609 ( .A1(n19002), .A2(n27951), .B(
        uart1_r_THOLD__14__0_), .C(n19104), .Y(n2260) );
  A2O1A1Ixp33_ASAP7_75t_SL U21610 ( .A1(uart1_r_IRQCNT__1_), .A2(n19002), .B(
        n29342), .C(n29338), .Y(n19291) );
  A2O1A1Ixp33_ASAP7_75t_SL U21611 ( .A1(n19002), .A2(n22433), .B(n32982), .C(
        n19089), .Y(n1711) );
  A2O1A1Ixp33_ASAP7_75t_SL U21612 ( .A1(dataout[15]), .A2(n19002), .B(n19287), 
        .C(n19002), .Y(n19288) );
  A2O1A1Ixp33_ASAP7_75t_SL U21613 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__29_), .A2(n19002), .B(n32565), .C(n19002), .Y(n19284) );
  A2O1A1Ixp33_ASAP7_75t_SL U21614 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[29]), 
        .A2(n19002), .B(n32593), .C(n19002), .Y(n19285) );
  O2A1O1Ixp33_ASAP7_75t_SL U21615 ( .A1(n32559), .A2(n19284), .B(n19002), .C(
        n19285), .Y(it_data[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21616 ( .A1(n32626), .A2(n19002), .B(n32543), .C(
        n19283), .Y(it_data[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21617 ( .A1(n18887), .A2(n32444), .B(n19279), .C(
        n19002), .Y(n19280) );
  A2O1A1Ixp33_ASAP7_75t_SL U21618 ( .A1(n33067), .A2(n19002), .B(n19280), .C(
        n19281), .Y(dc_address[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21619 ( .A1(n32640), .A2(n19002), .B(n32429), .C(
        n19002), .Y(n19271) );
  A2O1A1Ixp33_ASAP7_75t_SL U21620 ( .A1(n32379), .A2(n19002), .B(n32431), .C(
        n19002), .Y(n19272) );
  A2O1A1Ixp33_ASAP7_75t_SL U21621 ( .A1(dc_q[21]), .A2(n32385), .B(n19272), 
        .C(n19002), .Y(n19273) );
  A2O1A1Ixp33_ASAP7_75t_SL U21622 ( .A1(n32380), .A2(n19002), .B(n24543), .C(
        n19273), .Y(n19274) );
  A2O1A1Ixp33_ASAP7_75t_SL U21623 ( .A1(n19271), .A2(n19002), .B(n19274), .C(
        n19002), .Y(n19275) );
  A2O1A1Ixp33_ASAP7_75t_SL U21624 ( .A1(n32381), .A2(n19002), .B(n32408), .C(
        n19275), .Y(dc_data[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21625 ( .A1(n32214), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__17_), .B(n19269), .C(n19002), .Y(
        n19270) );
  A2O1A1Ixp33_ASAP7_75t_SL U21626 ( .A1(n32632), .A2(n19002), .B(n32217), .C(
        n19270), .Y(dt_data[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21627 ( .A1(n32162), .A2(n19002), .B(n33055), .C(
        n19002), .Y(n19264) );
  A2O1A1Ixp33_ASAP7_75t_SL U21628 ( .A1(n17278), .A2(n19002), .B(n19263), .C(
        n19002), .Y(n30801) );
  A2O1A1Ixp33_ASAP7_75t_SL U21629 ( .A1(n25568), .A2(n19002), .B(n19262), .C(
        n19002), .Y(n31876) );
  A2O1A1Ixp33_ASAP7_75t_SL U21630 ( .A1(n30224), .A2(n19002), .B(n22376), .C(
        n19002), .Y(n19261) );
  A2O1A1Ixp33_ASAP7_75t_SL U21631 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__29_), .B(n19261), .C(n19002), .Y(
        n29864) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21632 ( .A1(n28668), .A2(n28132), .B(n28133), 
        .C(n19002), .D(n19260), .Y(n32332) );
  A2O1A1Ixp33_ASAP7_75t_SL U21633 ( .A1(n23941), .A2(n19002), .B(n19243), .C(
        n19002), .Y(n19244) );
  A2O1A1Ixp33_ASAP7_75t_SL U21634 ( .A1(n19245), .A2(n19002), .B(n19246), .C(
        n19002), .Y(n19247) );
  A2O1A1Ixp33_ASAP7_75t_SL U21635 ( .A1(u0_0_leon3x0_p0_ici[59]), .A2(n19002), 
        .B(n19252), .C(n19002), .Y(n19253) );
  O2A1O1Ixp5_ASAP7_75t_SL U21636 ( .A1(n19244), .A2(n19254), .B(n19002), .C(
        n19249), .Y(n19255) );
  A2O1A1Ixp33_ASAP7_75t_SL U21637 ( .A1(n24903), .A2(n19241), .B(n24908), .C(
        n19002), .Y(n24904) );
  A2O1A1Ixp33_ASAP7_75t_SL U21638 ( .A1(n19238), .A2(n19002), .B(
        uart1_uarto_SCALER__11_), .C(n19002), .Y(n19239) );
  A2O1A1Ixp33_ASAP7_75t_SL U21639 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__0_), 
        .A2(n19002), .B(n19233), .C(n19002), .Y(n19234) );
  A2O1A1Ixp33_ASAP7_75t_SL U21640 ( .A1(n31423), .A2(n29731), .B(n19234), .C(
        n19002), .Y(n29476) );
  A2O1A1Ixp33_ASAP7_75t_SL U21641 ( .A1(n22376), .A2(n19002), .B(n30418), .C(
        n19232), .Y(n29680) );
  A2O1A1Ixp33_ASAP7_75t_SL U21642 ( .A1(u0_0_leon3x0_p0_divi[21]), .A2(n19002), 
        .B(n24631), .C(n19002), .Y(n19225) );
  A2O1A1Ixp33_ASAP7_75t_SL U21643 ( .A1(n28830), .A2(u0_0_leon3x0_p0_divi[21]), 
        .B(n28490), .C(n19002), .Y(n19227) );
  A2O1A1Ixp33_ASAP7_75t_SL U21644 ( .A1(n29150), .A2(n19002), .B(n19226), .C(
        n19227), .Y(n19228) );
  A2O1A1Ixp33_ASAP7_75t_SL U21645 ( .A1(u0_0_leon3x0_p0_divi[21]), .A2(n19002), 
        .B(n29148), .C(n19002), .Y(n19229) );
  A2O1A1Ixp33_ASAP7_75t_SL U21646 ( .A1(n22374), .A2(n19002), .B(n28347), .C(
        n19002), .Y(n19222) );
  A2O1A1Ixp33_ASAP7_75t_SL U21647 ( .A1(n18805), .A2(n19002), .B(n32616), .C(
        n19002), .Y(n19223) );
  A2O1A1Ixp33_ASAP7_75t_SL U21648 ( .A1(n22373), .A2(n19002), .B(n27127), .C(
        n19002), .Y(n19224) );
  O2A1O1Ixp5_ASAP7_75t_SL U21649 ( .A1(n19222), .A2(n19223), .B(n19002), .C(
        n19224), .Y(n27172) );
  A2O1A1Ixp33_ASAP7_75t_SL U21650 ( .A1(u0_0_leon3x0_p0_ici[30]), .A2(n19002), 
        .B(DP_OP_1196_128_7433_n452), .C(DP_OP_1196_128_7433_n357), .Y(n19220)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21651 ( .A1(n19219), .A2(n19002), .B(n19220), .C(
        n19002), .Y(n19221) );
  A2O1A1Ixp33_ASAP7_75t_SL U21652 ( .A1(u0_0_leon3x0_p0_ici[60]), .A2(n19218), 
        .B(n19221), .C(n19002), .Y(n32667) );
  A2O1A1Ixp33_ASAP7_75t_SL U21653 ( .A1(n22392), .A2(n19002), .B(n28725), .C(
        n19217), .Y(n28736) );
  A2O1A1Ixp33_ASAP7_75t_SL U21654 ( .A1(n19002), .A2(n28850), .B(n25463), .C(
        n19012), .Y(n19013) );
  A2O1A1Ixp33_ASAP7_75t_SL U21655 ( .A1(n28967), .A2(n26377), .B(n19013), .C(
        n19002), .Y(n19014) );
  A2O1A1Ixp33_ASAP7_75t_SL U21656 ( .A1(n28977), .A2(n19002), .B(n25464), .C(
        n19014), .Y(n26914) );
  A2O1A1Ixp33_ASAP7_75t_SL U21657 ( .A1(n19002), .A2(n22392), .B(n18299), .C(
        n19010), .Y(n26585) );
  A2O1A1Ixp33_ASAP7_75t_SL U21658 ( .A1(n29040), .A2(n19002), .B(n18876), .C(
        n19007), .Y(u0_0_leon3x0_p0_iu_fe_pc_22_) );
  A2O1A1Ixp33_ASAP7_75t_SL U21659 ( .A1(add_x_735_n92), .A2(n19002), .B(n19211), .C(n19002), .Y(add_x_735_n90) );
  A2O1A1Ixp33_ASAP7_75t_SL U21660 ( .A1(n28304), .A2(n19002), .B(n31660), .C(
        n19203), .Y(n19204) );
  A2O1A1Ixp33_ASAP7_75t_SL U21661 ( .A1(n28371), .A2(u0_0_leon3x0_p0_divo[26]), 
        .B(n19204), .C(n19002), .Y(n19205) );
  A2O1A1Ixp33_ASAP7_75t_SL U21662 ( .A1(n24040), .A2(n19002), .B(
        mult_x_1196_n2741), .C(n19002), .Y(n19192) );
  A2O1A1Ixp33_ASAP7_75t_SL U21663 ( .A1(n24041), .A2(n19002), .B(
        mult_x_1196_n2742), .C(n19002), .Y(n19193) );
  A2O1A1Ixp33_ASAP7_75t_SL U21664 ( .A1(n19192), .A2(n19002), .B(n19193), .C(
        n19002), .Y(n19194) );
  A2O1A1Ixp33_ASAP7_75t_SL U21665 ( .A1(n24034), .A2(n19002), .B(
        mult_x_1196_n2806), .C(n19002), .Y(n19198) );
  A2O1A1Ixp33_ASAP7_75t_SL U21666 ( .A1(n22251), .A2(n19002), .B(
        mult_x_1196_n2805), .C(n19002), .Y(n19199) );
  A2O1A1Ixp33_ASAP7_75t_SL U21667 ( .A1(n19194), .A2(n19002), .B(n19197), .C(
        n19200), .Y(n19201) );
  A2O1A1Ixp33_ASAP7_75t_SL U21668 ( .A1(n19002), .A2(n19198), .B(n19199), .C(
        n19002), .Y(n19200) );
  A2O1A1Ixp33_ASAP7_75t_SL U21669 ( .A1(n30805), .A2(n19002), .B(n19169), .C(
        n19170), .Y(n19171) );
  A2O1A1Ixp33_ASAP7_75t_SL U21670 ( .A1(n31248), .A2(irqctrl0_r_ILEVEL__13_), 
        .B(n19171), .C(n19002), .Y(n19172) );
  A2O1A1Ixp33_ASAP7_75t_SL U21671 ( .A1(n32004), .A2(n19002), .B(n30803), .C(
        n19002), .Y(n19177) );
  A2O1A1Ixp33_ASAP7_75t_SL U21672 ( .A1(n32008), .A2(n19176), .B(n19177), .C(
        n19002), .Y(n19178) );
  A2O1A1Ixp33_ASAP7_75t_SL U21673 ( .A1(n31323), .A2(n19002), .B(n30806), .C(
        n19178), .Y(n19179) );
  A2O1A1Ixp33_ASAP7_75t_SL U21674 ( .A1(n19175), .A2(n19002), .B(n19179), .C(
        n19002), .Y(n4662) );
  A2O1A1Ixp33_ASAP7_75t_SL U21675 ( .A1(n29517), .A2(n19002), .B(n19154), .C(
        n19002), .Y(n19155) );
  A2O1A1Ixp33_ASAP7_75t_SL U21676 ( .A1(n29516), .A2(n19002), .B(n28108), .C(
        n24694), .Y(n19156) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21677 ( .A1(n24628), .A2(n29521), .B(n19155), 
        .C(n19002), .D(n19156), .Y(n4369) );
  A2O1A1Ixp33_ASAP7_75t_SL U21678 ( .A1(n31448), .A2(n19002), .B(n19147), .C(
        n19002), .Y(n19148) );
  A2O1A1Ixp33_ASAP7_75t_SL U21679 ( .A1(n32197), .A2(n25014), .B(n31446), .C(
        n19002), .Y(n19149) );
  A2O1A1Ixp33_ASAP7_75t_SL U21680 ( .A1(n19148), .A2(n19002), .B(n19149), .C(
        n19002), .Y(n19150) );
  A2O1A1Ixp33_ASAP7_75t_SL U21681 ( .A1(n32443), .A2(n19002), .B(n19150), .C(
        n19002), .Y(n19151) );
  A2O1A1Ixp33_ASAP7_75t_SL U21682 ( .A1(n31001), .A2(n19002), .B(n31258), .C(
        n19002), .Y(n19152) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21683 ( .A1(n31262), .A2(n25399), .B(n22380), 
        .C(n19002), .D(n25586), .Y(n19153) );
  A2O1A1Ixp33_ASAP7_75t_SL U21684 ( .A1(n24291), .A2(mult_x_1196_n747), .B(
        mult_x_1196_n744), .C(n19002), .Y(n19142) );
  A2O1A1Ixp33_ASAP7_75t_SL U21685 ( .A1(n22427), .A2(n19002), .B(n19145), .C(
        n19146), .Y(n4293) );
  A2O1A1Ixp33_ASAP7_75t_SL U21686 ( .A1(n22428), .A2(n19002), .B(n29767), .C(
        n19141), .Y(n4125) );
  A2O1A1Ixp33_ASAP7_75t_SL U21687 ( .A1(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__31_), .A2(n19002), .B(n24654), .C(
        n19140), .Y(n4061) );
  A2O1A1Ixp33_ASAP7_75t_SL U21688 ( .A1(n24646), .A2(n19002), .B(n30473), .C(
        n19136), .Y(n3953) );
  A2O1A1Ixp33_ASAP7_75t_SL U21689 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_), .A2(n19002), .B(n24656), .C(
        n19134), .Y(n3747) );
  A2O1A1Ixp33_ASAP7_75t_SL U21690 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__8_), .A2(n19002), .B(n24495), .C(n19002), .Y(n19130) );
  A2O1A1Ixp33_ASAP7_75t_SL U21691 ( .A1(n23229), .A2(n19002), .B(
        u0_0_leon3x0_p0_iu_r_A__IMM__18_), .C(n19002), .Y(n19131) );
  A2O1A1Ixp33_ASAP7_75t_SL U21692 ( .A1(n24646), .A2(n19002), .B(n19126), .C(
        n19002), .Y(n19127) );
  A2O1A1Ixp33_ASAP7_75t_SL U21693 ( .A1(u0_0_leon3x0_p0_ici[53]), .A2(n19002), 
        .B(n24652), .C(n19125), .Y(n3406) );
  A2O1A1Ixp33_ASAP7_75t_SL U21694 ( .A1(u0_0_leon3x0_p0_ici[31]), .A2(n19002), 
        .B(n24651), .C(n19119), .Y(n3186) );
  A2O1A1Ixp33_ASAP7_75t_SL U21695 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__10_), 
        .A2(n19002), .B(n24653), .C(n19117), .Y(n3172) );
  A2O1A1Ixp33_ASAP7_75t_SL U21696 ( .A1(n31573), .A2(n19002), .B(n22396), .C(
        n19002), .Y(n19114) );
  A2O1A1Ixp33_ASAP7_75t_SL U21697 ( .A1(n31840), .A2(n19002), .B(apbi[17]), 
        .C(n19112), .Y(n2835) );
  A2O1A1Ixp33_ASAP7_75t_SL U21698 ( .A1(n31114), .A2(n19002), .B(n26126), .C(
        n19002), .Y(n19110) );
  A2O1A1Ixp33_ASAP7_75t_SL U21699 ( .A1(n31115), .A2(n19002), .B(n26127), .C(
        n19002), .Y(n19111) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21700 ( .A1(n31117), .A2(uart1_r_RHOLD__15__1_), 
        .B(n19110), .C(n19002), .D(n19111), .Y(n2451) );
  A2O1A1Ixp33_ASAP7_75t_SL U21701 ( .A1(n32040), .A2(n19002), .B(n31743), .C(
        n19002), .Y(n19109) );
  A2O1A1Ixp33_ASAP7_75t_SL U21702 ( .A1(sr1_r_SRHSEL_), .A2(n4722), .B(n19109), 
        .C(n19002), .Y(n2358) );
  A2O1A1Ixp33_ASAP7_75t_SL U21703 ( .A1(n32493), .A2(n19002), .B(n32512), .C(
        n19002), .Y(n19107) );
  A2O1A1Ixp33_ASAP7_75t_SL U21704 ( .A1(n32492), .A2(it_q[4]), .B(n19108), .C(
        n19002), .Y(n2288) );
  A2O1A1Ixp33_ASAP7_75t_SL U21705 ( .A1(uart1_r_TRADDR__3_), .A2(n27315), .B(
        n19103), .C(n19002), .Y(n2241) );
  A2O1A1Ixp33_ASAP7_75t_SL U21706 ( .A1(n32705), .A2(n19002), .B(n25412), .C(
        n19002), .Y(n19099) );
  A2O1A1Ixp33_ASAP7_75t_SL U21707 ( .A1(n22393), .A2(n19002), .B(n32998), .C(
        n19002), .Y(n19100) );
  A2O1A1Ixp33_ASAP7_75t_SL U21708 ( .A1(n19099), .A2(n19002), .B(n19100), .C(
        n19002), .Y(n1791) );
  A2O1A1Ixp33_ASAP7_75t_SL U21709 ( .A1(n31725), .A2(sr1_r_MCFG1__ROMWWS__2_), 
        .B(n19093), .C(n19002), .Y(n19094) );
  A2O1A1Ixp33_ASAP7_75t_SL U21710 ( .A1(dataout[7]), .A2(n19002), .B(n19087), 
        .C(n19002), .Y(n19088) );
  A2O1A1Ixp33_ASAP7_75t_SL U21711 ( .A1(n27279), .A2(n19002), .B(n30642), .C(
        n19002), .Y(n19078) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21712 ( .A1(n30644), .A2(n27275), .B(n19078), 
        .C(n19002), .D(n19081), .Y(n19082) );
  A2O1A1Ixp33_ASAP7_75t_SL U21713 ( .A1(n30645), .A2(n19002), .B(n27267), .C(
        n19082), .Y(n19083) );
  A2O1A1Ixp33_ASAP7_75t_SL U21714 ( .A1(n27263), .A2(n22432), .B(n19083), .C(
        n19002), .Y(n19084) );
  A2O1A1Ixp33_ASAP7_75t_SL U21715 ( .A1(n27257), .A2(n19002), .B(n22379), .C(
        n19002), .Y(n19086) );
  A2O1A1Ixp33_ASAP7_75t_SL U21716 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__27_), .A2(n19002), .B(n32565), .C(n19002), .Y(n19074) );
  A2O1A1Ixp33_ASAP7_75t_SL U21717 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[27]), 
        .A2(n19002), .B(n32593), .C(n19002), .Y(n19075) );
  O2A1O1Ixp33_ASAP7_75t_SL U21718 ( .A1(n32559), .A2(n19074), .B(n19002), .C(
        n19075), .Y(it_data[23]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21719 ( .A1(n32624), .A2(n19002), .B(n32543), .C(
        n19073), .Y(it_data[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21720 ( .A1(n32214), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__16_), .B(n19066), .C(n19002), .Y(
        n19067) );
  A2O1A1Ixp33_ASAP7_75t_SL U21721 ( .A1(n32630), .A2(n19002), .B(n32217), .C(
        n19067), .Y(dt_data[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21722 ( .A1(n29613), .A2(n19002), .B(n26522), .C(
        n19002), .Y(n19061) );
  A2O1A1Ixp33_ASAP7_75t_SL U21723 ( .A1(n18593), .A2(n19002), .B(n26329), .C(
        n19002), .Y(n19062) );
  A2O1A1Ixp33_ASAP7_75t_SL U21724 ( .A1(n25645), .A2(n19002), .B(n22375), .C(
        n19002), .Y(n19063) );
  A2O1A1Ixp33_ASAP7_75t_SL U21725 ( .A1(n19056), .A2(n19002), .B(n19057), .C(
        n19002), .Y(n19058) );
  A2O1A1Ixp33_ASAP7_75t_SL U21726 ( .A1(n28031), .A2(n19002), .B(n19059), .C(
        n19002), .Y(n19060) );
  A2O1A1Ixp33_ASAP7_75t_SL U21727 ( .A1(n31657), .A2(n19002), .B(n19052), .C(
        n19002), .Y(n19053) );
  A2O1A1Ixp33_ASAP7_75t_SL U21728 ( .A1(n22380), .A2(n19002), .B(n19053), .C(
        n19002), .Y(n24908) );
  A2O1A1Ixp33_ASAP7_75t_SL U21729 ( .A1(u0_0_leon3x0_p0_iu_de_icc_3_), .A2(
        n19002), .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_), .C(n19002), .Y(
        n19037) );
  A2O1A1Ixp33_ASAP7_75t_SL U21730 ( .A1(u0_0_leon3x0_p0_iu_de_icc_1_), .A2(
        n19002), .B(n30907), .C(n19002), .Y(n19038) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21731 ( .A1(u0_0_leon3x0_p0_iu_de_icc_2_), .A2(
        n30907), .B(u0_0_leon3x0_p0_iu_de_icc_0_), .C(n19002), .D(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_), .Y(n19039) );
  A2O1A1Ixp33_ASAP7_75t_SL U21732 ( .A1(n19040), .A2(n19002), .B(n19041), .C(
        n19002), .Y(n19042) );
  A2O1A1Ixp33_ASAP7_75t_SL U21733 ( .A1(n24873), .A2(n19002), .B(n30906), .C(
        n29173), .Y(n19043) );
  A2O1A1Ixp33_ASAP7_75t_SL U21734 ( .A1(n19037), .A2(n19002), .B(n19038), .C(
        n19002), .Y(n19046) );
  A2O1A1Ixp33_ASAP7_75t_SL U21735 ( .A1(n19046), .A2(n19002), .B(n19047), .C(
        n19002), .Y(n19048) );
  A2O1A1Ixp33_ASAP7_75t_SL U21736 ( .A1(n19039), .A2(n19002), .B(n19048), .C(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__27_), .Y(n19049) );
  A2O1A1Ixp33_ASAP7_75t_SL U21737 ( .A1(n19050), .A2(n19002), .B(n19045), .C(
        n19002), .Y(n19051) );
  A2O1A1Ixp33_ASAP7_75t_SL U21738 ( .A1(n23941), .A2(n19002), .B(n19029), .C(
        n19002), .Y(n19030) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21739 ( .A1(DP_OP_1196_128_7433_n234), .A2(
        DP_OP_1196_128_7433_n4), .B(n19030), .C(n19002), .D(
        DP_OP_1196_128_7433_n235), .Y(n19031) );
  A2O1A1Ixp33_ASAP7_75t_SL U21740 ( .A1(n24541), .A2(n19002), .B(n32119), .C(
        n19002), .Y(n19022) );
  A2O1A1Ixp33_ASAP7_75t_SL U21741 ( .A1(n29012), .A2(n30644), .B(n19025), .C(
        n19002), .Y(n19026) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21742 ( .A1(n31868), .A2(n31424), .B(n19022), 
        .C(n19002), .D(n19028), .Y(n29013) );
  A2O1A1Ixp33_ASAP7_75t_SL U21743 ( .A1(n32874), .A2(n19002), .B(n19020), .C(
        n19021), .Y(n32911) );
  A2O1A1Ixp33_ASAP7_75t_SL U21744 ( .A1(DP_OP_1196_128_7433_n168), .A2(n19002), 
        .B(n19008), .C(DP_OP_1196_128_7433_n161), .Y(n19009) );
  A2O1A1Ixp33_ASAP7_75t_SL U21745 ( .A1(n32142), .A2(n19002), .B(n32290), .C(
        n19002), .Y(n19003) );
  A2O1A1Ixp33_ASAP7_75t_SL U21746 ( .A1(n32290), .A2(u0_0_leon3x0_p0_dci[5]), 
        .B(n19003), .C(n19002), .Y(n32349) );
  O2A1O1Ixp33_ASAP7_75t_SL U21747 ( .A1(n19199), .A2(n19198), .B(n19002), .C(
        n19000), .Y(n19001) );
  A2O1A1Ixp33_ASAP7_75t_SL U21748 ( .A1(n21482), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n21483) );
  A2O1A1Ixp33_ASAP7_75t_SL U21749 ( .A1(n21504), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n21505) );
  O2A1O1Ixp33_ASAP7_75t_SL U21750 ( .A1(n31238), .A2(n21518), .B(n21519), .C(
        n18295), .Y(n21520) );
  A2O1A1Ixp33_ASAP7_75t_SL U21751 ( .A1(n20571), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n20572) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U21752 ( .A1(n32661), .A2(n32429), .B(n20576), 
        .C(n18295), .Y(n20577) );
  O2A1O1Ixp33_ASAP7_75t_SL U21753 ( .A1(n23941), .A2(n19447), .B(n19448), .C(
        n18295), .Y(n19449) );
  A2O1A1Ixp33_ASAP7_75t_SL U21754 ( .A1(n24622), .A2(n24621), .B(n18295), .C(
        n19002), .Y(n22198) );
  A2O1A1Ixp33_ASAP7_75t_SL U21755 ( .A1(timer0_r_SCALER__7_), .A2(n22198), .B(
        n18295), .C(n19002), .Y(n22199) );
  A2O1A1Ixp33_ASAP7_75t_SL U21756 ( .A1(n24622), .A2(n24621), .B(n18295), .C(
        n22200), .Y(n22201) );
  A2O1A1Ixp33_ASAP7_75t_SL U21757 ( .A1(n22199), .A2(n22201), .B(n18295), .C(
        n19002), .Y(n22202) );
  A2O1A1Ixp33_ASAP7_75t_SL U21758 ( .A1(n18845), .A2(n29884), .B(n18295), .C(
        n30687), .Y(n22192) );
  A2O1A1Ixp33_ASAP7_75t_SL U21759 ( .A1(n29881), .A2(n29882), .B(n18295), .C(
        n19002), .Y(n22195) );
  A2O1A1Ixp33_ASAP7_75t_SL U21760 ( .A1(n24648), .A2(
        u0_0_leon3x0_p0_iu_r_X__CTRL__TT__3_), .B(n18295), .C(n19002), .Y(
        n22196) );
  A2O1A1Ixp33_ASAP7_75t_SL U21761 ( .A1(n29885), .A2(n22195), .B(n18295), .C(
        n22196), .Y(n22197) );
  A2O1A1Ixp33_ASAP7_75t_SL U21762 ( .A1(n24665), .A2(n32574), .B(n18295), .C(
        n19002), .Y(n22190) );
  A2O1A1Ixp33_ASAP7_75t_SL U21763 ( .A1(n31639), .A2(n24694), .B(n18295), .C(
        n21968), .Y(n17243) );
  A2O1A1Ixp33_ASAP7_75t_SL U21764 ( .A1(n18295), .A2(n19002), .B(n21729), .C(
        n19002), .Y(n21730) );
  A2O1A1Ixp33_ASAP7_75t_SL U21765 ( .A1(n21963), .A2(n21964), .B(n18295), .C(
        n19002), .Y(n21965) );
  A2O1A1Ixp33_ASAP7_75t_SL U21766 ( .A1(n30640), .A2(rf_do_b[14]), .B(n18295), 
        .C(n19002), .Y(n22173) );
  A2O1A1Ixp33_ASAP7_75t_SL U21767 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__14_), .B(n18295), .C(n19002), .Y(n22174)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21768 ( .A1(n22173), .A2(n22174), .B(n18295), .C(
        n19002), .Y(n22175) );
  A2O1A1Ixp33_ASAP7_75t_SL U21769 ( .A1(n31542), .A2(n30491), .B(n18295), .C(
        n19002), .Y(n22163) );
  A2O1A1Ixp33_ASAP7_75t_SL U21770 ( .A1(n27242), .A2(n31054), .B(n18295), .C(
        n19002), .Y(n22164) );
  A2O1A1Ixp33_ASAP7_75t_SL U21771 ( .A1(n22163), .A2(n22164), .B(n18295), .C(
        n19002), .Y(n22165) );
  A2O1A1Ixp33_ASAP7_75t_SL U21772 ( .A1(n27240), .A2(n32114), .B(n18295), .C(
        n19002), .Y(n22166) );
  A2O1A1Ixp33_ASAP7_75t_SL U21773 ( .A1(n27241), .A2(n30492), .B(n18295), .C(
        n19002), .Y(n22167) );
  A2O1A1Ixp33_ASAP7_75t_SL U21774 ( .A1(n22166), .A2(n22167), .B(n18295), .C(
        n19002), .Y(n22168) );
  A2O1A1Ixp33_ASAP7_75t_SL U21775 ( .A1(n22165), .A2(n22168), .B(n18295), .C(
        n19002), .Y(n22169) );
  A2O1A1Ixp33_ASAP7_75t_SL U21776 ( .A1(n22427), .A2(n27243), .B(n18295), .C(
        n19002), .Y(n22170) );
  A2O1A1Ixp33_ASAP7_75t_SL U21777 ( .A1(n22169), .A2(n22170), .B(n18295), .C(
        n19002), .Y(n4639) );
  A2O1A1Ixp33_ASAP7_75t_SL U21778 ( .A1(n18295), .A2(n19002), .B(n21957), .C(
        n19002), .Y(n24509) );
  A2O1A1Ixp33_ASAP7_75t_SL U21779 ( .A1(n30248), .A2(n24678), .B(n18295), .C(
        n19002), .Y(n20832) );
  A2O1A1Ixp33_ASAP7_75t_SL U21780 ( .A1(u0_0_leon3x0_p0_divi[60]), .A2(n30430), 
        .B(n18295), .C(n19002), .Y(n22157) );
  A2O1A1Ixp33_ASAP7_75t_SL U21781 ( .A1(n22156), .A2(n22157), .B(n18295), .C(
        n19002), .Y(n22158) );
  A2O1A1Ixp33_ASAP7_75t_SL U21782 ( .A1(n29696), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), .B(n18295), .C(n19002), .Y(
        n22151) );
  A2O1A1Ixp33_ASAP7_75t_SL U21783 ( .A1(n29697), .A2(n29698), .B(n18295), .C(
        n19002), .Y(n22152) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U21784 ( .A1(n29874), .A2(n22151), .B(n18295), 
        .C(n22152), .D(n29875), .Y(n22153) );
  A2O1A1Ixp33_ASAP7_75t_SL U21785 ( .A1(n32618), .A2(n24663), .B(n18295), .C(
        n19002), .Y(n21441) );
  A2O1A1Ixp33_ASAP7_75t_SL U21786 ( .A1(n18295), .A2(n19002), .B(n20673), .C(
        n19002), .Y(n20674) );
  A2O1A1Ixp33_ASAP7_75t_SL U21787 ( .A1(n24668), .A2(n22147), .B(n18295), .C(
        n19002), .Y(n22148) );
  A2O1A1Ixp33_ASAP7_75t_SL U21788 ( .A1(n18295), .A2(n19002), .B(n21936), .C(
        n19002), .Y(n21937) );
  A2O1A1Ixp33_ASAP7_75t_SL U21789 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[32]), 
        .B(n18295), .C(n19002), .Y(n22145) );
  A2O1A1Ixp33_ASAP7_75t_SL U21790 ( .A1(n22144), .A2(n22145), .B(n18295), .C(
        n19002), .Y(n22146) );
  A2O1A1Ixp33_ASAP7_75t_SL U21791 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[39]), 
        .B(n18295), .C(n19002), .Y(n22141) );
  A2O1A1Ixp33_ASAP7_75t_SL U21792 ( .A1(n22140), .A2(n22141), .B(n18295), .C(
        n19002), .Y(n22142) );
  A2O1A1Ixp33_ASAP7_75t_SL U21793 ( .A1(n22396), .A2(n22137), .B(n18295), .C(
        n19002), .Y(n22138) );
  A2O1A1Ixp33_ASAP7_75t_SL U21794 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), 
        .A2(n31818), .B(n18295), .C(n19002), .Y(n22135) );
  A2O1A1Ixp33_ASAP7_75t_SL U21795 ( .A1(n26953), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n22134) );
  A2O1A1Ixp33_ASAP7_75t_SL U21796 ( .A1(n18295), .A2(n19002), .B(n21695), .C(
        n19002), .Y(n21696) );
  A2O1A1Ixp33_ASAP7_75t_SL U21797 ( .A1(n21696), .A2(n21697), .B(n18295), .C(
        n19002), .Y(n4374) );
  A2O1A1Ixp33_ASAP7_75t_SL U21798 ( .A1(n28522), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n21924) );
  A2O1A1Ixp33_ASAP7_75t_SL U21799 ( .A1(n30592), .A2(n24681), .B(n18295), .C(
        n19002), .Y(n22131) );
  A2O1A1Ixp33_ASAP7_75t_SL U21800 ( .A1(n29107), .A2(n24675), .B(n18295), .C(
        n19002), .Y(n21678) );
  A2O1A1Ixp33_ASAP7_75t_SL U21801 ( .A1(n24673), .A2(n25279), .B(n18295), .C(
        n19002), .Y(n22130) );
  A2O1A1Ixp33_ASAP7_75t_SL U21802 ( .A1(n24673), .A2(n25286), .B(n18295), .C(
        n19002), .Y(n22128) );
  A2O1A1Ixp33_ASAP7_75t_SL U21803 ( .A1(n24660), .A2(n21916), .B(n18295), .C(
        n19002), .Y(n21917) );
  A2O1A1Ixp33_ASAP7_75t_SL U21804 ( .A1(n24920), .A2(n24675), .B(n18295), .C(
        n19002), .Y(n21913) );
  A2O1A1Ixp33_ASAP7_75t_SL U21805 ( .A1(n32130), .A2(n24661), .B(n18295), .C(
        n19002), .Y(n21001) );
  A2O1A1Ixp33_ASAP7_75t_SL U21806 ( .A1(n22378), .A2(n32616), .B(n18295), .C(
        n19002), .Y(n22127) );
  A2O1A1Ixp33_ASAP7_75t_SL U21807 ( .A1(n24663), .A2(n32620), .B(n18295), .C(
        n19002), .Y(n22126) );
  A2O1A1Ixp33_ASAP7_75t_SL U21808 ( .A1(n23229), .A2(n29845), .B(n18295), .C(
        n19002), .Y(n21912) );
  A2O1A1Ixp33_ASAP7_75t_SL U21809 ( .A1(n29212), .A2(n24671), .B(n18295), .C(
        n19002), .Y(n21410) );
  A2O1A1Ixp33_ASAP7_75t_SL U21810 ( .A1(n24659), .A2(n21184), .B(n18295), .C(
        n19002), .Y(n21185) );
  A2O1A1Ixp33_ASAP7_75t_SL U21811 ( .A1(n24681), .A2(n29808), .B(n18295), .C(
        n19002), .Y(n21911) );
  A2O1A1Ixp33_ASAP7_75t_SL U21812 ( .A1(n25005), .A2(n24674), .B(n18295), .C(
        n19002), .Y(n20640) );
  A2O1A1Ixp33_ASAP7_75t_SL U21813 ( .A1(n24681), .A2(n30821), .B(n18295), .C(
        n19002), .Y(n21910) );
  A2O1A1Ixp33_ASAP7_75t_SL U21814 ( .A1(n24661), .A2(n29576), .B(n18295), .C(
        n19002), .Y(n22125) );
  A2O1A1Ixp33_ASAP7_75t_SL U21815 ( .A1(n31823), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n22124) );
  A2O1A1Ixp33_ASAP7_75t_SL U21816 ( .A1(n32606), .A2(n24661), .B(n18295), .C(
        n19002), .Y(n19880) );
  A2O1A1Ixp33_ASAP7_75t_SL U21817 ( .A1(n31018), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21904) );
  A2O1A1Ixp33_ASAP7_75t_SL U21818 ( .A1(n24681), .A2(n29693), .B(n18295), .C(
        n19002), .Y(n21170) );
  A2O1A1Ixp33_ASAP7_75t_SL U21819 ( .A1(n32562), .A2(n22122), .B(n18295), .C(
        n19002), .Y(n22123) );
  A2O1A1Ixp33_ASAP7_75t_SL U21820 ( .A1(n24674), .A2(n31962), .B(n18295), .C(
        n19002), .Y(n22121) );
  A2O1A1Ixp33_ASAP7_75t_SL U21821 ( .A1(n24681), .A2(n29907), .B(n18295), .C(
        n19002), .Y(n21169) );
  A2O1A1Ixp33_ASAP7_75t_SL U21822 ( .A1(n24681), .A2(n29795), .B(n18295), .C(
        n19002), .Y(n20638) );
  A2O1A1Ixp33_ASAP7_75t_SL U21823 ( .A1(n30224), .A2(n24676), .B(n18295), .C(
        n19002), .Y(n21900) );
  A2O1A1Ixp33_ASAP7_75t_SL U21824 ( .A1(n30610), .A2(n24662), .B(n18295), .C(
        n19002), .Y(n21899) );
  A2O1A1Ixp33_ASAP7_75t_SL U21825 ( .A1(n30458), .A2(n24673), .B(n18295), .C(
        n19002), .Y(n21897) );
  A2O1A1Ixp33_ASAP7_75t_SL U21826 ( .A1(n24681), .A2(n30412), .B(n18295), .C(
        n19002), .Y(n21398) );
  A2O1A1Ixp33_ASAP7_75t_SL U21827 ( .A1(n24681), .A2(n30391), .B(n18295), .C(
        n19002), .Y(n21653) );
  A2O1A1Ixp33_ASAP7_75t_SL U21828 ( .A1(n30382), .A2(n24673), .B(n18295), .C(
        n19002), .Y(n20986) );
  A2O1A1Ixp33_ASAP7_75t_SL U21829 ( .A1(n24681), .A2(n30376), .B(n18295), .C(
        n19002), .Y(n21896) );
  A2O1A1Ixp33_ASAP7_75t_SL U21830 ( .A1(n24681), .A2(n30366), .B(n18295), .C(
        n19002), .Y(n21895) );
  A2O1A1Ixp33_ASAP7_75t_SL U21831 ( .A1(n30350), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21652) );
  A2O1A1Ixp33_ASAP7_75t_SL U21832 ( .A1(n30338), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21396) );
  A2O1A1Ixp33_ASAP7_75t_SL U21833 ( .A1(n30327), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21651) );
  A2O1A1Ixp33_ASAP7_75t_SL U21834 ( .A1(n30320), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21894) );
  A2O1A1Ixp33_ASAP7_75t_SL U21835 ( .A1(n24681), .A2(n30291), .B(n18295), .C(
        n19002), .Y(n21893) );
  A2O1A1Ixp33_ASAP7_75t_SL U21836 ( .A1(n24670), .A2(n20455), .B(n18295), .C(
        n19002), .Y(n20456) );
  A2O1A1Ixp33_ASAP7_75t_SL U21837 ( .A1(n24664), .A2(n21882), .B(n18295), .C(
        n19002), .Y(n21883) );
  A2O1A1Ixp33_ASAP7_75t_SL U21838 ( .A1(n24663), .A2(n21880), .B(n18295), .C(
        n19002), .Y(n21881) );
  A2O1A1Ixp33_ASAP7_75t_SL U21839 ( .A1(n24665), .A2(n21878), .B(n18295), .C(
        n19002), .Y(n21879) );
  A2O1A1Ixp33_ASAP7_75t_SL U21840 ( .A1(n24668), .A2(n30927), .B(n18295), .C(
        n19002), .Y(n22119) );
  A2O1A1Ixp33_ASAP7_75t_SL U21841 ( .A1(n24674), .A2(n25152), .B(n18295), .C(
        n19002), .Y(n22118) );
  A2O1A1Ixp33_ASAP7_75t_SL U21842 ( .A1(n29481), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21381) );
  A2O1A1Ixp33_ASAP7_75t_SL U21843 ( .A1(n24665), .A2(n19705), .B(n18295), .C(
        n19002), .Y(n19706) );
  A2O1A1Ixp33_ASAP7_75t_SL U21844 ( .A1(n32577), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n20976) );
  A2O1A1Ixp33_ASAP7_75t_SL U21845 ( .A1(n32580), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21877) );
  A2O1A1Ixp33_ASAP7_75t_SL U21846 ( .A1(n30974), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21876) );
  A2O1A1Ixp33_ASAP7_75t_SL U21847 ( .A1(n29036), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21875) );
  A2O1A1Ixp33_ASAP7_75t_SL U21848 ( .A1(n31786), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21874) );
  A2O1A1Ixp33_ASAP7_75t_SL U21849 ( .A1(n30643), .A2(n24662), .B(n18295), .C(
        n19002), .Y(n21873) );
  A2O1A1Ixp33_ASAP7_75t_SL U21850 ( .A1(n24667), .A2(n20970), .B(n18295), .C(
        n19002), .Y(n20971) );
  A2O1A1Ixp33_ASAP7_75t_SL U21851 ( .A1(n24662), .A2(n21640), .B(n18295), .C(
        n19002), .Y(n21641) );
  A2O1A1Ixp33_ASAP7_75t_SL U21852 ( .A1(n31690), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21374) );
  A2O1A1Ixp33_ASAP7_75t_SL U21853 ( .A1(n22427), .A2(n20073), .B(n18295), .C(
        n19002), .Y(n20074) );
  A2O1A1Ixp33_ASAP7_75t_SL U21854 ( .A1(n29066), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21871) );
  A2O1A1Ixp33_ASAP7_75t_SL U21855 ( .A1(n31765), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21870) );
  A2O1A1Ixp33_ASAP7_75t_SL U21856 ( .A1(n30517), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21869) );
  A2O1A1Ixp33_ASAP7_75t_SL U21857 ( .A1(n30506), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21868) );
  A2O1A1Ixp33_ASAP7_75t_SL U21858 ( .A1(n32669), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21867) );
  A2O1A1Ixp33_ASAP7_75t_SL U21859 ( .A1(n24678), .A2(n22116), .B(n18295), .C(
        n19002), .Y(n22117) );
  A2O1A1Ixp33_ASAP7_75t_SL U21860 ( .A1(n28713), .A2(n24676), .B(n18295), .C(
        n19002), .Y(n21144) );
  A2O1A1Ixp33_ASAP7_75t_SL U21861 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__10_), .A2(
        n20308), .B(n18295), .C(n19002), .Y(n20309) );
  A2O1A1Ixp33_ASAP7_75t_SL U21862 ( .A1(n22396), .A2(n22114), .B(n18295), .C(
        n19002), .Y(n22115) );
  A2O1A1Ixp33_ASAP7_75t_SL U21863 ( .A1(n22396), .A2(n22112), .B(n18295), .C(
        n19002), .Y(n22113) );
  A2O1A1Ixp33_ASAP7_75t_SL U21864 ( .A1(n22396), .A2(n22110), .B(n18295), .C(
        n19002), .Y(n22111) );
  A2O1A1Ixp33_ASAP7_75t_SL U21865 ( .A1(n22396), .A2(n22108), .B(n18295), .C(
        n19002), .Y(n22109) );
  A2O1A1Ixp33_ASAP7_75t_SL U21866 ( .A1(n22396), .A2(n22106), .B(n18295), .C(
        n19002), .Y(n22107) );
  A2O1A1Ixp33_ASAP7_75t_SL U21867 ( .A1(n32219), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n21630) );
  A2O1A1Ixp33_ASAP7_75t_SL U21868 ( .A1(n32216), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n21860) );
  A2O1A1Ixp33_ASAP7_75t_SL U21869 ( .A1(n22396), .A2(n22104), .B(n18295), .C(
        n19002), .Y(n22105) );
  A2O1A1Ixp33_ASAP7_75t_SL U21870 ( .A1(n32213), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n21859) );
  A2O1A1Ixp33_ASAP7_75t_SL U21871 ( .A1(n22396), .A2(n22102), .B(n18295), .C(
        n19002), .Y(n22103) );
  A2O1A1Ixp33_ASAP7_75t_SL U21872 ( .A1(n22396), .A2(n22100), .B(n18295), .C(
        n19002), .Y(n22101) );
  A2O1A1Ixp33_ASAP7_75t_SL U21873 ( .A1(n22396), .A2(n22098), .B(n18295), .C(
        n19002), .Y(n22099) );
  A2O1A1Ixp33_ASAP7_75t_SL U21874 ( .A1(n32145), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n21852) );
  A2O1A1Ixp33_ASAP7_75t_SL U21875 ( .A1(n32148), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n21851) );
  A2O1A1Ixp33_ASAP7_75t_SL U21876 ( .A1(n32598), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n21359) );
  A2O1A1Ixp33_ASAP7_75t_SL U21877 ( .A1(n30169), .A2(n22094), .B(n18295), .C(
        n19002), .Y(n22095) );
  A2O1A1Ixp33_ASAP7_75t_SL U21878 ( .A1(n22095), .A2(n22097), .B(n18295), .C(
        n19002), .Y(n3050) );
  A2O1A1Ixp33_ASAP7_75t_SL U21879 ( .A1(n31501), .A2(n22088), .B(n18295), .C(
        n19002), .Y(n22089) );
  A2O1A1Ixp33_ASAP7_75t_SL U21880 ( .A1(n24603), .A2(n24602), .B(n18295), .C(
        n24594), .Y(n20778) );
  A2O1A1Ixp33_ASAP7_75t_SL U21881 ( .A1(n18295), .A2(n19002), .B(n21618), .C(
        n19002), .Y(n2863) );
  A2O1A1Ixp33_ASAP7_75t_SL U21882 ( .A1(n29383), .A2(n22084), .B(n18295), .C(
        n19002), .Y(n22085) );
  A2O1A1Ixp33_ASAP7_75t_SL U21883 ( .A1(n24661), .A2(n22082), .B(n18295), .C(
        n19002), .Y(n22083) );
  A2O1A1Ixp33_ASAP7_75t_SL U21884 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA2__4_), 
        .A2(n24661), .B(n18295), .C(n19002), .Y(n21833) );
  A2O1A1Ixp33_ASAP7_75t_SL U21885 ( .A1(n24681), .A2(n30445), .B(n18295), .C(
        n19002), .Y(n21831) );
  A2O1A1Ixp33_ASAP7_75t_SL U21886 ( .A1(n30487), .A2(n24663), .B(n18295), .C(
        n19002), .Y(n20769) );
  A2O1A1Ixp33_ASAP7_75t_SL U21887 ( .A1(n30489), .A2(n30488), .B(n18295), .C(
        n19002), .Y(n20770) );
  A2O1A1Ixp33_ASAP7_75t_SL U21888 ( .A1(n24666), .A2(n22078), .B(n18295), .C(
        n19002), .Y(n22079) );
  A2O1A1Ixp33_ASAP7_75t_SL U21889 ( .A1(n24677), .A2(n21825), .B(n18295), .C(
        n19002), .Y(n21826) );
  A2O1A1Ixp33_ASAP7_75t_SL U21890 ( .A1(n30540), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21822) );
  A2O1A1Ixp33_ASAP7_75t_SL U21891 ( .A1(n30828), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21818) );
  A2O1A1Ixp33_ASAP7_75t_SL U21892 ( .A1(n27009), .A2(n24671), .B(n18295), .C(
        n19002), .Y(n21817) );
  A2O1A1Ixp33_ASAP7_75t_SL U21893 ( .A1(n30270), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21816) );
  A2O1A1Ixp33_ASAP7_75t_SL U21894 ( .A1(n24678), .A2(n21814), .B(n18295), .C(
        n19002), .Y(n21815) );
  A2O1A1Ixp33_ASAP7_75t_SL U21895 ( .A1(n30251), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21813) );
  A2O1A1Ixp33_ASAP7_75t_SL U21896 ( .A1(n24676), .A2(n21811), .B(n18295), .C(
        n19002), .Y(n21812) );
  A2O1A1Ixp33_ASAP7_75t_SL U21897 ( .A1(n30590), .A2(n24663), .B(n18295), .C(
        n19002), .Y(n21810) );
  A2O1A1Ixp33_ASAP7_75t_SL U21898 ( .A1(n28108), .A2(n27947), .B(n18295), .C(
        n19002), .Y(n21805) );
  A2O1A1Ixp33_ASAP7_75t_SL U21899 ( .A1(n29383), .A2(n22070), .B(n18295), .C(
        n19002), .Y(n22071) );
  A2O1A1Ixp33_ASAP7_75t_SL U21900 ( .A1(n29350), .A2(n19685), .B(n18295), .C(
        n19002), .Y(n1764) );
  A2O1A1Ixp33_ASAP7_75t_SL U21901 ( .A1(n18295), .A2(n19002), .B(n21803), .C(
        n19002), .Y(n21804) );
  A2O1A1Ixp33_ASAP7_75t_SL U21902 ( .A1(n18295), .A2(n19002), .B(n21800), .C(
        n19002), .Y(n21801) );
  A2O1A1Ixp33_ASAP7_75t_SL U21903 ( .A1(n32660), .A2(n32653), .B(n18295), .C(
        n19002), .Y(n22069) );
  A2O1A1Ixp33_ASAP7_75t_SL U21904 ( .A1(n32660), .A2(n32629), .B(n18295), .C(
        n19002), .Y(n22068) );
  A2O1A1Ixp33_ASAP7_75t_SL U21905 ( .A1(n32660), .A2(n32623), .B(n18295), .C(
        n19002), .Y(n22067) );
  A2O1A1Ixp33_ASAP7_75t_SL U21906 ( .A1(n32603), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n21785) );
  A2O1A1Ixp33_ASAP7_75t_SL U21907 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__15_), .A2(n22065), .B(n18295), .C(n19002), .Y(n22066) );
  A2O1A1Ixp33_ASAP7_75t_SL U21908 ( .A1(n32433), .A2(n22061), .B(n18295), .C(
        n19002), .Y(n22062) );
  A2O1A1Ixp33_ASAP7_75t_SL U21909 ( .A1(n32611), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n22063) );
  A2O1A1Ixp33_ASAP7_75t_SL U21910 ( .A1(n32318), .A2(dc_q[7]), .B(n18295), .C(
        n19002), .Y(n22064) );
  A2O1A1Ixp33_ASAP7_75t_SL U21911 ( .A1(n22062), .A2(n22063), .B(n18295), .C(
        n22064), .Y(dc_data[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U21912 ( .A1(n32162), .A2(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__5_), .B(n18295), .C(n19002), .Y(
        n22060) );
  A2O1A1Ixp33_ASAP7_75t_SL U21913 ( .A1(n32162), .A2(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__4_), .B(n18295), .C(n19002), .Y(
        n22059) );
  A2O1A1Ixp33_ASAP7_75t_SL U21914 ( .A1(n29417), .A2(n22057), .B(n18295), .C(
        n19002), .Y(n22058) );
  A2O1A1Ixp33_ASAP7_75t_SL U21915 ( .A1(n22056), .A2(n22058), .B(n18295), .C(
        n19002), .Y(n29665) );
  A2O1A1Ixp33_ASAP7_75t_SL U21916 ( .A1(n31712), .A2(n21771), .B(n18295), .C(
        n19002), .Y(n31723) );
  A2O1A1Ixp33_ASAP7_75t_SL U21917 ( .A1(n24366), .A2(timer0_N65), .B(n18295), 
        .C(n19002), .Y(n21770) );
  A2O1A1Ixp33_ASAP7_75t_SL U21918 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[56]), 
        .B(n18295), .C(n19002), .Y(n22055) );
  A2O1A1Ixp33_ASAP7_75t_SL U21919 ( .A1(n18988), .A2(n22054), .B(n18295), .C(
        n19002), .Y(mult_x_1196_n247) );
  A2O1A1Ixp33_ASAP7_75t_SL U21920 ( .A1(mult_x_1196_n405), .A2(n22366), .B(
        n18295), .C(n22421), .Y(n21062) );
  A2O1A1Ixp33_ASAP7_75t_SL U21921 ( .A1(n21061), .A2(n21062), .B(n18295), .C(
        n19002), .Y(n23327) );
  A2O1A1Ixp33_ASAP7_75t_SL U21922 ( .A1(n25315), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21560) );
  A2O1A1Ixp33_ASAP7_75t_SL U21923 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__5_), .A2(n22052), .B(n18295), 
        .C(n19002), .Y(n31560) );
  A2O1A1Ixp33_ASAP7_75t_SL U21924 ( .A1(n32353), .A2(n32310), .B(n18295), .C(
        n19002), .Y(n20176) );
  A2O1A1Ixp33_ASAP7_75t_SL U21925 ( .A1(uart1_r_TRADDR__3_), .A2(n22047), .B(
        n18295), .C(n19002), .Y(n27408) );
  A2O1A1Ixp33_ASAP7_75t_SL U21926 ( .A1(rst0_r_3_), .A2(n22040), .B(n18295), 
        .C(n19002), .Y(n11537) );
  A2O1A1Ixp33_ASAP7_75t_SL U21927 ( .A1(n31246), .A2(uart1_r_BRATE__7_), .B(
        n18295), .C(n19002), .Y(n21979) );
  A2O1A1Ixp33_ASAP7_75t_SL U21928 ( .A1(n31247), .A2(irqctrl0_r_IPEND__7_), 
        .B(n18295), .C(n19002), .Y(n21980) );
  A2O1A1Ixp33_ASAP7_75t_SL U21929 ( .A1(uart1_r_LOOPB_), .A2(n31950), .B(
        n18295), .C(n19002), .Y(n21981) );
  A2O1A1Ixp33_ASAP7_75t_SL U21930 ( .A1(n21979), .A2(n21980), .B(n18295), .C(
        n21981), .Y(n21982) );
  A2O1A1Ixp33_ASAP7_75t_SL U21931 ( .A1(uart1_r_RHOLD__29__7_), .A2(n31217), 
        .B(n18295), .C(n19002), .Y(n21989) );
  A2O1A1Ixp33_ASAP7_75t_SL U21932 ( .A1(n31214), .A2(uart1_r_RHOLD__1__7_), 
        .B(n18295), .C(n19002), .Y(n21990) );
  A2O1A1Ixp33_ASAP7_75t_SL U21933 ( .A1(uart1_r_RHOLD__28__7_), .A2(n31215), 
        .B(n18295), .C(n19002), .Y(n21991) );
  A2O1A1Ixp33_ASAP7_75t_SL U21934 ( .A1(n21989), .A2(n21990), .B(n18295), .C(
        n21991), .Y(n21992) );
  A2O1A1Ixp33_ASAP7_75t_SL U21935 ( .A1(n31220), .A2(uart1_r_RHOLD__13__7_), 
        .B(n18295), .C(n19002), .Y(n21994) );
  A2O1A1Ixp33_ASAP7_75t_SL U21936 ( .A1(n31218), .A2(uart1_r_RHOLD__23__7_), 
        .B(n18295), .C(n19002), .Y(n21995) );
  A2O1A1Ixp33_ASAP7_75t_SL U21937 ( .A1(n31219), .A2(uart1_r_RHOLD__11__7_), 
        .B(n18295), .C(n19002), .Y(n21996) );
  A2O1A1Ixp33_ASAP7_75t_SL U21938 ( .A1(n21994), .A2(n21995), .B(n18295), .C(
        n21996), .Y(n21997) );
  A2O1A1Ixp33_ASAP7_75t_SL U21939 ( .A1(n31212), .A2(uart1_r_RHOLD__26__7_), 
        .B(n18295), .C(n19002), .Y(n21999) );
  A2O1A1Ixp33_ASAP7_75t_SL U21940 ( .A1(n31210), .A2(uart1_r_RHOLD__21__7_), 
        .B(n18295), .C(n19002), .Y(n22000) );
  A2O1A1Ixp33_ASAP7_75t_SL U21941 ( .A1(uart1_r_RHOLD__20__7_), .A2(n31211), 
        .B(n18295), .C(n19002), .Y(n22001) );
  A2O1A1Ixp33_ASAP7_75t_SL U21942 ( .A1(n21999), .A2(n22000), .B(n18295), .C(
        n22001), .Y(n22002) );
  A2O1A1Ixp33_ASAP7_75t_SL U21943 ( .A1(uart1_r_RHOLD__25__7_), .A2(n31209), 
        .B(n18295), .C(n19002), .Y(n22004) );
  A2O1A1Ixp33_ASAP7_75t_SL U21944 ( .A1(uart1_r_RHOLD__7__7_), .A2(n31207), 
        .B(n18295), .C(n19002), .Y(n22005) );
  A2O1A1Ixp33_ASAP7_75t_SL U21945 ( .A1(n31206), .A2(uart1_r_RHOLD__17__7_), 
        .B(n18295), .C(n19002), .Y(n22006) );
  A2O1A1Ixp33_ASAP7_75t_SL U21946 ( .A1(n22004), .A2(n22005), .B(n18295), .C(
        n22006), .Y(n22007) );
  A2O1A1Ixp33_ASAP7_75t_SL U21947 ( .A1(n31202), .A2(uart1_r_RHOLD__12__7_), 
        .B(n18295), .C(n19002), .Y(n22009) );
  A2O1A1Ixp33_ASAP7_75t_SL U21948 ( .A1(n22003), .A2(n22008), .B(n18295), .C(
        n22009), .Y(n22010) );
  A2O1A1Ixp33_ASAP7_75t_SL U21949 ( .A1(n31225), .A2(uart1_r_RHOLD__10__7_), 
        .B(n18295), .C(n19002), .Y(n22011) );
  A2O1A1Ixp33_ASAP7_75t_SL U21950 ( .A1(uart1_r_RHOLD__4__7_), .A2(n31224), 
        .B(n18295), .C(n19002), .Y(n22012) );
  A2O1A1Ixp33_ASAP7_75t_SL U21951 ( .A1(n31223), .A2(uart1_r_RHOLD__2__7_), 
        .B(n18295), .C(n19002), .Y(n22013) );
  A2O1A1Ixp33_ASAP7_75t_SL U21952 ( .A1(n22011), .A2(n22012), .B(n18295), .C(
        n22013), .Y(n22014) );
  A2O1A1Ixp33_ASAP7_75t_SL U21953 ( .A1(uart1_r_RHOLD__22__7_), .A2(n31229), 
        .B(n18295), .C(n19002), .Y(n22016) );
  A2O1A1Ixp33_ASAP7_75t_SL U21954 ( .A1(n31227), .A2(uart1_r_RHOLD__8__7_), 
        .B(n18295), .C(n19002), .Y(n22017) );
  A2O1A1Ixp33_ASAP7_75t_SL U21955 ( .A1(uart1_r_RHOLD__18__7_), .A2(n31228), 
        .B(n18295), .C(n19002), .Y(n22018) );
  A2O1A1Ixp33_ASAP7_75t_SL U21956 ( .A1(n22016), .A2(n22017), .B(n18295), .C(
        n22018), .Y(n22019) );
  A2O1A1Ixp33_ASAP7_75t_SL U21957 ( .A1(uart1_r_RHOLD__30__7_), .A2(n31201), 
        .B(n18295), .C(n19002), .Y(n22021) );
  A2O1A1Ixp33_ASAP7_75t_SL U21958 ( .A1(n31204), .A2(uart1_r_RHOLD__9__7_), 
        .B(n18295), .C(n19002), .Y(n22022) );
  A2O1A1Ixp33_ASAP7_75t_SL U21959 ( .A1(uart1_r_RHOLD__16__7_), .A2(n31205), 
        .B(n18295), .C(n19002), .Y(n22023) );
  A2O1A1Ixp33_ASAP7_75t_SL U21960 ( .A1(n22021), .A2(n22022), .B(n18295), .C(
        n22023), .Y(n22024) );
  A2O1A1Ixp33_ASAP7_75t_SL U21961 ( .A1(n22015), .A2(n22020), .B(n18295), .C(
        n22025), .Y(n22026) );
  A2O1A1Ixp33_ASAP7_75t_SL U21962 ( .A1(n21993), .A2(n21998), .B(n18295), .C(
        n22027), .Y(n22028) );
  A2O1A1Ixp33_ASAP7_75t_SL U21963 ( .A1(n31242), .A2(uart1_r_RHOLD__0__7_), 
        .B(n18295), .C(n19002), .Y(n22032) );
  A2O1A1Ixp33_ASAP7_75t_SL U21964 ( .A1(n21988), .A2(n22031), .B(n18295), .C(
        n22032), .Y(n22033) );
  A2O1A1Ixp33_ASAP7_75t_SL U21965 ( .A1(n21983), .A2(n22034), .B(n18295), .C(
        n19002), .Y(n22035) );
  A2O1A1Ixp33_ASAP7_75t_SL U21966 ( .A1(n21738), .A2(n21739), .B(n18295), .C(
        n19002), .Y(n4749) );
  A2O1A1Ixp33_ASAP7_75t_SL U21967 ( .A1(n28184), .A2(n28185), .B(n18295), .C(
        n21966), .Y(n4676) );
  A2O1A1Ixp33_ASAP7_75t_SL U21968 ( .A1(n31364), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__13_), .B(n18295), .C(n19002), .Y(
        n21963) );
  A2O1A1Ixp33_ASAP7_75t_SL U21969 ( .A1(n30024), .A2(n31043), .B(n18295), .C(
        n19002), .Y(n21964) );
  A2O1A1Ixp33_ASAP7_75t_SL U21970 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[45]), 
        .B(n18295), .C(n19002), .Y(n21960) );
  A2O1A1Ixp33_ASAP7_75t_SL U21971 ( .A1(n21959), .A2(n21960), .B(n18295), .C(
        n19002), .Y(n21961) );
  A2O1A1Ixp33_ASAP7_75t_SL U21972 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[59]), 
        .B(n18295), .C(n19002), .Y(n21950) );
  A2O1A1Ixp33_ASAP7_75t_SL U21973 ( .A1(n21949), .A2(n21950), .B(n18295), .C(
        n19002), .Y(n21951) );
  A2O1A1Ixp33_ASAP7_75t_SL U21974 ( .A1(n30640), .A2(rf_do_b[10]), .B(n18295), 
        .C(n19002), .Y(n21939) );
  A2O1A1Ixp33_ASAP7_75t_SL U21975 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__10_), .B(n18295), .C(n19002), .Y(n21940)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U21976 ( .A1(n21939), .A2(n21940), .B(n18295), .C(
        n19002), .Y(n21941) );
  A2O1A1Ixp33_ASAP7_75t_SL U21977 ( .A1(n21944), .A2(n30593), .B(n18295), .C(
        n19002), .Y(n21945) );
  A2O1A1Ixp33_ASAP7_75t_SL U21978 ( .A1(n24664), .A2(n19745), .B(n18295), .C(
        n19002), .Y(n19746) );
  A2O1A1Ixp33_ASAP7_75t_SL U21979 ( .A1(n24662), .A2(n32614), .B(n18295), .C(
        n19002), .Y(n21929) );
  A2O1A1Ixp33_ASAP7_75t_SL U21980 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[37]), 
        .B(n18295), .C(n19002), .Y(n21927) );
  A2O1A1Ixp33_ASAP7_75t_SL U21981 ( .A1(n21926), .A2(n21927), .B(n18295), .C(
        n19002), .Y(n21928) );
  A2O1A1Ixp33_ASAP7_75t_SL U21982 ( .A1(n32570), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n21421) );
  A2O1A1Ixp33_ASAP7_75t_SL U21983 ( .A1(n31687), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21694) );
  A2O1A1Ixp33_ASAP7_75t_SL U21984 ( .A1(n29817), .A2(n24666), .B(n18295), .C(
        n19002), .Y(n21923) );
  A2O1A1Ixp33_ASAP7_75t_SL U21985 ( .A1(n32126), .A2(n32127), .B(n18295), .C(
        n32128), .Y(n21922) );
  A2O1A1Ixp33_ASAP7_75t_SL U21986 ( .A1(n24669), .A2(n21679), .B(n18295), .C(
        n19002), .Y(n21680) );
  A2O1A1Ixp33_ASAP7_75t_SL U21987 ( .A1(n29105), .A2(n24675), .B(n18295), .C(
        n19002), .Y(n21418) );
  A2O1A1Ixp33_ASAP7_75t_SL U21988 ( .A1(n24673), .A2(n25280), .B(n18295), .C(
        n19002), .Y(n21921) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U21989 ( .A1(n24672), .A2(n25314), .B(n18295), 
        .C(n19002), .Y(n21919) );
  A2O1A1Ixp33_ASAP7_75t_SL U21990 ( .A1(n31980), .A2(n24659), .B(n18295), .C(
        n19002), .Y(n21674) );
  A2O1A1Ixp33_ASAP7_75t_SL U21991 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA1__0_), 
        .A2(n24660), .B(n18295), .C(n19002), .Y(n21914) );
  A2O1A1Ixp33_ASAP7_75t_SL U21992 ( .A1(n32176), .A2(n21914), .B(n18295), .C(
        n19002), .Y(n21915) );
  A2O1A1Ixp33_ASAP7_75t_SL U21993 ( .A1(n19002), .A2(n21915), .B(n18295), .C(
        n19002), .Y(n4169) );
  A2O1A1Ixp33_ASAP7_75t_SL U21994 ( .A1(n32608), .A2(n24667), .B(n18295), .C(
        n19002), .Y(n21411) );
  A2O1A1Ixp33_ASAP7_75t_SL U21995 ( .A1(n26753), .A2(n24673), .B(n18295), .C(
        n19002), .Y(n21671) );
  A2O1A1Ixp33_ASAP7_75t_SL U21996 ( .A1(n30920), .A2(n24668), .B(n18295), .C(
        n19002), .Y(n21409) );
  A2O1A1Ixp33_ASAP7_75t_SL U21997 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__18_), .A2(
        n21907), .B(n18295), .C(n19002), .Y(n21908) );
  A2O1A1Ixp33_ASAP7_75t_SL U21998 ( .A1(n28556), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n21906) );
  A2O1A1Ixp33_ASAP7_75t_SL U21999 ( .A1(n24663), .A2(n32612), .B(n18295), .C(
        n19002), .Y(n21905) );
  A2O1A1Ixp33_ASAP7_75t_SL U22000 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TT__4_), 
        .A2(n3916), .B(n18295), .C(n19002), .Y(n21901) );
  A2O1A1Ixp33_ASAP7_75t_SL U22001 ( .A1(n24659), .A2(n29741), .B(n18295), .C(
        n19002), .Y(n21903) );
  A2O1A1Ixp33_ASAP7_75t_SL U22002 ( .A1(n31815), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n21660) );
  A2O1A1Ixp33_ASAP7_75t_SL U22003 ( .A1(n24681), .A2(n30381), .B(n18295), .C(
        n19002), .Y(n21659) );
  A2O1A1Ixp33_ASAP7_75t_SL U22004 ( .A1(n24681), .A2(n28576), .B(n18295), .C(
        n19002), .Y(n21658) );
  A2O1A1Ixp33_ASAP7_75t_SL U22005 ( .A1(n24669), .A2(n26369), .B(n18295), .C(
        n19002), .Y(n21898) );
  A2O1A1Ixp33_ASAP7_75t_SL U22006 ( .A1(n24681), .A2(n30402), .B(n18295), .C(
        n19002), .Y(n21656) );
  A2O1A1Ixp33_ASAP7_75t_SL U22007 ( .A1(n30243), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21390) );
  A2O1A1Ixp33_ASAP7_75t_SL U22008 ( .A1(n30238), .A2(n24671), .B(n18295), .C(
        n19002), .Y(n21650) );
  A2O1A1Ixp33_ASAP7_75t_SL U22009 ( .A1(n24674), .A2(n21891), .B(n18295), .C(
        n19002), .Y(n21892) );
  A2O1A1Ixp33_ASAP7_75t_SL U22010 ( .A1(n24668), .A2(n21165), .B(n18295), .C(
        n19002), .Y(n21166) );
  A2O1A1Ixp33_ASAP7_75t_SL U22011 ( .A1(n24671), .A2(n21888), .B(n18295), .C(
        n19002), .Y(n21889) );
  A2O1A1Ixp33_ASAP7_75t_SL U22012 ( .A1(n19002), .A2(n24907), .B(n18295), .C(
        n19002), .Y(n21884) );
  A2O1A1Ixp33_ASAP7_75t_SL U22013 ( .A1(n24906), .A2(n21884), .B(n18295), .C(
        n19002), .Y(n21885) );
  A2O1A1Ixp33_ASAP7_75t_SL U22014 ( .A1(n21885), .A2(n21886), .B(n18295), .C(
        n19002), .Y(n21887) );
  A2O1A1Ixp33_ASAP7_75t_SL U22015 ( .A1(n23229), .A2(n31651), .B(n18295), .C(
        n19002), .Y(n21647) );
  A2O1A1Ixp33_ASAP7_75t_SL U22016 ( .A1(n30120), .A2(n24665), .B(n18295), .C(
        n19002), .Y(n21646) );
  A2O1A1Ixp33_ASAP7_75t_SL U22017 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA2__7_), 
        .A2(n24660), .B(n18295), .C(n19002), .Y(n21157) );
  A2O1A1Ixp33_ASAP7_75t_SL U22018 ( .A1(n32574), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21642) );
  A2O1A1Ixp33_ASAP7_75t_SL U22019 ( .A1(n24660), .A2(n29684), .B(n18295), .C(
        n19002), .Y(n21872) );
  A2O1A1Ixp33_ASAP7_75t_SL U22020 ( .A1(n32137), .A2(n32139), .B(n18295), .C(
        n32138), .Y(n20964) );
  A2O1A1Ixp33_ASAP7_75t_SL U22021 ( .A1(n32141), .A2(n20964), .B(n18295), .C(
        n19002), .Y(n20965) );
  A2O1A1Ixp33_ASAP7_75t_SL U22022 ( .A1(n22379), .A2(n20966), .B(n18295), .C(
        n19002), .Y(n20967) );
  A2O1A1Ixp33_ASAP7_75t_SL U22023 ( .A1(n24676), .A2(n21638), .B(n18295), .C(
        n19002), .Y(n21639) );
  A2O1A1Ixp33_ASAP7_75t_SL U22024 ( .A1(n28271), .A2(n22427), .B(n18295), .C(
        n19002), .Y(n20620) );
  A2O1A1Ixp33_ASAP7_75t_SL U22025 ( .A1(n24677), .A2(n19308), .B(n18295), .C(
        n19002), .Y(n19309) );
  A2O1A1Ixp33_ASAP7_75t_SL U22026 ( .A1(n32142), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n20785) );
  A2O1A1Ixp33_ASAP7_75t_SL U22027 ( .A1(n22396), .A2(n21861), .B(n18295), .C(
        n19002), .Y(n21862) );
  A2O1A1Ixp33_ASAP7_75t_SL U22028 ( .A1(n22396), .A2(n21857), .B(n18295), .C(
        n19002), .Y(n21858) );
  A2O1A1Ixp33_ASAP7_75t_SL U22029 ( .A1(n22396), .A2(n21855), .B(n18295), .C(
        n19002), .Y(n21856) );
  A2O1A1Ixp33_ASAP7_75t_SL U22030 ( .A1(n22396), .A2(n21853), .B(n18295), .C(
        n19002), .Y(n21854) );
  A2O1A1Ixp33_ASAP7_75t_SL U22031 ( .A1(n32592), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n21625) );
  A2O1A1Ixp33_ASAP7_75t_SL U22032 ( .A1(n30730), .A2(n24662), .B(n18295), .C(
        n19002), .Y(n21624) );
  A2O1A1Ixp33_ASAP7_75t_SL U22033 ( .A1(n19002), .A2(n21840), .B(n18295), .C(
        n19002), .Y(n32551) );
  A2O1A1Ixp33_ASAP7_75t_SL U22034 ( .A1(n31197), .A2(n31198), .B(n18295), .C(
        n19002), .Y(n21128) );
  A2O1A1Ixp33_ASAP7_75t_SL U22035 ( .A1(n24604), .A2(n24595), .B(n18295), .C(
        n19002), .Y(n21120) );
  A2O1A1Ixp33_ASAP7_75t_SL U22036 ( .A1(n24601), .A2(n24602), .B(n18295), .C(
        n21121), .Y(n21122) );
  A2O1A1Ixp33_ASAP7_75t_SL U22037 ( .A1(n30978), .A2(n24633), .B(n18295), .C(
        n19002), .Y(n21345) );
  A2O1A1Ixp33_ASAP7_75t_SL U22038 ( .A1(n30073), .A2(n24633), .B(n18295), .C(
        n19002), .Y(n21344) );
  A2O1A1Ixp33_ASAP7_75t_SL U22039 ( .A1(n29383), .A2(n21837), .B(n18295), .C(
        n19002), .Y(n21838) );
  A2O1A1Ixp33_ASAP7_75t_SL U22040 ( .A1(n23229), .A2(n32164), .B(n18295), .C(
        n19002), .Y(n21834) );
  A2O1A1Ixp33_ASAP7_75t_SL U22041 ( .A1(n21833), .A2(n21834), .B(n18295), .C(
        n19002), .Y(n21835) );
  A2O1A1Ixp33_ASAP7_75t_SL U22042 ( .A1(n19002), .A2(n21835), .B(n18295), .C(
        n19002), .Y(n2776) );
  A2O1A1Ixp33_ASAP7_75t_SL U22043 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA1__5_), 
        .A2(n24660), .B(n18295), .C(n19002), .Y(n21611) );
  A2O1A1Ixp33_ASAP7_75t_SL U22044 ( .A1(n24681), .A2(n30219), .B(n18295), .C(
        n19002), .Y(n21343) );
  A2O1A1Ixp33_ASAP7_75t_SL U22045 ( .A1(n30428), .A2(n24673), .B(n18295), .C(
        n19002), .Y(n21605) );
  A2O1A1Ixp33_ASAP7_75t_SL U22046 ( .A1(n24659), .A2(n21829), .B(n18295), .C(
        n19002), .Y(n21830) );
  A2O1A1Ixp33_ASAP7_75t_SL U22047 ( .A1(n24675), .A2(n21599), .B(n18295), .C(
        n19002), .Y(n21600) );
  A2O1A1Ixp33_ASAP7_75t_SL U22048 ( .A1(n24670), .A2(n28538), .B(n18295), .C(
        n19002), .Y(n21821) );
  A2O1A1Ixp33_ASAP7_75t_SL U22049 ( .A1(n27499), .A2(n27513), .B(n18295), .C(
        n19002), .Y(n21585) );
  A2O1A1Ixp33_ASAP7_75t_SL U22050 ( .A1(n19002), .A2(n21809), .B(n18295), .C(
        n19002), .Y(n32557) );
  A2O1A1Ixp33_ASAP7_75t_SL U22051 ( .A1(u0_0_leon3x0_p0_iu_r_X__ICC__0_), .A2(
        n20285), .B(n18295), .C(n19002), .Y(n20286) );
  A2O1A1Ixp33_ASAP7_75t_SL U22052 ( .A1(n26084), .A2(n19686), .B(n18295), .C(
        n19002), .Y(n19687) );
  A2O1A1Ixp33_ASAP7_75t_SL U22053 ( .A1(n26086), .A2(n26085), .B(n18295), .C(
        n19687), .Y(n2245) );
  A2O1A1Ixp33_ASAP7_75t_SL U22054 ( .A1(n24694), .A2(timer0_gpto_TICK__0_), 
        .B(n18295), .C(n18872), .Y(n24554) );
  A2O1A1Ixp33_ASAP7_75t_SL U22055 ( .A1(ahb0_r_HADDR__3_), .A2(n21798), .B(
        n18295), .C(n19002), .Y(n17273) );
  A2O1A1Ixp33_ASAP7_75t_SL U22056 ( .A1(n32583), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__5_), .B(n18295), .C(n19002), 
        .Y(n21793) );
  A2O1A1Ixp33_ASAP7_75t_SL U22057 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__10_), 
        .A2(n32584), .B(n18295), .C(n19002), .Y(n21794) );
  A2O1A1Ixp33_ASAP7_75t_SL U22058 ( .A1(n21793), .A2(n21794), .B(n18295), .C(
        n19002), .Y(n21795) );
  A2O1A1Ixp33_ASAP7_75t_SL U22059 ( .A1(n32587), .A2(n32588), .B(n18295), .C(
        n19002), .Y(n21797) );
  A2O1A1Ixp33_ASAP7_75t_SL U22060 ( .A1(n21796), .A2(n21797), .B(n18295), .C(
        n19002), .Y(ic_address[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22061 ( .A1(n32660), .A2(n32659), .B(n18295), .C(
        n19002), .Y(n21791) );
  A2O1A1Ixp33_ASAP7_75t_SL U22062 ( .A1(n32660), .A2(n32651), .B(n18295), .C(
        n19002), .Y(n21790) );
  A2O1A1Ixp33_ASAP7_75t_SL U22063 ( .A1(n32660), .A2(n32649), .B(n18295), .C(
        n19002), .Y(n21789) );
  A2O1A1Ixp33_ASAP7_75t_SL U22064 ( .A1(n32660), .A2(n32647), .B(n18295), .C(
        n19002), .Y(n21788) );
  A2O1A1Ixp33_ASAP7_75t_SL U22065 ( .A1(n32660), .A2(n32645), .B(n18295), .C(
        n19002), .Y(n21787) );
  A2O1A1Ixp33_ASAP7_75t_SL U22066 ( .A1(n32660), .A2(n32631), .B(n18295), .C(
        n19002), .Y(n21786) );
  A2O1A1Ixp33_ASAP7_75t_SL U22067 ( .A1(n32605), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n20428) );
  A2O1A1Ixp33_ASAP7_75t_SL U22068 ( .A1(n32601), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n21575) );
  A2O1A1Ixp33_ASAP7_75t_SL U22069 ( .A1(n32625), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n21780) );
  A2O1A1Ixp33_ASAP7_75t_SL U22070 ( .A1(n32344), .A2(dc_q[14]), .B(n18295), 
        .C(n19002), .Y(n21781) );
  A2O1A1Ixp33_ASAP7_75t_SL U22071 ( .A1(n21780), .A2(n21781), .B(n18295), .C(
        n19002), .Y(n21782) );
  A2O1A1Ixp33_ASAP7_75t_SL U22072 ( .A1(n32345), .A2(n32423), .B(n18295), .C(
        n19002), .Y(n21784) );
  A2O1A1Ixp33_ASAP7_75t_SL U22073 ( .A1(n21783), .A2(n21784), .B(n18295), .C(
        n19002), .Y(dc_data[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22074 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[30]), 
        .A2(n32231), .B(n18295), .C(n19002), .Y(n21778) );
  A2O1A1Ixp33_ASAP7_75t_SL U22075 ( .A1(n21777), .A2(n21778), .B(n18295), .C(
        n19002), .Y(dt_data[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22076 ( .A1(n24661), .A2(
        u0_0_leon3x0_p0_iu_r_A__RFA2__6_), .B(n18295), .C(n19002), .Y(n21775)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22077 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA2__5_), 
        .A2(n24661), .B(n18295), .C(n19002), .Y(n21568) );
  A2O1A1Ixp33_ASAP7_75t_SL U22078 ( .A1(n32162), .A2(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__6_), .B(n18295), .C(n19002), .Y(
        n21773) );
  A2O1A1Ixp33_ASAP7_75t_SL U22079 ( .A1(n29467), .A2(n30687), .B(n18295), .C(
        n19002), .Y(n19820) );
  A2O1A1Ixp33_ASAP7_75t_SL U22080 ( .A1(n31299), .A2(n21768), .B(n18295), .C(
        n19002), .Y(n31617) );
  A2O1A1Ixp33_ASAP7_75t_SL U22081 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[50]), 
        .B(n18295), .C(n19002), .Y(n21767) );
  A2O1A1Ixp33_ASAP7_75t_SL U22082 ( .A1(n32489), .A2(n32496), .B(n18295), .C(
        n19002), .Y(n21762) );
  A2O1A1Ixp33_ASAP7_75t_SL U22083 ( .A1(n32518), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__4_), .B(n18295), .C(n19002), 
        .Y(n21766) );
  A2O1A1Ixp33_ASAP7_75t_SL U22084 ( .A1(n21765), .A2(n21766), .B(n18295), .C(
        n19002), .Y(n32493) );
  A2O1A1Ixp33_ASAP7_75t_SL U22085 ( .A1(n24642), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[10]), .B(n18295), .C(n19002), .Y(n21760)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22086 ( .A1(mult_x_1196_n464), .A2(n22676), .B(
        n18295), .C(n21757), .Y(mult_x_1196_n357) );
  A2O1A1Ixp33_ASAP7_75t_SL U22087 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__0_), .B(n18295), .C(n19002), .Y(
        n21756) );
  A2O1A1Ixp33_ASAP7_75t_SL U22088 ( .A1(mult_x_1196_n317), .A2(n21755), .B(
        n18295), .C(n19002), .Y(mult_x_1196_n227) );
  A2O1A1Ixp33_ASAP7_75t_SL U22089 ( .A1(n31951), .A2(uart1_r_OVF_), .B(n18295), 
        .C(n19002), .Y(n21478) );
  A2O1A1Ixp33_ASAP7_75t_SL U22090 ( .A1(irqctrl0_r_ILEVEL__4_), .A2(n31248), 
        .B(n18295), .C(n19002), .Y(n21479) );
  A2O1A1Ixp33_ASAP7_75t_SL U22091 ( .A1(timer0_r_SCALER__4_), .A2(n31245), .B(
        n18295), .C(n19002), .Y(n21480) );
  A2O1A1Ixp33_ASAP7_75t_SL U22092 ( .A1(n21478), .A2(n21479), .B(n18295), .C(
        n21480), .Y(n21481) );
  A2O1A1Ixp33_ASAP7_75t_SL U22093 ( .A1(n30786), .A2(n30785), .B(n18295), .C(
        n19002), .Y(n21485) );
  A2O1A1Ixp33_ASAP7_75t_SL U22094 ( .A1(n30788), .A2(n30787), .B(n18295), .C(
        n19002), .Y(n21486) );
  A2O1A1Ixp33_ASAP7_75t_SL U22095 ( .A1(n31207), .A2(uart1_r_RHOLD__7__4_), 
        .B(n18295), .C(n19002), .Y(n21487) );
  A2O1A1Ixp33_ASAP7_75t_SL U22096 ( .A1(n31209), .A2(uart1_r_RHOLD__25__4_), 
        .B(n18295), .C(n19002), .Y(n21488) );
  A2O1A1Ixp33_ASAP7_75t_SL U22097 ( .A1(uart1_r_RHOLD__17__4_), .A2(n31206), 
        .B(n18295), .C(n19002), .Y(n21489) );
  A2O1A1Ixp33_ASAP7_75t_SL U22098 ( .A1(n21487), .A2(n21488), .B(n18295), .C(
        n21489), .Y(n21490) );
  A2O1A1Ixp33_ASAP7_75t_SL U22099 ( .A1(uart1_r_RHOLD__21__4_), .A2(n31210), 
        .B(n18295), .C(n19002), .Y(n21492) );
  A2O1A1Ixp33_ASAP7_75t_SL U22100 ( .A1(uart1_r_RHOLD__26__4_), .A2(n31212), 
        .B(n18295), .C(n19002), .Y(n21493) );
  A2O1A1Ixp33_ASAP7_75t_SL U22101 ( .A1(uart1_r_RHOLD__20__4_), .A2(n31211), 
        .B(n18295), .C(n19002), .Y(n21494) );
  A2O1A1Ixp33_ASAP7_75t_SL U22102 ( .A1(n21492), .A2(n21493), .B(n18295), .C(
        n21494), .Y(n21495) );
  A2O1A1Ixp33_ASAP7_75t_SL U22103 ( .A1(n31203), .A2(uart1_r_RHOLD__14__4_), 
        .B(n18295), .C(n19002), .Y(n21497) );
  A2O1A1Ixp33_ASAP7_75t_SL U22104 ( .A1(n21498), .A2(n21499), .B(n18295), .C(
        n19002), .Y(n21500) );
  A2O1A1Ixp33_ASAP7_75t_SL U22105 ( .A1(uart1_r_RHOLD__12__4_), .A2(n31202), 
        .B(n18295), .C(n19002), .Y(n21502) );
  A2O1A1Ixp33_ASAP7_75t_SL U22106 ( .A1(n21497), .A2(n21501), .B(n18295), .C(
        n21502), .Y(n21503) );
  A2O1A1Ixp33_ASAP7_75t_SL U22107 ( .A1(uart1_r_RHOLD__4__4_), .A2(n31224), 
        .B(n18295), .C(n19002), .Y(n21506) );
  A2O1A1Ixp33_ASAP7_75t_SL U22108 ( .A1(n31226), .A2(uart1_r_RHOLD__6__4_), 
        .B(n18295), .C(n19002), .Y(n21507) );
  A2O1A1Ixp33_ASAP7_75t_SL U22109 ( .A1(uart1_r_RHOLD__10__4_), .A2(n31225), 
        .B(n18295), .C(n19002), .Y(n21508) );
  A2O1A1Ixp33_ASAP7_75t_SL U22110 ( .A1(n30784), .A2(n21507), .B(n18295), .C(
        n21508), .Y(n21509) );
  A2O1A1Ixp33_ASAP7_75t_SL U22111 ( .A1(n21510), .A2(n21511), .B(n18295), .C(
        n19002), .Y(n21512) );
  A2O1A1Ixp33_ASAP7_75t_SL U22112 ( .A1(uart1_r_RHOLD__2__4_), .A2(n31223), 
        .B(n18295), .C(n19002), .Y(n21514) );
  A2O1A1Ixp33_ASAP7_75t_SL U22113 ( .A1(n21506), .A2(n21513), .B(n18295), .C(
        n21514), .Y(n21515) );
  A2O1A1Ixp33_ASAP7_75t_SL U22114 ( .A1(n21491), .A2(n21496), .B(n18295), .C(
        n21516), .Y(n21517) );
  A2O1A1Ixp33_ASAP7_75t_SL U22115 ( .A1(n21521), .A2(n21522), .B(n18295), .C(
        n19002), .Y(n21523) );
  A2O1A1Ixp33_ASAP7_75t_SL U22116 ( .A1(n31235), .A2(sr1_r_MCFG1__ROMWWS__0_), 
        .B(n18295), .C(n19002), .Y(n21525) );
  A2O1A1Ixp33_ASAP7_75t_SL U22117 ( .A1(irqctrl0_r_IMASK__0__4_), .A2(n31249), 
        .B(n18295), .C(n19002), .Y(n21528) );
  A2O1A1Ixp33_ASAP7_75t_SL U22118 ( .A1(sr1_r_MCFG2__RAMWIDTH__0_), .A2(n31250), .B(n18295), .C(n19002), .Y(n21531) );
  A2O1A1Ixp33_ASAP7_75t_SL U22119 ( .A1(n21525), .A2(n21530), .B(n18295), .C(
        n21531), .Y(n21532) );
  A2O1A1Ixp33_ASAP7_75t_SL U22120 ( .A1(n31240), .A2(n30782), .B(n18295), .C(
        n19002), .Y(n21536) );
  A2O1A1Ixp33_ASAP7_75t_SL U22121 ( .A1(n18295), .A2(n19002), .B(n21535), .C(
        n21536), .Y(n21537) );
  A2O1A1Ixp33_ASAP7_75t_SL U22122 ( .A1(n29659), .A2(n29660), .B(n18295), .C(
        n19002), .Y(n21740) );
  A2O1A1Ixp33_ASAP7_75t_SL U22123 ( .A1(n29665), .A2(n29660), .B(n18295), .C(
        n21743), .Y(n21744) );
  A2O1A1Ixp33_ASAP7_75t_SL U22124 ( .A1(n21742), .A2(n21744), .B(n18295), .C(
        n19002), .Y(n21745) );
  A2O1A1Ixp33_ASAP7_75t_SL U22125 ( .A1(n29664), .A2(n21745), .B(n18295), .C(
        n19002), .Y(n21746) );
  A2O1A1Ixp33_ASAP7_75t_SL U22126 ( .A1(n29666), .A2(n21746), .B(n18295), .C(
        n19002), .Y(irqctrl0_v_IRL__0__1_) );
  A2O1A1Ixp33_ASAP7_75t_SL U22127 ( .A1(n24681), .A2(n32568), .B(n18295), .C(
        n19002), .Y(n21738) );
  A2O1A1Ixp33_ASAP7_75t_SL U22128 ( .A1(n22428), .A2(n32567), .B(n18295), .C(
        n19002), .Y(n21739) );
  A2O1A1Ixp33_ASAP7_75t_SL U22129 ( .A1(u0_0_leon3x0_p0_c0mmu_icache0_r_BURST_), .A2(n32662), .B(n18295), .C(n19002), .Y(n21731) );
  A2O1A1Ixp33_ASAP7_75t_SL U22130 ( .A1(n32705), .A2(n32511), .B(n18295), .C(
        n31876), .Y(n21732) );
  A2O1A1Ixp33_ASAP7_75t_SL U22131 ( .A1(n32564), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__BURST_), .B(n18295), .C(n19002), 
        .Y(n21735) );
  A2O1A1Ixp33_ASAP7_75t_SL U22132 ( .A1(n31883), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_BURST_), .B(n18295), .C(n19002), .Y(
        n21736) );
  A2O1A1Ixp33_ASAP7_75t_SL U22133 ( .A1(n21244), .A2(n32749), .B(n18295), .C(
        n19002), .Y(n21245) );
  A2O1A1Ixp33_ASAP7_75t_SL U22134 ( .A1(n21464), .A2(n21465), .B(n18295), .C(
        n19002), .Y(n21466) );
  A2O1A1Ixp33_ASAP7_75t_SL U22135 ( .A1(n29618), .A2(n29617), .B(n18295), .C(
        n31542), .Y(n21724) );
  A2O1A1Ixp33_ASAP7_75t_SL U22136 ( .A1(n21723), .A2(n21724), .B(n18295), .C(
        n19002), .Y(n4658) );
  A2O1A1Ixp33_ASAP7_75t_SL U22137 ( .A1(n4832), .A2(n24694), .B(n18295), .C(
        n19002), .Y(n21720) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U22138 ( .A1(n32039), .A2(n32002), .B(n18295), 
        .C(n31803), .D(n21721), .Y(n4650) );
  A2O1A1Ixp33_ASAP7_75t_SL U22139 ( .A1(n21450), .A2(n21451), .B(n18295), .C(
        n19002), .Y(n21452) );
  A2O1A1Ixp33_ASAP7_75t_SL U22140 ( .A1(n21453), .A2(n21454), .B(n18295), .C(
        n19002), .Y(n21455) );
  A2O1A1Ixp33_ASAP7_75t_SL U22141 ( .A1(n23842), .A2(n24678), .B(n18295), .C(
        n19002), .Y(n21459) );
  A2O1A1Ixp33_ASAP7_75t_SL U22142 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[57]), 
        .B(n18295), .C(n19002), .Y(n21718) );
  A2O1A1Ixp33_ASAP7_75t_SL U22143 ( .A1(n21717), .A2(n21718), .B(n18295), .C(
        n19002), .Y(n21719) );
  A2O1A1Ixp33_ASAP7_75t_SL U22144 ( .A1(n24660), .A2(n21711), .B(n18295), .C(
        n19002), .Y(n21712) );
  A2O1A1Ixp33_ASAP7_75t_SL U22145 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[41]), 
        .B(n18295), .C(n19002), .Y(n21709) );
  A2O1A1Ixp33_ASAP7_75t_SL U22146 ( .A1(n21708), .A2(n21709), .B(n18295), .C(
        n19002), .Y(n21710) );
  A2O1A1Ixp33_ASAP7_75t_SL U22147 ( .A1(n22396), .A2(n21705), .B(n18295), .C(
        n19002), .Y(n21706) );
  A2O1A1Ixp33_ASAP7_75t_SL U22148 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), 
        .A2(u0_0_leon3x0_p0_iu_r_X__ICC__0_), .B(n18295), .C(n19002), .Y(
        n21434) );
  A2O1A1Ixp33_ASAP7_75t_SL U22149 ( .A1(n21436), .A2(n30953), .B(n18295), .C(
        n19002), .Y(n21437) );
  A2O1A1Ixp33_ASAP7_75t_SL U22150 ( .A1(n21426), .A2(n21433), .B(n18295), .C(
        n19002), .Y(n4467) );
  A2O1A1Ixp33_ASAP7_75t_SL U22151 ( .A1(n22408), .A2(n21698), .B(n18295), .C(
        n21699), .Y(n4389) );
  A2O1A1Ixp33_ASAP7_75t_SL U22152 ( .A1(n32610), .A2(n24663), .B(n18295), .C(
        n19002), .Y(n21697) );
  A2O1A1Ixp33_ASAP7_75t_SL U22153 ( .A1(n31457), .A2(n21685), .B(n18295), .C(
        n19002), .Y(n21686) );
  A2O1A1Ixp33_ASAP7_75t_SL U22154 ( .A1(n24684), .A2(n31459), .B(n18295), .C(
        n32292), .Y(n21689) );
  A2O1A1Ixp33_ASAP7_75t_SL U22155 ( .A1(n21688), .A2(n21690), .B(n18295), .C(
        n19002), .Y(n21691) );
  A2O1A1Ixp33_ASAP7_75t_SL U22156 ( .A1(n21692), .A2(n21693), .B(n18295), .C(
        n19002), .Y(u0_0_leon3x0_p0_c0mmu_dcache0_v_HOLDN_) );
  A2O1A1Ixp33_ASAP7_75t_SL U22157 ( .A1(n24673), .A2(n25281), .B(n18295), .C(
        n19002), .Y(n21677) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U22158 ( .A1(n24671), .A2(n25322), .B(n18295), 
        .C(n19002), .Y(n21676) );
  A2O1A1Ixp33_ASAP7_75t_SL U22159 ( .A1(n32640), .A2(n24666), .B(n18295), .C(
        n19002), .Y(n19737) );
  A2O1A1Ixp33_ASAP7_75t_SL U22160 ( .A1(n24673), .A2(n21672), .B(n18295), .C(
        n19002), .Y(n21673) );
  A2O1A1Ixp33_ASAP7_75t_SL U22161 ( .A1(n24665), .A2(n21669), .B(n18295), .C(
        n19002), .Y(n21670) );
  A2O1A1Ixp33_ASAP7_75t_SL U22162 ( .A1(n24661), .A2(n21407), .B(n18295), .C(
        n19002), .Y(n21408) );
  A2O1A1Ixp33_ASAP7_75t_SL U22163 ( .A1(n24663), .A2(n21405), .B(n18295), .C(
        n19002), .Y(n21406) );
  A2O1A1Ixp33_ASAP7_75t_SL U22164 ( .A1(n30370), .A2(n24666), .B(n18295), .C(
        n19002), .Y(n21404) );
  A2O1A1Ixp33_ASAP7_75t_SL U22165 ( .A1(n24669), .A2(n21667), .B(n18295), .C(
        n19002), .Y(n21668) );
  A2O1A1Ixp33_ASAP7_75t_SL U22166 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[36]), 
        .B(n18295), .C(n19002), .Y(n21663) );
  A2O1A1Ixp33_ASAP7_75t_SL U22167 ( .A1(n21662), .A2(n21663), .B(n18295), .C(
        n19002), .Y(n21664) );
  A2O1A1Ixp33_ASAP7_75t_SL U22168 ( .A1(n28273), .A2(n24681), .B(n18295), .C(
        n19002), .Y(n21657) );
  A2O1A1Ixp33_ASAP7_75t_SL U22169 ( .A1(n31680), .A2(n24666), .B(n18295), .C(
        n19002), .Y(n21399) );
  A2O1A1Ixp33_ASAP7_75t_SL U22170 ( .A1(n24681), .A2(n30393), .B(n18295), .C(
        n21654), .Y(n21655) );
  A2O1A1Ixp33_ASAP7_75t_SL U22171 ( .A1(n24681), .A2(n30312), .B(n18295), .C(
        n19002), .Y(n21395) );
  A2O1A1Ixp33_ASAP7_75t_SL U22172 ( .A1(n30296), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21394) );
  A2O1A1Ixp33_ASAP7_75t_SL U22173 ( .A1(n24681), .A2(n30282), .B(n18295), .C(
        n19002), .Y(n21393) );
  A2O1A1Ixp33_ASAP7_75t_SL U22174 ( .A1(n30262), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21392) );
  A2O1A1Ixp33_ASAP7_75t_SL U22175 ( .A1(n30247), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21391) );
  A2O1A1Ixp33_ASAP7_75t_SL U22176 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA1__1_), 
        .A2(n24660), .B(n18295), .C(n19002), .Y(n21648) );
  A2O1A1Ixp33_ASAP7_75t_SL U22177 ( .A1(n32177), .A2(n21648), .B(n18295), .C(
        n19002), .Y(n21649) );
  A2O1A1Ixp33_ASAP7_75t_SL U22178 ( .A1(n19002), .A2(n21649), .B(n18295), .C(
        n19002), .Y(n3758) );
  A2O1A1Ixp33_ASAP7_75t_SL U22179 ( .A1(n19002), .A2(n18295), .B(n20087), .C(
        n19002), .Y(n20088) );
  A2O1A1Ixp33_ASAP7_75t_SL U22180 ( .A1(n18295), .A2(n19002), .B(n21388), .C(
        n19002), .Y(n24508) );
  A2O1A1Ixp33_ASAP7_75t_SL U22181 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA2__3_), 
        .A2(n24661), .B(n18295), .C(n19002), .Y(n21382) );
  A2O1A1Ixp33_ASAP7_75t_SL U22182 ( .A1(n18295), .A2(n19002), .B(n19713), .C(
        n19002), .Y(n19714) );
  A2O1A1Ixp33_ASAP7_75t_SL U22183 ( .A1(n19712), .A2(n19714), .B(n18295), .C(
        n19002), .Y(n3532) );
  A2O1A1Ixp33_ASAP7_75t_SL U22184 ( .A1(n24660), .A2(n20624), .B(n18295), .C(
        n19002), .Y(n20625) );
  A2O1A1Ixp33_ASAP7_75t_SL U22185 ( .A1(n24677), .A2(n21377), .B(n18295), .C(
        n19002), .Y(n21378) );
  A2O1A1Ixp33_ASAP7_75t_SL U22186 ( .A1(n29032), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21373) );
  A2O1A1Ixp33_ASAP7_75t_SL U22187 ( .A1(n29034), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21372) );
  A2O1A1Ixp33_ASAP7_75t_SL U22188 ( .A1(n24678), .A2(n21636), .B(n18295), .C(
        n19002), .Y(n21637) );
  A2O1A1Ixp33_ASAP7_75t_SL U22189 ( .A1(n32586), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21369) );
  A2O1A1Ixp33_ASAP7_75t_SL U22190 ( .A1(u0_0_leon3x0_p0_muli[6]), .A2(n21633), 
        .B(n18295), .C(n19002), .Y(n21634) );
  A2O1A1Ixp33_ASAP7_75t_SL U22191 ( .A1(n22396), .A2(n21631), .B(n18295), .C(
        n19002), .Y(n21632) );
  A2O1A1Ixp33_ASAP7_75t_SL U22192 ( .A1(n22396), .A2(n21628), .B(n18295), .C(
        n19002), .Y(n21629) );
  A2O1A1Ixp33_ASAP7_75t_SL U22193 ( .A1(n22396), .A2(n21626), .B(n18295), .C(
        n19002), .Y(n21627) );
  A2O1A1Ixp33_ASAP7_75t_SL U22194 ( .A1(n22378), .A2(n28520), .B(n18295), .C(
        n19002), .Y(n21621) );
  A2O1A1Ixp33_ASAP7_75t_SL U22195 ( .A1(n29071), .A2(n22378), .B(n18295), .C(
        n19002), .Y(n21353) );
  A2O1A1Ixp33_ASAP7_75t_SL U22196 ( .A1(n26910), .A2(n24667), .B(n18295), .C(
        n19002), .Y(n21136) );
  A2O1A1Ixp33_ASAP7_75t_SL U22197 ( .A1(n19002), .A2(n28179), .B(n18295), .C(
        n19002), .Y(n21125) );
  A2O1A1Ixp33_ASAP7_75t_SL U22198 ( .A1(n21124), .A2(n21126), .B(n18295), .C(
        n19002), .Y(n21127) );
  A2O1A1Ixp33_ASAP7_75t_SL U22199 ( .A1(n30984), .A2(n29383), .B(n18295), .C(
        n19002), .Y(n20295) );
  A2O1A1Ixp33_ASAP7_75t_SL U22200 ( .A1(n23229), .A2(n32184), .B(n18295), .C(
        n19002), .Y(n21612) );
  A2O1A1Ixp33_ASAP7_75t_SL U22201 ( .A1(n21611), .A2(n21612), .B(n18295), .C(
        n19002), .Y(n21613) );
  A2O1A1Ixp33_ASAP7_75t_SL U22202 ( .A1(n19002), .A2(n21613), .B(n18295), .C(
        n19002), .Y(n2772) );
  A2O1A1Ixp33_ASAP7_75t_SL U22203 ( .A1(n24676), .A2(n21609), .B(n18295), .C(
        n19002), .Y(n21610) );
  A2O1A1Ixp33_ASAP7_75t_SL U22204 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__30_), .A2(
        n21606), .B(n18295), .C(n19002), .Y(n21607) );
  A2O1A1Ixp33_ASAP7_75t_SL U22205 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[34]), 
        .B(n18295), .C(n19002), .Y(n21603) );
  A2O1A1Ixp33_ASAP7_75t_SL U22206 ( .A1(n21602), .A2(n21603), .B(n18295), .C(
        n19002), .Y(n21604) );
  A2O1A1Ixp33_ASAP7_75t_SL U22207 ( .A1(n30524), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21335) );
  A2O1A1Ixp33_ASAP7_75t_SL U22208 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__13_), .A2(
        n21596), .B(n18295), .C(n19002), .Y(n21597) );
  A2O1A1Ixp33_ASAP7_75t_SL U22209 ( .A1(n30526), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21334) );
  A2O1A1Ixp33_ASAP7_75t_SL U22210 ( .A1(n30533), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21331) );
  A2O1A1Ixp33_ASAP7_75t_SL U22211 ( .A1(n24681), .A2(n27267), .B(n18295), .C(
        n19002), .Y(n21330) );
  A2O1A1Ixp33_ASAP7_75t_SL U22212 ( .A1(n31834), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21329) );
  A2O1A1Ixp33_ASAP7_75t_SL U22213 ( .A1(n24670), .A2(n28527), .B(n18295), .C(
        n19002), .Y(n21589) );
  A2O1A1Ixp33_ASAP7_75t_SL U22214 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__20_), .A2(
        n21586), .B(n18295), .C(n19002), .Y(n21587) );
  A2O1A1Ixp33_ASAP7_75t_SL U22215 ( .A1(n29043), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21328) );
  A2O1A1Ixp33_ASAP7_75t_SL U22216 ( .A1(n24681), .A2(n29081), .B(n18295), .C(
        n19002), .Y(n21327) );
  A2O1A1Ixp33_ASAP7_75t_SL U22217 ( .A1(n29040), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21326) );
  A2O1A1Ixp33_ASAP7_75t_SL U22218 ( .A1(n24681), .A2(n29768), .B(n18295), .C(
        n19002), .Y(n21325) );
  A2O1A1Ixp33_ASAP7_75t_SL U22219 ( .A1(n29773), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n21324) );
  A2O1A1Ixp33_ASAP7_75t_SL U22220 ( .A1(n27129), .A2(n24669), .B(n18295), .C(
        n19002), .Y(n20931) );
  A2O1A1Ixp33_ASAP7_75t_SL U22221 ( .A1(n28108), .A2(n27952), .B(n18295), .C(
        n19002), .Y(n21315) );
  A2O1A1Ixp33_ASAP7_75t_SL U22222 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__29_), .A2(
        n21581), .B(n18295), .C(n19002), .Y(n21582) );
  A2O1A1Ixp33_ASAP7_75t_SL U22223 ( .A1(n18295), .A2(n19002), .B(n21313), .C(
        n19002), .Y(n21314) );
  A2O1A1Ixp33_ASAP7_75t_SL U22224 ( .A1(n18295), .A2(n19002), .B(n21310), .C(
        n19002), .Y(n21311) );
  A2O1A1Ixp33_ASAP7_75t_SL U22225 ( .A1(n32660), .A2(n32657), .B(n18295), .C(
        n19002), .Y(n21580) );
  A2O1A1Ixp33_ASAP7_75t_SL U22226 ( .A1(n32660), .A2(n32637), .B(n18295), .C(
        n19002), .Y(n21579) );
  A2O1A1Ixp33_ASAP7_75t_SL U22227 ( .A1(n32660), .A2(n32635), .B(n18295), .C(
        n19002), .Y(n21578) );
  A2O1A1Ixp33_ASAP7_75t_SL U22228 ( .A1(n32660), .A2(n32633), .B(n18295), .C(
        n19002), .Y(n21577) );
  A2O1A1Ixp33_ASAP7_75t_SL U22229 ( .A1(n32660), .A2(n32625), .B(n18295), .C(
        n19002), .Y(n21576) );
  A2O1A1Ixp33_ASAP7_75t_SL U22230 ( .A1(n32599), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n21297) );
  A2O1A1Ixp33_ASAP7_75t_SL U22231 ( .A1(n32403), .A2(n21569), .B(n18295), .C(
        n19002), .Y(n21570) );
  A2O1A1Ixp33_ASAP7_75t_SL U22232 ( .A1(n32603), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n21571) );
  A2O1A1Ixp33_ASAP7_75t_SL U22233 ( .A1(n32318), .A2(dc_q[3]), .B(n18295), .C(
        n19002), .Y(n21572) );
  A2O1A1Ixp33_ASAP7_75t_SL U22234 ( .A1(n21570), .A2(n21571), .B(n18295), .C(
        n21572), .Y(dc_data[3]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22235 ( .A1(n23960), .A2(n28131), .B(n18295), .C(
        n19002), .Y(n21566) );
  A2O1A1Ixp33_ASAP7_75t_SL U22236 ( .A1(n29935), .A2(n21566), .B(n18295), .C(
        n19002), .Y(n21567) );
  A2O1A1Ixp33_ASAP7_75t_SL U22237 ( .A1(n29275), .A2(n21565), .B(n18295), .C(
        n19002), .Y(n29742) );
  A2O1A1Ixp33_ASAP7_75t_SL U22238 ( .A1(n24395), .A2(n24356), .B(n18295), .C(
        n19002), .Y(n21564) );
  A2O1A1Ixp33_ASAP7_75t_SL U22239 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[59]), 
        .B(n18295), .C(n19002), .Y(n21563) );
  A2O1A1Ixp33_ASAP7_75t_SL U22240 ( .A1(n31655), .A2(n21561), .B(n18295), .C(
        n21562), .Y(n31663) );
  A2O1A1Ixp33_ASAP7_75t_SL U22241 ( .A1(mult_x_1196_n591), .A2(n19002), .B(
        n18295), .C(n19002), .Y(n21277) );
  A2O1A1Ixp33_ASAP7_75t_SL U22242 ( .A1(n19002), .A2(n21278), .B(n18295), .C(
        n19002), .Y(mult_x_1196_n589) );
  A2O1A1Ixp33_ASAP7_75t_SL U22243 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[48]), 
        .B(n18295), .C(n19002), .Y(n21559) );
  A2O1A1Ixp33_ASAP7_75t_SL U22244 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[46]), 
        .B(n18295), .C(n19002), .Y(n21558) );
  A2O1A1Ixp33_ASAP7_75t_SL U22245 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__6_), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__5_), .B(n18295), .C(n19002), 
        .Y(n21555) );
  A2O1A1Ixp33_ASAP7_75t_SL U22246 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__0_), .A2(n31558), .B(n18295), 
        .C(n19002), .Y(n21556) );
  A2O1A1Ixp33_ASAP7_75t_SL U22247 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[53]), 
        .B(n18295), .C(n19002), .Y(n21554) );
  A2O1A1Ixp33_ASAP7_75t_SL U22248 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[55]), 
        .B(n18295), .C(n19002), .Y(n21553) );
  A2O1A1Ixp33_ASAP7_75t_SL U22249 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__3_), .B(n18295), .C(n19002), .Y(
        n21551) );
  A2O1A1Ixp33_ASAP7_75t_SL U22250 ( .A1(u0_0_leon3x0_p0_divi[62]), .A2(n22373), 
        .B(n18295), .C(n19002), .Y(n21261) );
  A2O1A1Ixp33_ASAP7_75t_SL U22251 ( .A1(n18295), .A2(n19002), .B(n20875), .C(
        n19002), .Y(n23224) );
  A2O1A1Ixp33_ASAP7_75t_SL U22252 ( .A1(mult_x_1196_n2225), .A2(
        mult_x_1196_n2535), .B(n18295), .C(n19002), .Y(n21542) );
  A2O1A1Ixp33_ASAP7_75t_SL U22253 ( .A1(n19002), .A2(n30783), .B(n18295), .C(
        n19002), .Y(n21476) );
  A2O1A1Ixp33_ASAP7_75t_SL U22254 ( .A1(uart1_r_RHOLD__24__4_), .A2(n21476), 
        .B(n18295), .C(n19002), .Y(n21477) );
  A2O1A1Ixp33_ASAP7_75t_SL U22255 ( .A1(n1630), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n21484) );
  A2O1A1Ixp33_ASAP7_75t_SL U22256 ( .A1(n31201), .A2(uart1_r_RHOLD__30__4_), 
        .B(n18295), .C(n19002), .Y(n21498) );
  A2O1A1Ixp33_ASAP7_75t_SL U22257 ( .A1(uart1_r_RHOLD__5__4_), .A2(n31200), 
        .B(n18295), .C(n19002), .Y(n21499) );
  A2O1A1Ixp33_ASAP7_75t_SL U22258 ( .A1(n31229), .A2(uart1_r_RHOLD__22__4_), 
        .B(n18295), .C(n19002), .Y(n21510) );
  A2O1A1Ixp33_ASAP7_75t_SL U22259 ( .A1(uart1_r_RHOLD__27__4_), .A2(n31230), 
        .B(n18295), .C(n19002), .Y(n21511) );
  A2O1A1Ixp33_ASAP7_75t_SL U22260 ( .A1(timer0_vtimers_1__IRQPEN_), .A2(n30790), .B(n18295), .C(n19002), .Y(n21519) );
  A2O1A1Ixp33_ASAP7_75t_SL U22261 ( .A1(uart1_r_BRATE__4_), .A2(n31246), .B(
        n18295), .C(n19002), .Y(n21521) );
  A2O1A1Ixp33_ASAP7_75t_SL U22262 ( .A1(timer0_r_RELOAD__4_), .A2(n31237), .B(
        n18295), .C(n19002), .Y(n21522) );
  A2O1A1Ixp33_ASAP7_75t_SL U22263 ( .A1(n19002), .A2(n31023), .B(n18295), .C(
        n19002), .Y(n21526) );
  A2O1A1Ixp33_ASAP7_75t_SL U22264 ( .A1(irqctrl0_r_IPEND__4_), .A2(n21526), 
        .B(n18295), .C(n19002), .Y(n21527) );
  A2O1A1Ixp33_ASAP7_75t_SL U22265 ( .A1(n21527), .A2(n21528), .B(n18295), .C(
        n19002), .Y(n21529) );
  A2O1A1Ixp33_ASAP7_75t_SL U22266 ( .A1(n21524), .A2(n21533), .B(n18295), .C(
        n19002), .Y(n21534) );
  A2O1A1Ixp33_ASAP7_75t_SL U22267 ( .A1(n21477), .A2(n21538), .B(n18295), .C(
        n19002), .Y(n21539) );
  A2O1A1Ixp33_ASAP7_75t_SL U22268 ( .A1(n29631), .A2(n20864), .B(n18295), .C(
        n19002), .Y(n20865) );
  A2O1A1Ixp33_ASAP7_75t_SL U22269 ( .A1(n31877), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[0]), .B(n18295), .C(
        u0_0_leon3x0_p0_c0mmu_icache0_r_BURST_), .Y(n21473) );
  A2O1A1Ixp33_ASAP7_75t_SL U22270 ( .A1(n32786), .A2(n31698), .B(n18295), .C(
        n19002), .Y(n21475) );
  A2O1A1Ixp33_ASAP7_75t_SL U22271 ( .A1(n31720), .A2(sr1_r_MCFG1__IOWS__3_), 
        .B(n18295), .C(n19002), .Y(n21468) );
  A2O1A1Ixp33_ASAP7_75t_SL U22272 ( .A1(n31725), .A2(sr1_r_MCFG1__ROMWWS__3_), 
        .B(n18295), .C(n19002), .Y(n21469) );
  A2O1A1Ixp33_ASAP7_75t_SL U22273 ( .A1(n31726), .A2(sr1_r_MCFG1__ROMRWS__3_), 
        .B(n18295), .C(n19002), .Y(n21470) );
  A2O1A1Ixp33_ASAP7_75t_SL U22274 ( .A1(n21468), .A2(n21469), .B(n18295), .C(
        n21470), .Y(n21471) );
  A2O1A1Ixp33_ASAP7_75t_SL U22275 ( .A1(uart1_r_TSHIFT__9_), .A2(n29951), .B(
        n18295), .C(n19002), .Y(n21464) );
  A2O1A1Ixp33_ASAP7_75t_SL U22276 ( .A1(uart1_r_TSHIFT__8_), .A2(n29954), .B(
        n18295), .C(n19002), .Y(n21465) );
  A2O1A1Ixp33_ASAP7_75t_SL U22277 ( .A1(n24663), .A2(n32626), .B(n18295), .C(
        n19002), .Y(n21462) );
  A2O1A1Ixp33_ASAP7_75t_SL U22278 ( .A1(n32577), .A2(n24662), .B(n18295), .C(
        n19002), .Y(n21235) );
  A2O1A1Ixp33_ASAP7_75t_SL U22279 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__25_), 
        .A2(n30641), .B(n18295), .C(n19002), .Y(n21450) );
  A2O1A1Ixp33_ASAP7_75t_SL U22280 ( .A1(rf_do_b[25]), .A2(n30640), .B(n18295), 
        .C(n19002), .Y(n21451) );
  A2O1A1Ixp33_ASAP7_75t_SL U22281 ( .A1(u0_0_leon3x0_p0_iu_r_W__RESULT__25_), 
        .A2(n29863), .B(n18295), .C(n19002), .Y(n21454) );
  A2O1A1Ixp33_ASAP7_75t_SL U22282 ( .A1(n29804), .A2(n21446), .B(n18295), .C(
        n19002), .Y(n21447) );
  A2O1A1Ixp33_ASAP7_75t_SL U22283 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[60]), 
        .B(n18295), .C(n19002), .Y(n21444) );
  A2O1A1Ixp33_ASAP7_75t_SL U22284 ( .A1(n21443), .A2(n21444), .B(n18295), .C(
        n19002), .Y(n21445) );
  A2O1A1Ixp33_ASAP7_75t_SL U22285 ( .A1(n26746), .A2(n24669), .B(n18295), .C(
        n19002), .Y(n21426) );
  A2O1A1Ixp33_ASAP7_75t_SL U22286 ( .A1(n30626), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n21427) );
  A2O1A1Ixp33_ASAP7_75t_SL U22287 ( .A1(n31415), .A2(n21427), .B(n18295), .C(
        n19002), .Y(n21428) );
  A2O1A1Ixp33_ASAP7_75t_SL U22288 ( .A1(n21428), .A2(n21432), .B(n18295), .C(
        n19002), .Y(n21433) );
  A2O1A1Ixp33_ASAP7_75t_SL U22289 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[42]), 
        .B(n18295), .C(n19002), .Y(n21424) );
  A2O1A1Ixp33_ASAP7_75t_SL U22290 ( .A1(n21423), .A2(n21424), .B(n18295), .C(
        n19002), .Y(n21425) );
  A2O1A1Ixp33_ASAP7_75t_SL U22291 ( .A1(n24670), .A2(n21419), .B(n18295), .C(
        n19002), .Y(n21420) );
  A2O1A1Ixp33_ASAP7_75t_SL U22292 ( .A1(mult_x_1196_n765), .A2(
        mult_x_1196_n766), .B(n18295), .C(n21415), .Y(n21416) );
  A2O1A1Ixp33_ASAP7_75t_SL U22293 ( .A1(n24673), .A2(n25284), .B(n18295), .C(
        n19002), .Y(n21414) );
  A2O1A1Ixp33_ASAP7_75t_SL U22294 ( .A1(n24666), .A2(n32138), .B(n18295), .C(
        n19002), .Y(n21412) );
  A2O1A1Ixp33_ASAP7_75t_SL U22295 ( .A1(n24648), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__6_), .B(n18295), .C(n19002), .Y(
        n20469) );
  A2O1A1Ixp33_ASAP7_75t_SL U22296 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[38]), 
        .B(n18295), .C(n19002), .Y(n21402) );
  A2O1A1Ixp33_ASAP7_75t_SL U22297 ( .A1(n21401), .A2(n21402), .B(n18295), .C(
        n19002), .Y(n21403) );
  A2O1A1Ixp33_ASAP7_75t_SL U22298 ( .A1(n24660), .A2(n20801), .B(n18295), .C(
        n19002), .Y(n20802) );
  A2O1A1Ixp33_ASAP7_75t_SL U22299 ( .A1(n24681), .A2(n29932), .B(n18295), .C(
        n19002), .Y(n21168) );
  A2O1A1Ixp33_ASAP7_75t_SL U22300 ( .A1(n30417), .A2(n24673), .B(n18295), .C(
        n19002), .Y(n20987) );
  A2O1A1Ixp33_ASAP7_75t_SL U22301 ( .A1(n30234), .A2(n24671), .B(n18295), .C(
        n19002), .Y(n21167) );
  A2O1A1Ixp33_ASAP7_75t_SL U22302 ( .A1(n18295), .A2(n19002), .B(n20090), .C(
        n19002), .Y(n20091) );
  A2O1A1Ixp33_ASAP7_75t_SL U22303 ( .A1(n20091), .A2(n20092), .B(n18295), .C(
        n19002), .Y(n3737) );
  A2O1A1Ixp33_ASAP7_75t_SL U22304 ( .A1(n24670), .A2(n21162), .B(n18295), .C(
        n19002), .Y(n21163) );
  A2O1A1Ixp33_ASAP7_75t_SL U22305 ( .A1(n22421), .A2(DP_OP_1196_128_7433_n455), 
        .B(n18295), .C(n19002), .Y(n21383) );
  A2O1A1Ixp33_ASAP7_75t_SL U22306 ( .A1(n21382), .A2(n21383), .B(n18295), .C(
        n19002), .Y(n21384) );
  A2O1A1Ixp33_ASAP7_75t_SL U22307 ( .A1(n19002), .A2(n21384), .B(n18295), .C(
        n19002), .Y(n3552) );
  A2O1A1Ixp33_ASAP7_75t_SL U22308 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA1__2_), 
        .A2(n24660), .B(n18295), .C(n19002), .Y(n21154) );
  A2O1A1Ixp33_ASAP7_75t_SL U22309 ( .A1(n22378), .A2(n20797), .B(n18295), .C(
        n19002), .Y(n20798) );
  A2O1A1Ixp33_ASAP7_75t_SL U22310 ( .A1(n24665), .A2(n21379), .B(n18295), .C(
        n19002), .Y(n21380) );
  A2O1A1Ixp33_ASAP7_75t_SL U22311 ( .A1(n29736), .A2(n29737), .B(n18295), .C(
        n19002), .Y(n20794) );
  A2O1A1Ixp33_ASAP7_75t_SL U22312 ( .A1(n24677), .A2(n21370), .B(n18295), .C(
        n19002), .Y(n21371) );
  A2O1A1Ixp33_ASAP7_75t_SL U22313 ( .A1(n28585), .A2(n22378), .B(n18295), .C(
        n19002), .Y(n20619) );
  A2O1A1Ixp33_ASAP7_75t_SL U22314 ( .A1(n32677), .A2(n18830), .B(n18295), .C(
        n19002), .Y(n21145) );
  A2O1A1Ixp33_ASAP7_75t_SL U22315 ( .A1(n31596), .A2(n31584), .B(n18295), .C(
        n21362), .Y(n21363) );
  A2O1A1Ixp33_ASAP7_75t_SL U22316 ( .A1(n31588), .A2(n21363), .B(n18295), .C(
        n21364), .Y(n18101) );
  A2O1A1Ixp33_ASAP7_75t_SL U22317 ( .A1(n22396), .A2(n21360), .B(n18295), .C(
        n19002), .Y(n21361) );
  A2O1A1Ixp33_ASAP7_75t_SL U22318 ( .A1(n30182), .A2(n21354), .B(n18295), .C(
        n19002), .Y(n21355) );
  A2O1A1Ixp33_ASAP7_75t_SL U22319 ( .A1(n21356), .A2(n21357), .B(n18295), .C(
        n19002), .Y(n21358) );
  A2O1A1Ixp33_ASAP7_75t_SL U22320 ( .A1(n21355), .A2(n21358), .B(n18295), .C(
        n19002), .Y(u0_0_leon3x0_p0_c0mmu_dcache0_v_FADDR__6_) );
  A2O1A1Ixp33_ASAP7_75t_SL U22321 ( .A1(n28952), .A2(n24676), .B(n18295), .C(
        n19002), .Y(n21137) );
  A2O1A1Ixp33_ASAP7_75t_SL U22322 ( .A1(n19002), .A2(n21350), .B(n18295), .C(
        n19002), .Y(n32548) );
  A2O1A1Ixp33_ASAP7_75t_SL U22323 ( .A1(n28042), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n21346) );
  A2O1A1Ixp33_ASAP7_75t_SL U22324 ( .A1(n24694), .A2(n21346), .B(n18295), .C(
        n19002), .Y(n21347) );
  A2O1A1Ixp33_ASAP7_75t_SL U22325 ( .A1(n29374), .A2(n21347), .B(n18295), .C(
        n19002), .Y(n21348) );
  A2O1A1Ixp33_ASAP7_75t_SL U22326 ( .A1(n31021), .A2(n31840), .B(n18295), .C(
        n19002), .Y(n20776) );
  A2O1A1Ixp33_ASAP7_75t_SL U22327 ( .A1(u0_0_leon3x0_p0_muli[3]), .A2(n21340), 
        .B(n18295), .C(n19002), .Y(n21341) );
  A2O1A1Ixp33_ASAP7_75t_SL U22328 ( .A1(n30429), .A2(n24661), .B(n18295), .C(
        n19002), .Y(n20771) );
  A2O1A1Ixp33_ASAP7_75t_SL U22329 ( .A1(n24681), .A2(n27172), .B(n18295), .C(
        n19002), .Y(n21095) );
  A2O1A1Ixp33_ASAP7_75t_SL U22330 ( .A1(n21094), .A2(n29350), .B(n18295), .C(
        n19002), .Y(n1761) );
  A2O1A1Ixp33_ASAP7_75t_SL U22331 ( .A1(n32583), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__4_), .B(n18295), .C(n19002), 
        .Y(n21303) );
  A2O1A1Ixp33_ASAP7_75t_SL U22332 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__9_), 
        .A2(n32584), .B(n18295), .C(n19002), .Y(n21304) );
  A2O1A1Ixp33_ASAP7_75t_SL U22333 ( .A1(n21303), .A2(n21304), .B(n18295), .C(
        n19002), .Y(n21305) );
  A2O1A1Ixp33_ASAP7_75t_SL U22334 ( .A1(n32581), .A2(n32588), .B(n18295), .C(
        n19002), .Y(n21307) );
  A2O1A1Ixp33_ASAP7_75t_SL U22335 ( .A1(n21306), .A2(n21307), .B(n18295), .C(
        n19002), .Y(ic_address[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22336 ( .A1(n32660), .A2(n32655), .B(n18295), .C(
        n19002), .Y(n21301) );
  A2O1A1Ixp33_ASAP7_75t_SL U22337 ( .A1(n32660), .A2(n32643), .B(n18295), .C(
        n19002), .Y(n21300) );
  A2O1A1Ixp33_ASAP7_75t_SL U22338 ( .A1(n32660), .A2(n32639), .B(n18295), .C(
        n19002), .Y(n21299) );
  A2O1A1Ixp33_ASAP7_75t_SL U22339 ( .A1(n32660), .A2(n32627), .B(n18295), .C(
        n19002), .Y(n21298) );
  A2O1A1Ixp33_ASAP7_75t_SL U22340 ( .A1(n32619), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n20921) );
  A2O1A1Ixp33_ASAP7_75t_SL U22341 ( .A1(n32600), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n20046) );
  A2O1A1Ixp33_ASAP7_75t_SL U22342 ( .A1(n32653), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n21292) );
  A2O1A1Ixp33_ASAP7_75t_SL U22343 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__6_), 
        .A2(n30723), .B(n18295), .C(n19002), .Y(n20563) );
  A2O1A1Ixp33_ASAP7_75t_SL U22344 ( .A1(n28805), .A2(n32162), .B(n18295), .C(
        n19002), .Y(n20564) );
  A2O1A1Ixp33_ASAP7_75t_SL U22345 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__6_), 
        .A2(n30726), .B(n18295), .C(n19002), .Y(n20565) );
  A2O1A1Ixp33_ASAP7_75t_SL U22346 ( .A1(u0_0_leon3x0_p0_ici[3]), .A2(n30722), 
        .B(n18295), .C(n19002), .Y(n20566) );
  A2O1A1Ixp33_ASAP7_75t_SL U22347 ( .A1(n20564), .A2(n20565), .B(n18295), .C(
        n20566), .Y(n20567) );
  A2O1A1Ixp33_ASAP7_75t_SL U22348 ( .A1(u0_0_leon3x0_p0_ici[34]), .A2(n30724), 
        .B(n18295), .C(n19002), .Y(n20569) );
  A2O1A1Ixp33_ASAP7_75t_SL U22349 ( .A1(n20563), .A2(n20568), .B(n18295), .C(
        n20569), .Y(rf_di_w[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22350 ( .A1(n31392), .A2(
        u0_0_leon3x0_p0_iu_r_W__RESULT__30_), .B(n18295), .C(n19002), .Y(
        n21287) );
  A2O1A1Ixp33_ASAP7_75t_SL U22351 ( .A1(rf_do_a[30]), .A2(n31391), .B(n18295), 
        .C(n19002), .Y(n21288) );
  A2O1A1Ixp33_ASAP7_75t_SL U22352 ( .A1(n21287), .A2(n21288), .B(n18295), .C(
        n19002), .Y(n21289) );
  A2O1A1Ixp33_ASAP7_75t_SL U22353 ( .A1(n24393), .A2(n24361), .B(n18295), .C(
        n19002), .Y(n21285) );
  A2O1A1Ixp33_ASAP7_75t_SL U22354 ( .A1(n18580), .A2(n21277), .B(n18295), .C(
        n19002), .Y(n21278) );
  A2O1A1Ixp33_ASAP7_75t_SL U22355 ( .A1(n24600), .A2(n24587), .B(n18295), .C(
        n19002), .Y(n19235) );
  A2O1A1Ixp33_ASAP7_75t_SL U22356 ( .A1(n24600), .A2(n24587), .B(n18295), .C(
        n19002), .Y(n19238) );
  A2O1A1Ixp33_ASAP7_75t_SL U22357 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[35]), 
        .B(n18295), .C(n19002), .Y(n21267) );
  A2O1A1Ixp33_ASAP7_75t_SL U22358 ( .A1(n31537), .A2(n24987), .B(n18295), .C(
        n19002), .Y(n20184) );
  A2O1A1Ixp33_ASAP7_75t_SL U22359 ( .A1(n31737), .A2(n32801), .B(n18295), .C(
        n19002), .Y(n21266) );
  A2O1A1Ixp33_ASAP7_75t_SL U22360 ( .A1(n32917), .A2(n21265), .B(n18295), .C(
        n19002), .Y(n32979) );
  A2O1A1Ixp33_ASAP7_75t_SL U22361 ( .A1(mult_x_1196_n391), .A2(
        mult_x_1196_n787), .B(n18295), .C(n23769), .Y(n21262) );
  A2O1A1Ixp33_ASAP7_75t_SL U22362 ( .A1(n21252), .A2(n21253), .B(n18295), .C(
        n19002), .Y(n21255) );
  A2O1A1Ixp33_ASAP7_75t_SL U22363 ( .A1(n21254), .A2(n21255), .B(n18295), .C(
        n19002), .Y(mult_x_1196_n849) );
  A2O1A1Ixp33_ASAP7_75t_SL U22364 ( .A1(n22408), .A2(n21241), .B(n18295), .C(
        n19002), .Y(n21242) );
  A2O1A1Ixp33_ASAP7_75t_SL U22365 ( .A1(n31213), .A2(n27496), .B(n18295), .C(
        n19002), .Y(n21041) );
  A2O1A1Ixp33_ASAP7_75t_SL U22366 ( .A1(n21038), .A2(n21039), .B(n18295), .C(
        n19002), .Y(n21040) );
  A2O1A1Ixp33_ASAP7_75t_SL U22367 ( .A1(n25600), .A2(n31806), .B(n18295), .C(
        n21238), .Y(n4649) );
  A2O1A1Ixp33_ASAP7_75t_SL U22368 ( .A1(n20686), .A2(n20688), .B(n18295), .C(
        n19002), .Y(n4648) );
  A2O1A1Ixp33_ASAP7_75t_SL U22369 ( .A1(n30640), .A2(rf_do_b[26]), .B(n18295), 
        .C(n19002), .Y(n21226) );
  A2O1A1Ixp33_ASAP7_75t_SL U22370 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__26_), .B(n18295), .C(n19002), .Y(n21227)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22371 ( .A1(n21226), .A2(n21227), .B(n18295), .C(
        n19002), .Y(n21228) );
  A2O1A1Ixp33_ASAP7_75t_SL U22372 ( .A1(n28802), .A2(n21231), .B(n18295), .C(
        n19002), .Y(n21232) );
  A2O1A1Ixp33_ASAP7_75t_SL U22373 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[56]), 
        .B(n18295), .C(n19002), .Y(n21222) );
  A2O1A1Ixp33_ASAP7_75t_SL U22374 ( .A1(n21221), .A2(n21222), .B(n18295), .C(
        n19002), .Y(n21223) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U22375 ( .A1(n29614), .A2(n29615), .B(n18295), 
        .C(n31054), .D(n21217), .Y(n21218) );
  A2O1A1Ixp33_ASAP7_75t_SL U22376 ( .A1(n31542), .A2(n28279), .B(n18295), .C(
        n19002), .Y(n21219) );
  A2O1A1Ixp33_ASAP7_75t_SL U22377 ( .A1(n21219), .A2(n21218), .B(n18295), .C(
        n19002), .Y(n4587) );
  A2O1A1Ixp33_ASAP7_75t_SL U22378 ( .A1(u0_0_leon3x0_p0_divi[43]), .A2(n30430), 
        .B(n18295), .C(n19002), .Y(n21205) );
  A2O1A1Ixp33_ASAP7_75t_SL U22379 ( .A1(n21204), .A2(n21205), .B(n18295), .C(
        n19002), .Y(n21206) );
  A2O1A1Ixp33_ASAP7_75t_SL U22380 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[46]), 
        .B(n18295), .C(n19002), .Y(n21201) );
  A2O1A1Ixp33_ASAP7_75t_SL U22381 ( .A1(n21200), .A2(n21201), .B(n18295), .C(
        n19002), .Y(n21202) );
  A2O1A1Ixp33_ASAP7_75t_SL U22382 ( .A1(n18295), .A2(n19002), .B(n21005), .C(
        n19002), .Y(n21006) );
  A2O1A1Ixp33_ASAP7_75t_SL U22383 ( .A1(n24668), .A2(n26752), .B(n18295), .C(
        n19002), .Y(n21191) );
  A2O1A1Ixp33_ASAP7_75t_SL U22384 ( .A1(n24673), .A2(n25285), .B(n18295), .C(
        n19002), .Y(n21188) );
  A2O1A1Ixp33_ASAP7_75t_SL U22385 ( .A1(n24661), .A2(n21186), .B(n18295), .C(
        n19002), .Y(n21187) );
  A2O1A1Ixp33_ASAP7_75t_SL U22386 ( .A1(n32624), .A2(n24669), .B(n18295), .C(
        n19002), .Y(n21000) );
  A2O1A1Ixp33_ASAP7_75t_SL U22387 ( .A1(n24664), .A2(n20471), .B(n18295), .C(
        n19002), .Y(n20472) );
  A2O1A1Ixp33_ASAP7_75t_SL U22388 ( .A1(n31352), .A2(n31451), .B(n18295), .C(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DFRZ_), .Y(n21181) );
  A2O1A1Ixp33_ASAP7_75t_SL U22389 ( .A1(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DCS__1_), .A2(n21181), .B(n18295), 
        .C(n19002), .Y(n21182) );
  A2O1A1Ixp33_ASAP7_75t_SL U22390 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[33]), 
        .B(n18295), .C(n19002), .Y(n21173) );
  A2O1A1Ixp33_ASAP7_75t_SL U22391 ( .A1(n21172), .A2(n21173), .B(n18295), .C(
        n19002), .Y(n21174) );
  A2O1A1Ixp33_ASAP7_75t_SL U22392 ( .A1(n24674), .A2(n20810), .B(n18295), .C(
        n19002), .Y(n20811) );
  A2O1A1Ixp33_ASAP7_75t_SL U22393 ( .A1(n24681), .A2(n30496), .B(n18295), .C(
        n19002), .Y(n20988) );
  A2O1A1Ixp33_ASAP7_75t_SL U22394 ( .A1(u0_0_leon3x0_p0_div0_r_CNT__3_), .A2(
        n24904), .B(n18295), .C(n19002), .Y(n21164) );
  A2O1A1Ixp33_ASAP7_75t_SL U22395 ( .A1(n30817), .A2(n24663), .B(n18295), .C(
        n19002), .Y(n19521) );
  A2O1A1Ixp33_ASAP7_75t_SL U22396 ( .A1(n30818), .A2(n31872), .B(n18295), .C(
        n19002), .Y(n19522) );
  A2O1A1Ixp33_ASAP7_75t_SL U22397 ( .A1(n23229), .A2(n32171), .B(n18295), .C(
        n19002), .Y(n21158) );
  A2O1A1Ixp33_ASAP7_75t_SL U22398 ( .A1(n21157), .A2(n21158), .B(n18295), .C(
        n19002), .Y(n21159) );
  A2O1A1Ixp33_ASAP7_75t_SL U22399 ( .A1(n19002), .A2(n21159), .B(n18295), .C(
        n19002), .Y(n3550) );
  A2O1A1Ixp33_ASAP7_75t_SL U22400 ( .A1(n24671), .A2(n19517), .B(n18295), .C(
        n19002), .Y(n19518) );
  A2O1A1Ixp33_ASAP7_75t_SL U22401 ( .A1(n22421), .A2(n32178), .B(n18295), .C(
        n19002), .Y(n21155) );
  A2O1A1Ixp33_ASAP7_75t_SL U22402 ( .A1(n21154), .A2(n21155), .B(n18295), .C(
        n19002), .Y(n21156) );
  A2O1A1Ixp33_ASAP7_75t_SL U22403 ( .A1(n19002), .A2(n21156), .B(n18295), .C(
        n19002), .Y(n3501) );
  A2O1A1Ixp33_ASAP7_75t_SL U22404 ( .A1(n24677), .A2(n21152), .B(n18295), .C(
        n19002), .Y(n21153) );
  A2O1A1Ixp33_ASAP7_75t_SL U22405 ( .A1(n32567), .A2(n18829), .B(n18295), .C(
        n19002), .Y(n20979) );
  A2O1A1Ixp33_ASAP7_75t_SL U22406 ( .A1(n22378), .A2(n19871), .B(n18295), .C(
        n19002), .Y(n19872) );
  A2O1A1Ixp33_ASAP7_75t_SL U22407 ( .A1(n24677), .A2(n21150), .B(n18295), .C(
        n19002), .Y(n21151) );
  A2O1A1Ixp33_ASAP7_75t_SL U22408 ( .A1(n24663), .A2(n21148), .B(n18295), .C(
        n19002), .Y(n21149) );
  A2O1A1Ixp33_ASAP7_75t_SL U22409 ( .A1(n24677), .A2(n21146), .B(n18295), .C(
        n19002), .Y(n21147) );
  A2O1A1Ixp33_ASAP7_75t_SL U22410 ( .A1(n22396), .A2(n21138), .B(n18295), .C(
        n19002), .Y(n21139) );
  A2O1A1Ixp33_ASAP7_75t_SL U22411 ( .A1(uart1_r_BRATE__8_), .A2(n21125), .B(
        n18295), .C(n19002), .Y(n21126) );
  A2O1A1Ixp33_ASAP7_75t_SL U22412 ( .A1(n30780), .A2(n24633), .B(n18295), .C(
        n19002), .Y(n20941) );
  A2O1A1Ixp33_ASAP7_75t_SL U22413 ( .A1(n29383), .A2(n21118), .B(n18295), .C(
        n19002), .Y(n21119) );
  A2O1A1Ixp33_ASAP7_75t_SL U22414 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__31_), .A2(
        n21115), .B(n18295), .C(n19002), .Y(n21116) );
  A2O1A1Ixp33_ASAP7_75t_SL U22415 ( .A1(n22420), .A2(n31422), .B(n18295), .C(
        n19002), .Y(n20057) );
  A2O1A1Ixp33_ASAP7_75t_SL U22416 ( .A1(n20058), .A2(n20059), .B(n18295), .C(
        n19002), .Y(n20060) );
  A2O1A1Ixp33_ASAP7_75t_SL U22417 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[35]), 
        .B(n18295), .C(n19002), .Y(n21113) );
  A2O1A1Ixp33_ASAP7_75t_SL U22418 ( .A1(n21112), .A2(n21113), .B(n18295), .C(
        n19002), .Y(n21114) );
  A2O1A1Ixp33_ASAP7_75t_SL U22419 ( .A1(n24677), .A2(n21107), .B(n18295), .C(
        n19002), .Y(n21108) );
  A2O1A1Ixp33_ASAP7_75t_SL U22420 ( .A1(n28552), .A2(n22427), .B(n18295), .C(
        n19002), .Y(n20937) );
  A2O1A1Ixp33_ASAP7_75t_SL U22421 ( .A1(n27279), .A2(n22427), .B(n18295), .C(
        n19002), .Y(n20936) );
  A2O1A1Ixp33_ASAP7_75t_SL U22422 ( .A1(n24681), .A2(n27030), .B(n18295), .C(
        n19002), .Y(n20935) );
  A2O1A1Ixp33_ASAP7_75t_SL U22423 ( .A1(n24678), .A2(n21099), .B(n18295), .C(
        n19002), .Y(n21100) );
  A2O1A1Ixp33_ASAP7_75t_SL U22424 ( .A1(n29782), .A2(n24667), .B(n18295), .C(
        n19002), .Y(n20932) );
  A2O1A1Ixp33_ASAP7_75t_SL U22425 ( .A1(ahb0_r_HADDR__10_), .A2(
        ahb0_r_HADDR__8_), .B(n18295), .C(n19002), .Y(n20595) );
  A2O1A1Ixp33_ASAP7_75t_SL U22426 ( .A1(ahb0_r_HADDR__7_), .A2(
        ahb0_r_HADDR__6_), .B(n18295), .C(n19002), .Y(n20596) );
  A2O1A1Ixp33_ASAP7_75t_SL U22427 ( .A1(n28108), .A2(n27926), .B(n18295), .C(
        n19002), .Y(n19849) );
  A2O1A1Ixp33_ASAP7_75t_SL U22428 ( .A1(n28108), .A2(n27948), .B(n18295), .C(
        n19002), .Y(n19848) );
  A2O1A1Ixp33_ASAP7_75t_SL U22429 ( .A1(n18295), .A2(n19002), .B(n20924), .C(
        n19002), .Y(n20925) );
  A2O1A1Ixp33_ASAP7_75t_SL U22430 ( .A1(n18295), .A2(n19002), .B(n20758), .C(
        n19002), .Y(n20759) );
  A2O1A1Ixp33_ASAP7_75t_SL U22431 ( .A1(n24420), .A2(n24389), .B(n18295), .C(
        n21090), .Y(n21091) );
  A2O1A1Ixp33_ASAP7_75t_SL U22432 ( .A1(n24389), .A2(n24420), .B(n18295), .C(
        n19002), .Y(n21092) );
  A2O1A1Ixp33_ASAP7_75t_SL U22433 ( .A1(n32583), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__2_), .B(n18295), .C(n19002), 
        .Y(n21085) );
  A2O1A1Ixp33_ASAP7_75t_SL U22434 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__7_), 
        .A2(n32584), .B(n18295), .C(n19002), .Y(n21086) );
  A2O1A1Ixp33_ASAP7_75t_SL U22435 ( .A1(n21085), .A2(n21086), .B(n18295), .C(
        n19002), .Y(n21087) );
  A2O1A1Ixp33_ASAP7_75t_SL U22436 ( .A1(n32575), .A2(n32588), .B(n18295), .C(
        n19002), .Y(n21089) );
  A2O1A1Ixp33_ASAP7_75t_SL U22437 ( .A1(n21088), .A2(n21089), .B(n18295), .C(
        n19002), .Y(ic_address[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22438 ( .A1(n32660), .A2(n32641), .B(n18295), .C(
        n19002), .Y(n21083) );
  A2O1A1Ixp33_ASAP7_75t_SL U22439 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__9_), 
        .A2(n32447), .B(n18295), .C(n19002), .Y(n19475) );
  A2O1A1Ixp33_ASAP7_75t_SL U22440 ( .A1(n32446), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[42]), .B(n18295), .C(n19002), .Y(n19476) );
  A2O1A1Ixp33_ASAP7_75t_SL U22441 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[9]), .A2(
        n32448), .B(n18295), .C(n19002), .Y(n19477) );
  A2O1A1Ixp33_ASAP7_75t_SL U22442 ( .A1(n19475), .A2(n19476), .B(n18295), .C(
        n19477), .Y(n19478) );
  A2O1A1Ixp33_ASAP7_75t_SL U22443 ( .A1(n33067), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__4_), .B(n18295), .C(n19002), 
        .Y(n19480) );
  A2O1A1Ixp33_ASAP7_75t_SL U22444 ( .A1(n18295), .A2(n19002), .B(n20574), .C(
        n19002), .Y(n20575) );
  A2O1A1Ixp33_ASAP7_75t_SL U22445 ( .A1(n20575), .A2(n20581), .B(n18295), .C(
        n19002), .Y(dc_data[31]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22446 ( .A1(n32215), .A2(n32234), .B(n18295), .C(
        n19002), .Y(n20741) );
  A2O1A1Ixp33_ASAP7_75t_SL U22447 ( .A1(n24622), .A2(n24621), .B(n18295), .C(
        n19002), .Y(n21082) );
  A2O1A1Ixp33_ASAP7_75t_SL U22448 ( .A1(n29629), .A2(n21081), .B(n18295), .C(
        n19002), .Y(n29662) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U22449 ( .A1(n29504), .A2(n30007), .B(n18295), 
        .C(n29505), .D(n29503), .Y(n21080) );
  A2O1A1Ixp33_ASAP7_75t_SL U22450 ( .A1(n31392), .A2(
        u0_0_leon3x0_p0_iu_r_W__RESULT__23_), .B(n18295), .C(n19002), .Y(
        n21076) );
  A2O1A1Ixp33_ASAP7_75t_SL U22451 ( .A1(rf_do_a[23]), .A2(n31391), .B(n18295), 
        .C(n19002), .Y(n21077) );
  A2O1A1Ixp33_ASAP7_75t_SL U22452 ( .A1(n21076), .A2(n21077), .B(n18295), .C(
        n19002), .Y(n21078) );
  A2O1A1Ixp33_ASAP7_75t_SL U22453 ( .A1(n24397), .A2(n24351), .B(n18295), .C(
        n19002), .Y(n21069) );
  A2O1A1Ixp33_ASAP7_75t_SL U22454 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[58]), 
        .B(n18295), .C(n19002), .Y(n21068) );
  A2O1A1Ixp33_ASAP7_75t_SL U22455 ( .A1(n31392), .A2(
        u0_0_leon3x0_p0_iu_r_W__RESULT__18_), .B(n18295), .C(n19002), .Y(
        n21065) );
  A2O1A1Ixp33_ASAP7_75t_SL U22456 ( .A1(rf_do_a[18]), .A2(n31391), .B(n18295), 
        .C(n19002), .Y(n21066) );
  A2O1A1Ixp33_ASAP7_75t_SL U22457 ( .A1(n21065), .A2(n21066), .B(n18295), .C(
        n19002), .Y(n21067) );
  A2O1A1Ixp33_ASAP7_75t_SL U22458 ( .A1(add_x_746_n12), .A2(
        u0_0_leon3x0_p0_iu_fe_pc_30_), .B(n18295), .C(n19002), .Y(n21063) );
  A2O1A1Ixp33_ASAP7_75t_SL U22459 ( .A1(n25307), .A2(n24672), .B(n18295), .C(
        n19002), .Y(n21061) );
  A2O1A1Ixp33_ASAP7_75t_SL U22460 ( .A1(mult_x_1196_n348), .A2(n21060), .B(
        n18295), .C(n19002), .Y(mult_x_1196_n230) );
  A2O1A1Ixp33_ASAP7_75t_SL U22461 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[47]), 
        .B(n18295), .C(n19002), .Y(n21058) );
  A2O1A1Ixp33_ASAP7_75t_SL U22462 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[45]), 
        .B(n18295), .C(n19002), .Y(n21057) );
  A2O1A1Ixp33_ASAP7_75t_SL U22463 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[36]), 
        .B(n18295), .C(n19002), .Y(n21055) );
  A2O1A1Ixp33_ASAP7_75t_SL U22464 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__9_), 
        .A2(n29060), .B(n18295), .C(n19002), .Y(n20523) );
  A2O1A1Ixp33_ASAP7_75t_SL U22465 ( .A1(n18532), .A2(
        u0_0_leon3x0_p0_iu_r_E__SHCNT__4_), .B(n18295), .C(n19002), .Y(n21050)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22466 ( .A1(n21050), .A2(n28820), .B(n18295), .C(
        n19002), .Y(n26139) );
  A2O1A1Ixp33_ASAP7_75t_SL U22467 ( .A1(n29881), .A2(irqi_0__IRL__0_), .B(
        n18295), .C(n19002), .Y(n21045) );
  A2O1A1Ixp33_ASAP7_75t_SL U22468 ( .A1(n24649), .A2(
        u0_0_leon3x0_p0_iu_r_X__CTRL__TT__0_), .B(n18295), .C(n19002), .Y(
        n21046) );
  A2O1A1Ixp33_ASAP7_75t_SL U22469 ( .A1(n29642), .A2(n21045), .B(n18295), .C(
        n21046), .Y(n21047) );
  O2A1O1Ixp33_ASAP7_75t_SL U22470 ( .A1(n18295), .A2(n20851), .B(n19002), .C(
        n20852), .Y(n20853) );
  A2O1A1Ixp33_ASAP7_75t_SL U22471 ( .A1(sr1_r_MCFG1__ROMRWS__1_), .A2(n31726), 
        .B(n18295), .C(n19002), .Y(n20856) );
  A2O1A1Ixp33_ASAP7_75t_SL U22472 ( .A1(uart1_r_TSHIFT__7_), .A2(n29951), .B(
        n18295), .C(n19002), .Y(n21038) );
  A2O1A1Ixp33_ASAP7_75t_SL U22473 ( .A1(uart1_r_TSHIFT__6_), .A2(n29954), .B(
        n18295), .C(n19002), .Y(n21039) );
  A2O1A1Ixp33_ASAP7_75t_SL U22474 ( .A1(u0_0_leon3x0_p0_divi[57]), .A2(n30430), 
        .B(n18295), .C(n19002), .Y(n21030) );
  A2O1A1Ixp33_ASAP7_75t_SL U22475 ( .A1(n21029), .A2(n21030), .B(n18295), .C(
        n19002), .Y(n21031) );
  A2O1A1Ixp33_ASAP7_75t_SL U22476 ( .A1(n30640), .A2(rf_do_b[28]), .B(n18295), 
        .C(n19002), .Y(n21019) );
  A2O1A1Ixp33_ASAP7_75t_SL U22477 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__28_), .B(n18295), .C(n19002), .Y(n21020)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22478 ( .A1(n21019), .A2(n21020), .B(n18295), .C(
        n19002), .Y(n21021) );
  A2O1A1Ixp33_ASAP7_75t_SL U22479 ( .A1(n23833), .A2(n22427), .B(n18295), .C(
        n19002), .Y(n21026) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U22480 ( .A1(n29614), .A2(n29615), .B(n18295), 
        .C(n31542), .D(n21015), .Y(n21016) );
  A2O1A1Ixp33_ASAP7_75t_SL U22481 ( .A1(n30600), .A2(n30599), .B(n18295), .C(
        n31054), .Y(n21017) );
  A2O1A1Ixp33_ASAP7_75t_SL U22482 ( .A1(n21016), .A2(n21017), .B(n18295), .C(
        n19002), .Y(n4583) );
  A2O1A1Ixp33_ASAP7_75t_SL U22483 ( .A1(n24669), .A2(n32580), .B(n18295), .C(
        n19002), .Y(n21014) );
  A2O1A1Ixp33_ASAP7_75t_SL U22484 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[54]), 
        .B(n18295), .C(n19002), .Y(n21009) );
  A2O1A1Ixp33_ASAP7_75t_SL U22485 ( .A1(n21008), .A2(n21009), .B(n18295), .C(
        n19002), .Y(n21010) );
  A2O1A1Ixp33_ASAP7_75t_SL U22486 ( .A1(n24684), .A2(n24666), .B(n18295), .C(
        n19002), .Y(n21002) );
  A2O1A1Ixp33_ASAP7_75t_SL U22487 ( .A1(n24675), .A2(n29106), .B(n18295), .C(
        n19002), .Y(n20655) );
  A2O1A1Ixp33_ASAP7_75t_SL U22488 ( .A1(n24663), .A2(n20996), .B(n18295), .C(
        n19002), .Y(n20997) );
  A2O1A1Ixp33_ASAP7_75t_SL U22489 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[43]), 
        .B(n18295), .C(n19002), .Y(n20994) );
  A2O1A1Ixp33_ASAP7_75t_SL U22490 ( .A1(n20993), .A2(n20994), .B(n18295), .C(
        n19002), .Y(n20995) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U22491 ( .A1(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__IFRZ_), .A2(n31352), .B(n18295), 
        .C(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__0_), .D(n32461), .Y(n20989)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22492 ( .A1(n32120), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[1]), .B(n18295), .C(n19002), .Y(n20990)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22493 ( .A1(n32124), .A2(n32127), .B(n18295), .C(
        n19002), .Y(n20805) );
  A2O1A1Ixp33_ASAP7_75t_SL U22494 ( .A1(n24684), .A2(n32676), .B(n18295), .C(
        u0_0_leon3x0_p0_c0mmu_icache0_r_UNDERRUN_), .Y(n20806) );
  A2O1A1Ixp33_ASAP7_75t_SL U22495 ( .A1(n20804), .A2(n20807), .B(n18295), .C(
        n19002), .Y(n3895) );
  A2O1A1Ixp33_ASAP7_75t_SL U22496 ( .A1(n26755), .A2(n24671), .B(n18295), .C(
        n19002), .Y(n20803) );
  A2O1A1Ixp33_ASAP7_75t_SL U22497 ( .A1(n30407), .A2(n24677), .B(n18295), .C(
        n19002), .Y(n20800) );
  A2O1A1Ixp33_ASAP7_75t_SL U22498 ( .A1(n24681), .A2(n30385), .B(n18295), .C(
        n19002), .Y(n20799) );
  A2O1A1Ixp33_ASAP7_75t_SL U22499 ( .A1(n24674), .A2(n20984), .B(n18295), .C(
        n19002), .Y(n20985) );
  A2O1A1Ixp33_ASAP7_75t_SL U22500 ( .A1(n24665), .A2(n20453), .B(n18295), .C(
        n19002), .Y(n20454) );
  A2O1A1Ixp33_ASAP7_75t_SL U22501 ( .A1(n24675), .A2(n20980), .B(n18295), .C(
        n19002), .Y(n20981) );
  A2O1A1Ixp33_ASAP7_75t_SL U22502 ( .A1(n24665), .A2(n20977), .B(n18295), .C(
        n19002), .Y(n20978) );
  A2O1A1Ixp33_ASAP7_75t_SL U22503 ( .A1(n24677), .A2(n20974), .B(n18295), .C(
        n19002), .Y(n20975) );
  A2O1A1Ixp33_ASAP7_75t_SL U22504 ( .A1(n24678), .A2(n20972), .B(n18295), .C(
        n19002), .Y(n20973) );
  A2O1A1Ixp33_ASAP7_75t_SL U22505 ( .A1(n24666), .A2(n20968), .B(n18295), .C(
        n19002), .Y(n20969) );
  A2O1A1Ixp33_ASAP7_75t_SL U22506 ( .A1(n32140), .A2(n20965), .B(n18295), .C(
        n19002), .Y(n20966) );
  A2O1A1Ixp33_ASAP7_75t_SL U22507 ( .A1(n31945), .A2(n20960), .B(n18295), .C(
        n19002), .Y(n20961) );
  A2O1A1Ixp33_ASAP7_75t_SL U22508 ( .A1(n24677), .A2(n20958), .B(n18295), .C(
        n19002), .Y(n20959) );
  A2O1A1Ixp33_ASAP7_75t_SL U22509 ( .A1(u0_0_leon3x0_p0_muli[7]), .A2(n20615), 
        .B(n18295), .C(n19002), .Y(n20616) );
  A2O1A1Ixp33_ASAP7_75t_SL U22510 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__8_), .A2(
        n20953), .B(n18295), .C(n19002), .Y(n20954) );
  A2O1A1Ixp33_ASAP7_75t_SL U22511 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__21_), .A2(
        n20948), .B(n18295), .C(n19002), .Y(n20949) );
  A2O1A1Ixp33_ASAP7_75t_SL U22512 ( .A1(n31198), .A2(n30978), .B(n18295), .C(
        n19002), .Y(n20064) );
  A2O1A1Ixp33_ASAP7_75t_SL U22513 ( .A1(n28056), .A2(n20942), .B(n18295), .C(
        n19002), .Y(n20943) );
  A2O1A1Ixp33_ASAP7_75t_SL U22514 ( .A1(n19002), .A2(n28179), .B(n18295), .C(
        n19002), .Y(n20781) );
  A2O1A1Ixp33_ASAP7_75t_SL U22515 ( .A1(n20780), .A2(n20782), .B(n18295), .C(
        n19002), .Y(n20783) );
  A2O1A1Ixp33_ASAP7_75t_SL U22516 ( .A1(n29510), .A2(n24633), .B(n18295), .C(
        n19002), .Y(n20777) );
  A2O1A1Ixp33_ASAP7_75t_SL U22517 ( .A1(n24666), .A2(n30439), .B(n18295), .C(
        n19002), .Y(n20938) );
  A2O1A1Ixp33_ASAP7_75t_SL U22518 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA1__3_), 
        .A2(n24660), .B(n18295), .C(n19002), .Y(n20762) );
  A2O1A1Ixp33_ASAP7_75t_SL U22519 ( .A1(n24678), .A2(n20933), .B(n18295), .C(
        n19002), .Y(n20934) );
  A2O1A1Ixp33_ASAP7_75t_SL U22520 ( .A1(u0_0_leon3x0_p0_iu_r_X__ICC__3_), .A2(
        n20601), .B(n18295), .C(n19002), .Y(n20602) );
  A2O1A1Ixp33_ASAP7_75t_SL U22521 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__9_), .A2(
        n20928), .B(n18295), .C(n19002), .Y(n20929) );
  A2O1A1Ixp33_ASAP7_75t_SL U22522 ( .A1(n18295), .A2(n19002), .B(n20587), .C(
        n19002), .Y(n20588) );
  A2O1A1Ixp33_ASAP7_75t_SL U22523 ( .A1(n32613), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n20584) );
  A2O1A1Ixp33_ASAP7_75t_SL U22524 ( .A1(n32660), .A2(n32611), .B(n18295), .C(
        n19002), .Y(n20920) );
  A2O1A1Ixp33_ASAP7_75t_SL U22525 ( .A1(n32607), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n20754) );
  A2O1A1Ixp33_ASAP7_75t_SL U22526 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__21_), .A2(n20916), .B(n18295), .C(n19002), .Y(n20917) );
  A2O1A1Ixp33_ASAP7_75t_SL U22527 ( .A1(n32647), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n20911) );
  A2O1A1Ixp33_ASAP7_75t_SL U22528 ( .A1(n32212), .A2(n32234), .B(n18295), .C(
        n19002), .Y(n20260) );
  A2O1A1Ixp33_ASAP7_75t_SL U22529 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__27_), 
        .A2(n30723), .B(n18295), .C(n19002), .Y(n20734) );
  A2O1A1Ixp33_ASAP7_75t_SL U22530 ( .A1(n26950), .A2(n32162), .B(n18295), .C(
        n19002), .Y(n20735) );
  A2O1A1Ixp33_ASAP7_75t_SL U22531 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__27_), 
        .A2(n30726), .B(n18295), .C(n19002), .Y(n20736) );
  A2O1A1Ixp33_ASAP7_75t_SL U22532 ( .A1(u0_0_leon3x0_p0_ici[24]), .A2(n30722), 
        .B(n18295), .C(n19002), .Y(n20737) );
  A2O1A1Ixp33_ASAP7_75t_SL U22533 ( .A1(n20735), .A2(n20736), .B(n18295), .C(
        n20737), .Y(n20738) );
  A2O1A1Ixp33_ASAP7_75t_SL U22534 ( .A1(u0_0_leon3x0_p0_ici[55]), .A2(n30724), 
        .B(n18295), .C(n19002), .Y(n20740) );
  A2O1A1Ixp33_ASAP7_75t_SL U22535 ( .A1(n20734), .A2(n20739), .B(n18295), .C(
        n20740), .Y(rf_di_w[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22536 ( .A1(apbi[46]), .A2(n20904), .B(n18295), 
        .C(n19002), .Y(n20905) );
  A2O1A1Ixp33_ASAP7_75t_SL U22537 ( .A1(u0_0_leon3x0_p0_dci[37]), .A2(
        u0_0_leon3x0_p0_dci[38]), .B(n18295), .C(n19002), .Y(n20899) );
  A2O1A1Ixp33_ASAP7_75t_SL U22538 ( .A1(n18295), .A2(n19002), .B(n19456), .C(
        n19002), .Y(n19457) );
  A2O1A1Ixp33_ASAP7_75t_SL U22539 ( .A1(n19457), .A2(n19458), .B(n18295), .C(
        n19002), .Y(n30678) );
  A2O1A1Ixp33_ASAP7_75t_SL U22540 ( .A1(DP_OP_1196_128_7433_n8), .A2(n20888), 
        .B(n18295), .C(n19002), .Y(n20889) );
  A2O1A1Ixp33_ASAP7_75t_SL U22541 ( .A1(DP_OP_1196_128_7433_n7), .A2(n20888), 
        .B(n18295), .C(n19002), .Y(n20891) );
  A2O1A1Ixp33_ASAP7_75t_SL U22542 ( .A1(DP_OP_1196_128_7433_n67), .A2(n20891), 
        .B(n18295), .C(n19002), .Y(n20892) );
  A2O1A1Ixp33_ASAP7_75t_SL U22543 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__15_), 
        .A2(n29060), .B(n18295), .C(n19002), .Y(n20001) );
  A2O1A1Ixp33_ASAP7_75t_SL U22544 ( .A1(n19002), .A2(n18888), .B(n18295), .C(
        n19002), .Y(n20876) );
  A2O1A1Ixp33_ASAP7_75t_SL U22545 ( .A1(add_x_735_n168), .A2(n20876), .B(
        n18295), .C(n19002), .Y(n20877) );
  A2O1A1Ixp33_ASAP7_75t_SL U22546 ( .A1(add_x_735_n163), .A2(n20877), .B(
        n18295), .C(n19002), .Y(add_x_735_n159) );
  A2O1A1Ixp33_ASAP7_75t_SL U22547 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[60]), 
        .B(n18295), .C(n19002), .Y(n20366) );
  A2O1A1Ixp33_ASAP7_75t_SL U22548 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__29_), .B(n18295), .C(n19002), .Y(n20367) );
  A2O1A1Ixp33_ASAP7_75t_SL U22549 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[61]), 
        .B(n18295), .C(n19002), .Y(n20370) );
  A2O1A1Ixp33_ASAP7_75t_SL U22550 ( .A1(n20366), .A2(n20369), .B(n18295), .C(
        n20370), .Y(u0_0_leon3x0_p0_div0_vaddin1[30]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22551 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[49]), 
        .B(n18295), .C(n19002), .Y(n20509) );
  A2O1A1Ixp33_ASAP7_75t_SL U22552 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__17_), .B(n18295), .C(n19002), .Y(n20510) );
  A2O1A1Ixp33_ASAP7_75t_SL U22553 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[48]), 
        .B(n18295), .C(n19002), .Y(n20513) );
  A2O1A1Ixp33_ASAP7_75t_SL U22554 ( .A1(n20509), .A2(n20512), .B(n18295), .C(
        n20513), .Y(u0_0_leon3x0_p0_div0_vaddin1[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22555 ( .A1(n20872), .A2(mult_x_1196_n844), .B(
        n18295), .C(n19002), .Y(n20874) );
  A2O1A1Ixp33_ASAP7_75t_SL U22556 ( .A1(n20873), .A2(n20874), .B(n18295), .C(
        n19002), .Y(mult_x_1196_n842) );
  A2O1A1Ixp33_ASAP7_75t_SL U22557 ( .A1(n18295), .A2(n19002), .B(n20695), .C(
        n19002), .Y(n20696) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U22558 ( .A1(n20853), .A2(n20855), .B(n18295), 
        .C(n20856), .D(n18295), .Y(n20857) );
  A2O1A1Ixp33_ASAP7_75t_SL U22559 ( .A1(apbi[39]), .A2(apbi[38]), .B(n18295), 
        .C(n19002), .Y(n20843) );
  A2O1A1Ixp33_ASAP7_75t_SL U22560 ( .A1(apbi[42]), .A2(apbi[41]), .B(n18295), 
        .C(apbi[40]), .Y(n20844) );
  A2O1A1Ixp33_ASAP7_75t_SL U22561 ( .A1(apbi[44]), .A2(n20845), .B(n18295), 
        .C(n19002), .Y(n17252) );
  A2O1A1Ixp33_ASAP7_75t_SL U22562 ( .A1(n29954), .A2(uart1_r_TSHIFT__4_), .B(
        n18295), .C(n19002), .Y(n20840) );
  A2O1A1Ixp33_ASAP7_75t_SL U22563 ( .A1(uart1_r_TSHIFT__5_), .A2(n29951), .B(
        n18295), .C(n19002), .Y(n20841) );
  A2O1A1Ixp33_ASAP7_75t_SL U22564 ( .A1(n20840), .A2(n20841), .B(n18295), .C(
        n19002), .Y(n20842) );
  A2O1A1Ixp33_ASAP7_75t_SL U22565 ( .A1(n30244), .A2(n30394), .B(n18295), .C(
        n19002), .Y(n20836) );
  A2O1A1Ixp33_ASAP7_75t_SL U22566 ( .A1(n20835), .A2(n20836), .B(n18295), .C(
        n19002), .Y(n20837) );
  A2O1A1Ixp33_ASAP7_75t_SL U22567 ( .A1(n24665), .A2(n30245), .B(n18295), .C(
        n19002), .Y(n20838) );
  A2O1A1Ixp33_ASAP7_75t_SL U22568 ( .A1(n30640), .A2(rf_do_b[29]), .B(n18295), 
        .C(n19002), .Y(n20822) );
  A2O1A1Ixp33_ASAP7_75t_SL U22569 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__29_), .B(n18295), .C(n19002), .Y(n20823)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22570 ( .A1(n20822), .A2(n20823), .B(n18295), .C(
        n19002), .Y(n20824) );
  A2O1A1Ixp33_ASAP7_75t_SL U22571 ( .A1(n29866), .A2(n31868), .B(n18295), .C(
        n19002), .Y(n20826) );
  A2O1A1Ixp33_ASAP7_75t_SL U22572 ( .A1(n20825), .A2(n20826), .B(n18295), .C(
        n19002), .Y(n20827) );
  A2O1A1Ixp33_ASAP7_75t_SL U22573 ( .A1(n29072), .A2(n29073), .B(n18295), .C(
        n31054), .Y(n20682) );
  A2O1A1Ixp33_ASAP7_75t_SL U22574 ( .A1(n20681), .A2(n20682), .B(n18295), .C(
        n19002), .Y(n4577) );
  A2O1A1Ixp33_ASAP7_75t_SL U22575 ( .A1(n33000), .A2(n22408), .B(n18295), .C(
        n19002), .Y(n20501) );
  A2O1A1Ixp33_ASAP7_75t_SL U22576 ( .A1(n22919), .A2(n20665), .B(n18295), .C(
        n19002), .Y(n20666) );
  A2O1A1Ixp33_ASAP7_75t_SL U22577 ( .A1(n24430), .A2(
        u0_0_leon3x0_p0_div0_r_X__30_), .B(n18295), .C(n19002), .Y(n20668) );
  A2O1A1Ixp33_ASAP7_75t_SL U22578 ( .A1(n24662), .A2(n30677), .B(n18295), .C(
        n19002), .Y(n20102) );
  A2O1A1Ixp33_ASAP7_75t_SL U22579 ( .A1(mult_x_1196_n770), .A2(n24254), .B(
        n18295), .C(n20650), .Y(n20651) );
  A2O1A1Ixp33_ASAP7_75t_SL U22580 ( .A1(n24254), .A2(mult_x_1196_n770), .B(
        n18295), .C(n19002), .Y(n20652) );
  A2O1A1Ixp33_ASAP7_75t_SL U22581 ( .A1(n18384), .A2(n20652), .B(n18295), .C(
        n19002), .Y(n20653) );
  A2O1A1Ixp33_ASAP7_75t_SL U22582 ( .A1(n20651), .A2(n20653), .B(n18295), .C(
        n19002), .Y(n20654) );
  A2O1A1Ixp33_ASAP7_75t_SL U22583 ( .A1(n24664), .A2(n32734), .B(n18295), .C(
        n19002), .Y(n20817) );
  A2O1A1Ixp33_ASAP7_75t_SL U22584 ( .A1(n32630), .A2(n24667), .B(n18295), .C(
        n19002), .Y(n20649) );
  A2O1A1Ixp33_ASAP7_75t_SL U22585 ( .A1(n24674), .A2(n20815), .B(n18295), .C(
        n19002), .Y(n20816) );
  A2O1A1Ixp33_ASAP7_75t_SL U22586 ( .A1(n22393), .A2(ahb0_r_HTRANS__1_), .B(
        n18295), .C(n19002), .Y(n20808) );
  A2O1A1Ixp33_ASAP7_75t_SL U22587 ( .A1(n32036), .A2(n20808), .B(n18295), .C(
        n19002), .Y(n20809) );
  A2O1A1Ixp33_ASAP7_75t_SL U22588 ( .A1(n24694), .A2(n20809), .B(n18295), .C(
        n19002), .Y(n3900) );
  A2O1A1Ixp33_ASAP7_75t_SL U22589 ( .A1(n32126), .A2(n32128), .B(n18295), .C(
        n19002), .Y(n20804) );
  A2O1A1Ixp33_ASAP7_75t_SL U22590 ( .A1(n20805), .A2(n20806), .B(n18295), .C(
        n19002), .Y(n20807) );
  A2O1A1Ixp33_ASAP7_75t_SL U22591 ( .A1(n24670), .A2(n20083), .B(n18295), .C(
        n19002), .Y(n20084) );
  A2O1A1Ixp33_ASAP7_75t_SL U22592 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA2__1_), 
        .A2(n24662), .B(n18295), .C(n19002), .Y(n20628) );
  A2O1A1Ixp33_ASAP7_75t_SL U22593 ( .A1(n24675), .A2(n20626), .B(n18295), .C(
        n19002), .Y(n20627) );
  A2O1A1Ixp33_ASAP7_75t_SL U22594 ( .A1(n24677), .A2(n20795), .B(n18295), .C(
        n19002), .Y(n20796) );
  A2O1A1Ixp33_ASAP7_75t_SL U22595 ( .A1(n28400), .A2(n22378), .B(n18295), .C(
        n19002), .Y(n20450) );
  A2O1A1Ixp33_ASAP7_75t_SL U22596 ( .A1(n22427), .A2(n20792), .B(n18295), .C(
        n19002), .Y(n20793) );
  A2O1A1Ixp33_ASAP7_75t_SL U22597 ( .A1(n24663), .A2(n32677), .B(n18295), .C(
        n19002), .Y(n20791) );
  A2O1A1Ixp33_ASAP7_75t_SL U22598 ( .A1(n19002), .A2(n31583), .B(n18295), .C(
        n19002), .Y(n20786) );
  A2O1A1Ixp33_ASAP7_75t_SL U22599 ( .A1(n13499), .A2(n20786), .B(n18295), .C(
        n19002), .Y(n20787) );
  A2O1A1Ixp33_ASAP7_75t_SL U22600 ( .A1(n31596), .A2(n31582), .B(n18295), .C(
        n20787), .Y(n20788) );
  A2O1A1Ixp33_ASAP7_75t_SL U22601 ( .A1(n19002), .A2(n20788), .B(n18295), .C(
        n19002), .Y(n18102) );
  A2O1A1Ixp33_ASAP7_75t_SL U22602 ( .A1(n24665), .A2(n29898), .B(n18295), .C(
        n19002), .Y(n20784) );
  A2O1A1Ixp33_ASAP7_75t_SL U22603 ( .A1(n28572), .A2(n24677), .B(n18295), .C(
        n19002), .Y(n20612) );
  A2O1A1Ixp33_ASAP7_75t_SL U22604 ( .A1(n29851), .A2(n31198), .B(n18295), .C(
        n19002), .Y(n20610) );
  A2O1A1Ixp33_ASAP7_75t_SL U22605 ( .A1(uart1_r_BRATE__7_), .A2(n20781), .B(
        n18295), .C(n19002), .Y(n20782) );
  A2O1A1Ixp33_ASAP7_75t_SL U22606 ( .A1(n24681), .A2(n20774), .B(n18295), .C(
        n19002), .Y(n20775) );
  A2O1A1Ixp33_ASAP7_75t_SL U22607 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__12_), .A2(
        n20606), .B(n18295), .C(n19002), .Y(n20607) );
  A2O1A1Ixp33_ASAP7_75t_SL U22608 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[44]), 
        .B(n18295), .C(n19002), .Y(n20767) );
  A2O1A1Ixp33_ASAP7_75t_SL U22609 ( .A1(n20766), .A2(n20767), .B(n18295), .C(
        n19002), .Y(n20768) );
  A2O1A1Ixp33_ASAP7_75t_SL U22610 ( .A1(n28593), .A2(n24677), .B(n18295), .C(
        n19002), .Y(n20604) );
  A2O1A1Ixp33_ASAP7_75t_SL U22611 ( .A1(n22421), .A2(n32179), .B(n18295), .C(
        n19002), .Y(n20763) );
  A2O1A1Ixp33_ASAP7_75t_SL U22612 ( .A1(n20762), .A2(n20763), .B(n18295), .C(
        n19002), .Y(n20764) );
  A2O1A1Ixp33_ASAP7_75t_SL U22613 ( .A1(n19002), .A2(n20764), .B(n18295), .C(
        n19002), .Y(n2567) );
  A2O1A1Ixp33_ASAP7_75t_SL U22614 ( .A1(n24678), .A2(n20760), .B(n18295), .C(
        n19002), .Y(n20761) );
  A2O1A1Ixp33_ASAP7_75t_SL U22615 ( .A1(n18295), .A2(n19002), .B(n20590), .C(
        n19002), .Y(n20591) );
  A2O1A1Ixp33_ASAP7_75t_SL U22616 ( .A1(n25239), .A2(n25243), .B(n18295), .C(
        n20756), .Y(n17270) );
  A2O1A1Ixp33_ASAP7_75t_SL U22617 ( .A1(n32660), .A2(n32621), .B(n18295), .C(
        n19002), .Y(n20755) );
  A2O1A1Ixp33_ASAP7_75t_SL U22618 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__19_), .A2(n20750), .B(n18295), .C(n19002), .Y(n20751) );
  A2O1A1Ixp33_ASAP7_75t_SL U22619 ( .A1(n32651), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n20745) );
  A2O1A1Ixp33_ASAP7_75t_SL U22620 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__21_), 
        .A2(n32214), .B(n18295), .C(n19002), .Y(n20742) );
  A2O1A1Ixp33_ASAP7_75t_SL U22621 ( .A1(n20741), .A2(n20742), .B(n18295), .C(
        n19002), .Y(n20743) );
  A2O1A1Ixp33_ASAP7_75t_SL U22622 ( .A1(n19002), .A2(n20743), .B(n18295), .C(
        n19002), .Y(n20744) );
  A2O1A1Ixp33_ASAP7_75t_SL U22623 ( .A1(n30726), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__9_), .B(n18295), .C(n19002), .Y(
        n20727) );
  A2O1A1Ixp33_ASAP7_75t_SL U22624 ( .A1(n27169), .A2(n32162), .B(n18295), .C(
        n19002), .Y(n20728) );
  A2O1A1Ixp33_ASAP7_75t_SL U22625 ( .A1(n30722), .A2(u0_0_leon3x0_p0_ici[6]), 
        .B(n18295), .C(n19002), .Y(n20729) );
  A2O1A1Ixp33_ASAP7_75t_SL U22626 ( .A1(n20727), .A2(n20728), .B(n18295), .C(
        n20729), .Y(n20730) );
  A2O1A1Ixp33_ASAP7_75t_SL U22627 ( .A1(n30723), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__9_), .B(n18295), .C(n19002), .Y(
        n20732) );
  A2O1A1Ixp33_ASAP7_75t_SL U22628 ( .A1(n30724), .A2(u0_0_leon3x0_p0_ici[37]), 
        .B(n18295), .C(n19002), .Y(n20733) );
  A2O1A1Ixp33_ASAP7_75t_SL U22629 ( .A1(n20731), .A2(n20732), .B(n18295), .C(
        n20733), .Y(rf_di_w[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22630 ( .A1(u0_0_leon3x0_p0_iu_fe_pc_17_), .A2(
        u0_0_leon3x0_p0_iu_fe_pc_16_), .B(n18295), .C(n19002), .Y(n20720) );
  A2O1A1Ixp33_ASAP7_75t_SL U22631 ( .A1(add_x_746_n103), .A2(n20721), .B(
        n18295), .C(n19002), .Y(n20722) );
  A2O1A1Ixp33_ASAP7_75t_SL U22632 ( .A1(n28403), .A2(n29778), .B(n18295), .C(
        n19002), .Y(n20716) );
  A2O1A1Ixp33_ASAP7_75t_SL U22633 ( .A1(n22375), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__24_), .B(n18295), .C(n19002), .Y(n20717)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22634 ( .A1(n23002), .A2(n28402), .B(n18295), .C(
        n19002), .Y(n20718) );
  A2O1A1Ixp33_ASAP7_75t_SL U22635 ( .A1(n20716), .A2(n20717), .B(n18295), .C(
        n20718), .Y(n20719) );
  A2O1A1Ixp33_ASAP7_75t_SL U22636 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[33]), 
        .B(n18295), .C(n19002), .Y(n20712) );
  A2O1A1Ixp33_ASAP7_75t_SL U22637 ( .A1(n32786), .A2(n20704), .B(n18295), .C(
        n19002), .Y(n32809) );
  A2O1A1Ixp33_ASAP7_75t_SL U22638 ( .A1(n32353), .A2(n32339), .B(n18295), .C(
        n19002), .Y(n20703) );
  A2O1A1Ixp33_ASAP7_75t_SL U22639 ( .A1(n32353), .A2(n32302), .B(n18295), .C(
        n19002), .Y(n20702) );
  A2O1A1Ixp33_ASAP7_75t_SL U22640 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[41]), 
        .B(n18295), .C(n19002), .Y(n20701) );
  A2O1A1Ixp33_ASAP7_75t_SL U22641 ( .A1(DP_OP_1196_128_7433_n264), .A2(
        DP_OP_1196_128_7433_n291), .B(n18295), .C(n19002), .Y(n20514) );
  A2O1A1Ixp33_ASAP7_75t_SL U22642 ( .A1(n19002), .A2(n20515), .B(n18295), .C(
        n19002), .Y(DP_OP_1196_128_7433_n263) );
  A2O1A1Ixp33_ASAP7_75t_SL U22643 ( .A1(n28193), .A2(uart1_r_RWADDR__2_), .B(
        n18295), .C(n19002), .Y(n20698) );
  A2O1A1Ixp33_ASAP7_75t_SL U22644 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[54]), 
        .B(n18295), .C(n19002), .Y(n19985) );
  A2O1A1Ixp33_ASAP7_75t_SL U22645 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__23_), .B(n18295), .C(n19002), .Y(n19986) );
  A2O1A1Ixp33_ASAP7_75t_SL U22646 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[55]), 
        .B(n18295), .C(n19002), .Y(n19989) );
  A2O1A1Ixp33_ASAP7_75t_SL U22647 ( .A1(n19985), .A2(n19988), .B(n18295), .C(
        n19989), .Y(u0_0_leon3x0_p0_div0_vaddin1[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22648 ( .A1(mult_x_1196_n867), .A2(n20697), .B(
        n18295), .C(n19002), .Y(mult_x_1196_n339) );
  A2O1A1Ixp33_ASAP7_75t_SL U22649 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[49]), 
        .B(n18295), .C(n19002), .Y(n20157) );
  A2O1A1Ixp33_ASAP7_75t_SL U22650 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__18_), .B(n18295), .C(n19002), .Y(n20158) );
  A2O1A1Ixp33_ASAP7_75t_SL U22651 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[50]), 
        .B(n18295), .C(n19002), .Y(n20161) );
  A2O1A1Ixp33_ASAP7_75t_SL U22652 ( .A1(n20157), .A2(n20160), .B(n18295), .C(
        n20161), .Y(u0_0_leon3x0_p0_div0_vaddin1[19]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22653 ( .A1(n18295), .A2(n19002), .B(n20505), .C(
        n19002), .Y(n20506) );
  A2O1A1Ixp33_ASAP7_75t_SL U22654 ( .A1(n4742), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n20693) );
  A2O1A1Ixp33_ASAP7_75t_SL U22655 ( .A1(n30030), .A2(n20693), .B(n18295), .C(
        n19002), .Y(n20694) );
  A2O1A1Ixp33_ASAP7_75t_SL U22656 ( .A1(n20694), .A2(n20696), .B(n18295), .C(
        n19002), .Y(n17722) );
  A2O1A1Ixp33_ASAP7_75t_SL U22657 ( .A1(sr1_r_MCFG1__IOWS__0_), .A2(n31720), 
        .B(n18295), .C(n19002), .Y(n20140) );
  A2O1A1Ixp33_ASAP7_75t_SL U22658 ( .A1(sr1_r_MCFG1__ROMWWS__0_), .A2(n31725), 
        .B(n18295), .C(n19002), .Y(n20150) );
  A2O1A1Ixp33_ASAP7_75t_SL U22659 ( .A1(n20140), .A2(n20149), .B(n18295), .C(
        n20150), .Y(n20151) );
  A2O1A1Ixp33_ASAP7_75t_SL U22660 ( .A1(n24694), .A2(n20151), .B(n18295), .C(
        n19002), .Y(n4723) );
  A2O1A1Ixp33_ASAP7_75t_SL U22661 ( .A1(n29954), .A2(uart1_r_TSHIFT__2_), .B(
        n18295), .C(n19002), .Y(n20359) );
  A2O1A1Ixp33_ASAP7_75t_SL U22662 ( .A1(n18845), .A2(n20687), .B(n18295), .C(
        n19002), .Y(n20688) );
  A2O1A1Ixp33_ASAP7_75t_SL U22663 ( .A1(n22408), .A2(n20683), .B(n18295), .C(
        n19002), .Y(n20684) );
  A2O1A1Ixp33_ASAP7_75t_SL U22664 ( .A1(n31043), .A2(n31357), .B(n18295), .C(
        n19002), .Y(n20677) );
  A2O1A1Ixp33_ASAP7_75t_SL U22665 ( .A1(n31364), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__9_), .B(n18295), .C(n19002), .Y(
        n20678) );
  A2O1A1Ixp33_ASAP7_75t_SL U22666 ( .A1(n20677), .A2(n20678), .B(n18295), .C(
        n19002), .Y(n20679) );
  A2O1A1Ixp33_ASAP7_75t_SL U22667 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_div0_r_NEG_), .B(n18295), .C(n19002), .Y(n20665) );
  A2O1A1Ixp33_ASAP7_75t_SL U22668 ( .A1(n31674), .A2(n20666), .B(n18295), .C(
        n19002), .Y(n20667) );
  A2O1A1Ixp33_ASAP7_75t_SL U22669 ( .A1(n19002), .A2(n20669), .B(n18295), .C(
        n19002), .Y(n20670) );
  A2O1A1Ixp33_ASAP7_75t_SL U22670 ( .A1(n20667), .A2(n20670), .B(n18295), .C(
        n19002), .Y(n20671) );
  A2O1A1Ixp33_ASAP7_75t_SL U22671 ( .A1(n30640), .A2(rf_do_b[30]), .B(n18295), 
        .C(n19002), .Y(n20657) );
  A2O1A1Ixp33_ASAP7_75t_SL U22672 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__30_), .B(n18295), .C(n19002), .Y(n20658)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22673 ( .A1(n20657), .A2(n20658), .B(n18295), .C(
        n19002), .Y(n20659) );
  A2O1A1Ixp33_ASAP7_75t_SL U22674 ( .A1(n20662), .A2(n30593), .B(n18295), .C(
        n19002), .Y(n20663) );
  A2O1A1Ixp33_ASAP7_75t_SL U22675 ( .A1(u0_0_leon3x0_p0_divi[42]), .A2(n19352), 
        .B(n18295), .C(n19002), .Y(n19353) );
  A2O1A1Ixp33_ASAP7_75t_SL U22676 ( .A1(n30390), .A2(n24664), .B(n18295), .C(
        n19002), .Y(n19357) );
  A2O1A1Ixp33_ASAP7_75t_SL U22677 ( .A1(n31981), .A2(n24659), .B(n18295), .C(
        n19002), .Y(n20474) );
  A2O1A1Ixp33_ASAP7_75t_SL U22678 ( .A1(n27521), .A2(n31940), .B(n18295), .C(
        n19002), .Y(n20641) );
  A2O1A1Ixp33_ASAP7_75t_SL U22679 ( .A1(n20641), .A2(n20642), .B(n18295), .C(
        n19002), .Y(n20643) );
  A2O1A1Ixp33_ASAP7_75t_SL U22680 ( .A1(n29980), .A2(n27523), .B(n18295), .C(
        n20643), .Y(n20644) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U22681 ( .A1(n29980), .A2(n27523), .B(n18295), 
        .C(n20643), .D(n20646), .Y(n20647) );
  A2O1A1Ixp33_ASAP7_75t_SL U22682 ( .A1(n24648), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PV_), .B(n18295), .C(n19002), .Y(n19732)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22683 ( .A1(n24674), .A2(n25170), .B(n18295), .C(
        n19002), .Y(n20639) );
  A2O1A1Ixp33_ASAP7_75t_SL U22684 ( .A1(n31339), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n20462) );
  A2O1A1Ixp33_ASAP7_75t_SL U22685 ( .A1(n24673), .A2(n25689), .B(n18295), .C(
        n19002), .Y(n20637) );
  A2O1A1Ixp33_ASAP7_75t_SL U22686 ( .A1(n24667), .A2(n23835), .B(n18295), .C(
        n19002), .Y(n20634) );
  A2O1A1Ixp33_ASAP7_75t_SL U22687 ( .A1(n23229), .A2(DP_OP_1196_128_7433_n453), 
        .B(n18295), .C(n19002), .Y(n20629) );
  A2O1A1Ixp33_ASAP7_75t_SL U22688 ( .A1(n20628), .A2(n20629), .B(n18295), .C(
        n19002), .Y(n20630) );
  A2O1A1Ixp33_ASAP7_75t_SL U22689 ( .A1(n19002), .A2(n20630), .B(n18295), .C(
        n19002), .Y(n3540) );
  A2O1A1Ixp33_ASAP7_75t_SL U22690 ( .A1(n24659), .A2(n20621), .B(n18295), .C(
        n19002), .Y(n20622) );
  A2O1A1Ixp33_ASAP7_75t_SL U22691 ( .A1(n24676), .A2(n20448), .B(n18295), .C(
        n19002), .Y(n20449) );
  A2O1A1Ixp33_ASAP7_75t_SL U22692 ( .A1(n24677), .A2(n32586), .B(n18295), .C(
        n19002), .Y(n20618) );
  A2O1A1Ixp33_ASAP7_75t_SL U22693 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA1__7_), 
        .A2(n24659), .B(n18295), .C(n19002), .Y(n20311) );
  A2O1A1Ixp33_ASAP7_75t_SL U22694 ( .A1(n3135), .A2(n32562), .B(n18295), .C(
        n19002), .Y(n19507) );
  A2O1A1Ixp33_ASAP7_75t_SL U22695 ( .A1(n22396), .A2(n20613), .B(n18295), .C(
        n19002), .Y(n20614) );
  A2O1A1Ixp33_ASAP7_75t_SL U22696 ( .A1(n28699), .A2(n24677), .B(n18295), .C(
        n19002), .Y(n20438) );
  A2O1A1Ixp33_ASAP7_75t_SL U22697 ( .A1(n24604), .A2(n24603), .B(n18295), .C(
        n24595), .Y(n20297) );
  A2O1A1Ixp33_ASAP7_75t_SL U22698 ( .A1(n29568), .A2(n24633), .B(n18295), .C(
        n19002), .Y(n20061) );
  A2O1A1Ixp33_ASAP7_75t_SL U22699 ( .A1(n31423), .A2(n24665), .B(n18295), .C(
        n19002), .Y(n20437) );
  A2O1A1Ixp33_ASAP7_75t_SL U22700 ( .A1(n24677), .A2(n30361), .B(n18295), .C(
        n19002), .Y(n20605) );
  A2O1A1Ixp33_ASAP7_75t_SL U22701 ( .A1(n32786), .A2(n32834), .B(n18295), .C(
        n19002), .Y(n20600) );
  A2O1A1Ixp33_ASAP7_75t_SL U22702 ( .A1(n29356), .A2(n24694), .B(n18295), .C(
        n19002), .Y(n20593) );
  A2O1A1Ixp33_ASAP7_75t_SL U22703 ( .A1(n27357), .A2(n20593), .B(n18295), .C(
        n19002), .Y(n20594) );
  A2O1A1Ixp33_ASAP7_75t_SL U22704 ( .A1(n32617), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n20430) );
  A2O1A1Ixp33_ASAP7_75t_SL U22705 ( .A1(n32609), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n20429) );
  A2O1A1Ixp33_ASAP7_75t_SL U22706 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__18_), .A2(n20582), .B(n18295), .C(n19002), .Y(n20583) );
  A2O1A1Ixp33_ASAP7_75t_SL U22707 ( .A1(n33069), .A2(dc_q[31]), .B(n18295), 
        .C(n19002), .Y(n20576) );
  A2O1A1Ixp33_ASAP7_75t_SL U22708 ( .A1(DP_OP_5187J1_124_3275_n213), .A2(
        DP_OP_5187J1_124_3275_n231), .B(n18295), .C(n19002), .Y(n20557) );
  A2O1A1Ixp33_ASAP7_75t_SL U22709 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[57]), 
        .B(n18295), .C(n19002), .Y(n20556) );
  A2O1A1Ixp33_ASAP7_75t_SL U22710 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__27_), .B(n18295), .C(n19002), .Y(
        n20188) );
  A2O1A1Ixp33_ASAP7_75t_SL U22711 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__21_), .B(n18295), .C(n19002), .Y(
        n20551) );
  A2O1A1Ixp33_ASAP7_75t_SL U22712 ( .A1(n23914), .A2(mult_x_1196_n524), .B(
        n18295), .C(n19002), .Y(n20547) );
  A2O1A1Ixp33_ASAP7_75t_SL U22713 ( .A1(n22274), .A2(add_x_735_n272), .B(
        n18295), .C(n20384), .Y(n20385) );
  A2O1A1Ixp33_ASAP7_75t_SL U22714 ( .A1(n22274), .A2(add_x_735_n272), .B(
        n18295), .C(n19002), .Y(n20386) );
  A2O1A1Ixp33_ASAP7_75t_SL U22715 ( .A1(n20386), .A2(
        u0_0_leon3x0_p0_iu_r_E__ALUCIN_), .B(n18295), .C(n19002), .Y(n20387)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22716 ( .A1(n20385), .A2(n20387), .B(n18295), .C(
        n19002), .Y(u0_0_leon3x0_p0_dci[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22717 ( .A1(n19642), .A2(n19643), .B(n18295), .C(
        n19002), .Y(n19644) );
  A2O1A1Ixp33_ASAP7_75t_SL U22718 ( .A1(n19645), .A2(n19646), .B(n18295), .C(
        n19002), .Y(n19647) );
  A2O1A1Ixp33_ASAP7_75t_SL U22719 ( .A1(n20537), .A2(n20538), .B(n18295), .C(
        n19002), .Y(n20539) );
  A2O1A1Ixp33_ASAP7_75t_SL U22720 ( .A1(n20539), .A2(n20540), .B(n18295), .C(
        n19002), .Y(n29694) );
  A2O1A1Ixp33_ASAP7_75t_SL U22721 ( .A1(DP_OP_1196_128_7433_n91), .A2(n20536), 
        .B(n18295), .C(n19002), .Y(DP_OP_1196_128_7433_n14) );
  A2O1A1Ixp33_ASAP7_75t_SL U22722 ( .A1(uart1_r_TXCLK__1_), .A2(n20531), .B(
        n18295), .C(n19002), .Y(n26086) );
  A2O1A1Ixp33_ASAP7_75t_SL U22723 ( .A1(n2388), .A2(n20527), .B(n18295), .C(
        n19002), .Y(n27446) );
  A2O1A1Ixp33_ASAP7_75t_SL U22724 ( .A1(n29059), .A2(u0_0_leon3x0_p0_ici[37]), 
        .B(n18295), .C(n19002), .Y(n20524) );
  A2O1A1Ixp33_ASAP7_75t_SL U22725 ( .A1(n20523), .A2(n20524), .B(n18295), .C(
        n19002), .Y(n20525) );
  A2O1A1Ixp33_ASAP7_75t_SL U22726 ( .A1(n19002), .A2(n20525), .B(n18295), .C(
        n19002), .Y(n20526) );
  A2O1A1Ixp33_ASAP7_75t_SL U22727 ( .A1(n28847), .A2(n28966), .B(n18295), .C(
        n19002), .Y(n20518) );
  A2O1A1Ixp33_ASAP7_75t_SL U22728 ( .A1(n26293), .A2(n24575), .B(n18295), .C(
        n19002), .Y(n20519) );
  A2O1A1Ixp33_ASAP7_75t_SL U22729 ( .A1(n20518), .A2(n20519), .B(n18295), .C(
        n19002), .Y(n20520) );
  A2O1A1Ixp33_ASAP7_75t_SL U22730 ( .A1(n27098), .A2(n26552), .B(n18295), .C(
        n19002), .Y(n20522) );
  A2O1A1Ixp33_ASAP7_75t_SL U22731 ( .A1(n20521), .A2(n20522), .B(n18295), .C(
        n19002), .Y(n28741) );
  A2O1A1Ixp33_ASAP7_75t_SL U22732 ( .A1(n19002), .A2(n22406), .B(n18295), .C(
        n19002), .Y(n20516) );
  A2O1A1Ixp33_ASAP7_75t_SL U22733 ( .A1(n23768), .A2(n20516), .B(n18295), .C(
        n19002), .Y(n20517) );
  A2O1A1Ixp33_ASAP7_75t_SL U22734 ( .A1(mult_x_1196_n355), .A2(n20517), .B(
        n18295), .C(n19002), .Y(n23671) );
  A2O1A1Ixp33_ASAP7_75t_SL U22735 ( .A1(DP_OP_1196_128_7433_n267), .A2(n20514), 
        .B(n18295), .C(n19002), .Y(n20515) );
  A2O1A1Ixp33_ASAP7_75t_SL U22736 ( .A1(uart1_r_RWADDR__2_), .A2(
        uart1_r_RWADDR__0_), .B(n18295), .C(n19002), .Y(n20371) );
  A2O1A1Ixp33_ASAP7_75t_SL U22737 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[53]), 
        .B(n18295), .C(n19002), .Y(n19783) );
  A2O1A1Ixp33_ASAP7_75t_SL U22738 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__21_), .B(n18295), .C(n19002), .Y(n19784) );
  A2O1A1Ixp33_ASAP7_75t_SL U22739 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[52]), 
        .B(n18295), .C(n19002), .Y(n19787) );
  A2O1A1Ixp33_ASAP7_75t_SL U22740 ( .A1(n19783), .A2(n19786), .B(n18295), .C(
        n19787), .Y(u0_0_leon3x0_p0_div0_vaddin1[22]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22741 ( .A1(mult_x_1196_n849), .A2(n20506), .B(
        n18295), .C(n20507), .Y(n20508) );
  A2O1A1Ixp33_ASAP7_75t_SL U22742 ( .A1(n19002), .A2(n28028), .B(n18295), .C(
        n19002), .Y(n20360) );
  A2O1A1Ixp33_ASAP7_75t_SL U22743 ( .A1(n20359), .A2(n20361), .B(n18295), .C(
        n19002), .Y(n20362) );
  A2O1A1Ixp33_ASAP7_75t_SL U22744 ( .A1(n18295), .A2(n19002), .B(n20124), .C(
        n19002), .Y(n20125) );
  A2O1A1Ixp33_ASAP7_75t_SL U22745 ( .A1(n30733), .A2(n31542), .B(n18295), .C(
        n19002), .Y(n20126) );
  A2O1A1Ixp33_ASAP7_75t_SL U22746 ( .A1(n27175), .A2(n24647), .B(n18295), .C(
        n19002), .Y(n20127) );
  A2O1A1Ixp33_ASAP7_75t_SL U22747 ( .A1(n20125), .A2(n20126), .B(n18295), .C(
        n20127), .Y(n4555) );
  A2O1A1Ixp33_ASAP7_75t_SL U22748 ( .A1(n30640), .A2(rf_do_b[31]), .B(n18295), 
        .C(n19002), .Y(n20490) );
  A2O1A1Ixp33_ASAP7_75t_SL U22749 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__31_), .B(n18295), .C(n19002), .Y(n20491)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22750 ( .A1(n20490), .A2(n20491), .B(n18295), .C(
        n19002), .Y(n20492) );
  A2O1A1Ixp33_ASAP7_75t_SL U22751 ( .A1(n31681), .A2(n31868), .B(n18295), .C(
        n19002), .Y(n20494) );
  A2O1A1Ixp33_ASAP7_75t_SL U22752 ( .A1(n20493), .A2(n20494), .B(n18295), .C(
        n19002), .Y(n20495) );
  A2O1A1Ixp33_ASAP7_75t_SL U22753 ( .A1(u0_0_leon3x0_p0_divi[40]), .A2(n30430), 
        .B(n18295), .C(n19002), .Y(n20484) );
  A2O1A1Ixp33_ASAP7_75t_SL U22754 ( .A1(n20483), .A2(n20484), .B(n18295), .C(
        n19002), .Y(n20485) );
  A2O1A1Ixp33_ASAP7_75t_SL U22755 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[58]), 
        .B(n18295), .C(n19002), .Y(n20477) );
  A2O1A1Ixp33_ASAP7_75t_SL U22756 ( .A1(n20476), .A2(n20477), .B(n18295), .C(
        n19002), .Y(n20478) );
  A2O1A1Ixp33_ASAP7_75t_SL U22757 ( .A1(n29104), .A2(n24675), .B(n18295), .C(
        n19002), .Y(n20335) );
  A2O1A1Ixp33_ASAP7_75t_SL U22758 ( .A1(n24663), .A2(n32636), .B(n18295), .C(
        n19002), .Y(n20473) );
  A2O1A1Ixp33_ASAP7_75t_SL U22759 ( .A1(n19002), .A2(n26808), .B(n18295), .C(
        n19002), .Y(n20466) );
  A2O1A1Ixp33_ASAP7_75t_SL U22760 ( .A1(n26811), .A2(n20466), .B(n18295), .C(
        n19002), .Y(n20467) );
  A2O1A1Ixp33_ASAP7_75t_SL U22761 ( .A1(n26810), .A2(n20467), .B(n18295), .C(
        n19002), .Y(n20468) );
  A2O1A1Ixp33_ASAP7_75t_SL U22762 ( .A1(n22379), .A2(n30464), .B(n18295), .C(
        n19002), .Y(n19725) );
  A2O1A1Ixp33_ASAP7_75t_SL U22763 ( .A1(n24675), .A2(n25670), .B(n18295), .C(
        n19002), .Y(n20463) );
  A2O1A1Ixp33_ASAP7_75t_SL U22764 ( .A1(n25553), .A2(n24670), .B(n18295), .C(
        n19002), .Y(n19135) );
  A2O1A1Ixp33_ASAP7_75t_SL U22765 ( .A1(n24670), .A2(n19315), .B(n18295), .C(
        n19002), .Y(n19316) );
  A2O1A1Ixp33_ASAP7_75t_SL U22766 ( .A1(n24661), .A2(n19715), .B(n18295), .C(
        n19002), .Y(n19716) );
  A2O1A1Ixp33_ASAP7_75t_SL U22767 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA2__2_), 
        .A2(n24662), .B(n18295), .C(n19002), .Y(n20451) );
  A2O1A1Ixp33_ASAP7_75t_SL U22768 ( .A1(n32163), .A2(n20451), .B(n18295), .C(
        n19002), .Y(n20452) );
  A2O1A1Ixp33_ASAP7_75t_SL U22769 ( .A1(n19002), .A2(n20452), .B(n18295), .C(
        n19002), .Y(n3536) );
  A2O1A1Ixp33_ASAP7_75t_SL U22770 ( .A1(n24675), .A2(n19707), .B(n18295), .C(
        n19002), .Y(n19708) );
  A2O1A1Ixp33_ASAP7_75t_SL U22771 ( .A1(n32150), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n20305) );
  A2O1A1Ixp33_ASAP7_75t_SL U22772 ( .A1(n22396), .A2(n20444), .B(n18295), .C(
        n19002), .Y(n20445) );
  A2O1A1Ixp33_ASAP7_75t_SL U22773 ( .A1(n31299), .A2(n24684), .B(n18295), .C(
        n20442), .Y(n20443) );
  A2O1A1Ixp33_ASAP7_75t_SL U22774 ( .A1(n24661), .A2(n20303), .B(n18295), .C(
        n19002), .Y(n20304) );
  A2O1A1Ixp33_ASAP7_75t_SL U22775 ( .A1(n19002), .A2(n28179), .B(n18295), .C(
        n19002), .Y(n20300) );
  A2O1A1Ixp33_ASAP7_75t_SL U22776 ( .A1(n20299), .A2(n20301), .B(n18295), .C(
        n19002), .Y(n20302) );
  A2O1A1Ixp33_ASAP7_75t_SL U22777 ( .A1(n29851), .A2(n24633), .B(n18295), .C(
        n19002), .Y(n20296) );
  A2O1A1Ixp33_ASAP7_75t_SL U22778 ( .A1(n28509), .A2(n24678), .B(n18295), .C(
        n19002), .Y(n20290) );
  A2O1A1Ixp33_ASAP7_75t_SL U22779 ( .A1(n18295), .A2(n19002), .B(n20053), .C(
        n19002), .Y(n20054) );
  A2O1A1Ixp33_ASAP7_75t_SL U22780 ( .A1(n29356), .A2(n20054), .B(n18295), .C(
        n19002), .Y(n20055) );
  A2O1A1Ixp33_ASAP7_75t_SL U22781 ( .A1(n18295), .A2(n19002), .B(n20280), .C(
        n19002), .Y(n20281) );
  A2O1A1Ixp33_ASAP7_75t_SL U22782 ( .A1(n18295), .A2(n19002), .B(n20277), .C(
        n19002), .Y(n20278) );
  A2O1A1Ixp33_ASAP7_75t_SL U22783 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__17_), .A2(n20426), .B(n18295), .C(n19002), .Y(n20427) );
  A2O1A1Ixp33_ASAP7_75t_SL U22784 ( .A1(n32414), .A2(n32400), .B(n18295), .C(
        n19002), .Y(n20425) );
  A2O1A1Ixp33_ASAP7_75t_SL U22785 ( .A1(n20424), .A2(n20425), .B(n18295), .C(
        n19002), .Y(dc_data[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22786 ( .A1(n32396), .A2(n20415), .B(n18295), .C(
        n19002), .Y(n20416) );
  A2O1A1Ixp33_ASAP7_75t_SL U22787 ( .A1(n32600), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n20417) );
  A2O1A1Ixp33_ASAP7_75t_SL U22788 ( .A1(n32318), .A2(dc_q[1]), .B(n18295), .C(
        n19002), .Y(n20418) );
  A2O1A1Ixp33_ASAP7_75t_SL U22789 ( .A1(n20416), .A2(n20417), .B(n18295), .C(
        n20418), .Y(dc_data[1]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22790 ( .A1(n32211), .A2(n32234), .B(n18295), .C(
        n19002), .Y(n19660) );
  A2O1A1Ixp33_ASAP7_75t_SL U22791 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__15_), 
        .A2(n30723), .B(n18295), .C(n19002), .Y(n20253) );
  A2O1A1Ixp33_ASAP7_75t_SL U22792 ( .A1(n28574), .A2(n32162), .B(n18295), .C(
        n19002), .Y(n20254) );
  A2O1A1Ixp33_ASAP7_75t_SL U22793 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__15_), 
        .A2(n30726), .B(n18295), .C(n19002), .Y(n20255) );
  A2O1A1Ixp33_ASAP7_75t_SL U22794 ( .A1(u0_0_leon3x0_p0_ici[12]), .A2(n30722), 
        .B(n18295), .C(n19002), .Y(n20256) );
  A2O1A1Ixp33_ASAP7_75t_SL U22795 ( .A1(n20254), .A2(n20255), .B(n18295), .C(
        n20256), .Y(n20257) );
  A2O1A1Ixp33_ASAP7_75t_SL U22796 ( .A1(u0_0_leon3x0_p0_ici[43]), .A2(n30724), 
        .B(n18295), .C(n19002), .Y(n20259) );
  A2O1A1Ixp33_ASAP7_75t_SL U22797 ( .A1(n20253), .A2(n20258), .B(n18295), .C(
        n20259), .Y(rf_di_w[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22798 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__14_), .B(n18295), .C(n19002), .Y(
        n20414) );
  A2O1A1Ixp33_ASAP7_75t_SL U22799 ( .A1(n28403), .A2(n29783), .B(n18295), .C(
        n19002), .Y(n20411) );
  A2O1A1Ixp33_ASAP7_75t_SL U22800 ( .A1(n18606), .A2(n28402), .B(n18295), .C(
        n19002), .Y(n20412) );
  A2O1A1Ixp33_ASAP7_75t_SL U22801 ( .A1(n28419), .A2(n20411), .B(n18295), .C(
        n20412), .Y(n20413) );
  A2O1A1Ixp33_ASAP7_75t_SL U22802 ( .A1(n31392), .A2(
        u0_0_leon3x0_p0_iu_r_W__RESULT__21_), .B(n18295), .C(n19002), .Y(
        n20403) );
  A2O1A1Ixp33_ASAP7_75t_SL U22803 ( .A1(n31391), .A2(rf_do_a[21]), .B(n18295), 
        .C(n19002), .Y(n20404) );
  A2O1A1Ixp33_ASAP7_75t_SL U22804 ( .A1(n20403), .A2(n20404), .B(n18295), .C(
        n19002), .Y(n20405) );
  A2O1A1Ixp33_ASAP7_75t_SL U22805 ( .A1(n31545), .A2(n31342), .B(n18295), .C(
        n19002), .Y(n20407) );
  A2O1A1Ixp33_ASAP7_75t_SL U22806 ( .A1(n20406), .A2(n20407), .B(n18295), .C(
        n19002), .Y(n31543) );
  A2O1A1Ixp33_ASAP7_75t_SL U22807 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[42]), 
        .B(n18295), .C(n19002), .Y(n20401) );
  A2O1A1Ixp33_ASAP7_75t_SL U22808 ( .A1(DP_OP_5187J1_124_3275_n231), .A2(
        n20392), .B(n18295), .C(n19002), .Y(n20393) );
  A2O1A1Ixp33_ASAP7_75t_SL U22809 ( .A1(DP_OP_5187J1_124_3275_n214), .A2(
        n20395), .B(n18295), .C(n19002), .Y(n20396) );
  A2O1A1Ixp33_ASAP7_75t_SL U22810 ( .A1(DP_OP_5187J1_124_3275_n209), .A2(
        n20396), .B(n18295), .C(n19002), .Y(n20397) );
  A2O1A1Ixp33_ASAP7_75t_SL U22811 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[54]), 
        .B(n18295), .C(n19002), .Y(n20390) );
  A2O1A1Ixp33_ASAP7_75t_SL U22812 ( .A1(u0_0_leon3x0_p0_ici[55]), .A2(n29059), 
        .B(n18295), .C(n19002), .Y(n20187) );
  A2O1A1Ixp33_ASAP7_75t_SL U22813 ( .A1(n19002), .A2(n20189), .B(n18295), .C(
        n19002), .Y(n20190) );
  A2O1A1Ixp33_ASAP7_75t_SL U22814 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__6_), .B(n18295), .C(n19002), .Y(
        n20389) );
  A2O1A1Ixp33_ASAP7_75t_SL U22815 ( .A1(n24681), .A2(n20388), .B(n18295), .C(
        n19002), .Y(n32176) );
  A2O1A1Ixp33_ASAP7_75t_SL U22816 ( .A1(n31609), .A2(n20376), .B(n18295), .C(
        n19002), .Y(n31313) );
  A2O1A1Ixp33_ASAP7_75t_SL U22817 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__13_), 
        .A2(n29060), .B(n18295), .C(n19002), .Y(n20180) );
  A2O1A1Ixp33_ASAP7_75t_SL U22818 ( .A1(n2387), .A2(n20373), .B(n18295), .C(
        n19002), .Y(n27451) );
  A2O1A1Ixp33_ASAP7_75t_SL U22819 ( .A1(u0_0_leon3x0_p0_iu_fe_pc_8_), .A2(
        n20372), .B(n18295), .C(n19002), .Y(add_x_746_n131) );
  A2O1A1Ixp33_ASAP7_75t_SL U22820 ( .A1(n22214), .A2(mult_x_1196_n229), .B(
        n18295), .C(n22421), .Y(n23210) );
  A2O1A1Ixp33_ASAP7_75t_SL U22821 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[50]), 
        .B(n18295), .C(n19002), .Y(n19619) );
  A2O1A1Ixp33_ASAP7_75t_SL U22822 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__19_), .B(n18295), .C(n19002), .Y(n19620) );
  A2O1A1Ixp33_ASAP7_75t_SL U22823 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[51]), 
        .B(n18295), .C(n19002), .Y(n19623) );
  A2O1A1Ixp33_ASAP7_75t_SL U22824 ( .A1(n19619), .A2(n19622), .B(n18295), .C(
        n19623), .Y(u0_0_leon3x0_p0_div0_vaddin1[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22825 ( .A1(n31727), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n20144) );
  A2O1A1Ixp33_ASAP7_75t_SL U22826 ( .A1(n19002), .A2(n20145), .B(n18295), .C(
        n19002), .Y(n20146) );
  A2O1A1Ixp33_ASAP7_75t_SL U22827 ( .A1(uart1_r_TSHIFT__3_), .A2(n20360), .B(
        n18295), .C(n19002), .Y(n20361) );
  A2O1A1Ixp33_ASAP7_75t_SL U22828 ( .A1(n19002), .A2(n29727), .B(n18295), .C(
        n19002), .Y(n20354) );
  A2O1A1Ixp33_ASAP7_75t_SL U22829 ( .A1(n30708), .A2(n20354), .B(n18295), .C(
        n19002), .Y(n20355) );
  A2O1A1Ixp33_ASAP7_75t_SL U22830 ( .A1(n20355), .A2(n29886), .B(n18295), .C(
        n19002), .Y(n20356) );
  A2O1A1Ixp33_ASAP7_75t_SL U22831 ( .A1(n22408), .A2(n32998), .B(n18295), .C(
        n19002), .Y(n20353) );
  A2O1A1Ixp33_ASAP7_75t_SL U22832 ( .A1(n30640), .A2(rf_do_b[11]), .B(n18295), 
        .C(n19002), .Y(n20343) );
  A2O1A1Ixp33_ASAP7_75t_SL U22833 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__11_), .B(n18295), .C(n19002), .Y(n20344)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22834 ( .A1(n20343), .A2(n20344), .B(n18295), .C(
        n19002), .Y(n20345) );
  A2O1A1Ixp33_ASAP7_75t_SL U22835 ( .A1(n19157), .A2(n19162), .B(n18295), .C(
        n19002), .Y(n19163) );
  A2O1A1Ixp33_ASAP7_75t_SL U22836 ( .A1(n24665), .A2(n30265), .B(n18295), .C(
        n19002), .Y(n19164) );
  A2O1A1Ixp33_ASAP7_75t_SL U22837 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[52]), 
        .B(n18295), .C(n19002), .Y(n20338) );
  A2O1A1Ixp33_ASAP7_75t_SL U22838 ( .A1(n20337), .A2(n20338), .B(n18295), .C(
        n19002), .Y(n20339) );
  A2O1A1Ixp33_ASAP7_75t_SL U22839 ( .A1(mult_x_1196_n761), .A2(n22624), .B(
        n18295), .C(n20332), .Y(n20333) );
  A2O1A1Ixp33_ASAP7_75t_SL U22840 ( .A1(n32638), .A2(n24678), .B(n18295), .C(
        n19002), .Y(n20097) );
  A2O1A1Ixp33_ASAP7_75t_SL U22841 ( .A1(n31959), .A2(n24659), .B(n18295), .C(
        n19002), .Y(n19532) );
  A2O1A1Ixp33_ASAP7_75t_SL U22842 ( .A1(n30935), .A2(n24668), .B(n18295), .C(
        n19002), .Y(n19137) );
  A2O1A1Ixp33_ASAP7_75t_SL U22843 ( .A1(n32037), .A2(n24694), .B(n18295), .C(
        n20330), .Y(n20331) );
  A2O1A1Ixp33_ASAP7_75t_SL U22844 ( .A1(n24659), .A2(n19878), .B(n18295), .C(
        n19002), .Y(n19879) );
  A2O1A1Ixp33_ASAP7_75t_SL U22845 ( .A1(n32054), .A2(n32055), .B(n18295), .C(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), .Y(n19317) );
  A2O1A1Ixp33_ASAP7_75t_SL U22846 ( .A1(n31811), .A2(n19322), .B(n18295), .C(
        n19002), .Y(n19323) );
  A2O1A1Ixp33_ASAP7_75t_SL U22847 ( .A1(n19319), .A2(n19325), .B(n18295), .C(
        n19002), .Y(n19326) );
  A2O1A1Ixp33_ASAP7_75t_SL U22848 ( .A1(n24670), .A2(n20328), .B(n18295), .C(
        n19002), .Y(n20329) );
  A2O1A1Ixp33_ASAP7_75t_SL U22849 ( .A1(n31658), .A2(n24684), .B(n18295), .C(
        n24680), .Y(n20327) );
  A2O1A1Ixp33_ASAP7_75t_SL U22850 ( .A1(n20323), .A2(n20324), .B(n18295), .C(
        n19002), .Y(n24497) );
  A2O1A1Ixp33_ASAP7_75t_SL U22851 ( .A1(n24661), .A2(n29575), .B(n18295), .C(
        n19002), .Y(n20320) );
  A2O1A1Ixp33_ASAP7_75t_SL U22852 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__2_), .A2(
        n24648), .B(n18295), .C(n19002), .Y(n19519) );
  A2O1A1Ixp33_ASAP7_75t_SL U22853 ( .A1(n24495), .A2(n19520), .B(n18295), .C(
        n19002), .Y(n3544) );
  A2O1A1Ixp33_ASAP7_75t_SL U22854 ( .A1(n24660), .A2(n20318), .B(n18295), .C(
        n19002), .Y(n20319) );
  A2O1A1Ixp33_ASAP7_75t_SL U22855 ( .A1(n24661), .A2(n20316), .B(n18295), .C(
        n19002), .Y(n20317) );
  A2O1A1Ixp33_ASAP7_75t_SL U22856 ( .A1(n24662), .A2(n20314), .B(n18295), .C(
        n19002), .Y(n20315) );
  A2O1A1Ixp33_ASAP7_75t_SL U22857 ( .A1(n24676), .A2(n20071), .B(n18295), .C(
        n19002), .Y(n20072) );
  A2O1A1Ixp33_ASAP7_75t_SL U22858 ( .A1(n22421), .A2(n32186), .B(n18295), .C(
        n19002), .Y(n20312) );
  A2O1A1Ixp33_ASAP7_75t_SL U22859 ( .A1(n20311), .A2(n20312), .B(n18295), .C(
        n19002), .Y(n20313) );
  A2O1A1Ixp33_ASAP7_75t_SL U22860 ( .A1(n19002), .A2(n20313), .B(n18295), .C(
        n19002), .Y(n3160) );
  A2O1A1Ixp33_ASAP7_75t_SL U22861 ( .A1(n31258), .A2(n31259), .B(n18295), .C(
        n19002), .Y(n20306) );
  A2O1A1Ixp33_ASAP7_75t_SL U22862 ( .A1(n31573), .A2(n20307), .B(n18295), .C(
        n19002), .Y(n3131) );
  A2O1A1Ixp33_ASAP7_75t_SL U22863 ( .A1(uart1_r_BRATE__6_), .A2(n20300), .B(
        n18295), .C(n19002), .Y(n20301) );
  A2O1A1Ixp33_ASAP7_75t_SL U22864 ( .A1(n27308), .A2(n24694), .B(n18295), .C(
        n19002), .Y(n20283) );
  A2O1A1Ixp33_ASAP7_75t_SL U22865 ( .A1(n27327), .A2(n20283), .B(n18295), .C(
        n19002), .Y(n20284) );
  A2O1A1Ixp33_ASAP7_75t_SL U22866 ( .A1(n32591), .A2(n20273), .B(n18295), .C(
        n19002), .Y(n20274) );
  A2O1A1Ixp33_ASAP7_75t_SL U22867 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__10_), 
        .A2(n32447), .B(n18295), .C(n19002), .Y(n19672) );
  A2O1A1Ixp33_ASAP7_75t_SL U22868 ( .A1(n32446), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[43]), .B(n18295), .C(n19002), .Y(n19673) );
  A2O1A1Ixp33_ASAP7_75t_SL U22869 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[10]), 
        .A2(n32448), .B(n18295), .C(n19002), .Y(n19674) );
  A2O1A1Ixp33_ASAP7_75t_SL U22870 ( .A1(n19672), .A2(n19673), .B(n18295), .C(
        n19674), .Y(n19675) );
  A2O1A1Ixp33_ASAP7_75t_SL U22871 ( .A1(n33067), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__5_), .B(n18295), .C(n19002), 
        .Y(n19677) );
  A2O1A1Ixp33_ASAP7_75t_SL U22872 ( .A1(n32385), .A2(dc_q[22]), .B(n18295), 
        .C(n19002), .Y(n20268) );
  A2O1A1Ixp33_ASAP7_75t_SL U22873 ( .A1(n20267), .A2(n20268), .B(n18295), .C(
        n19002), .Y(n20269) );
  A2O1A1Ixp33_ASAP7_75t_SL U22874 ( .A1(n32386), .A2(n32423), .B(n18295), .C(
        n19002), .Y(n20271) );
  A2O1A1Ixp33_ASAP7_75t_SL U22875 ( .A1(n20270), .A2(n20271), .B(n18295), .C(
        n19002), .Y(dc_data[22]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22876 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__19_), 
        .A2(n32214), .B(n18295), .C(n19002), .Y(n20261) );
  A2O1A1Ixp33_ASAP7_75t_SL U22877 ( .A1(n20260), .A2(n20261), .B(n18295), .C(
        n19002), .Y(n20262) );
  A2O1A1Ixp33_ASAP7_75t_SL U22878 ( .A1(n19002), .A2(n20262), .B(n18295), .C(
        n19002), .Y(n20263) );
  A2O1A1Ixp33_ASAP7_75t_SL U22879 ( .A1(n28001), .A2(uart1_r_THOLD__21__7_), 
        .B(n18295), .C(n19002), .Y(n20207) );
  A2O1A1Ixp33_ASAP7_75t_SL U22880 ( .A1(n27998), .A2(uart1_r_THOLD__25__7_), 
        .B(n18295), .C(n19002), .Y(n20208) );
  A2O1A1Ixp33_ASAP7_75t_SL U22881 ( .A1(n27999), .A2(uart1_r_THOLD__17__7_), 
        .B(n18295), .C(n19002), .Y(n20209) );
  A2O1A1Ixp33_ASAP7_75t_SL U22882 ( .A1(n20207), .A2(n20208), .B(n18295), .C(
        n20209), .Y(n20210) );
  A2O1A1Ixp33_ASAP7_75t_SL U22883 ( .A1(n28003), .A2(uart1_r_THOLD__1__7_), 
        .B(n18295), .C(n19002), .Y(n20212) );
  A2O1A1Ixp33_ASAP7_75t_SL U22884 ( .A1(n27996), .A2(uart1_r_THOLD__29__7_), 
        .B(n18295), .C(n19002), .Y(n20213) );
  A2O1A1Ixp33_ASAP7_75t_SL U22885 ( .A1(n27997), .A2(uart1_r_THOLD__13__7_), 
        .B(n18295), .C(n19002), .Y(n20214) );
  A2O1A1Ixp33_ASAP7_75t_SL U22886 ( .A1(n20212), .A2(n20213), .B(n18295), .C(
        n20214), .Y(n20215) );
  A2O1A1Ixp33_ASAP7_75t_SL U22887 ( .A1(n20211), .A2(n20216), .B(n18295), .C(
        n19002), .Y(n20217) );
  A2O1A1Ixp33_ASAP7_75t_SL U22888 ( .A1(n28011), .A2(uart1_r_THOLD__20__7_), 
        .B(n18295), .C(n19002), .Y(n20219) );
  A2O1A1Ixp33_ASAP7_75t_SL U22889 ( .A1(uart1_r_THOLD__12__7_), .A2(n20220), 
        .B(n18295), .C(n19002), .Y(n20221) );
  A2O1A1Ixp33_ASAP7_75t_SL U22890 ( .A1(n20218), .A2(n20219), .B(n18295), .C(
        n20221), .Y(n20222) );
  A2O1A1Ixp33_ASAP7_75t_SL U22891 ( .A1(n28008), .A2(uart1_r_THOLD__0__7_), 
        .B(n18295), .C(n19002), .Y(n20224) );
  A2O1A1Ixp33_ASAP7_75t_SL U22892 ( .A1(n28015), .A2(uart1_r_THOLD__4__7_), 
        .B(n18295), .C(n19002), .Y(n20225) );
  A2O1A1Ixp33_ASAP7_75t_SL U22893 ( .A1(n28009), .A2(uart1_r_THOLD__8__7_), 
        .B(n18295), .C(n19002), .Y(n20226) );
  A2O1A1Ixp33_ASAP7_75t_SL U22894 ( .A1(n20224), .A2(n20225), .B(n18295), .C(
        n20226), .Y(n20227) );
  A2O1A1Ixp33_ASAP7_75t_SL U22895 ( .A1(n20223), .A2(n20228), .B(n18295), .C(
        n19002), .Y(n20229) );
  A2O1A1Ixp33_ASAP7_75t_SL U22896 ( .A1(n27999), .A2(uart1_r_THOLD__19__7_), 
        .B(n18295), .C(n19002), .Y(n20230) );
  A2O1A1Ixp33_ASAP7_75t_SL U22897 ( .A1(n27996), .A2(uart1_r_THOLD__31__7_), 
        .B(n18295), .C(n19002), .Y(n20231) );
  A2O1A1Ixp33_ASAP7_75t_SL U22898 ( .A1(n27997), .A2(uart1_r_THOLD__15__7_), 
        .B(n18295), .C(n19002), .Y(n20232) );
  A2O1A1Ixp33_ASAP7_75t_SL U22899 ( .A1(n20230), .A2(n20231), .B(n18295), .C(
        n20232), .Y(n20233) );
  A2O1A1Ixp33_ASAP7_75t_SL U22900 ( .A1(n28003), .A2(uart1_r_THOLD__3__7_), 
        .B(n18295), .C(n19002), .Y(n20235) );
  A2O1A1Ixp33_ASAP7_75t_SL U22901 ( .A1(n28001), .A2(uart1_r_THOLD__23__7_), 
        .B(n18295), .C(n19002), .Y(n20236) );
  A2O1A1Ixp33_ASAP7_75t_SL U22902 ( .A1(n28000), .A2(uart1_r_THOLD__11__7_), 
        .B(n18295), .C(n19002), .Y(n20237) );
  A2O1A1Ixp33_ASAP7_75t_SL U22903 ( .A1(n20235), .A2(n20236), .B(n18295), .C(
        n20237), .Y(n20238) );
  A2O1A1Ixp33_ASAP7_75t_SL U22904 ( .A1(n20234), .A2(n20239), .B(n18295), .C(
        n19002), .Y(n20240) );
  A2O1A1Ixp33_ASAP7_75t_SL U22905 ( .A1(uart1_r_THOLD__14__7_), .A2(n20220), 
        .B(n18295), .C(n19002), .Y(n20242) );
  A2O1A1Ixp33_ASAP7_75t_SL U22906 ( .A1(n28015), .A2(uart1_r_THOLD__6__7_), 
        .B(n18295), .C(n19002), .Y(n20243) );
  A2O1A1Ixp33_ASAP7_75t_SL U22907 ( .A1(n20241), .A2(n20242), .B(n18295), .C(
        n20243), .Y(n20244) );
  A2O1A1Ixp33_ASAP7_75t_SL U22908 ( .A1(n28010), .A2(uart1_r_THOLD__18__7_), 
        .B(n18295), .C(n19002), .Y(n20246) );
  A2O1A1Ixp33_ASAP7_75t_SL U22909 ( .A1(n28011), .A2(uart1_r_THOLD__22__7_), 
        .B(n18295), .C(n19002), .Y(n20247) );
  A2O1A1Ixp33_ASAP7_75t_SL U22910 ( .A1(n20245), .A2(n20246), .B(n18295), .C(
        n20247), .Y(n20248) );
  A2O1A1Ixp33_ASAP7_75t_SL U22911 ( .A1(n28008), .A2(uart1_r_THOLD__2__7_), 
        .B(n18295), .C(n19002), .Y(n20250) );
  A2O1A1Ixp33_ASAP7_75t_SL U22912 ( .A1(n28009), .A2(uart1_r_THOLD__10__7_), 
        .B(n18295), .C(n19002), .Y(n20251) );
  A2O1A1Ixp33_ASAP7_75t_SL U22913 ( .A1(n20249), .A2(n20250), .B(n18295), .C(
        n20251), .Y(n20252) );
  A2O1A1Ixp33_ASAP7_75t_SL U22914 ( .A1(n31392), .A2(
        u0_0_leon3x0_p0_iu_r_W__RESULT__16_), .B(n18295), .C(n19002), .Y(
        n20204) );
  A2O1A1Ixp33_ASAP7_75t_SL U22915 ( .A1(rf_do_a[16]), .A2(n31391), .B(n18295), 
        .C(n19002), .Y(n20205) );
  A2O1A1Ixp33_ASAP7_75t_SL U22916 ( .A1(n20204), .A2(n20205), .B(n18295), .C(
        n19002), .Y(n20206) );
  A2O1A1Ixp33_ASAP7_75t_SL U22917 ( .A1(DP_OP_1196_128_7433_n95), .A2(
        DP_OP_1196_128_7433_n98), .B(n18295), .C(n20201), .Y(n20202) );
  A2O1A1Ixp33_ASAP7_75t_SL U22918 ( .A1(add_x_735_A_2_), .A2(n28131), .B(
        n18295), .C(n19002), .Y(n20195) );
  A2O1A1Ixp33_ASAP7_75t_SL U22919 ( .A1(n27489), .A2(n30639), .B(n18295), .C(
        n20195), .Y(n20196) );
  A2O1A1Ixp33_ASAP7_75t_SL U22920 ( .A1(n18593), .A2(n22418), .B(n18295), .C(
        n19002), .Y(n20194) );
  A2O1A1Ixp33_ASAP7_75t_SL U22921 ( .A1(DP_OP_5187J1_124_3275_n301), .A2(
        n24317), .B(n18295), .C(n20192), .Y(n20193) );
  A2O1A1Ixp33_ASAP7_75t_SL U22922 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[32]), 
        .B(n18295), .C(n19002), .Y(n20191) );
  A2O1A1Ixp33_ASAP7_75t_SL U22923 ( .A1(n20187), .A2(n20188), .B(n18295), .C(
        n19002), .Y(n20189) );
  A2O1A1Ixp33_ASAP7_75t_SL U22924 ( .A1(n22373), .A2(u0_0_leon3x0_p0_divi[31]), 
        .B(n18295), .C(n19002), .Y(n20186) );
  A2O1A1Ixp33_ASAP7_75t_SL U22925 ( .A1(n31458), .A2(n30199), .B(n18295), .C(
        n19002), .Y(n20185) );
  A2O1A1Ixp33_ASAP7_75t_SL U22926 ( .A1(n29059), .A2(u0_0_leon3x0_p0_ici[41]), 
        .B(n18295), .C(n19002), .Y(n20181) );
  A2O1A1Ixp33_ASAP7_75t_SL U22927 ( .A1(n20180), .A2(n20181), .B(n18295), .C(
        n19002), .Y(n20182) );
  A2O1A1Ixp33_ASAP7_75t_SL U22928 ( .A1(n19002), .A2(n20182), .B(n18295), .C(
        n19002), .Y(n20183) );
  A2O1A1Ixp33_ASAP7_75t_SL U22929 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__13_), .B(n18295), .C(n19002), .Y(
        n20179) );
  A2O1A1Ixp33_ASAP7_75t_SL U22930 ( .A1(n32808), .A2(n20178), .B(n18295), .C(
        n19002), .Y(n32796) );
  A2O1A1Ixp33_ASAP7_75t_SL U22931 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[45]), 
        .B(n18295), .C(n19002), .Y(n19793) );
  A2O1A1Ixp33_ASAP7_75t_SL U22932 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__13_), .B(n18295), .C(n19002), .Y(n19794) );
  A2O1A1Ixp33_ASAP7_75t_SL U22933 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[44]), 
        .B(n18295), .C(n19002), .Y(n19797) );
  A2O1A1Ixp33_ASAP7_75t_SL U22934 ( .A1(n19793), .A2(n19796), .B(n18295), .C(
        n19797), .Y(u0_0_leon3x0_p0_div0_vaddin1[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22935 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__25_), .B(n18295), .C(n19002), .Y(n20167) );
  A2O1A1Ixp33_ASAP7_75t_SL U22936 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[57]), 
        .B(n18295), .C(n19002), .Y(n20170) );
  A2O1A1Ixp33_ASAP7_75t_SL U22937 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[56]), 
        .B(n18295), .C(n19002), .Y(n20171) );
  A2O1A1Ixp33_ASAP7_75t_SL U22938 ( .A1(n20169), .A2(n20170), .B(n18295), .C(
        n20171), .Y(u0_0_leon3x0_p0_div0_vaddin1[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22939 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__28_), .B(n18295), .C(n19002), .Y(n20162) );
  A2O1A1Ixp33_ASAP7_75t_SL U22940 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[60]), 
        .B(n18295), .C(n19002), .Y(n20165) );
  A2O1A1Ixp33_ASAP7_75t_SL U22941 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[59]), 
        .B(n18295), .C(n19002), .Y(n20166) );
  A2O1A1Ixp33_ASAP7_75t_SL U22942 ( .A1(n20164), .A2(n20165), .B(n18295), .C(
        n20166), .Y(u0_0_leon3x0_p0_div0_vaddin1[29]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22943 ( .A1(n24046), .A2(n22642), .B(n18295), .C(
        n19002), .Y(n20155) );
  A2O1A1Ixp33_ASAP7_75t_SL U22944 ( .A1(n20154), .A2(n20155), .B(n18295), .C(
        n19002), .Y(n20156) );
  A2O1A1Ixp33_ASAP7_75t_SL U22945 ( .A1(n19002), .A2(n20156), .B(n18295), .C(
        n19002), .Y(mult_x_1196_n844) );
  A2O1A1Ixp33_ASAP7_75t_SL U22946 ( .A1(sr1_r_MCFG2__RAMRWS__0_), .A2(n20144), 
        .B(n18295), .C(n19002), .Y(n20145) );
  A2O1A1Ixp33_ASAP7_75t_SL U22947 ( .A1(n29948), .A2(n20137), .B(n18295), .C(
        n19002), .Y(n20138) );
  A2O1A1Ixp33_ASAP7_75t_SL U22948 ( .A1(n30205), .A2(n32195), .B(n18295), .C(
        n19002), .Y(n20120) );
  A2O1A1Ixp33_ASAP7_75t_SL U22949 ( .A1(n30208), .A2(n30209), .B(n18295), .C(
        n19002), .Y(n20123) );
  A2O1A1Ixp33_ASAP7_75t_SL U22950 ( .A1(n30640), .A2(rf_do_b[23]), .B(n18295), 
        .C(n19002), .Y(n20111) );
  A2O1A1Ixp33_ASAP7_75t_SL U22951 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__23_), .B(n18295), .C(n19002), .Y(n20112)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U22952 ( .A1(n20111), .A2(n20112), .B(n18295), .C(
        n19002), .Y(n20113) );
  A2O1A1Ixp33_ASAP7_75t_SL U22953 ( .A1(n20116), .A2(n30593), .B(n18295), .C(
        n19002), .Y(n20117) );
  A2O1A1Ixp33_ASAP7_75t_SL U22954 ( .A1(u0_0_leon3x0_p0_divi[59]), .A2(n30430), 
        .B(n18295), .C(n19002), .Y(n20106) );
  A2O1A1Ixp33_ASAP7_75t_SL U22955 ( .A1(n20105), .A2(n20106), .B(n18295), .C(
        n19002), .Y(n20107) );
  A2O1A1Ixp33_ASAP7_75t_SL U22956 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[61]), 
        .B(n18295), .C(n19002), .Y(n20100) );
  A2O1A1Ixp33_ASAP7_75t_SL U22957 ( .A1(n20099), .A2(n20100), .B(n18295), .C(
        n19002), .Y(n20101) );
  A2O1A1Ixp33_ASAP7_75t_SL U22958 ( .A1(n24669), .A2(n26285), .B(n18295), .C(
        n19002), .Y(n19743) );
  A2O1A1Ixp33_ASAP7_75t_SL U22959 ( .A1(n24675), .A2(n19889), .B(n18295), .C(
        n19002), .Y(n19890) );
  A2O1A1Ixp33_ASAP7_75t_SL U22960 ( .A1(n31626), .A2(n20095), .B(n18295), .C(
        n20096), .Y(n10972) );
  A2O1A1Ixp33_ASAP7_75t_SL U22961 ( .A1(n30684), .A2(n24662), .B(n18295), .C(
        n19002), .Y(n19531) );
  A2O1A1Ixp33_ASAP7_75t_SL U22962 ( .A1(n24668), .A2(n20093), .B(n18295), .C(
        n19002), .Y(n20094) );
  A2O1A1Ixp33_ASAP7_75t_SL U22963 ( .A1(n24670), .A2(n19722), .B(n18295), .C(
        n19002), .Y(n19723) );
  A2O1A1Ixp33_ASAP7_75t_SL U22964 ( .A1(n19002), .A2(n24908), .B(n18295), .C(
        n19002), .Y(n20085) );
  A2O1A1Ixp33_ASAP7_75t_SL U22965 ( .A1(u0_0_leon3x0_p0_div0_r_CNT__0_), .A2(
        n20085), .B(n18295), .C(n19002), .Y(n20086) );
  A2O1A1Ixp33_ASAP7_75t_SL U22966 ( .A1(n19002), .A2(n20086), .B(n18295), .C(
        n19002), .Y(n20087) );
  A2O1A1Ixp33_ASAP7_75t_SL U22967 ( .A1(n19002), .A2(n24646), .B(n18295), .C(
        n19002), .Y(n20080) );
  A2O1A1Ixp33_ASAP7_75t_SL U22968 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__6_), .A2(n20080), .B(n18295), .C(n19002), .Y(n20081) );
  A2O1A1Ixp33_ASAP7_75t_SL U22969 ( .A1(n19002), .A2(n20081), .B(n18295), .C(
        n19002), .Y(n20082) );
  A2O1A1Ixp33_ASAP7_75t_SL U22970 ( .A1(n24674), .A2(n20078), .B(n18295), .C(
        n19002), .Y(n20079) );
  A2O1A1Ixp33_ASAP7_75t_SL U22971 ( .A1(n24668), .A2(n26819), .B(n18295), .C(
        n19002), .Y(n19712) );
  A2O1A1Ixp33_ASAP7_75t_SL U22972 ( .A1(u0_0_leon3x0_p0_iu_r_A__RFA2__0_), 
        .A2(n24662), .B(n18295), .C(n19002), .Y(n19709) );
  A2O1A1Ixp33_ASAP7_75t_SL U22973 ( .A1(n24660), .A2(n20076), .B(n18295), .C(
        n19002), .Y(n20077) );
  A2O1A1Ixp33_ASAP7_75t_SL U22974 ( .A1(n31347), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n20075) );
  A2O1A1Ixp33_ASAP7_75t_SL U22975 ( .A1(n31260), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n19702) );
  A2O1A1Ixp33_ASAP7_75t_SL U22976 ( .A1(n19002), .A2(n20068), .B(n18295), .C(
        n19002), .Y(n20069) );
  A2O1A1Ixp33_ASAP7_75t_SL U22977 ( .A1(n19002), .A2(n20070), .B(n18295), .C(
        n19002), .Y(n30914) );
  A2O1A1Ixp33_ASAP7_75t_SL U22978 ( .A1(n24592), .A2(n24607), .B(n18295), .C(
        n19002), .Y(n19861) );
  A2O1A1Ixp33_ASAP7_75t_SL U22979 ( .A1(n24604), .A2(n24605), .B(n18295), .C(
        n19862), .Y(n19863) );
  A2O1A1Ixp33_ASAP7_75t_SL U22980 ( .A1(u0_0_leon3x0_p0_divi[31]), .A2(n31662), 
        .B(n18295), .C(n19002), .Y(n20059) );
  A2O1A1Ixp33_ASAP7_75t_SL U22981 ( .A1(n18295), .A2(n19002), .B(n19683), .C(
        n19002), .Y(n19684) );
  A2O1A1Ixp33_ASAP7_75t_SL U22982 ( .A1(n18295), .A2(n19002), .B(n19844), .C(
        n19002), .Y(n19845) );
  A2O1A1Ixp33_ASAP7_75t_SL U22983 ( .A1(n32583), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__3_), .B(n18295), .C(n19002), 
        .Y(n20048) );
  A2O1A1Ixp33_ASAP7_75t_SL U22984 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__8_), 
        .A2(n32584), .B(n18295), .C(n19002), .Y(n20049) );
  A2O1A1Ixp33_ASAP7_75t_SL U22985 ( .A1(n20048), .A2(n20049), .B(n18295), .C(
        n19002), .Y(n20050) );
  A2O1A1Ixp33_ASAP7_75t_SL U22986 ( .A1(n32578), .A2(n32588), .B(n18295), .C(
        n19002), .Y(n20052) );
  A2O1A1Ixp33_ASAP7_75t_SL U22987 ( .A1(n20051), .A2(n20052), .B(n18295), .C(
        n19002), .Y(ic_address[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22988 ( .A1(n32615), .A2(n32660), .B(n18295), .C(
        n19002), .Y(n19831) );
  A2O1A1Ixp33_ASAP7_75t_SL U22989 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[28]), 
        .A2(n32231), .B(n18295), .C(n19002), .Y(n20040) );
  A2O1A1Ixp33_ASAP7_75t_SL U22990 ( .A1(n20039), .A2(n20040), .B(n18295), .C(
        n19002), .Y(dt_data[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22991 ( .A1(n30726), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__22_), .B(n18295), .C(n19002), .Y(
        n20031) );
  A2O1A1Ixp33_ASAP7_75t_SL U22992 ( .A1(n29074), .A2(n32162), .B(n18295), .C(
        n19002), .Y(n20032) );
  A2O1A1Ixp33_ASAP7_75t_SL U22993 ( .A1(n30722), .A2(u0_0_leon3x0_p0_ici[19]), 
        .B(n18295), .C(n19002), .Y(n20033) );
  A2O1A1Ixp33_ASAP7_75t_SL U22994 ( .A1(n20031), .A2(n20032), .B(n18295), .C(
        n20033), .Y(n20034) );
  A2O1A1Ixp33_ASAP7_75t_SL U22995 ( .A1(n30723), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__22_), .B(n18295), .C(n19002), .Y(
        n20036) );
  A2O1A1Ixp33_ASAP7_75t_SL U22996 ( .A1(n30724), .A2(u0_0_leon3x0_p0_ici[50]), 
        .B(n18295), .C(n19002), .Y(n20037) );
  A2O1A1Ixp33_ASAP7_75t_SL U22997 ( .A1(n20035), .A2(n20036), .B(n18295), .C(
        n20037), .Y(rf_di_w[22]) );
  A2O1A1Ixp33_ASAP7_75t_SL U22998 ( .A1(n31392), .A2(
        u0_0_leon3x0_p0_iu_r_W__RESULT__15_), .B(n18295), .C(n19002), .Y(
        n20028) );
  A2O1A1Ixp33_ASAP7_75t_SL U22999 ( .A1(rf_do_a[15]), .A2(n31391), .B(n18295), 
        .C(n19002), .Y(n20029) );
  A2O1A1Ixp33_ASAP7_75t_SL U23000 ( .A1(n20028), .A2(n20029), .B(n18295), .C(
        n19002), .Y(n20030) );
  A2O1A1Ixp33_ASAP7_75t_SL U23001 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__25_), .B(n18295), .C(n19002), .Y(
        n20026) );
  A2O1A1Ixp33_ASAP7_75t_SL U23002 ( .A1(DP_OP_5187J1_124_3275_n249), .A2(
        DP_OP_5187J1_124_3275_n329), .B(n18295), .C(n19002), .Y(n20019) );
  A2O1A1Ixp33_ASAP7_75t_SL U23003 ( .A1(DP_OP_5187J1_124_3275_n250), .A2(
        DP_OP_5187J1_124_3275_n329), .B(n18295), .C(n19002), .Y(n20021) );
  A2O1A1Ixp33_ASAP7_75t_SL U23004 ( .A1(DP_OP_5187J1_124_3275_n245), .A2(
        n20021), .B(n18295), .C(n19002), .Y(n20022) );
  A2O1A1Ixp33_ASAP7_75t_SL U23005 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__11_), .B(n18295), .C(n19002), .Y(
        n20018) );
  A2O1A1Ixp33_ASAP7_75t_SL U23006 ( .A1(DP_OP_1196_128_7433_n8), .A2(
        DP_OP_1196_128_7433_n84), .B(n18295), .C(n19002), .Y(n20014) );
  A2O1A1Ixp33_ASAP7_75t_SL U23007 ( .A1(n32176), .A2(n32177), .B(n18295), .C(
        n19002), .Y(n20009) );
  A2O1A1Ixp33_ASAP7_75t_SL U23008 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__29_), 
        .A2(n29060), .B(n18295), .C(n19002), .Y(n19033) );
  A2O1A1Ixp33_ASAP7_75t_SL U23009 ( .A1(n29059), .A2(u0_0_leon3x0_p0_ici[43]), 
        .B(n18295), .C(n19002), .Y(n20002) );
  A2O1A1Ixp33_ASAP7_75t_SL U23010 ( .A1(n20001), .A2(n20002), .B(n18295), .C(
        n19002), .Y(n20003) );
  A2O1A1Ixp33_ASAP7_75t_SL U23011 ( .A1(n19002), .A2(n20003), .B(n18295), .C(
        n19002), .Y(n20004) );
  A2O1A1Ixp33_ASAP7_75t_SL U23012 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__24_), .B(n18295), .C(n19002), .Y(
        n19439) );
  A2O1A1Ixp33_ASAP7_75t_SL U23013 ( .A1(n24931), .A2(n19019), .B(n18295), .C(
        n19002), .Y(n24964) );
  A2O1A1Ixp33_ASAP7_75t_SL U23014 ( .A1(n28977), .A2(n25469), .B(n18295), .C(
        n19002), .Y(n19995) );
  A2O1A1Ixp33_ASAP7_75t_SL U23015 ( .A1(n26423), .A2(n24575), .B(n18295), .C(
        n19002), .Y(n19996) );
  A2O1A1Ixp33_ASAP7_75t_SL U23016 ( .A1(n19995), .A2(n19996), .B(n18295), .C(
        n19002), .Y(n19997) );
  A2O1A1Ixp33_ASAP7_75t_SL U23017 ( .A1(n28967), .A2(n25470), .B(n18295), .C(
        n19002), .Y(n19999) );
  A2O1A1Ixp33_ASAP7_75t_SL U23018 ( .A1(n19998), .A2(n19999), .B(n18295), .C(
        n19002), .Y(n26937) );
  A2O1A1Ixp33_ASAP7_75t_SL U23019 ( .A1(n19998), .A2(n19999), .B(n18295), .C(
        n19002), .Y(n18794) );
  A2O1A1Ixp33_ASAP7_75t_SL U23020 ( .A1(n26023), .A2(uart1_r_RWADDR__0_), .B(
        n18295), .C(n19002), .Y(n19990) );
  A2O1A1Ixp33_ASAP7_75t_SL U23021 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__15_), .B(n18295), .C(n19002), .Y(n19980) );
  A2O1A1Ixp33_ASAP7_75t_SL U23022 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[46]), 
        .B(n18295), .C(n19002), .Y(n19983) );
  A2O1A1Ixp33_ASAP7_75t_SL U23023 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[47]), 
        .B(n18295), .C(n19002), .Y(n19984) );
  A2O1A1Ixp33_ASAP7_75t_SL U23024 ( .A1(n19982), .A2(n19983), .B(n18295), .C(
        n19984), .Y(u0_0_leon3x0_p0_div0_vaddin1[16]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23025 ( .A1(n32696), .A2(n32704), .B(n18295), .C(
        n24694), .Y(n19975) );
  A2O1A1Ixp33_ASAP7_75t_SL U23026 ( .A1(n31199), .A2(apb0_r_CFGSEL_), .B(
        n18295), .C(n19002), .Y(n19917) );
  A2O1A1Ixp33_ASAP7_75t_SL U23027 ( .A1(n31249), .A2(irqctrl0_r_IMASK__0__6_), 
        .B(n18295), .C(n19002), .Y(n19921) );
  A2O1A1Ixp33_ASAP7_75t_SL U23028 ( .A1(n31247), .A2(irqctrl0_r_IPEND__6_), 
        .B(n18295), .C(n19002), .Y(n19922) );
  A2O1A1Ixp33_ASAP7_75t_SL U23029 ( .A1(n19920), .A2(n19921), .B(n18295), .C(
        n19922), .Y(n19923) );
  A2O1A1Ixp33_ASAP7_75t_SL U23030 ( .A1(timer0_r_SCALER__6_), .A2(n31245), .B(
        n18295), .C(n19002), .Y(n19924) );
  A2O1A1Ixp33_ASAP7_75t_SL U23031 ( .A1(uart1_r_FRAME_), .A2(n31951), .B(
        n18295), .C(n19002), .Y(n19925) );
  A2O1A1Ixp33_ASAP7_75t_SL U23032 ( .A1(n31246), .A2(uart1_r_BRATE__6_), .B(
        n18295), .C(n19002), .Y(n19926) );
  A2O1A1Ixp33_ASAP7_75t_SL U23033 ( .A1(n19924), .A2(n19925), .B(n18295), .C(
        n19926), .Y(n19927) );
  A2O1A1Ixp33_ASAP7_75t_SL U23034 ( .A1(n31250), .A2(sr1_r_MCFG2__RMW_), .B(
        n18295), .C(n19002), .Y(n19929) );
  A2O1A1Ixp33_ASAP7_75t_SL U23035 ( .A1(n31251), .A2(irqctrl0_r_IFORCE__0__6_), 
        .B(n18295), .C(n19002), .Y(n19930) );
  A2O1A1Ixp33_ASAP7_75t_SL U23036 ( .A1(n19928), .A2(n19929), .B(n18295), .C(
        n19930), .Y(n19931) );
  A2O1A1Ixp33_ASAP7_75t_SL U23037 ( .A1(n31233), .A2(n31234), .B(n18295), .C(
        n19002), .Y(n19933) );
  A2O1A1Ixp33_ASAP7_75t_SL U23038 ( .A1(n31231), .A2(n31232), .B(n18295), .C(
        n19002), .Y(n19934) );
  A2O1A1Ixp33_ASAP7_75t_SL U23039 ( .A1(n31209), .A2(uart1_r_RHOLD__25__6_), 
        .B(n18295), .C(n19002), .Y(n19935) );
  A2O1A1Ixp33_ASAP7_75t_SL U23040 ( .A1(n31206), .A2(uart1_r_RHOLD__17__6_), 
        .B(n18295), .C(n19002), .Y(n19936) );
  A2O1A1Ixp33_ASAP7_75t_SL U23041 ( .A1(n31207), .A2(uart1_r_RHOLD__7__6_), 
        .B(n18295), .C(n19002), .Y(n19937) );
  A2O1A1Ixp33_ASAP7_75t_SL U23042 ( .A1(n19935), .A2(n19936), .B(n18295), .C(
        n19937), .Y(n19938) );
  A2O1A1Ixp33_ASAP7_75t_SL U23043 ( .A1(n31213), .A2(uart1_r_RHOLD__15__6_), 
        .B(n18295), .C(n19002), .Y(n19940) );
  A2O1A1Ixp33_ASAP7_75t_SL U23044 ( .A1(n31210), .A2(uart1_r_RHOLD__21__6_), 
        .B(n18295), .C(n19002), .Y(n19941) );
  A2O1A1Ixp33_ASAP7_75t_SL U23045 ( .A1(n31211), .A2(uart1_r_RHOLD__20__6_), 
        .B(n18295), .C(n19002), .Y(n19942) );
  A2O1A1Ixp33_ASAP7_75t_SL U23046 ( .A1(n19940), .A2(n19941), .B(n18295), .C(
        n19942), .Y(n19943) );
  A2O1A1Ixp33_ASAP7_75t_SL U23047 ( .A1(n31200), .A2(uart1_r_RHOLD__5__6_), 
        .B(n18295), .C(n19002), .Y(n19945) );
  A2O1A1Ixp33_ASAP7_75t_SL U23048 ( .A1(n31201), .A2(uart1_r_RHOLD__30__6_), 
        .B(n18295), .C(n19002), .Y(n19946) );
  A2O1A1Ixp33_ASAP7_75t_SL U23049 ( .A1(n19945), .A2(n19946), .B(n18295), .C(
        n19002), .Y(n19947) );
  A2O1A1Ixp33_ASAP7_75t_SL U23050 ( .A1(n31202), .A2(uart1_r_RHOLD__12__6_), 
        .B(n18295), .C(n19002), .Y(n19949) );
  A2O1A1Ixp33_ASAP7_75t_SL U23051 ( .A1(n31203), .A2(uart1_r_RHOLD__14__6_), 
        .B(n18295), .C(n19002), .Y(n19950) );
  A2O1A1Ixp33_ASAP7_75t_SL U23052 ( .A1(n19948), .A2(n19949), .B(n18295), .C(
        n19950), .Y(n19951) );
  A2O1A1Ixp33_ASAP7_75t_SL U23053 ( .A1(n31218), .A2(uart1_r_RHOLD__23__6_), 
        .B(n18295), .C(n19002), .Y(n19952) );
  A2O1A1Ixp33_ASAP7_75t_SL U23054 ( .A1(n31219), .A2(uart1_r_RHOLD__11__6_), 
        .B(n18295), .C(n19002), .Y(n19953) );
  A2O1A1Ixp33_ASAP7_75t_SL U23055 ( .A1(n19952), .A2(n19953), .B(n18295), .C(
        n19002), .Y(n19954) );
  A2O1A1Ixp33_ASAP7_75t_SL U23056 ( .A1(n31216), .A2(uart1_r_RHOLD__3__6_), 
        .B(n18295), .C(n19002), .Y(n19955) );
  A2O1A1Ixp33_ASAP7_75t_SL U23057 ( .A1(n31217), .A2(uart1_r_RHOLD__29__6_), 
        .B(n18295), .C(n19002), .Y(n19956) );
  A2O1A1Ixp33_ASAP7_75t_SL U23058 ( .A1(n31222), .A2(n19955), .B(n18295), .C(
        n19956), .Y(n19957) );
  A2O1A1Ixp33_ASAP7_75t_SL U23059 ( .A1(n31214), .A2(uart1_r_RHOLD__1__6_), 
        .B(n18295), .C(n19002), .Y(n19959) );
  A2O1A1Ixp33_ASAP7_75t_SL U23060 ( .A1(n31215), .A2(uart1_r_RHOLD__28__6_), 
        .B(n18295), .C(n19002), .Y(n19960) );
  A2O1A1Ixp33_ASAP7_75t_SL U23061 ( .A1(n19958), .A2(n19959), .B(n18295), .C(
        n19960), .Y(n19961) );
  A2O1A1Ixp33_ASAP7_75t_SL U23062 ( .A1(n19939), .A2(n19944), .B(n18295), .C(
        n19962), .Y(n19963) );
  A2O1A1Ixp33_ASAP7_75t_SL U23063 ( .A1(n31235), .A2(sr1_r_MCFG1__ROMWWS__2_), 
        .B(n18295), .C(n19002), .Y(n19965) );
  A2O1A1Ixp33_ASAP7_75t_SL U23064 ( .A1(n31236), .A2(n19965), .B(n18295), .C(
        n19002), .Y(n19966) );
  A2O1A1Ixp33_ASAP7_75t_SL U23065 ( .A1(uart1_r_RHOLD__0__6_), .A2(n31242), 
        .B(n18295), .C(n19002), .Y(n19970) );
  A2O1A1Ixp33_ASAP7_75t_SL U23066 ( .A1(n19969), .A2(n19970), .B(n18295), .C(
        n19002), .Y(n19971) );
  A2O1A1Ixp33_ASAP7_75t_SL U23067 ( .A1(n19932), .A2(n19972), .B(n18295), .C(
        n19002), .Y(n19973) );
  A2O1A1Ixp33_ASAP7_75t_SL U23068 ( .A1(n19760), .A2(n19761), .B(n18295), .C(
        n19002), .Y(n19762) );
  A2O1A1Ixp33_ASAP7_75t_SL U23069 ( .A1(n19763), .A2(n19764), .B(n18295), .C(
        n19002), .Y(n19765) );
  A2O1A1Ixp33_ASAP7_75t_SL U23070 ( .A1(n31670), .A2(n31669), .B(n18295), .C(
        n19002), .Y(n19766) );
  A2O1A1Ixp33_ASAP7_75t_SL U23071 ( .A1(n31672), .A2(n31671), .B(n18295), .C(
        n19002), .Y(n19767) );
  A2O1A1Ixp33_ASAP7_75t_SL U23072 ( .A1(n31666), .A2(n31665), .B(n18295), .C(
        n19768), .Y(n19769) );
  A2O1A1Ixp33_ASAP7_75t_SL U23073 ( .A1(n19771), .A2(n19772), .B(n18295), .C(
        n19002), .Y(n19773) );
  A2O1A1Ixp33_ASAP7_75t_SL U23074 ( .A1(n19774), .A2(n19775), .B(n18295), .C(
        n19002), .Y(n19776) );
  A2O1A1Ixp33_ASAP7_75t_SL U23075 ( .A1(n22379), .A2(n19750), .B(n18295), .C(
        n19002), .Y(n19751) );
  A2O1A1Ixp33_ASAP7_75t_SL U23076 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__9_), 
        .A2(n19752), .B(n18295), .C(n19002), .Y(n19753) );
  A2O1A1Ixp33_ASAP7_75t_SL U23077 ( .A1(n19746), .A2(n19756), .B(n18295), .C(
        n19002), .Y(n4443) );
  A2O1A1Ixp33_ASAP7_75t_SL U23078 ( .A1(n31478), .A2(n30024), .B(n18295), .C(
        n19002), .Y(n19907) );
  A2O1A1Ixp33_ASAP7_75t_SL U23079 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__5_), 
        .A2(n31364), .B(n18295), .C(n19002), .Y(n19908) );
  A2O1A1Ixp33_ASAP7_75t_SL U23080 ( .A1(n19907), .A2(n19908), .B(n18295), .C(
        n19002), .Y(n19909) );
  A2O1A1Ixp33_ASAP7_75t_SL U23081 ( .A1(n31479), .A2(n30025), .B(n18295), .C(
        n19002), .Y(n19911) );
  A2O1A1Ixp33_ASAP7_75t_SL U23082 ( .A1(n19910), .A2(n19911), .B(n18295), .C(
        n19002), .Y(n19912) );
  A2O1A1Ixp33_ASAP7_75t_SL U23083 ( .A1(n30640), .A2(rf_do_b[21]), .B(n18295), 
        .C(n19002), .Y(n19892) );
  A2O1A1Ixp33_ASAP7_75t_SL U23084 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__21_), .B(n18295), .C(n19002), .Y(n19893)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U23085 ( .A1(n19892), .A2(n19893), .B(n18295), .C(
        n19002), .Y(n19894) );
  A2O1A1Ixp33_ASAP7_75t_SL U23086 ( .A1(n19897), .A2(n30593), .B(n18295), .C(
        n19002), .Y(n19898) );
  A2O1A1Ixp33_ASAP7_75t_SL U23087 ( .A1(mult_x_1196_n752), .A2(n24272), .B(
        n18295), .C(n19738), .Y(n19739) );
  A2O1A1Ixp33_ASAP7_75t_SL U23088 ( .A1(n24272), .A2(mult_x_1196_n752), .B(
        n18295), .C(n19002), .Y(n19740) );
  A2O1A1Ixp33_ASAP7_75t_SL U23089 ( .A1(n22664), .A2(n19740), .B(n18295), .C(
        n19002), .Y(n19741) );
  A2O1A1Ixp33_ASAP7_75t_SL U23090 ( .A1(n19739), .A2(n19741), .B(n18295), .C(
        n19002), .Y(n19742) );
  A2O1A1Ixp33_ASAP7_75t_SL U23091 ( .A1(n32642), .A2(n24677), .B(n18295), .C(
        n19002), .Y(n19533) );
  A2O1A1Ixp33_ASAP7_75t_SL U23092 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[50]), 
        .B(n18295), .C(n19002), .Y(n19887) );
  A2O1A1Ixp33_ASAP7_75t_SL U23093 ( .A1(n19886), .A2(n19887), .B(n18295), .C(
        n19002), .Y(n19888) );
  A2O1A1Ixp33_ASAP7_75t_SL U23094 ( .A1(n19730), .A2(n30683), .B(n18295), .C(
        n19002), .Y(n19731) );
  A2O1A1Ixp33_ASAP7_75t_SL U23095 ( .A1(n19002), .A2(n19733), .B(n18295), .C(
        n19002), .Y(n4024) );
  A2O1A1Ixp33_ASAP7_75t_SL U23096 ( .A1(n31444), .A2(n24665), .B(n18295), .C(
        n19002), .Y(n19528) );
  A2O1A1Ixp33_ASAP7_75t_SL U23097 ( .A1(n24901), .A2(n24902), .B(n18295), .C(
        n19002), .Y(n19719) );
  A2O1A1Ixp33_ASAP7_75t_SL U23098 ( .A1(n24675), .A2(n19876), .B(n18295), .C(
        n19002), .Y(n19877) );
  A2O1A1Ixp33_ASAP7_75t_SL U23099 ( .A1(n29695), .A2(n24684), .B(n18295), .C(
        n19002), .Y(n19122) );
  A2O1A1Ixp33_ASAP7_75t_SL U23100 ( .A1(n29694), .A2(n24681), .B(n18295), .C(
        n19122), .Y(n19123) );
  A2O1A1Ixp33_ASAP7_75t_SL U23101 ( .A1(n22378), .A2(n19869), .B(n18295), .C(
        n19002), .Y(n19870) );
  A2O1A1Ixp33_ASAP7_75t_SL U23102 ( .A1(n24676), .A2(n19703), .B(n18295), .C(
        n19002), .Y(n19704) );
  A2O1A1Ixp33_ASAP7_75t_SL U23103 ( .A1(n19002), .A2(n28179), .B(n18295), .C(
        n19002), .Y(n19865) );
  A2O1A1Ixp33_ASAP7_75t_SL U23104 ( .A1(uart1_r_BRATE__5_), .A2(n19865), .B(
        n18295), .C(n19002), .Y(n19866) );
  A2O1A1Ixp33_ASAP7_75t_SL U23105 ( .A1(n19866), .A2(n19867), .B(n18295), .C(
        n19002), .Y(n19868) );
  A2O1A1Ixp33_ASAP7_75t_SL U23106 ( .A1(n30774), .A2(n30068), .B(n18295), .C(
        n19860), .Y(n2862) );
  A2O1A1Ixp33_ASAP7_75t_SL U23107 ( .A1(n29428), .A2(n29383), .B(n18295), .C(
        n19002), .Y(n19693) );
  A2O1A1Ixp33_ASAP7_75t_SL U23108 ( .A1(n31437), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n19859) );
  A2O1A1Ixp33_ASAP7_75t_SL U23109 ( .A1(n27517), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n19855) );
  A2O1A1Ixp33_ASAP7_75t_SL U23110 ( .A1(n19854), .A2(n19855), .B(n18295), .C(
        n19002), .Y(n19856) );
  A2O1A1Ixp33_ASAP7_75t_SL U23111 ( .A1(n29981), .A2(n27509), .B(n18295), .C(
        n19856), .Y(n19857) );
  A2O1A1Ixp33_ASAP7_75t_SL U23112 ( .A1(n19002), .A2(n19857), .B(n18295), .C(
        n19002), .Y(n19858) );
  A2O1A1Ixp33_ASAP7_75t_SL U23113 ( .A1(n30547), .A2(n24633), .B(n18295), .C(
        n19002), .Y(n19688) );
  A2O1A1Ixp33_ASAP7_75t_SL U23114 ( .A1(n18295), .A2(n19002), .B(n19487), .C(
        n19002), .Y(n19488) );
  A2O1A1Ixp33_ASAP7_75t_SL U23115 ( .A1(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_), .A2(n31961), .B(n18295), .C(
        n19840), .Y(n19841) );
  A2O1A1Ixp33_ASAP7_75t_SL U23116 ( .A1(n24681), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_), .B(n18295), .C(n19841), .Y(
        n19842) );
  A2O1A1Ixp33_ASAP7_75t_SL U23117 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__6_), .A2(n32590), .B(n18295), 
        .C(n19002), .Y(n19836) );
  A2O1A1Ixp33_ASAP7_75t_SL U23118 ( .A1(n19835), .A2(n19836), .B(n18295), .C(
        n19002), .Y(n19837) );
  A2O1A1Ixp33_ASAP7_75t_SL U23119 ( .A1(u0_0_leon3x0_p0_ici[64]), .A2(n32594), 
        .B(n18295), .C(n19002), .Y(n19839) );
  A2O1A1Ixp33_ASAP7_75t_SL U23120 ( .A1(n19838), .A2(n19839), .B(n18295), .C(
        n19002), .Y(ic_address[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23121 ( .A1(n32623), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n19826) );
  A2O1A1Ixp33_ASAP7_75t_SL U23122 ( .A1(n32344), .A2(dc_q[13]), .B(n18295), 
        .C(n19002), .Y(n19827) );
  A2O1A1Ixp33_ASAP7_75t_SL U23123 ( .A1(n19826), .A2(n19827), .B(n18295), .C(
        n19002), .Y(n19828) );
  A2O1A1Ixp33_ASAP7_75t_SL U23124 ( .A1(n32413), .A2(n32340), .B(n18295), .C(
        n19002), .Y(n19830) );
  A2O1A1Ixp33_ASAP7_75t_SL U23125 ( .A1(n19829), .A2(n19830), .B(n18295), .C(
        n19002), .Y(dc_data[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23126 ( .A1(n32233), .A2(n32234), .B(n18295), .C(
        n19002), .Y(n19824) );
  A2O1A1Ixp33_ASAP7_75t_SL U23127 ( .A1(n19823), .A2(n19824), .B(n18295), .C(
        n19002), .Y(dt_data[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23128 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__26_), .B(n18295), .C(n19002), .Y(
        n19819) );
  A2O1A1Ixp33_ASAP7_75t_SL U23129 ( .A1(n19242), .A2(DP_OP_1196_128_7433_n8), 
        .B(n18295), .C(n19002), .Y(n19243) );
  A2O1A1Ixp33_ASAP7_75t_SL U23130 ( .A1(n19247), .A2(n19248), .B(n18295), .C(
        n19002), .Y(n19249) );
  A2O1A1Ixp33_ASAP7_75t_SL U23131 ( .A1(n23965), .A2(n29146), .B(n18295), .C(
        n19002), .Y(n19807) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U23132 ( .A1(n24579), .A2(
        u0_0_leon3x0_p0_divi[16]), .B(n18295), .C(n19808), .D(n19812), .Y(
        n30326) );
  A2O1A1Ixp33_ASAP7_75t_SL U23133 ( .A1(uart1_r_RXSTATE__0_), .A2(n2867), .B(
        n18295), .C(n19002), .Y(n19799) );
  A2O1A1Ixp33_ASAP7_75t_SL U23134 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__9_), .B(n18295), .C(n19002), .Y(
        n19798) );
  A2O1A1Ixp33_ASAP7_75t_SL U23135 ( .A1(n22392), .A2(n29837), .B(n18295), .C(
        n19002), .Y(n19792) );
  A2O1A1Ixp33_ASAP7_75t_SL U23136 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__15_), .A2(n24796), .B(n18295), .C(
        n19002), .Y(n19427) );
  A2O1A1Ixp33_ASAP7_75t_SL U23137 ( .A1(DP_OP_1196_128_7433_n235), .A2(
        DP_OP_1196_128_7433_n208), .B(n18295), .C(n19002), .Y(n19789) );
  A2O1A1Ixp33_ASAP7_75t_SL U23138 ( .A1(DP_OP_1196_128_7433_n211), .A2(n19789), 
        .B(n18295), .C(n19002), .Y(n19790) );
  A2O1A1Ixp33_ASAP7_75t_SL U23139 ( .A1(n19002), .A2(n19790), .B(n18295), .C(
        n19002), .Y(DP_OP_1196_128_7433_n207) );
  A2O1A1Ixp33_ASAP7_75t_SL U23140 ( .A1(n32296), .A2(n19788), .B(n18295), .C(
        n19002), .Y(n32389) );
  A2O1A1Ixp33_ASAP7_75t_SL U23141 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[55]), 
        .B(n18295), .C(n19002), .Y(n19624) );
  A2O1A1Ixp33_ASAP7_75t_SL U23142 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__24_), .B(n18295), .C(n19002), .Y(n19625) );
  A2O1A1Ixp33_ASAP7_75t_SL U23143 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[56]), 
        .B(n18295), .C(n19002), .Y(n19628) );
  A2O1A1Ixp33_ASAP7_75t_SL U23144 ( .A1(n19624), .A2(n19627), .B(n18295), .C(
        n19628), .Y(u0_0_leon3x0_p0_div0_vaddin1[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23145 ( .A1(n27534), .A2(n19183), .B(n18295), .C(
        n19002), .Y(n19184) );
  A2O1A1Ixp33_ASAP7_75t_SL U23146 ( .A1(uart1_v_RXDB__1_), .A2(
        uart1_r_RCNT__5_), .B(n18295), .C(n19002), .Y(n19185) );
  A2O1A1Ixp33_ASAP7_75t_SL U23147 ( .A1(n27538), .A2(n27537), .B(n18295), .C(
        n19002), .Y(n19187) );
  A2O1A1Ixp33_ASAP7_75t_SL U23148 ( .A1(n28251), .A2(n28250), .B(n18295), .C(
        n19002), .Y(n19556) );
  A2O1A1Ixp33_ASAP7_75t_SL U23149 ( .A1(n19557), .A2(n19558), .B(n18295), .C(
        n19002), .Y(n19559) );
  A2O1A1Ixp33_ASAP7_75t_SL U23150 ( .A1(uart1_r_RHOLD__21__3_), .A2(n31210), 
        .B(n18295), .C(n19002), .Y(n19562) );
  A2O1A1Ixp33_ASAP7_75t_SL U23151 ( .A1(uart1_r_RHOLD__26__3_), .A2(n31212), 
        .B(n18295), .C(n19002), .Y(n19563) );
  A2O1A1Ixp33_ASAP7_75t_SL U23152 ( .A1(uart1_r_RHOLD__20__3_), .A2(n31211), 
        .B(n18295), .C(n19002), .Y(n19564) );
  A2O1A1Ixp33_ASAP7_75t_SL U23153 ( .A1(n19562), .A2(n19563), .B(n18295), .C(
        n19564), .Y(n19565) );
  A2O1A1Ixp33_ASAP7_75t_SL U23154 ( .A1(uart1_r_RHOLD__7__3_), .A2(n31207), 
        .B(n18295), .C(n19002), .Y(n19567) );
  A2O1A1Ixp33_ASAP7_75t_SL U23155 ( .A1(uart1_r_RHOLD__25__3_), .A2(n31209), 
        .B(n18295), .C(n19002), .Y(n19568) );
  A2O1A1Ixp33_ASAP7_75t_SL U23156 ( .A1(uart1_r_RHOLD__17__3_), .A2(n31206), 
        .B(n18295), .C(n19002), .Y(n19569) );
  A2O1A1Ixp33_ASAP7_75t_SL U23157 ( .A1(n19567), .A2(n19568), .B(n18295), .C(
        n19569), .Y(n19570) );
  A2O1A1Ixp33_ASAP7_75t_SL U23158 ( .A1(n19566), .A2(n19571), .B(n18295), .C(
        n19002), .Y(n19572) );
  A2O1A1Ixp33_ASAP7_75t_SL U23159 ( .A1(uart1_r_RHOLD__4__3_), .A2(n31224), 
        .B(n18295), .C(n19002), .Y(n19573) );
  A2O1A1Ixp33_ASAP7_75t_SL U23160 ( .A1(uart1_r_RHOLD__10__3_), .A2(n31225), 
        .B(n18295), .C(n19002), .Y(n19574) );
  A2O1A1Ixp33_ASAP7_75t_SL U23161 ( .A1(uart1_r_RHOLD__2__3_), .A2(n31223), 
        .B(n18295), .C(n19002), .Y(n19575) );
  A2O1A1Ixp33_ASAP7_75t_SL U23162 ( .A1(n19573), .A2(n19574), .B(n18295), .C(
        n19575), .Y(n19576) );
  A2O1A1Ixp33_ASAP7_75t_SL U23163 ( .A1(uart1_r_RHOLD__14__3_), .A2(n31203), 
        .B(n18295), .C(n19002), .Y(n19578) );
  A2O1A1Ixp33_ASAP7_75t_SL U23164 ( .A1(n19579), .A2(n19580), .B(n18295), .C(
        n19002), .Y(n19581) );
  A2O1A1Ixp33_ASAP7_75t_SL U23165 ( .A1(uart1_r_RHOLD__12__3_), .A2(n31202), 
        .B(n18295), .C(n19002), .Y(n19583) );
  A2O1A1Ixp33_ASAP7_75t_SL U23166 ( .A1(n19578), .A2(n19582), .B(n18295), .C(
        n19583), .Y(n19584) );
  A2O1A1Ixp33_ASAP7_75t_SL U23167 ( .A1(uart1_r_RHOLD__8__3_), .A2(n31227), 
        .B(n18295), .C(n19002), .Y(n19586) );
  A2O1A1Ixp33_ASAP7_75t_SL U23168 ( .A1(uart1_r_RHOLD__22__3_), .A2(n31229), 
        .B(n18295), .C(n19002), .Y(n19587) );
  A2O1A1Ixp33_ASAP7_75t_SL U23169 ( .A1(uart1_r_RHOLD__18__3_), .A2(n31228), 
        .B(n18295), .C(n19002), .Y(n19588) );
  A2O1A1Ixp33_ASAP7_75t_SL U23170 ( .A1(n19586), .A2(n19587), .B(n18295), .C(
        n19588), .Y(n19589) );
  A2O1A1Ixp33_ASAP7_75t_SL U23171 ( .A1(n19577), .A2(n19585), .B(n18295), .C(
        n19590), .Y(n19591) );
  A2O1A1Ixp33_ASAP7_75t_SL U23172 ( .A1(n19595), .A2(n19596), .B(n18295), .C(
        n19002), .Y(n19597) );
  A2O1A1Ixp33_ASAP7_75t_SL U23173 ( .A1(n19598), .A2(n19599), .B(n18295), .C(
        n19002), .Y(n19600) );
  A2O1A1Ixp33_ASAP7_75t_SL U23174 ( .A1(n31951), .A2(uart1_r_BREAK_), .B(
        n18295), .C(n19002), .Y(n19602) );
  A2O1A1Ixp33_ASAP7_75t_SL U23175 ( .A1(uart1_r_BRATE__3_), .A2(n31246), .B(
        n18295), .C(n19002), .Y(n19603) );
  A2O1A1Ixp33_ASAP7_75t_SL U23176 ( .A1(n19601), .A2(n19602), .B(n18295), .C(
        n19603), .Y(n19604) );
  A2O1A1Ixp33_ASAP7_75t_SL U23177 ( .A1(timer0_r_SCALER__3_), .A2(n31245), .B(
        n18295), .C(n19002), .Y(n19609) );
  A2O1A1Ixp33_ASAP7_75t_SL U23178 ( .A1(irqctrl0_r_IPEND__3_), .A2(n31247), 
        .B(n18295), .C(n19002), .Y(n19610) );
  A2O1A1Ixp33_ASAP7_75t_SL U23179 ( .A1(timer0_vtimers_1__IRQEN_), .A2(n30790), 
        .B(n18295), .C(n19002), .Y(n19611) );
  A2O1A1Ixp33_ASAP7_75t_SL U23180 ( .A1(n19609), .A2(n19610), .B(n18295), .C(
        n19611), .Y(n19612) );
  A2O1A1Ixp33_ASAP7_75t_SL U23181 ( .A1(n19613), .A2(n19614), .B(n18295), .C(
        n19002), .Y(n19615) );
  A2O1A1Ixp33_ASAP7_75t_SL U23182 ( .A1(n19002), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__24_), .B(n18295), .C(n19002), .Y(n19552)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U23183 ( .A1(n19551), .A2(n19553), .B(n18295), .C(
        n19002), .Y(n4509) );
  A2O1A1Ixp33_ASAP7_75t_SL U23184 ( .A1(n19759), .A2(n19778), .B(n18295), .C(
        n19002), .Y(n4508) );
  A2O1A1Ixp33_ASAP7_75t_SL U23185 ( .A1(n19002), .A2(n30389), .B(n18295), .C(
        n19002), .Y(n19747) );
  A2O1A1Ixp33_ASAP7_75t_SL U23186 ( .A1(n31415), .A2(n19747), .B(n18295), .C(
        n19002), .Y(n19748) );
  A2O1A1Ixp33_ASAP7_75t_SL U23187 ( .A1(n19002), .A2(n24638), .B(n18295), .C(
        n19002), .Y(n19752) );
  A2O1A1Ixp33_ASAP7_75t_SL U23188 ( .A1(n19748), .A2(n19755), .B(n18295), .C(
        n19002), .Y(n19756) );
  A2O1A1Ixp33_ASAP7_75t_SL U23189 ( .A1(n24681), .A2(n19734), .B(n18295), .C(
        n19735), .Y(n19736) );
  A2O1A1Ixp33_ASAP7_75t_SL U23190 ( .A1(n31958), .A2(n24659), .B(n18295), .C(
        n19002), .Y(n19327) );
  A2O1A1Ixp33_ASAP7_75t_SL U23191 ( .A1(n19731), .A2(n19732), .B(n18295), .C(
        n19002), .Y(n19733) );
  A2O1A1Ixp33_ASAP7_75t_SL U23192 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[47]), 
        .B(n18295), .C(n19002), .Y(n19728) );
  A2O1A1Ixp33_ASAP7_75t_SL U23193 ( .A1(n19727), .A2(n19728), .B(n18295), .C(
        n19002), .Y(n19729) );
  A2O1A1Ixp33_ASAP7_75t_SL U23194 ( .A1(n31968), .A2(n19720), .B(n18295), .C(
        n19002), .Y(n19721) );
  A2O1A1Ixp33_ASAP7_75t_SL U23195 ( .A1(n28562), .A2(n19718), .B(n18295), .C(
        n19002), .Y(n3640) );
  A2O1A1Ixp33_ASAP7_75t_SL U23196 ( .A1(n22421), .A2(DP_OP_1196_128_7433_n452), 
        .B(n18295), .C(n19002), .Y(n19710) );
  A2O1A1Ixp33_ASAP7_75t_SL U23197 ( .A1(n19709), .A2(n19710), .B(n18295), .C(
        n19002), .Y(n19711) );
  A2O1A1Ixp33_ASAP7_75t_SL U23198 ( .A1(n19002), .A2(n19711), .B(n18295), .C(
        n19002), .Y(n3474) );
  A2O1A1Ixp33_ASAP7_75t_SL U23199 ( .A1(u0_0_leon3x0_p0_dci[2]), .A2(n30199), 
        .B(n18295), .C(n19002), .Y(n19696) );
  A2O1A1Ixp33_ASAP7_75t_SL U23200 ( .A1(n19697), .A2(n19698), .B(n18295), .C(
        n19002), .Y(n19699) );
  A2O1A1Ixp33_ASAP7_75t_SL U23201 ( .A1(n19700), .A2(n31600), .B(n18295), .C(
        n19002), .Y(n19701) );
  A2O1A1Ixp33_ASAP7_75t_SL U23202 ( .A1(n29383), .A2(n19694), .B(n18295), .C(
        n19002), .Y(n19695) );
  A2O1A1Ixp33_ASAP7_75t_SL U23203 ( .A1(n24664), .A2(n19302), .B(n18295), .C(
        n19002), .Y(n19303) );
  A2O1A1Ixp33_ASAP7_75t_SL U23204 ( .A1(n31730), .A2(n19689), .B(n18295), .C(
        n19002), .Y(n19690) );
  A2O1A1Ixp33_ASAP7_75t_SL U23205 ( .A1(n28108), .A2(n27968), .B(n18295), .C(
        n19002), .Y(n19490) );
  A2O1A1Ixp33_ASAP7_75t_SL U23206 ( .A1(n28108), .A2(n27929), .B(n18295), .C(
        n19002), .Y(n19489) );
  A2O1A1Ixp33_ASAP7_75t_SL U23207 ( .A1(n32566), .A2(n19679), .B(n18295), .C(
        n19002), .Y(n19680) );
  A2O1A1Ixp33_ASAP7_75t_SL U23208 ( .A1(n32385), .A2(dc_q[23]), .B(n18295), 
        .C(n19002), .Y(n19668) );
  A2O1A1Ixp33_ASAP7_75t_SL U23209 ( .A1(n19667), .A2(n19668), .B(n18295), .C(
        n19002), .Y(n19669) );
  A2O1A1Ixp33_ASAP7_75t_SL U23210 ( .A1(n32386), .A2(n32433), .B(n18295), .C(
        n19002), .Y(n19671) );
  A2O1A1Ixp33_ASAP7_75t_SL U23211 ( .A1(n19670), .A2(n19671), .B(n18295), .C(
        n19002), .Y(dc_data[23]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23212 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__18_), 
        .A2(n32214), .B(n18295), .C(n19002), .Y(n19661) );
  A2O1A1Ixp33_ASAP7_75t_SL U23213 ( .A1(n19660), .A2(n19661), .B(n18295), .C(
        n19002), .Y(n19662) );
  A2O1A1Ixp33_ASAP7_75t_SL U23214 ( .A1(n19002), .A2(n19662), .B(n18295), .C(
        n19002), .Y(n19663) );
  A2O1A1Ixp33_ASAP7_75t_SL U23215 ( .A1(n29723), .A2(n19659), .B(n18295), .C(
        n19002), .Y(n29639) );
  A2O1A1Ixp33_ASAP7_75t_SL U23216 ( .A1(n24574), .A2(ahb0_r_HRDATAS__13_), .B(
        n18295), .C(n19002), .Y(n19655) );
  A2O1A1Ixp33_ASAP7_75t_SL U23217 ( .A1(n30001), .A2(ahb0_r_HRDATAM__13_), .B(
        n18295), .C(n19002), .Y(n19656) );
  A2O1A1Ixp33_ASAP7_75t_SL U23218 ( .A1(n30002), .A2(ahbso_1__HRDATA__13_), 
        .B(n18295), .C(n19002), .Y(n19657) );
  A2O1A1Ixp33_ASAP7_75t_SL U23219 ( .A1(n19655), .A2(n19656), .B(n18295), .C(
        n19657), .Y(n19658) );
  A2O1A1Ixp33_ASAP7_75t_SL U23220 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__10_), .B(n18295), .C(n19002), .Y(
        n19654) );
  A2O1A1Ixp33_ASAP7_75t_SL U23221 ( .A1(n19650), .A2(n19651), .B(n18295), .C(
        n19002), .Y(n19652) );
  A2O1A1Ixp33_ASAP7_75t_SL U23222 ( .A1(DP_OP_1196_128_7433_n8), .A2(n19446), 
        .B(n18295), .C(n19002), .Y(n19447) );
  A2O1A1Ixp33_ASAP7_75t_SL U23223 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__3_), .A2(
        n30641), .B(n18295), .C(n19002), .Y(n19642) );
  A2O1A1Ixp33_ASAP7_75t_SL U23224 ( .A1(rf_do_b[3]), .A2(n30640), .B(n18295), 
        .C(n19002), .Y(n19643) );
  A2O1A1Ixp33_ASAP7_75t_SL U23225 ( .A1(u0_0_leon3x0_p0_iu_r_W__RESULT__3_), 
        .A2(n29863), .B(n18295), .C(n19002), .Y(n19646) );
  A2O1A1Ixp33_ASAP7_75t_SL U23226 ( .A1(n29731), .A2(
        u0_0_leon3x0_p0_iu_r_X__RESULT__5_), .B(n18295), .C(n19002), .Y(n19640) );
  A2O1A1Ixp33_ASAP7_75t_SL U23227 ( .A1(u0_0_leon3x0_p0_ici[52]), .A2(n29059), 
        .B(n18295), .C(n19002), .Y(n19438) );
  A2O1A1Ixp33_ASAP7_75t_SL U23228 ( .A1(n19002), .A2(n19440), .B(n18295), .C(
        n19002), .Y(n19441) );
  A2O1A1Ixp33_ASAP7_75t_SL U23229 ( .A1(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__1_), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_HIT_), .B(n18295), .C(n19002), .Y(
        n19632) );
  A2O1A1Ixp33_ASAP7_75t_SL U23230 ( .A1(n31352), .A2(n19629), .B(n18295), .C(
        n19002), .Y(n29328) );
  A2O1A1Ixp33_ASAP7_75t_SL U23231 ( .A1(n19002), .A2(n19182), .B(n18295), .C(
        n19002), .Y(n19183) );
  A2O1A1Ixp33_ASAP7_75t_SL U23232 ( .A1(n29336), .A2(n19188), .B(n18295), .C(
        n19002), .Y(n19189) );
  A2O1A1Ixp33_ASAP7_75t_SL U23233 ( .A1(n29973), .A2(n19189), .B(n18295), .C(
        n19002), .Y(n19190) );
  A2O1A1Ixp33_ASAP7_75t_SL U23234 ( .A1(uart1_r_RHOLD__13__3_), .A2(n31220), 
        .B(n18295), .C(n19002), .Y(n19557) );
  A2O1A1Ixp33_ASAP7_75t_SL U23235 ( .A1(uart1_r_RHOLD__31__3_), .A2(n31221), 
        .B(n18295), .C(n19002), .Y(n19558) );
  A2O1A1Ixp33_ASAP7_75t_SL U23236 ( .A1(n28252), .A2(n19560), .B(n18295), .C(
        n19002), .Y(n19561) );
  A2O1A1Ixp33_ASAP7_75t_SL U23237 ( .A1(uart1_r_RHOLD__30__3_), .A2(n31201), 
        .B(n18295), .C(n19002), .Y(n19579) );
  A2O1A1Ixp33_ASAP7_75t_SL U23238 ( .A1(n31200), .A2(uart1_r_RHOLD__5__3_), 
        .B(n18295), .C(n19002), .Y(n19580) );
  A2O1A1Ixp33_ASAP7_75t_SL U23239 ( .A1(timer0_r_RELOAD__3_), .A2(n31237), .B(
        n18295), .C(n19002), .Y(n19593) );
  A2O1A1Ixp33_ASAP7_75t_SL U23240 ( .A1(irqctrl0_r_IMASK__0__3_), .A2(n31249), 
        .B(n18295), .C(n19002), .Y(n19595) );
  A2O1A1Ixp33_ASAP7_75t_SL U23241 ( .A1(irqctrl0_r_IFORCE__0__3_), .A2(n31251), 
        .B(n18295), .C(n19002), .Y(n19596) );
  A2O1A1Ixp33_ASAP7_75t_SL U23242 ( .A1(n31235), .A2(sr1_r_MCFG1__ROMRWS__3_), 
        .B(n18295), .C(n19002), .Y(n19599) );
  A2O1A1Ixp33_ASAP7_75t_SL U23243 ( .A1(n19002), .A2(n30783), .B(n18295), .C(
        n19002), .Y(n19607) );
  A2O1A1Ixp33_ASAP7_75t_SL U23244 ( .A1(uart1_r_RHOLD__24__3_), .A2(n19607), 
        .B(n18295), .C(n19002), .Y(n19608) );
  A2O1A1Ixp33_ASAP7_75t_SL U23245 ( .A1(uart1_r_TIRQEN_), .A2(n31950), .B(
        n18295), .C(n19002), .Y(n19614) );
  A2O1A1Ixp33_ASAP7_75t_SL U23246 ( .A1(n19606), .A2(n19608), .B(n18295), .C(
        n19616), .Y(n19617) );
  A2O1A1Ixp33_ASAP7_75t_SL U23247 ( .A1(n24667), .A2(n19552), .B(n18295), .C(
        n19002), .Y(n19553) );
  A2O1A1Ixp33_ASAP7_75t_SL U23248 ( .A1(n19002), .A2(n31757), .B(n18295), .C(
        n19002), .Y(n19547) );
  A2O1A1Ixp33_ASAP7_75t_SL U23249 ( .A1(n31758), .A2(n19547), .B(n18295), .C(
        n19002), .Y(n19548) );
  A2O1A1Ixp33_ASAP7_75t_SL U23250 ( .A1(n31756), .A2(n19548), .B(n18295), .C(
        n19002), .Y(n4483) );
  A2O1A1Ixp33_ASAP7_75t_SL U23251 ( .A1(n31043), .A2(n31044), .B(n18295), .C(
        n19002), .Y(n19544) );
  A2O1A1Ixp33_ASAP7_75t_SL U23252 ( .A1(n31364), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__10_), .B(n18295), .C(n19002), .Y(
        n19545) );
  A2O1A1Ixp33_ASAP7_75t_SL U23253 ( .A1(n19544), .A2(n19545), .B(n18295), .C(
        n19002), .Y(n19546) );
  A2O1A1Ixp33_ASAP7_75t_SL U23254 ( .A1(n30264), .A2(n30453), .B(n18295), .C(
        n19002), .Y(n19157) );
  A2O1A1Ixp33_ASAP7_75t_SL U23255 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__23_), 
        .A2(n19159), .B(n18295), .C(n19002), .Y(n19160) );
  A2O1A1Ixp33_ASAP7_75t_SL U23256 ( .A1(n19158), .A2(n19160), .B(n18295), .C(
        n19002), .Y(n19161) );
  A2O1A1Ixp33_ASAP7_75t_SL U23257 ( .A1(n30640), .A2(rf_do_b[27]), .B(n18295), 
        .C(n19002), .Y(n19535) );
  A2O1A1Ixp33_ASAP7_75t_SL U23258 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__27_), .B(n18295), .C(n19002), .Y(n19536)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U23259 ( .A1(n19535), .A2(n19536), .B(n18295), .C(
        n19002), .Y(n19537) );
  A2O1A1Ixp33_ASAP7_75t_SL U23260 ( .A1(n23843), .A2(n24667), .B(n18295), .C(
        n19002), .Y(n19542) );
  A2O1A1Ixp33_ASAP7_75t_SL U23261 ( .A1(n19329), .A2(n19334), .B(n18295), .C(
        n19002), .Y(n4295) );
  A2O1A1Ixp33_ASAP7_75t_SL U23262 ( .A1(n32042), .A2(n19529), .B(n18295), .C(
        n19002), .Y(n19530) );
  A2O1A1Ixp33_ASAP7_75t_SL U23263 ( .A1(n24666), .A2(n19526), .B(n18295), .C(
        n19002), .Y(n19527) );
  A2O1A1Ixp33_ASAP7_75t_SL U23264 ( .A1(n24678), .A2(n19524), .B(n18295), .C(
        n19002), .Y(n19525) );
  A2O1A1Ixp33_ASAP7_75t_SL U23265 ( .A1(n24670), .A2(n25881), .B(n18295), .C(
        n19002), .Y(n19523) );
  A2O1A1Ixp33_ASAP7_75t_SL U23266 ( .A1(n32163), .A2(n19519), .B(n18295), .C(
        n19002), .Y(n19520) );
  A2O1A1Ixp33_ASAP7_75t_SL U23267 ( .A1(n24676), .A2(n19312), .B(n18295), .C(
        n19002), .Y(n19313) );
  A2O1A1Ixp33_ASAP7_75t_SL U23268 ( .A1(n31438), .A2(n22379), .B(n18295), .C(
        n19002), .Y(n19516) );
  A2O1A1Ixp33_ASAP7_75t_SL U23269 ( .A1(n30701), .A2(n30700), .B(n18295), .C(
        n19002), .Y(n19515) );
  A2O1A1Ixp33_ASAP7_75t_SL U23270 ( .A1(n24662), .A2(n19513), .B(n18295), .C(
        n19002), .Y(n19514) );
  A2O1A1Ixp33_ASAP7_75t_SL U23271 ( .A1(n22427), .A2(n19511), .B(n18295), .C(
        n19002), .Y(n19512) );
  A2O1A1Ixp33_ASAP7_75t_SL U23272 ( .A1(n24676), .A2(n19509), .B(n18295), .C(
        n19002), .Y(n19510) );
  A2O1A1Ixp33_ASAP7_75t_SL U23273 ( .A1(n29383), .A2(n19505), .B(n18295), .C(
        n19002), .Y(n19506) );
  A2O1A1Ixp33_ASAP7_75t_SL U23274 ( .A1(n26619), .A2(n31840), .B(n18295), .C(
        n19002), .Y(n19307) );
  A2O1A1Ixp33_ASAP7_75t_SL U23275 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[48]), 
        .B(n18295), .C(n19002), .Y(n19499) );
  A2O1A1Ixp33_ASAP7_75t_SL U23276 ( .A1(n19498), .A2(n19499), .B(n18295), .C(
        n19002), .Y(n19500) );
  A2O1A1Ixp33_ASAP7_75t_SL U23277 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[40]), 
        .B(n18295), .C(n19002), .Y(n19493) );
  A2O1A1Ixp33_ASAP7_75t_SL U23278 ( .A1(n19492), .A2(n19493), .B(n18295), .C(
        n19002), .Y(n19494) );
  A2O1A1Ixp33_ASAP7_75t_SL U23279 ( .A1(n30139), .A2(n24633), .B(n18295), .C(
        n19002), .Y(n19292) );
  A2O1A1Ixp33_ASAP7_75t_SL U23280 ( .A1(n18295), .A2(n19002), .B(n19288), .C(
        n19002), .Y(n19289) );
  A2O1A1Ixp33_ASAP7_75t_SL U23281 ( .A1(n22386), .A2(n19484), .B(n18295), .C(
        n19002), .Y(n19485) );
  A2O1A1Ixp33_ASAP7_75t_SL U23282 ( .A1(ahb0_r_HADDR__2_), .A2(n19483), .B(
        n18295), .C(n19002), .Y(n17288) );
  A2O1A1Ixp33_ASAP7_75t_SL U23283 ( .A1(n22379), .A2(n32119), .B(n18295), .C(
        n19002), .Y(n19286) );
  A2O1A1Ixp33_ASAP7_75t_SL U23284 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__16_), .A2(n19481), .B(n18295), .C(n19002), .Y(n19482) );
  A2O1A1Ixp33_ASAP7_75t_SL U23285 ( .A1(n29405), .A2(n19469), .B(n18295), .C(
        n19002), .Y(n29658) );
  A2O1A1Ixp33_ASAP7_75t_SL U23286 ( .A1(n30640), .A2(rf_do_b[1]), .B(n18295), 
        .C(n19002), .Y(n19463) );
  A2O1A1Ixp33_ASAP7_75t_SL U23287 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__1_), .B(n18295), .C(n19002), .Y(n19464)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U23288 ( .A1(n19463), .A2(n19464), .B(n18295), .C(
        n19002), .Y(n19465) );
  A2O1A1Ixp33_ASAP7_75t_SL U23289 ( .A1(DP_OP_1196_128_7433_n7), .A2(n19446), 
        .B(n18295), .C(n19002), .Y(n19448) );
  A2O1A1Ixp33_ASAP7_75t_SL U23290 ( .A1(n19451), .A2(DP_OP_1196_128_7433_n51), 
        .B(n18295), .C(n19002), .Y(n19452) );
  A2O1A1Ixp33_ASAP7_75t_SL U23291 ( .A1(DP_OP_1196_128_7433_n51), .A2(n19453), 
        .B(n18295), .C(n19002), .Y(n19454) );
  A2O1A1Ixp33_ASAP7_75t_SL U23292 ( .A1(DP_OP_5187J1_124_3275_n297), .A2(
        DP_OP_5187J1_124_3275_n298), .B(n18295), .C(n19444), .Y(n19445) );
  A2O1A1Ixp33_ASAP7_75t_SL U23293 ( .A1(n29731), .A2(
        u0_0_leon3x0_p0_iu_r_X__RESULT__2_), .B(n18295), .C(n19002), .Y(n19443) );
  A2O1A1Ixp33_ASAP7_75t_SL U23294 ( .A1(n19237), .A2(n19239), .B(n18295), .C(
        n19002), .Y(n19240) );
  A2O1A1Ixp33_ASAP7_75t_SL U23295 ( .A1(n19236), .A2(n19240), .B(n18295), .C(
        n19002), .Y(uart1_scaler_11_) );
  A2O1A1Ixp33_ASAP7_75t_SL U23296 ( .A1(n19438), .A2(n19439), .B(n18295), .C(
        n19002), .Y(n19440) );
  A2O1A1Ixp33_ASAP7_75t_SL U23297 ( .A1(n31833), .A2(n19437), .B(n18295), .C(
        n19002), .Y(n32665) );
  A2O1A1Ixp33_ASAP7_75t_SL U23298 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__5_), .B(n18295), .C(n19002), .Y(n19432) );
  A2O1A1Ixp33_ASAP7_75t_SL U23299 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[37]), 
        .B(n18295), .C(n19002), .Y(n19435) );
  A2O1A1Ixp33_ASAP7_75t_SL U23300 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[36]), 
        .B(n18295), .C(n19002), .Y(n19436) );
  A2O1A1Ixp33_ASAP7_75t_SL U23301 ( .A1(n19434), .A2(n19435), .B(n18295), .C(
        n19436), .Y(u0_0_leon3x0_p0_div0_vaddin1[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23302 ( .A1(n32202), .A2(n19429), .B(n18295), .C(
        n19002), .Y(n32203) );
  A2O1A1Ixp33_ASAP7_75t_SL U23303 ( .A1(n28602), .A2(n22392), .B(n18295), .C(
        n19002), .Y(n19011) );
  A2O1A1Ixp33_ASAP7_75t_SL U23304 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[43]), 
        .B(n18295), .C(n19002), .Y(n19212) );
  A2O1A1Ixp33_ASAP7_75t_SL U23305 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__12_), .B(n18295), .C(n19002), .Y(n19213) );
  A2O1A1Ixp33_ASAP7_75t_SL U23306 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[44]), 
        .B(n18295), .C(n19002), .Y(n19216) );
  A2O1A1Ixp33_ASAP7_75t_SL U23307 ( .A1(n19212), .A2(n19215), .B(n18295), .C(
        n19216), .Y(u0_0_leon3x0_p0_div0_vaddin1[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23308 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__27_), .B(n18295), .C(n19002), .Y(n19422) );
  A2O1A1Ixp33_ASAP7_75t_SL U23309 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[59]), 
        .B(n18295), .C(n19002), .Y(n19425) );
  A2O1A1Ixp33_ASAP7_75t_SL U23310 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[58]), 
        .B(n18295), .C(n19002), .Y(n19426) );
  A2O1A1Ixp33_ASAP7_75t_SL U23311 ( .A1(n19424), .A2(n19425), .B(n18295), .C(
        n19426), .Y(u0_0_leon3x0_p0_div0_vaddin1[28]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23312 ( .A1(n29336), .A2(n19180), .B(n18295), .C(
        n19002), .Y(n19181) );
  A2O1A1Ixp33_ASAP7_75t_SL U23313 ( .A1(n29973), .A2(n19181), .B(n18295), .C(
        n19002), .Y(n19182) );
  A2O1A1Ixp33_ASAP7_75t_SL U23314 ( .A1(n19002), .A2(n27536), .B(n18295), .C(
        n19002), .Y(n19188) );
  A2O1A1Ixp33_ASAP7_75t_SL U23315 ( .A1(n31249), .A2(irqctrl0_r_IMASK__0__2_), 
        .B(n18295), .C(n19002), .Y(n19359) );
  A2O1A1Ixp33_ASAP7_75t_SL U23316 ( .A1(irqctrl0_r_IFORCE__0__2_), .A2(n31251), 
        .B(n18295), .C(n19002), .Y(n19360) );
  A2O1A1Ixp33_ASAP7_75t_SL U23317 ( .A1(n31235), .A2(sr1_r_MCFG1__ROMRWS__2_), 
        .B(n18295), .C(n19002), .Y(n19361) );
  A2O1A1Ixp33_ASAP7_75t_SL U23318 ( .A1(n19359), .A2(n19360), .B(n18295), .C(
        n19361), .Y(n19362) );
  A2O1A1Ixp33_ASAP7_75t_SL U23319 ( .A1(timer0_r_SCALER__2_), .A2(n31245), .B(
        n18295), .C(n19002), .Y(n19364) );
  A2O1A1Ixp33_ASAP7_75t_SL U23320 ( .A1(n19363), .A2(n19364), .B(n18295), .C(
        n19002), .Y(n19365) );
  A2O1A1Ixp33_ASAP7_75t_SL U23321 ( .A1(n31226), .A2(uart1_r_RHOLD__6__2_), 
        .B(n18295), .C(n19002), .Y(n19368) );
  A2O1A1Ixp33_ASAP7_75t_SL U23322 ( .A1(uart1_r_RHOLD__2__2_), .A2(n31223), 
        .B(n18295), .C(n19002), .Y(n19369) );
  A2O1A1Ixp33_ASAP7_75t_SL U23323 ( .A1(n31224), .A2(uart1_r_RHOLD__4__2_), 
        .B(n18295), .C(n19002), .Y(n19370) );
  A2O1A1Ixp33_ASAP7_75t_SL U23324 ( .A1(n19368), .A2(n19369), .B(n18295), .C(
        n19370), .Y(n19371) );
  A2O1A1Ixp33_ASAP7_75t_SL U23325 ( .A1(n31230), .A2(uart1_r_RHOLD__27__2_), 
        .B(n18295), .C(n19002), .Y(n19373) );
  A2O1A1Ixp33_ASAP7_75t_SL U23326 ( .A1(n31227), .A2(uart1_r_RHOLD__8__2_), 
        .B(n18295), .C(n19002), .Y(n19374) );
  A2O1A1Ixp33_ASAP7_75t_SL U23327 ( .A1(n31228), .A2(uart1_r_RHOLD__18__2_), 
        .B(n18295), .C(n19002), .Y(n19375) );
  A2O1A1Ixp33_ASAP7_75t_SL U23328 ( .A1(n19373), .A2(n19374), .B(n18295), .C(
        n19375), .Y(n19376) );
  A2O1A1Ixp33_ASAP7_75t_SL U23329 ( .A1(n31213), .A2(uart1_r_RHOLD__15__2_), 
        .B(n18295), .C(n19002), .Y(n19378) );
  A2O1A1Ixp33_ASAP7_75t_SL U23330 ( .A1(n31210), .A2(uart1_r_RHOLD__21__2_), 
        .B(n18295), .C(n19002), .Y(n19379) );
  A2O1A1Ixp33_ASAP7_75t_SL U23331 ( .A1(n31211), .A2(uart1_r_RHOLD__20__2_), 
        .B(n18295), .C(n19002), .Y(n19380) );
  A2O1A1Ixp33_ASAP7_75t_SL U23332 ( .A1(n19378), .A2(n19379), .B(n18295), .C(
        n19380), .Y(n19381) );
  A2O1A1Ixp33_ASAP7_75t_SL U23333 ( .A1(n31209), .A2(uart1_r_RHOLD__25__2_), 
        .B(n18295), .C(n19002), .Y(n19383) );
  A2O1A1Ixp33_ASAP7_75t_SL U23334 ( .A1(n31206), .A2(uart1_r_RHOLD__17__2_), 
        .B(n18295), .C(n19002), .Y(n19384) );
  A2O1A1Ixp33_ASAP7_75t_SL U23335 ( .A1(n31207), .A2(uart1_r_RHOLD__7__2_), 
        .B(n18295), .C(n19002), .Y(n19385) );
  A2O1A1Ixp33_ASAP7_75t_SL U23336 ( .A1(n19383), .A2(n19384), .B(n18295), .C(
        n19385), .Y(n19386) );
  A2O1A1Ixp33_ASAP7_75t_SL U23337 ( .A1(n31203), .A2(uart1_r_RHOLD__14__2_), 
        .B(n18295), .C(n19002), .Y(n19388) );
  A2O1A1Ixp33_ASAP7_75t_SL U23338 ( .A1(n19382), .A2(n19387), .B(n18295), .C(
        n19388), .Y(n19389) );
  A2O1A1Ixp33_ASAP7_75t_SL U23339 ( .A1(n31201), .A2(uart1_r_RHOLD__30__2_), 
        .B(n18295), .C(n19002), .Y(n19390) );
  A2O1A1Ixp33_ASAP7_75t_SL U23340 ( .A1(n31204), .A2(uart1_r_RHOLD__9__2_), 
        .B(n18295), .C(n19002), .Y(n19391) );
  A2O1A1Ixp33_ASAP7_75t_SL U23341 ( .A1(n31205), .A2(uart1_r_RHOLD__16__2_), 
        .B(n18295), .C(n19002), .Y(n19392) );
  A2O1A1Ixp33_ASAP7_75t_SL U23342 ( .A1(n19390), .A2(n19391), .B(n18295), .C(
        n19392), .Y(n19393) );
  A2O1A1Ixp33_ASAP7_75t_SL U23343 ( .A1(n31217), .A2(uart1_r_RHOLD__29__2_), 
        .B(n18295), .C(n19002), .Y(n19395) );
  A2O1A1Ixp33_ASAP7_75t_SL U23344 ( .A1(n31214), .A2(uart1_r_RHOLD__1__2_), 
        .B(n18295), .C(n19002), .Y(n19396) );
  A2O1A1Ixp33_ASAP7_75t_SL U23345 ( .A1(uart1_r_RHOLD__28__2_), .A2(n31215), 
        .B(n18295), .C(n19002), .Y(n19397) );
  A2O1A1Ixp33_ASAP7_75t_SL U23346 ( .A1(n19395), .A2(n19396), .B(n18295), .C(
        n19397), .Y(n19398) );
  A2O1A1Ixp33_ASAP7_75t_SL U23347 ( .A1(n31221), .A2(uart1_r_RHOLD__31__2_), 
        .B(n18295), .C(n19002), .Y(n19400) );
  A2O1A1Ixp33_ASAP7_75t_SL U23348 ( .A1(n31218), .A2(uart1_r_RHOLD__23__2_), 
        .B(n18295), .C(n19002), .Y(n19401) );
  A2O1A1Ixp33_ASAP7_75t_SL U23349 ( .A1(uart1_r_RHOLD__11__2_), .A2(n31219), 
        .B(n18295), .C(n19002), .Y(n19402) );
  A2O1A1Ixp33_ASAP7_75t_SL U23350 ( .A1(n19400), .A2(n19401), .B(n18295), .C(
        n19402), .Y(n19403) );
  A2O1A1Ixp33_ASAP7_75t_SL U23351 ( .A1(n19394), .A2(n19399), .B(n18295), .C(
        n19404), .Y(n19405) );
  A2O1A1Ixp33_ASAP7_75t_SL U23352 ( .A1(n19372), .A2(n19377), .B(n18295), .C(
        n19406), .Y(n19407) );
  A2O1A1Ixp33_ASAP7_75t_SL U23353 ( .A1(n31237), .A2(timer0_r_RELOAD__2_), .B(
        n18295), .C(n19002), .Y(n19408) );
  A2O1A1Ixp33_ASAP7_75t_SL U23354 ( .A1(n31246), .A2(uart1_r_BRATE__2_), .B(
        n18295), .C(n19002), .Y(n19409) );
  A2O1A1Ixp33_ASAP7_75t_SL U23355 ( .A1(n19408), .A2(n19409), .B(n18295), .C(
        n19002), .Y(n19410) );
  A2O1A1Ixp33_ASAP7_75t_SL U23356 ( .A1(n31247), .A2(irqctrl0_r_IPEND__2_), 
        .B(n18295), .C(n19002), .Y(n19411) );
  A2O1A1Ixp33_ASAP7_75t_SL U23357 ( .A1(n31248), .A2(irqctrl0_r_ILEVEL__2_), 
        .B(n18295), .C(n19002), .Y(n19412) );
  A2O1A1Ixp33_ASAP7_75t_SL U23358 ( .A1(n19411), .A2(n19412), .B(n18295), .C(
        n19002), .Y(n19413) );
  A2O1A1Ixp33_ASAP7_75t_SL U23359 ( .A1(n31950), .A2(uart1_r_RIRQEN_), .B(
        n18295), .C(n19002), .Y(n19415) );
  A2O1A1Ixp33_ASAP7_75t_SL U23360 ( .A1(n29558), .A2(n31951), .B(n18295), .C(
        n19002), .Y(n19416) );
  A2O1A1Ixp33_ASAP7_75t_SL U23361 ( .A1(n19414), .A2(n19415), .B(n18295), .C(
        n19416), .Y(n19417) );
  A2O1A1Ixp33_ASAP7_75t_SL U23362 ( .A1(n31956), .A2(
        timer0_vtimers_1__RELOAD__2_), .B(n18295), .C(n19002), .Y(n19419) );
  A2O1A1Ixp33_ASAP7_75t_SL U23363 ( .A1(n30790), .A2(timer0_vtimers_1__LOAD_), 
        .B(n18295), .C(n19002), .Y(n19420) );
  A2O1A1Ixp33_ASAP7_75t_SL U23364 ( .A1(n19418), .A2(n19419), .B(n18295), .C(
        n19420), .Y(n19421) );
  A2O1A1Ixp33_ASAP7_75t_SL U23365 ( .A1(n31542), .A2(n27087), .B(n18295), .C(
        n19002), .Y(n19165) );
  A2O1A1Ixp33_ASAP7_75t_SL U23366 ( .A1(n18295), .A2(n19002), .B(n19166), .C(
        n19002), .Y(n19167) );
  A2O1A1Ixp33_ASAP7_75t_SL U23367 ( .A1(n24647), .A2(n27088), .B(n18295), .C(
        n19002), .Y(n19168) );
  A2O1A1Ixp33_ASAP7_75t_SL U23368 ( .A1(n19165), .A2(n19167), .B(n18295), .C(
        n19168), .Y(n4501) );
  A2O1A1Ixp33_ASAP7_75t_SL U23369 ( .A1(n24638), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n19350) );
  A2O1A1Ixp33_ASAP7_75t_SL U23370 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__Y__10_), 
        .A2(n19350), .B(n18295), .C(n19002), .Y(n19351) );
  A2O1A1Ixp33_ASAP7_75t_SL U23371 ( .A1(n19351), .A2(n19353), .B(n18295), .C(
        n19002), .Y(n19354) );
  A2O1A1Ixp33_ASAP7_75t_SL U23372 ( .A1(n31043), .A2(n30573), .B(n18295), .C(
        n19002), .Y(n19346) );
  A2O1A1Ixp33_ASAP7_75t_SL U23373 ( .A1(n31364), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__14_), .B(n18295), .C(n19002), .Y(
        n19347) );
  A2O1A1Ixp33_ASAP7_75t_SL U23374 ( .A1(n19346), .A2(n19347), .B(n18295), .C(
        n19002), .Y(n19348) );
  A2O1A1Ixp33_ASAP7_75t_SL U23375 ( .A1(n30640), .A2(rf_do_b[6]), .B(n18295), 
        .C(n19002), .Y(n19335) );
  A2O1A1Ixp33_ASAP7_75t_SL U23376 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__6_), .B(n18295), .C(n19002), .Y(n19336)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U23377 ( .A1(n19335), .A2(n19336), .B(n18295), .C(
        n19002), .Y(n19337) );
  A2O1A1Ixp33_ASAP7_75t_SL U23378 ( .A1(n29863), .A2(
        u0_0_leon3x0_p0_iu_r_W__RESULT__6_), .B(n18295), .C(n19002), .Y(n19339) );
  A2O1A1Ixp33_ASAP7_75t_SL U23379 ( .A1(n19338), .A2(n19339), .B(n18295), .C(
        n19002), .Y(n19340) );
  A2O1A1Ixp33_ASAP7_75t_SL U23380 ( .A1(n23847), .A2(n24676), .B(n18295), .C(
        n19002), .Y(n19344) );
  A2O1A1Ixp33_ASAP7_75t_SL U23381 ( .A1(n29101), .A2(n24678), .B(n18295), .C(
        n19002), .Y(n19329) );
  A2O1A1Ixp33_ASAP7_75t_SL U23382 ( .A1(n24291), .A2(n19332), .B(n18295), .C(
        n19002), .Y(n19333) );
  A2O1A1Ixp33_ASAP7_75t_SL U23383 ( .A1(n19331), .A2(n19333), .B(n18295), .C(
        n19002), .Y(n19334) );
  A2O1A1Ixp33_ASAP7_75t_SL U23384 ( .A1(n24666), .A2(n32644), .B(n18295), .C(
        n19002), .Y(n19328) );
  A2O1A1Ixp33_ASAP7_75t_SL U23385 ( .A1(n30685), .A2(n24664), .B(n18295), .C(
        n19002), .Y(n19138) );
  A2O1A1Ixp33_ASAP7_75t_SL U23386 ( .A1(n18295), .A2(n19002), .B(n19132), .C(
        n19002), .Y(n24507) );
  A2O1A1Ixp33_ASAP7_75t_SL U23387 ( .A1(n24666), .A2(n32152), .B(n18295), .C(
        n19002), .Y(n19314) );
  A2O1A1Ixp33_ASAP7_75t_SL U23388 ( .A1(n24677), .A2(n19310), .B(n18295), .C(
        n19002), .Y(n19311) );
  A2O1A1Ixp33_ASAP7_75t_SL U23389 ( .A1(n32681), .A2(n22396), .B(n18295), .C(
        n19002), .Y(n19115) );
  A2O1A1Ixp33_ASAP7_75t_SL U23390 ( .A1(n29416), .A2(n29383), .B(n18295), .C(
        n19002), .Y(n19113) );
  A2O1A1Ixp33_ASAP7_75t_SL U23391 ( .A1(n30965), .A2(n24681), .B(n18295), .C(
        n19002), .Y(n19301) );
  A2O1A1Ixp33_ASAP7_75t_SL U23392 ( .A1(n31662), .A2(u0_0_leon3x0_p0_divi[49]), 
        .B(n18295), .C(n19002), .Y(n19299) );
  A2O1A1Ixp33_ASAP7_75t_SL U23393 ( .A1(n19298), .A2(n19299), .B(n18295), .C(
        n19002), .Y(n19300) );
  A2O1A1Ixp33_ASAP7_75t_SL U23394 ( .A1(n32786), .A2(n32835), .B(n18295), .C(
        n19002), .Y(n19296) );
  A2O1A1Ixp33_ASAP7_75t_SL U23395 ( .A1(n28108), .A2(n27946), .B(n18295), .C(
        n19002), .Y(n19105) );
  A2O1A1Ixp33_ASAP7_75t_SL U23396 ( .A1(n28108), .A2(n27951), .B(n18295), .C(
        n19002), .Y(n19104) );
  A2O1A1Ixp33_ASAP7_75t_SL U23397 ( .A1(n26085), .A2(n19293), .B(n18295), .C(
        n19002), .Y(n19294) );
  A2O1A1Ixp33_ASAP7_75t_SL U23398 ( .A1(n18295), .A2(n19002), .B(n19088), .C(
        n19002), .Y(n19089) );
  A2O1A1Ixp33_ASAP7_75t_SL U23399 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__14_), .A2(n19282), .B(n18295), .C(n19002), .Y(n19283) );
  A2O1A1Ixp33_ASAP7_75t_SL U23400 ( .A1(n32446), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[41]), .B(n18295), .C(n19002), .Y(n19276) );
  A2O1A1Ixp33_ASAP7_75t_SL U23401 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__8_), 
        .A2(n32447), .B(n18295), .C(n19002), .Y(n19277) );
  A2O1A1Ixp33_ASAP7_75t_SL U23402 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[8]), .A2(
        n32448), .B(n18295), .C(n19002), .Y(n19278) );
  A2O1A1Ixp33_ASAP7_75t_SL U23403 ( .A1(n19276), .A2(n19277), .B(n18295), .C(
        n19278), .Y(n19279) );
  A2O1A1Ixp33_ASAP7_75t_SL U23404 ( .A1(n33067), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__3_), .B(n18295), .C(n19002), 
        .Y(n19281) );
  A2O1A1Ixp33_ASAP7_75t_SL U23405 ( .A1(n32210), .A2(n32234), .B(n18295), .C(
        n19002), .Y(n19268) );
  A2O1A1Ixp33_ASAP7_75t_SL U23406 ( .A1(n19264), .A2(n19265), .B(n18295), .C(
        n19002), .Y(n19266) );
  A2O1A1Ixp33_ASAP7_75t_SL U23407 ( .A1(n32161), .A2(
        u0_0_leon3x0_p0_iu_r_X__CTRL__WREG_), .B(n18295), .C(n19002), .Y(
        n19267) );
  A2O1A1Ixp33_ASAP7_75t_SL U23408 ( .A1(n19266), .A2(n19267), .B(n18295), .C(
        n19002), .Y(rf_we_w) );
  A2O1A1Ixp33_ASAP7_75t_SL U23409 ( .A1(n25240), .A2(n25241), .B(n18295), .C(
        n19002), .Y(n19263) );
  A2O1A1Ixp33_ASAP7_75t_SL U23410 ( .A1(n3897), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[0]), .B(n18295), .C(n19002), .Y(n19262) );
  A2O1A1Ixp33_ASAP7_75t_SL U23411 ( .A1(n23091), .A2(n28131), .B(n18295), .C(
        n19002), .Y(n19258) );
  NAND2xp5_ASAP7_75t_SL U23412 ( .A(n22375), .B(
        u0_0_leon3x0_p0_iu_r_E__OP1__11_), .Y(n19259) );
  A2O1A1Ixp33_ASAP7_75t_SL U23413 ( .A1(n19258), .A2(n19259), .B(n18295), .C(
        n19002), .Y(n19260) );
  A2O1A1Ixp33_ASAP7_75t_SL U23414 ( .A1(n19242), .A2(DP_OP_1196_128_7433_n7), 
        .B(n18295), .C(n19002), .Y(n19248) );
  A2O1A1Ixp33_ASAP7_75t_SL U23415 ( .A1(n30909), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n19250) );
  A2O1A1Ixp33_ASAP7_75t_SL U23416 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_), .A2(n19250), .B(n18295), .C(
        n19002), .Y(n19251) );
  A2O1A1Ixp33_ASAP7_75t_SL U23417 ( .A1(n30908), .A2(n19251), .B(n18295), .C(
        n19002), .Y(n19252) );
  A2O1A1Ixp33_ASAP7_75t_SL U23418 ( .A1(n19002), .A2(uart1_uarto_SCALER__10_), 
        .B(n18295), .C(n19002), .Y(n19237) );
  A2O1A1Ixp33_ASAP7_75t_SL U23419 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__5_), .B(n18295), .C(n19002), .Y(
        n19232) );
  A2O1A1Ixp33_ASAP7_75t_SL U23420 ( .A1(n19228), .A2(n19230), .B(n18295), .C(
        n19002), .Y(n19231) );
  A2O1A1Ixp33_ASAP7_75t_SL U23421 ( .A1(n22392), .A2(n30721), .B(n18295), .C(
        n19002), .Y(n19217) );
  A2O1A1Ixp33_ASAP7_75t_SL U23422 ( .A1(n28847), .A2(n26376), .B(n18295), .C(
        n19002), .Y(n19012) );
  A2O1A1Ixp33_ASAP7_75t_SL U23423 ( .A1(n28574), .A2(n22392), .B(n18295), .C(
        n19002), .Y(n19010) );
  A2O1A1Ixp33_ASAP7_75t_SL U23424 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__22_), 
        .A2(n29060), .B(n18295), .C(n19002), .Y(n19004) );
  A2O1A1Ixp33_ASAP7_75t_SL U23425 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__26_), .B(n18295), .C(n19002), .Y(n19203) );
  A2O1A1Ixp33_ASAP7_75t_SL U23426 ( .A1(n28367), .A2(u0_0_leon3x0_p0_divi[57]), 
        .B(n18295), .C(n19002), .Y(n19206) );
  A2O1A1Ixp33_ASAP7_75t_SL U23427 ( .A1(n28378), .A2(u0_0_leon3x0_p0_divi[58]), 
        .B(n18295), .C(n19002), .Y(n19207) );
  A2O1A1Ixp33_ASAP7_75t_SL U23428 ( .A1(n19205), .A2(n19206), .B(n18295), .C(
        n19207), .Y(u0_0_leon3x0_p0_div0_vaddin1[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23429 ( .A1(n19194), .A2(n19197), .B(n18295), .C(
        n19002), .Y(n19202) );
  A2O1A1Ixp33_ASAP7_75t_SL U23430 ( .A1(n19201), .A2(n19202), .B(n18295), .C(
        n19002), .Y(mult_x_1196_n873) );
  A2O1A1Ixp33_ASAP7_75t_SL U23431 ( .A1(n19002), .A2(n27536), .B(n18295), .C(
        n19002), .Y(n19180) );
  A2O1A1Ixp33_ASAP7_75t_SL U23432 ( .A1(n31251), .A2(irqctrl0_r_IFORCE__0__13_), .B(n18295), .C(n19002), .Y(n19170) );
  A2O1A1Ixp33_ASAP7_75t_SL U23433 ( .A1(n31247), .A2(irqctrl0_r_IPEND__13_), 
        .B(n18295), .C(n19002), .Y(n19173) );
  A2O1A1Ixp33_ASAP7_75t_SL U23434 ( .A1(n31950), .A2(n30804), .B(n18295), .C(
        n19002), .Y(n19174) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U23435 ( .A1(n19172), .A2(n19173), .B(n18295), 
        .C(n19174), .D(apb0_r_CFGSEL_), .Y(n19175) );
  A2O1A1Ixp33_ASAP7_75t_SL U23436 ( .A1(n24638), .A2(n19002), .B(n18295), .C(
        n19002), .Y(n19159) );
  A2O1A1Ixp33_ASAP7_75t_SL U23437 ( .A1(n25014), .A2(n32197), .B(n18295), .C(
        n19002), .Y(n19147) );
  A2O1A1Ixp33_ASAP7_75t_SL U23438 ( .A1(n22378), .A2(n29100), .B(n18295), .C(
        n19002), .Y(n19146) );
  A2O1A1Ixp33_ASAP7_75t_SL U23439 ( .A1(n24659), .A2(n32646), .B(n18295), .C(
        n19002), .Y(n19141) );
  A2O1A1Ixp33_ASAP7_75t_SL U23440 ( .A1(n24659), .A2(n19139), .B(n18295), .C(
        n19002), .Y(n19140) );
  A2O1A1Ixp33_ASAP7_75t_SL U23441 ( .A1(n24663), .A2(n32602), .B(n18295), .C(
        n19002), .Y(n19136) );
  A2O1A1Ixp33_ASAP7_75t_SL U23442 ( .A1(n24660), .A2(n19133), .B(n18295), .C(
        n19002), .Y(n19134) );
  A2O1A1Ixp33_ASAP7_75t_SL U23443 ( .A1(n24674), .A2(n26783), .B(n18295), .C(
        n19002), .Y(n19129) );
  A2O1A1Ixp33_ASAP7_75t_SL U23444 ( .A1(n22378), .A2(n19124), .B(n18295), .C(
        n19002), .Y(n19125) );
  A2O1A1Ixp33_ASAP7_75t_SL U23445 ( .A1(u0_0_leon3x0_p0_iu_v_E__ET_), .A2(
        n19002), .B(n18295), .C(n19002), .Y(n19120) );
  A2O1A1Ixp33_ASAP7_75t_SL U23446 ( .A1(n24660), .A2(n19120), .B(n18295), .C(
        n19002), .Y(n19121) );
  A2O1A1Ixp33_ASAP7_75t_SL U23447 ( .A1(n19121), .A2(n19123), .B(n18295), .C(
        n19002), .Y(n3374) );
  A2O1A1Ixp33_ASAP7_75t_SL U23448 ( .A1(n22378), .A2(n19118), .B(n18295), .C(
        n19002), .Y(n19119) );
  A2O1A1Ixp33_ASAP7_75t_SL U23449 ( .A1(n24676), .A2(n19116), .B(n18295), .C(
        n19002), .Y(n19117) );
  A2O1A1Ixp33_ASAP7_75t_SL U23450 ( .A1(n31840), .A2(n26550), .B(n18295), .C(
        n19002), .Y(n19112) );
  A2O1A1Ixp33_ASAP7_75t_SL U23451 ( .A1(n27314), .A2(n19101), .B(n18295), .C(
        n19002), .Y(n19102) );
  A2O1A1Ixp33_ASAP7_75t_SL U23452 ( .A1(n31720), .A2(sr1_r_MCFG1__IOWS__2_), 
        .B(n18295), .C(n19002), .Y(n19090) );
  A2O1A1Ixp33_ASAP7_75t_SL U23453 ( .A1(sr1_r_WS__2_), .A2(n31760), .B(n18295), 
        .C(n19002), .Y(n19091) );
  A2O1A1Ixp33_ASAP7_75t_SL U23454 ( .A1(n19090), .A2(n19091), .B(n18295), .C(
        n19092), .Y(n19093) );
  A2O1A1Ixp33_ASAP7_75t_SL U23455 ( .A1(n31726), .A2(sr1_r_MCFG1__ROMRWS__2_), 
        .B(n18295), .C(n19002), .Y(n19095) );
  A2O1A1Ixp33_ASAP7_75t_SL U23456 ( .A1(n19094), .A2(n19095), .B(n18295), .C(
        n19002), .Y(n19096) );
  A2O1A1Ixp33_ASAP7_75t_SL U23457 ( .A1(n24694), .A2(n19096), .B(n18295), .C(
        n19002), .Y(n1725) );
  A2O1A1Ixp33_ASAP7_75t_SL U23458 ( .A1(n30640), .A2(rf_do_b[17]), .B(n18295), 
        .C(n19002), .Y(n19079) );
  A2O1A1Ixp33_ASAP7_75t_SL U23459 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__17_), .B(n18295), .C(n19002), .Y(n19080)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U23460 ( .A1(n19079), .A2(n19080), .B(n18295), .C(
        n19002), .Y(n19081) );
  A2O1A1Ixp33_ASAP7_75t_SL U23461 ( .A1(n19084), .A2(n30593), .B(n18295), .C(
        n19002), .Y(n19085) );
  A2O1A1Ixp33_ASAP7_75t_SL U23462 ( .A1(u0_0_leon3x0_p0_div0_r_NEG_), .A2(
        n29109), .B(n18295), .C(n29110), .Y(n19076) );
  A2O1A1Ixp33_ASAP7_75t_SL U23463 ( .A1(n22431), .A2(n19077), .B(n18295), .C(
        n19002), .Y(n29018) );
  A2O1A1Ixp33_ASAP7_75t_SL U23464 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__13_), .A2(n19072), .B(n18295), .C(n19002), .Y(n19073) );
  A2O1A1Ixp33_ASAP7_75t_SL U23465 ( .A1(n32423), .A2(n19068), .B(n18295), .C(
        n19002), .Y(n19069) );
  A2O1A1Ixp33_ASAP7_75t_SL U23466 ( .A1(n32609), .A2(n24643), .B(n18295), .C(
        n19002), .Y(n19070) );
  A2O1A1Ixp33_ASAP7_75t_SL U23467 ( .A1(n32318), .A2(dc_q[6]), .B(n18295), .C(
        n19002), .Y(n19071) );
  A2O1A1Ixp33_ASAP7_75t_SL U23468 ( .A1(n19069), .A2(n19070), .B(n18295), .C(
        n19071), .Y(dc_data[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U23469 ( .A1(n32209), .A2(n32234), .B(n18295), .C(
        n19002), .Y(n19065) );
  A2O1A1Ixp33_ASAP7_75t_SL U23470 ( .A1(uart1_r_TSHIFT__2_), .A2(
        uart1_r_TSHIFT__4_), .B(n18295), .C(n19002), .Y(n19056) );
  A2O1A1Ixp33_ASAP7_75t_SL U23471 ( .A1(uart1_r_TSHIFT__9_), .A2(
        uart1_r_TSHIFT__3_), .B(n18295), .C(n19002), .Y(n19057) );
  A2O1A1Ixp33_ASAP7_75t_SL U23472 ( .A1(n19058), .A2(uart1_r_TSHIFT__6_), .B(
        n18295), .C(uart1_r_TSHIFT__5_), .Y(n19059) );
  A2O1A1Ixp33_ASAP7_75t_SL U23473 ( .A1(uart1_r_TSHIFT__8_), .A2(
        uart1_r_TSHIFT__7_), .B(n18295), .C(n19060), .Y(n28037) );
  A2O1A1Ixp33_ASAP7_75t_SL U23474 ( .A1(add_x_735_n267), .A2(n18892), .B(
        n18295), .C(n19054), .Y(n19055) );
  A2O1A1Ixp33_ASAP7_75t_SL U23475 ( .A1(n28371), .A2(n24681), .B(n18295), .C(
        n19002), .Y(n19052) );
  A2O1A1Ixp33_ASAP7_75t_SL U23476 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_), .B(n18295), .C(n24873), .Y(
        n19044) );
  A2O1A1Ixp33_ASAP7_75t_SL U23477 ( .A1(n25234), .A2(n19049), .B(n18295), .C(
        n19002), .Y(n19050) );
  A2O1A1Ixp33_ASAP7_75t_SL U23478 ( .A1(n29059), .A2(u0_0_leon3x0_p0_ici[57]), 
        .B(n18295), .C(n19002), .Y(n19034) );
  A2O1A1Ixp33_ASAP7_75t_SL U23479 ( .A1(n19033), .A2(n19034), .B(n18295), .C(
        n19002), .Y(n19035) );
  A2O1A1Ixp33_ASAP7_75t_SL U23480 ( .A1(n19002), .A2(n19035), .B(n18295), .C(
        n19002), .Y(n19036) );
  A2O1A1Ixp33_ASAP7_75t_SL U23481 ( .A1(DP_OP_1196_128_7433_n6), .A2(
        DP_OP_1196_128_7433_n234), .B(n18295), .C(n19002), .Y(n19029) );
  A2O1A1Ixp33_ASAP7_75t_SL U23482 ( .A1(n30640), .A2(rf_do_b[0]), .B(n18295), 
        .C(n19002), .Y(n19023) );
  A2O1A1Ixp33_ASAP7_75t_SL U23483 ( .A1(n30641), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__0_), .B(n18295), .C(n19002), .Y(n19024)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U23484 ( .A1(n19023), .A2(n19024), .B(n18295), .C(
        n19002), .Y(n19025) );
  A2O1A1Ixp33_ASAP7_75t_SL U23485 ( .A1(n29863), .A2(
        u0_0_leon3x0_p0_iu_r_W__RESULT__0_), .B(n18295), .C(n19002), .Y(n19027) );
  A2O1A1Ixp33_ASAP7_75t_SL U23486 ( .A1(n19026), .A2(n19027), .B(n18295), .C(
        n19002), .Y(n19028) );
  A2O1A1Ixp33_ASAP7_75t_SL U23487 ( .A1(n32871), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[12]), .B(n18295), .C(n19002), .Y(n19021) );
  A2O1A1Ixp33_ASAP7_75t_SL U23488 ( .A1(n25659), .A2(n25676), .B(n18295), .C(
        n19002), .Y(n19019) );
  A2O1A1Ixp33_ASAP7_75t_SL U23489 ( .A1(DP_OP_1196_128_7433_n348), .A2(n19015), 
        .B(n18295), .C(n19002), .Y(n19016) );
  A2O1A1Ixp33_ASAP7_75t_SL U23490 ( .A1(n19002), .A2(n19009), .B(n18295), .C(
        n19002), .Y(DP_OP_1196_128_7433_n157) );
  A2O1A1Ixp33_ASAP7_75t_SL U23491 ( .A1(n29059), .A2(u0_0_leon3x0_p0_ici[50]), 
        .B(n18295), .C(n19002), .Y(n19005) );
  A2O1A1Ixp33_ASAP7_75t_SL U23492 ( .A1(n19004), .A2(n19005), .B(n18295), .C(
        n19002), .Y(n19006) );
  A2O1A1Ixp33_ASAP7_75t_SL U23493 ( .A1(n19002), .A2(n19006), .B(n18295), .C(
        n19002), .Y(n19007) );
  HB1xp67_ASAP7_75t_SL U23494 ( .A(n23089), .Y(n18296) );
  HB1xp67_ASAP7_75t_SL U23495 ( .A(u0_0_leon3x0_p0_muli[21]), .Y(n18297) );
  XNOR2x1_ASAP7_75t_SL U23496 ( .A(n22653), .B(n24302), .Y(n18721) );
  XNOR2x1_ASAP7_75t_SL U23497 ( .A(n24050), .B(n18394), .Y(mult_x_1196_n3151)
         );
  BUFx2_ASAP7_75t_SL U23498 ( .A(mult_x_1196_n1963), .Y(n18298) );
  INVx5_ASAP7_75t_SL U23499 ( .A(add_x_735_A_22_), .Y(n23968) );
  INVx2_ASAP7_75t_SL U23500 ( .A(n23661), .Y(n23659) );
  BUFx5_ASAP7_75t_SL U23501 ( .A(n23963), .Y(n18299) );
  INVx4_ASAP7_75t_SRAM U23502 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__9_), .Y(
        n27110) );
  NOR2x1p5_ASAP7_75t_SL U23503 ( .A(n18300), .B(n18702), .Y(mult_x_1196_n1133)
         );
  NOR2x1p5_ASAP7_75t_SL U23504 ( .A(mult_x_1196_n2884), .B(n23708), .Y(n18300)
         );
  XNOR2xp5_ASAP7_75t_SL U23505 ( .A(n23750), .B(n18301), .Y(mult_x_1196_n1787)
         );
  XNOR2xp5_ASAP7_75t_SL U23506 ( .A(n18302), .B(n22292), .Y(n18301) );
  INVx1_ASAP7_75t_SL U23507 ( .A(mult_x_1196_n2364), .Y(n18302) );
  BUFx2_ASAP7_75t_SL U23508 ( .A(n24256), .Y(n18303) );
  BUFx2_ASAP7_75t_SL U23509 ( .A(mult_x_1196_n2136), .Y(n18304) );
  BUFx2_ASAP7_75t_SL U23510 ( .A(n23536), .Y(n22720) );
  XNOR2x1_ASAP7_75t_SL U23511 ( .A(n24048), .B(n22448), .Y(mult_x_1196_n3115)
         );
  BUFx2_ASAP7_75t_SL U23512 ( .A(n24025), .Y(n18305) );
  XOR2x2_ASAP7_75t_SL U23513 ( .A(n23513), .B(n23596), .Y(n23512) );
  HB1xp67_ASAP7_75t_SL U23514 ( .A(n24072), .Y(n18306) );
  INVx8_ASAP7_75t_SL U23515 ( .A(n26917), .Y(n24048) );
  XOR2xp5_ASAP7_75t_SL U23516 ( .A(n22834), .B(n22835), .Y(mult_x_1196_n1793)
         );
  OAI22xp5_ASAP7_75t_SL U23517 ( .A1(mult_x_1196_n3224), .A2(n22953), .B1(
        mult_x_1196_n3223), .B2(n23984), .Y(n22834) );
  HB1xp67_ASAP7_75t_SL U23518 ( .A(n22395), .Y(n18307) );
  BUFx10_ASAP7_75t_SL U23519 ( .A(u0_0_leon3x0_p0_muli[19]), .Y(n24067) );
  XNOR2x2_ASAP7_75t_SL U23520 ( .A(n22589), .B(n18970), .Y(mult_x_1196_n1520)
         );
  NAND2x1_ASAP7_75t_SL U23521 ( .A(mult_x_1196_n328), .B(n22443), .Y(n23601)
         );
  NAND3x1_ASAP7_75t_SL U23522 ( .A(n23601), .B(n23237), .C(n23236), .Y(n23234)
         );
  OAI21xp5_ASAP7_75t_SL U23523 ( .A1(mult_x_1196_n225), .A2(mult_x_1196_n296), 
        .B(n23229), .Y(n21675) );
  OAI21xp5_ASAP7_75t_SL U23524 ( .A1(n22258), .A2(mult_x_1196_n297), .B(
        mult_x_1196_n298), .Y(mult_x_1196_n296) );
  XOR2x2_ASAP7_75t_SL U23525 ( .A(n23694), .B(mult_x_1196_n1088), .Y(
        mult_x_1196_n1062) );
  NAND2x1p5_ASAP7_75t_SL U23526 ( .A(mult_x_1196_n932), .B(n22221), .Y(
        mult_x_1196_n377) );
  NAND2xp5_ASAP7_75t_SL U23527 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__19_), .B(
        n18910), .Y(n23531) );
  HB1xp67_ASAP7_75t_SL U23528 ( .A(n24012), .Y(n18308) );
  HB1xp67_ASAP7_75t_SL U23529 ( .A(n24031), .Y(n18309) );
  INVx2_ASAP7_75t_SL U23530 ( .A(n23981), .Y(n18310) );
  INVx2_ASAP7_75t_SL U23531 ( .A(n18754), .Y(n18311) );
  NAND2x1p5_ASAP7_75t_SL U23532 ( .A(n18311), .B(n18310), .Y(n18753) );
  INVx2_ASAP7_75t_SL U23533 ( .A(n18312), .Y(u0_0_leon3x0_p0_muli[13]) );
  AOI21x1_ASAP7_75t_SL U23534 ( .A1(n18997), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__2_), .B(n30604), .Y(n18312) );
  XOR2x2_ASAP7_75t_SL U23535 ( .A(mult_x_1196_n2531), .B(n23271), .Y(n24265)
         );
  OAI22xp5_ASAP7_75t_SL U23536 ( .A1(mult_x_1196_n3107), .A2(n23100), .B1(
        n24002), .B2(mult_x_1196_n3106), .Y(mult_x_1196_n2531) );
  OAI21xp5_ASAP7_75t_SL U23537 ( .A1(n23831), .A2(n28904), .B(n18313), .Y(
        u0_0_leon3x0_p0_muli[14]) );
  NAND2x1_ASAP7_75t_SL U23538 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__3_), .B(
        n23831), .Y(n18313) );
  BUFx3_ASAP7_75t_SL U23539 ( .A(mult_x_1196_n1350), .Y(n18400) );
  OAI22x1_ASAP7_75t_SL U23540 ( .A1(n18654), .A2(mult_x_1196_n3108), .B1(
        mult_x_1196_n3107), .B2(n24002), .Y(n23500) );
  BUFx5_ASAP7_75t_SL U23541 ( .A(n23956), .Y(n18314) );
  BUFx3_ASAP7_75t_SL U23542 ( .A(mult_x_1196_n1522), .Y(n18315) );
  HB1xp67_ASAP7_75t_SL U23543 ( .A(u0_0_leon3x0_p0_muli[22]), .Y(n18316) );
  BUFx12f_ASAP7_75t_SL U23544 ( .A(n24018), .Y(n23141) );
  NAND2x1p5_ASAP7_75t_SL U23545 ( .A(n25140), .B(n25139), .Y(
        u0_0_leon3x0_p0_muli[48]) );
  INVx5_ASAP7_75t_SL U23546 ( .A(u0_0_leon3x0_p0_muli[48]), .Y(n22424) );
  MAJIxp5_ASAP7_75t_SL U23547 ( .A(mult_x_1196_n2555), .B(mult_x_1196_n2587), 
        .C(n23517), .Y(n23591) );
  OAI21xp5_ASAP7_75t_SL U23548 ( .A1(mult_x_1196_n3131), .A2(n18397), .B(
        n18317), .Y(mult_x_1196_n2555) );
  INVx1_ASAP7_75t_SL U23549 ( .A(n18318), .Y(n18317) );
  NOR2x1_ASAP7_75t_SL U23550 ( .A(n23996), .B(mult_x_1196_n3130), .Y(n18318)
         );
  XNOR2x2_ASAP7_75t_SL U23551 ( .A(n24072), .B(n23089), .Y(mult_x_1196_n2901)
         );
  OAI22x1_ASAP7_75t_SL U23552 ( .A1(mult_x_1196_n2895), .A2(n23116), .B1(
        n24025), .B2(mult_x_1196_n2894), .Y(mult_x_1196_n2323) );
  XNOR2x2_ASAP7_75t_SL U23553 ( .A(n23089), .B(n24065), .Y(mult_x_1196_n2894)
         );
  NOR2x1p5_ASAP7_75t_SL U23554 ( .A(n23387), .B(mult_x_1196_n387), .Y(n23386)
         );
  NAND2x1_ASAP7_75t_SL U23555 ( .A(n23386), .B(n23385), .Y(mult_x_1196_n308)
         );
  BUFx2_ASAP7_75t_SL U23556 ( .A(n23982), .Y(n18319) );
  NAND2xp5_ASAP7_75t_SL U23557 ( .A(mult_x_1196_n794), .B(mult_x_1196_n472), 
        .Y(n22491) );
  NAND2x1_ASAP7_75t_SL U23558 ( .A(mult_x_1196_n299), .B(mult_x_1196_n464), 
        .Y(mult_x_1196_n297) );
  XNOR2x1_ASAP7_75t_SL U23559 ( .A(n24073), .B(n22926), .Y(n18720) );
  INVx5_ASAP7_75t_SL U23560 ( .A(n18466), .Y(n24060) );
  XNOR2x1_ASAP7_75t_SL U23561 ( .A(n18320), .B(n22513), .Y(n22325) );
  XNOR2x1_ASAP7_75t_SL U23562 ( .A(n22608), .B(mult_x_1196_n1928), .Y(n18320)
         );
  NAND2x1_ASAP7_75t_SL U23563 ( .A(n22332), .B(n18321), .Y(mult_x_1196_n706)
         );
  INVx1_ASAP7_75t_SL U23564 ( .A(mult_x_1196_n1989), .Y(n18321) );
  XNOR2xp5_ASAP7_75t_SL U23565 ( .A(n23039), .B(n23037), .Y(mult_x_1196_n1989)
         );
  OAI21xp5_ASAP7_75t_SL U23566 ( .A1(n24247), .A2(n23740), .B(
        mult_x_1196_n1063), .Y(n24249) );
  INVx1_ASAP7_75t_SL U23567 ( .A(mult_x_1196_n1046), .Y(n24247) );
  XNOR2xp5_ASAP7_75t_SL U23568 ( .A(n18322), .B(n18417), .Y(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N54) );
  INVx1_ASAP7_75t_SL U23569 ( .A(n18418), .Y(n18322) );
  XNOR2xp5_ASAP7_75t_SL U23570 ( .A(n18324), .B(n18323), .Y(mult_x_1196_n933)
         );
  XOR2xp5_ASAP7_75t_SL U23571 ( .A(n22340), .B(mult_x_1196_n949), .Y(n18323)
         );
  INVx1_ASAP7_75t_SL U23572 ( .A(n22633), .Y(n18324) );
  XOR2x2_ASAP7_75t_SL U23573 ( .A(n23614), .B(n22600), .Y(mult_x_1196_n1434)
         );
  OAI22x1_ASAP7_75t_SL U23574 ( .A1(mult_x_1196_n3069), .A2(n23637), .B1(
        mult_x_1196_n3068), .B2(n24005), .Y(n23169) );
  HB1xp67_ASAP7_75t_SL U23575 ( .A(n23957), .Y(n18325) );
  HB1xp67_ASAP7_75t_SL U23576 ( .A(mult_x_1196_n2417), .Y(n18326) );
  HB1xp67_ASAP7_75t_SL U23577 ( .A(u0_0_leon3x0_p0_muli[27]), .Y(n18327) );
  INVx1_ASAP7_75t_SL U23578 ( .A(mult_x_1196_n1561), .Y(n18703) );
  INVx13_ASAP7_75t_SL U23579 ( .A(n22427), .Y(n23229) );
  BUFx2_ASAP7_75t_SL U23580 ( .A(mult_x_1196_n2379), .Y(n23940) );
  OAI22x1_ASAP7_75t_SL U23581 ( .A1(n22792), .A2(mult_x_1196_n3066), .B1(
        n24005), .B2(mult_x_1196_n3065), .Y(n18663) );
  XNOR2x1_ASAP7_75t_SL U23582 ( .A(n24074), .B(n22926), .Y(mult_x_1196_n2767)
         );
  NOR2x1_ASAP7_75t_SL U23583 ( .A(mult_x_1196_n2767), .B(n24041), .Y(n18715)
         );
  OAI22x1_ASAP7_75t_SL U23584 ( .A1(mult_x_1196_n3130), .A2(n24000), .B1(
        n23996), .B2(n18958), .Y(mult_x_1196_n2554) );
  NAND2x1p5_ASAP7_75t_SL U23585 ( .A(n25196), .B(n25195), .Y(add_x_735_A_14_)
         );
  NAND2xp33_ASAP7_75t_SRAM U23586 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__12_), 
        .B(n18910), .Y(n25100) );
  OAI22xp5_ASAP7_75t_SL U23587 ( .A1(mult_x_1196_n2926), .A2(n24022), .B1(
        n24020), .B2(mult_x_1196_n2925), .Y(mult_x_1196_n2354) );
  OAI22xp5_ASAP7_75t_SL U23588 ( .A1(n22251), .A2(mult_x_1196_n2818), .B1(
        mult_x_1196_n2819), .B2(n24034), .Y(mult_x_1196_n2253) );
  XNOR2xp5_ASAP7_75t_SL U23589 ( .A(n22395), .B(n22442), .Y(mult_x_1196_n2818)
         );
  OAI21xp5_ASAP7_75t_SL U23590 ( .A1(mult_x_1196_n760), .A2(n24262), .B(
        mult_x_1196_n761), .Y(mult_x_1196_n759) );
  NOR2x1_ASAP7_75t_SL U23591 ( .A(n18329), .B(n18328), .Y(n24262) );
  NOR2x1_ASAP7_75t_SL U23592 ( .A(mult_x_1196_n764), .B(mult_x_1196_n766), .Y(
        n18328) );
  INVx1_ASAP7_75t_SL U23593 ( .A(mult_x_1196_n765), .Y(n18329) );
  BUFx5_ASAP7_75t_SL U23594 ( .A(mult_x_1196_n1141), .Y(n18330) );
  MAJIxp5_ASAP7_75t_SL U23595 ( .A(n18331), .B(mult_x_1196_n2405), .C(
        mult_x_1196_n2341), .Y(mult_x_1196_n1052) );
  INVx1_ASAP7_75t_SL U23596 ( .A(n18333), .Y(n18331) );
  XNOR2xp5_ASAP7_75t_SL U23597 ( .A(n18333), .B(n18332), .Y(mult_x_1196_n1053)
         );
  XNOR2xp5_ASAP7_75t_SL U23598 ( .A(mult_x_1196_n2405), .B(mult_x_1196_n2341), 
        .Y(n18332) );
  NOR2x1_ASAP7_75t_SL U23599 ( .A(n18335), .B(n18334), .Y(n18333) );
  NOR2x1_ASAP7_75t_SL U23600 ( .A(mult_x_1196_n2849), .B(n23449), .Y(n18334)
         );
  NOR2x1_ASAP7_75t_SL U23601 ( .A(mult_x_1196_n2848), .B(n24030), .Y(n18335)
         );
  XNOR2x1_ASAP7_75t_SL U23602 ( .A(mult_x_1196_n1386), .B(n23852), .Y(n23058)
         );
  XNOR2x1_ASAP7_75t_SL U23603 ( .A(n23742), .B(n22557), .Y(mult_x_1196_n1386)
         );
  NAND3xp33_ASAP7_75t_SL U23604 ( .A(n18502), .B(n18504), .C(n18336), .Y(n4191) );
  NAND2xp5_ASAP7_75t_SL U23605 ( .A(n18338), .B(n18337), .Y(n18336) );
  NAND2xp5_ASAP7_75t_SL U23606 ( .A(mult_x_1196_n328), .B(n18343), .Y(n18337)
         );
  NOR2x1_ASAP7_75t_SL U23607 ( .A(n18506), .B(n18508), .Y(n18338) );
  OR2x2_ASAP7_75t_SL U23608 ( .A(mult_x_1196_n1844), .B(n18477), .Y(
        mult_x_1196_n815) );
  XNOR2xp5_ASAP7_75t_SL U23609 ( .A(n22886), .B(n18939), .Y(n18477) );
  BUFx5_ASAP7_75t_SL U23610 ( .A(n23073), .Y(n18339) );
  OAI22x1_ASAP7_75t_SL U23611 ( .A1(mult_x_1196_n2917), .A2(n22781), .B1(
        mult_x_1196_n2916), .B2(n24020), .Y(mult_x_1196_n2345) );
  XOR2xp5_ASAP7_75t_SL U23612 ( .A(mult_x_1196_n2281), .B(n18340), .Y(
        mult_x_1196_n1011) );
  XNOR2xp5_ASAP7_75t_SL U23613 ( .A(mult_x_1196_n2339), .B(n22995), .Y(n18340)
         );
  MAJIxp5_ASAP7_75t_SL U23614 ( .A(mult_x_1196_n2473), .B(mult_x_1196_n2377), 
        .C(mult_x_1196_n2409), .Y(mult_x_1196_n1156) );
  OAI22xp5_ASAP7_75t_SL U23615 ( .A1(mult_x_1196_n2949), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2948), .Y(mult_x_1196_n2377) );
  OAI21x1_ASAP7_75t_SL U23616 ( .A1(n24097), .A2(n24096), .B(mult_x_1196_n1113), .Y(n24099) );
  NAND2x1p5_ASAP7_75t_SL U23617 ( .A(n24098), .B(n24099), .Y(mult_x_1196_n1086) );
  BUFx5_ASAP7_75t_SL U23618 ( .A(n22509), .Y(n18341) );
  NAND2xp5_ASAP7_75t_SL U23619 ( .A(n18344), .B(n18343), .Y(n18975) );
  NAND3xp33_ASAP7_75t_SL U23620 ( .A(n18343), .B(n18344), .C(n18342), .Y(
        n18972) );
  INVx1_ASAP7_75t_SL U23621 ( .A(n18345), .Y(n18342) );
  INVxp67_ASAP7_75t_SL U23622 ( .A(n22258), .Y(n18343) );
  NOR2xp67_ASAP7_75t_SL U23623 ( .A(mult_x_1196_n294), .B(mult_x_1196_n297), 
        .Y(n18344) );
  INVx1_ASAP7_75t_SL U23624 ( .A(n18980), .Y(n18345) );
  HB1xp67_ASAP7_75t_SL U23625 ( .A(n24030), .Y(n18346) );
  XNOR2x1_ASAP7_75t_SL U23626 ( .A(n24056), .B(n18926), .Y(mult_x_1196_n3259)
         );
  XNOR2xp5_ASAP7_75t_SL U23627 ( .A(mult_x_1196_n1346), .B(mult_x_1196_n1352), 
        .Y(n22594) );
  MAJIxp5_ASAP7_75t_SL U23628 ( .A(n23137), .B(mult_x_1196_n2168), .C(
        mult_x_1196_n2509), .Y(mult_x_1196_n1352) );
  XNOR2x1_ASAP7_75t_SL U23629 ( .A(n23408), .B(mult_x_1196_n2471), .Y(n18690)
         );
  AO21x1_ASAP7_75t_SL U23630 ( .A1(n24007), .A2(n18550), .B(mult_x_1196_n3043), 
        .Y(mult_x_1196_n2471) );
  AOI21xp33_ASAP7_75t_SL U23631 ( .A1(n18932), .A2(n22676), .B(n23926), .Y(
        mult_x_1196_n430) );
  MAJIxp5_ASAP7_75t_SL U23632 ( .A(mult_x_1196_n984), .B(mult_x_1196_n986), 
        .C(mult_x_1196_n970), .Y(mult_x_1196_n965) );
  XNOR2xp5_ASAP7_75t_SL U23633 ( .A(n18347), .B(n22590), .Y(mult_x_1196_n964)
         );
  INVx1_ASAP7_75t_SL U23634 ( .A(mult_x_1196_n966), .Y(n18347) );
  XNOR2xp5_ASAP7_75t_SL U23635 ( .A(mult_x_1196_n970), .B(n18348), .Y(
        mult_x_1196_n966) );
  XNOR2xp5_ASAP7_75t_SL U23636 ( .A(n18349), .B(mult_x_1196_n984), .Y(n18348)
         );
  INVx1_ASAP7_75t_SL U23637 ( .A(mult_x_1196_n986), .Y(n18349) );
  BUFx2_ASAP7_75t_SL U23638 ( .A(n22206), .Y(n18394) );
  BUFx5_ASAP7_75t_SL U23639 ( .A(mult_x_1196_n496), .Y(n18350) );
  NAND2x1_ASAP7_75t_SL U23640 ( .A(n18352), .B(n18351), .Y(n18408) );
  INVx2_ASAP7_75t_SL U23641 ( .A(mult_x_1196_n2859), .Y(n18351) );
  INVx2_ASAP7_75t_SL U23642 ( .A(n24031), .Y(n18352) );
  INVx1_ASAP7_75t_SL U23643 ( .A(n18353), .Y(n21758) );
  HB1xp67_ASAP7_75t_SL U23644 ( .A(mult_x_1196_n534), .Y(n18353) );
  NOR2x1p5_ASAP7_75t_SL U23645 ( .A(mult_x_1196_n1820), .B(mult_x_1196_n1797), 
        .Y(mult_x_1196_n651) );
  INVx2_ASAP7_75t_SL U23646 ( .A(n23706), .Y(n23705) );
  HB1xp67_ASAP7_75t_SL U23647 ( .A(mult_x_1196_n1685), .Y(n18354) );
  BUFx2_ASAP7_75t_SL U23648 ( .A(n24008), .Y(n22540) );
  MAJIxp5_ASAP7_75t_SL U23649 ( .A(mult_x_1196_n1940), .B(n22307), .C(
        mult_x_1196_n1957), .Y(mult_x_1196_n1934) );
  XOR2xp5_ASAP7_75t_SL U23650 ( .A(n18355), .B(n22555), .Y(mult_x_1196_n1940)
         );
  INVx1_ASAP7_75t_SL U23651 ( .A(n23715), .Y(n18355) );
  BUFx8_ASAP7_75t_SL U23652 ( .A(u0_0_leon3x0_p0_muli[29]), .Y(n24055) );
  BUFx6f_ASAP7_75t_SL U23653 ( .A(n24000), .Y(n18397) );
  NOR2x1_ASAP7_75t_SL U23654 ( .A(mult_x_1196_n1597), .B(mult_x_1196_n1627), 
        .Y(n22855) );
  AO21x2_ASAP7_75t_SL U23655 ( .A1(n22856), .A2(mult_x_1196_n1624), .B(n22855), 
        .Y(mult_x_1196_n1586) );
  NAND2x2_ASAP7_75t_SL U23656 ( .A(mult_x_1196_n464), .B(mult_x_1196_n385), 
        .Y(mult_x_1196_n379) );
  INVx2_ASAP7_75t_SL U23657 ( .A(mult_x_1196_n1064), .Y(n22511) );
  AOI21xp5_ASAP7_75t_SL U23658 ( .A1(n23212), .A2(mult_x_1196_n360), .B(n23211), .Y(n22368) );
  MAJIxp5_ASAP7_75t_SL U23659 ( .A(mult_x_1196_n2308), .B(mult_x_1196_n2244), 
        .C(n18358), .Y(mult_x_1196_n927) );
  XNOR2xp5_ASAP7_75t_SL U23660 ( .A(n18357), .B(n18356), .Y(mult_x_1196_n928)
         );
  INVx1_ASAP7_75t_SL U23661 ( .A(mult_x_1196_n2308), .Y(n18356) );
  XNOR2xp5_ASAP7_75t_SL U23662 ( .A(n18358), .B(mult_x_1196_n2244), .Y(n18357)
         );
  OAI22xp5_ASAP7_75t_SL U23663 ( .A1(n18346), .A2(mult_x_1196_n2841), .B1(
        n18309), .B2(mult_x_1196_n2842), .Y(n18358) );
  NAND2x1p5_ASAP7_75t_SL U23664 ( .A(mult_x_1196_n1081), .B(mult_x_1196_n1084), 
        .Y(mult_x_1196_n482) );
  INVx4_ASAP7_75t_SL U23665 ( .A(n24689), .Y(n23559) );
  XNOR2xp5_ASAP7_75t_SL U23666 ( .A(mult_x_1196_n240), .B(n18359), .Y(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N50) );
  OAI21xp5_ASAP7_75t_SL U23667 ( .A1(mult_x_1196_n466), .A2(n22533), .B(
        mult_x_1196_n467), .Y(n18359) );
  OAI21x1_ASAP7_75t_SL U23668 ( .A1(mult_x_1196_n3099), .A2(n18654), .B(n18360), .Y(n23104) );
  NAND2x1p5_ASAP7_75t_SL U23669 ( .A(n22582), .B(n22583), .Y(n18360) );
  OAI22xp5_ASAP7_75t_SL U23670 ( .A1(n23839), .A2(n23831), .B1(n27110), .B2(
        n24689), .Y(u0_0_leon3x0_p0_muli[19]) );
  BUFx6f_ASAP7_75t_SL U23671 ( .A(u0_0_leon3x0_p0_muli[25]), .Y(n24059) );
  BUFx5_ASAP7_75t_SL U23672 ( .A(mult_x_1196_n464), .Y(n18361) );
  XNOR2x2_ASAP7_75t_SL U23673 ( .A(n22532), .B(n18362), .Y(mult_x_1196_n1013)
         );
  XNOR2xp5_ASAP7_75t_SL U23674 ( .A(mult_x_1196_n2156), .B(n22531), .Y(n18362)
         );
  INVx3_ASAP7_75t_SL U23675 ( .A(n23491), .Y(u0_0_leon3x0_p0_muli[45]) );
  INVx6_ASAP7_75t_SL U23676 ( .A(n23529), .Y(add_x_735_A_20_) );
  BUFx2_ASAP7_75t_SL U23677 ( .A(n23989), .Y(n18528) );
  XNOR2xp5_ASAP7_75t_SL U23678 ( .A(mult_x_1196_n1921), .B(mult_x_1196_n1902), 
        .Y(n23264) );
  XNOR2xp5_ASAP7_75t_SL U23679 ( .A(n23270), .B(n22625), .Y(mult_x_1196_n1902)
         );
  BUFx5_ASAP7_75t_SL U23680 ( .A(n23182), .Y(n18363) );
  XNOR2xp5_ASAP7_75t_SL U23681 ( .A(mult_x_1196_n1569), .B(mult_x_1196_n1571), 
        .Y(n23015) );
  MAJIxp5_ASAP7_75t_SL U23682 ( .A(mult_x_1196_n2577), .B(mult_x_1196_n2609), 
        .C(n23384), .Y(mult_x_1196_n1571) );
  OAI22x1_ASAP7_75t_SL U23683 ( .A1(n24007), .A2(mult_x_1196_n3052), .B1(
        n24005), .B2(mult_x_1196_n3051), .Y(mult_x_1196_n2480) );
  XNOR2xp5_ASAP7_75t_SL U23684 ( .A(n24081), .B(n24052), .Y(mult_x_1196_n3051)
         );
  BUFx3_ASAP7_75t_SL U23685 ( .A(n24029), .Y(n18390) );
  BUFx6f_ASAP7_75t_SL U23686 ( .A(u0_0_leon3x0_p0_muli[12]), .Y(n24075) );
  XOR2x2_ASAP7_75t_SL U23687 ( .A(n23616), .B(n23617), .Y(mult_x_1196_n1355)
         );
  HB1xp67_ASAP7_75t_SL U23688 ( .A(n24041), .Y(n18364) );
  HB1xp67_ASAP7_75t_SL U23689 ( .A(n23983), .Y(n18365) );
  BUFx2_ASAP7_75t_SL U23690 ( .A(n24226), .Y(n18366) );
  INVx5_ASAP7_75t_SL U23691 ( .A(add_x_735_A_14_), .Y(n23962) );
  XNOR2x1_ASAP7_75t_SL U23692 ( .A(n18605), .B(n18367), .Y(mult_x_1196_n1493)
         );
  XNOR2x1_ASAP7_75t_SL U23693 ( .A(mult_x_1196_n2451), .B(n24280), .Y(n18367)
         );
  INVx6_ASAP7_75t_SL U23694 ( .A(n18789), .Y(n24050) );
  XNOR2xp5_ASAP7_75t_SL U23695 ( .A(mult_x_1196_n2663), .B(n23400), .Y(n23399)
         );
  MAJIxp5_ASAP7_75t_SL U23696 ( .A(mult_x_1196_n1066), .B(mult_x_1196_n1068), 
        .C(n18369), .Y(mult_x_1196_n1042) );
  XOR2xp5_ASAP7_75t_SL U23697 ( .A(n18368), .B(mult_x_1196_n1066), .Y(
        mult_x_1196_n1043) );
  XNOR2xp5_ASAP7_75t_SL U23698 ( .A(mult_x_1196_n1068), .B(n18369), .Y(n18368)
         );
  XNOR2xp5_ASAP7_75t_SL U23699 ( .A(n18370), .B(n22611), .Y(n18369) );
  INVx1_ASAP7_75t_SL U23700 ( .A(mult_x_1196_n1049), .Y(n18370) );
  NAND2x2_ASAP7_75t_SL U23701 ( .A(n18956), .B(n24257), .Y(n24182) );
  BUFx8_ASAP7_75t_SL U23702 ( .A(u0_0_leon3x0_p0_muli[30]), .Y(n24054) );
  OAI22xp5_ASAP7_75t_SL U23703 ( .A1(n23843), .A2(n23831), .B1(n24689), .B2(
        n26889), .Y(u0_0_leon3x0_p0_muli[34]) );
  XNOR2x1_ASAP7_75t_SL U23704 ( .A(n24052), .B(n23952), .Y(mult_x_1196_n3255)
         );
  MAJIxp5_ASAP7_75t_SL U23705 ( .A(mult_x_1196_n1780), .B(mult_x_1196_n1810), 
        .C(mult_x_1196_n1791), .Y(mult_x_1196_n1781) );
  NAND2x1p5_ASAP7_75t_SL U23706 ( .A(n22830), .B(n18592), .Y(add_x_735_A_22_)
         );
  INVx2_ASAP7_75t_SL U23707 ( .A(n18529), .Y(n24291) );
  BUFx5_ASAP7_75t_SL U23708 ( .A(n24259), .Y(n18371) );
  MAJIxp5_ASAP7_75t_SL U23709 ( .A(n18373), .B(mult_x_1196_n2455), .C(
        mult_x_1196_n2391), .Y(mult_x_1196_n1638) );
  XNOR2xp5_ASAP7_75t_SL U23710 ( .A(n18373), .B(n18372), .Y(mult_x_1196_n1639)
         );
  XOR2xp5_ASAP7_75t_SL U23711 ( .A(mult_x_1196_n2391), .B(mult_x_1196_n2455), 
        .Y(n18372) );
  OAI22xp5_ASAP7_75t_SL U23712 ( .A1(n24039), .A2(mult_x_1196_n2803), .B1(
        mult_x_1196_n2802), .B2(n22391), .Y(n18373) );
  XNOR2xp5_ASAP7_75t_SL U23713 ( .A(mult_x_1196_n2010), .B(mult_x_1196_n2012), 
        .Y(n22804) );
  HB1xp67_ASAP7_75t_SL U23714 ( .A(n26683), .Y(n18374) );
  HB1xp67_ASAP7_75t_SL U23715 ( .A(n23071), .Y(n18375) );
  HB1xp67_ASAP7_75t_SL U23716 ( .A(n18633), .Y(n18376) );
  INVx1_ASAP7_75t_SL U23717 ( .A(mult_x_1196_n723), .Y(mult_x_1196_n721) );
  NAND2xp5_ASAP7_75t_SL U23718 ( .A(mult_x_1196_n2043), .B(mult_x_1196_n2030), 
        .Y(mult_x_1196_n723) );
  INVx1_ASAP7_75t_SL U23719 ( .A(n18971), .Y(mult_x_1196_n1535) );
  XOR2xp5_ASAP7_75t_SL U23720 ( .A(n18377), .B(n22435), .Y(n18971) );
  INVx1_ASAP7_75t_SL U23721 ( .A(mult_x_1196_n2608), .Y(n18377) );
  MAJIxp5_ASAP7_75t_SL U23722 ( .A(mult_x_1196_n1385), .B(n23306), .C(
        mult_x_1196_n1379), .Y(mult_x_1196_n1341) );
  MAJIxp5_ASAP7_75t_SL U23723 ( .A(mult_x_1196_n2604), .B(mult_x_1196_n2262), 
        .C(n23742), .Y(mult_x_1196_n1385) );
  MAJIxp5_ASAP7_75t_SL U23724 ( .A(n18379), .B(mult_x_1196_n971), .C(
        mult_x_1196_n957), .Y(mult_x_1196_n951) );
  XOR2xp5_ASAP7_75t_SL U23725 ( .A(n18379), .B(n18378), .Y(mult_x_1196_n952)
         );
  XNOR2xp5_ASAP7_75t_SL U23726 ( .A(mult_x_1196_n971), .B(mult_x_1196_n957), 
        .Y(n18378) );
  XNOR2xp5_ASAP7_75t_SL U23727 ( .A(mult_x_1196_n2246), .B(n22762), .Y(n18379)
         );
  HB1xp67_ASAP7_75t_SL U23728 ( .A(n25491), .Y(n18380) );
  BUFx5_ASAP7_75t_SL U23729 ( .A(n24205), .Y(n18381) );
  MAJIxp5_ASAP7_75t_SL U23730 ( .A(mult_x_1196_n2380), .B(n18383), .C(
        mult_x_1196_n2165), .Y(mult_x_1196_n1246) );
  XOR2xp5_ASAP7_75t_SL U23731 ( .A(n18382), .B(mult_x_1196_n2380), .Y(
        mult_x_1196_n1247) );
  XNOR2xp5_ASAP7_75t_SL U23732 ( .A(n18383), .B(mult_x_1196_n2165), .Y(n18382)
         );
  OAI22xp5_ASAP7_75t_SL U23733 ( .A1(mult_x_1196_n2920), .A2(n24022), .B1(
        mult_x_1196_n2919), .B2(n24020), .Y(n18383) );
  BUFx5_ASAP7_75t_SL U23734 ( .A(mult_x_1196_n771), .Y(n18384) );
  OAI22xp5_ASAP7_75t_SL U23735 ( .A1(n24030), .A2(n18622), .B1(n24031), .B2(
        mult_x_1196_n2870), .Y(n18772) );
  XNOR2x1_ASAP7_75t_SL U23736 ( .A(n24074), .B(n18385), .Y(n18622) );
  INVx3_ASAP7_75t_SL U23737 ( .A(n18771), .Y(n18385) );
  NAND2xp5_ASAP7_75t_SL U23738 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__13_), .B(
        n24685), .Y(n25196) );
  XNOR2x1_ASAP7_75t_SL U23739 ( .A(n24227), .B(n18386), .Y(mult_x_1196_n1497)
         );
  XNOR2x1_ASAP7_75t_SL U23740 ( .A(mult_x_1196_n2233), .B(n22714), .Y(n18386)
         );
  INVx1_ASAP7_75t_SRAM U23741 ( .A(n18932), .Y(mult_x_1196_n467) );
  OAI22x1_ASAP7_75t_SL U23742 ( .A1(mult_x_1196_n2890), .A2(n23116), .B1(
        n22983), .B2(mult_x_1196_n2889), .Y(mult_x_1196_n2318) );
  XNOR2xp5_ASAP7_75t_SL U23743 ( .A(n23089), .B(n24061), .Y(mult_x_1196_n2890)
         );
  BUFx2_ASAP7_75t_SL U23744 ( .A(n23439), .Y(n22565) );
  NOR2x2_ASAP7_75t_SL U23745 ( .A(mult_x_1196_n3167), .B(n23992), .Y(n23277)
         );
  XNOR2xp5_ASAP7_75t_SL U23746 ( .A(n18387), .B(n23510), .Y(n23509) );
  INVx1_ASAP7_75t_SL U23747 ( .A(mult_x_1196_n1147), .Y(n18387) );
  OAI22x1_ASAP7_75t_SL U23748 ( .A1(n23072), .A2(mult_x_1196_n3209), .B1(
        mult_x_1196_n3208), .B2(n24106), .Y(mult_x_1196_n2633) );
  BUFx5_ASAP7_75t_SL U23749 ( .A(n25644), .Y(n18388) );
  XNOR2x1_ASAP7_75t_SL U23750 ( .A(mult_x_1196_n2419), .B(n22932), .Y(n23648)
         );
  NOR2x1p5_ASAP7_75t_SL U23751 ( .A(n18716), .B(n18715), .Y(n22932) );
  XNOR2x1_ASAP7_75t_SL U23752 ( .A(n24181), .B(n18389), .Y(mult_x_1196_n1288)
         );
  XNOR2x1_ASAP7_75t_SL U23753 ( .A(n23856), .B(n23428), .Y(n18389) );
  BUFx5_ASAP7_75t_SL U23754 ( .A(n23303), .Y(n18391) );
  XNOR2xp5_ASAP7_75t_SL U23755 ( .A(n18392), .B(mult_x_1196_n1863), .Y(n23590)
         );
  INVx1_ASAP7_75t_SL U23756 ( .A(mult_x_1196_n1832), .Y(n18392) );
  NOR2x1_ASAP7_75t_SL U23757 ( .A(n22950), .B(n22951), .Y(mult_x_1196_n1832)
         );
  BUFx5_ASAP7_75t_SL U23758 ( .A(add_x_735_A_4_), .Y(n18393) );
  AOI21x1_ASAP7_75t_SL U23759 ( .A1(mult_x_1196_n668), .A2(n23451), .B(n18395), 
        .Y(mult_x_1196_n648) );
  OAI21x1_ASAP7_75t_SL U23760 ( .A1(mult_x_1196_n651), .A2(mult_x_1196_n655), 
        .B(mult_x_1196_n652), .Y(n18395) );
  BUFx5_ASAP7_75t_SL U23761 ( .A(mult_x_1196_n1596), .Y(n18396) );
  INVx1_ASAP7_75t_SL U23762 ( .A(add_x_735_A_22_), .Y(n24421) );
  NOR2x1p5_ASAP7_75t_SL U23763 ( .A(n18545), .B(n18544), .Y(n23746) );
  NOR2x1_ASAP7_75t_SL U23764 ( .A(n23224), .B(mult_x_1196_n411), .Y(n23223) );
  NOR2x1_ASAP7_75t_SL U23765 ( .A(n18398), .B(mult_x_1196_n418), .Y(
        mult_x_1196_n411) );
  INVx1_ASAP7_75t_SL U23766 ( .A(n18446), .Y(n18398) );
  BUFx3_ASAP7_75t_SL U23767 ( .A(mult_x_1196_n1807), .Y(n18415) );
  AND2x2_ASAP7_75t_SL U23768 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__10_), .B(n22434), .Y(n18544) );
  XNOR2x1_ASAP7_75t_SL U23769 ( .A(n23149), .B(n18986), .Y(mult_x_1196_n1486)
         );
  NAND2xp5_ASAP7_75t_SL U23770 ( .A(n18470), .B(n18579), .Y(n18577) );
  XNOR2xp5_ASAP7_75t_SL U23771 ( .A(n18578), .B(n23789), .Y(n18470) );
  XNOR2x1_ASAP7_75t_SL U23772 ( .A(n22978), .B(n18732), .Y(n18735) );
  XNOR2x1_ASAP7_75t_SL U23773 ( .A(n18736), .B(n22483), .Y(n22978) );
  XOR2xp5_ASAP7_75t_SL U23774 ( .A(mult_x_1196_n1879), .B(mult_x_1196_n1877), 
        .Y(n18722) );
  BUFx5_ASAP7_75t_SL U23775 ( .A(mult_x_1196_n785), .Y(n18399) );
  MAJIxp5_ASAP7_75t_SL U23776 ( .A(mult_x_1196_n1076), .B(mult_x_1196_n1097), 
        .C(mult_x_1196_n1099), .Y(mult_x_1196_n1068) );
  XOR2xp5_ASAP7_75t_SL U23777 ( .A(n23023), .B(mult_x_1196_n1080), .Y(
        mult_x_1196_n1076) );
  INVx2_ASAP7_75t_SL U23778 ( .A(n18361), .Y(mult_x_1196_n466) );
  NAND2x1_ASAP7_75t_SL U23779 ( .A(n23228), .B(n23226), .Y(n23218) );
  NAND2xp33_ASAP7_75t_SL U23780 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__6_), .B(
        n24685), .Y(n25113) );
  BUFx2_ASAP7_75t_SL U23781 ( .A(n18747), .Y(n18401) );
  XNOR2x1_ASAP7_75t_SL U23782 ( .A(n24074), .B(n23089), .Y(mult_x_1196_n2903)
         );
  XOR2x2_ASAP7_75t_SL U23783 ( .A(n23608), .B(mult_x_1196_n1712), .Y(
        mult_x_1196_n1690) );
  HB1xp67_ASAP7_75t_SL U23784 ( .A(n22251), .Y(n18402) );
  NAND3xp33_ASAP7_75t_SL U23785 ( .A(n18974), .B(n18972), .C(n18973), .Y(n4183) );
  HB1xp67_ASAP7_75t_SL U23786 ( .A(n22584), .Y(n18403) );
  INVx3_ASAP7_75t_SL U23787 ( .A(n18404), .Y(n24086) );
  NOR2x1p5_ASAP7_75t_SL U23788 ( .A(n22356), .B(mult_x_1196_n1648), .Y(n18404)
         );
  XNOR2xp5_ASAP7_75t_SL U23789 ( .A(n23778), .B(n18405), .Y(mult_x_1196_n1351)
         );
  XOR2xp5_ASAP7_75t_SL U23790 ( .A(mult_x_1196_n2571), .B(mult_x_1196_n2319), 
        .Y(n18405) );
  NOR2x1p5_ASAP7_75t_SL U23791 ( .A(n22251), .B(n18676), .Y(n23791) );
  INVx4_ASAP7_75t_SL U23792 ( .A(n18910), .Y(n18862) );
  BUFx5_ASAP7_75t_SL U23793 ( .A(n18374), .Y(n18406) );
  INVx1_ASAP7_75t_SL U23794 ( .A(n23137), .Y(n23139) );
  NAND2xp5_ASAP7_75t_SL U23795 ( .A(n18408), .B(n18407), .Y(n23137) );
  INVx1_ASAP7_75t_SL U23796 ( .A(n23140), .Y(n18407) );
  OAI22xp5_ASAP7_75t_SL U23797 ( .A1(n22743), .A2(mult_x_1196_n2852), .B1(
        mult_x_1196_n2853), .B2(n24031), .Y(n23913) );
  XNOR2xp5_ASAP7_75t_SL U23798 ( .A(n22897), .B(n22442), .Y(mult_x_1196_n2852)
         );
  OAI22x1_ASAP7_75t_SL U23799 ( .A1(mult_x_1196_n2752), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2751), .Y(n23824) );
  XNOR2x1_ASAP7_75t_SL U23800 ( .A(n23824), .B(mult_x_1196_n2157), .Y(n23823)
         );
  OAI21xp5_ASAP7_75t_SL U23801 ( .A1(n24646), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N59), .B(n25312), .Y(n4197) );
  INVx2_ASAP7_75t_SL U23802 ( .A(mult_x_1196_n2225), .Y(n23739) );
  INVx6_ASAP7_75t_SL U23803 ( .A(n24681), .Y(n22377) );
  NOR2x1_ASAP7_75t_SL U23804 ( .A(mult_x_1196_n2826), .B(n24035), .Y(n23790)
         );
  XNOR2xp5_ASAP7_75t_SL U23805 ( .A(n22395), .B(n24065), .Y(mult_x_1196_n2826)
         );
  NAND2xp5_ASAP7_75t_SL U23806 ( .A(n24112), .B(n18409), .Y(n24278) );
  OAI21xp5_ASAP7_75t_SL U23807 ( .A1(n22262), .A2(n24077), .B(
        mult_x_1196_n1801), .Y(n18409) );
  INVx8_ASAP7_75t_SL U23808 ( .A(n23619), .Y(n24046) );
  INVx2_ASAP7_75t_SL U23809 ( .A(mult_x_1196_n407), .Y(mult_x_1196_n405) );
  AOI21x1_ASAP7_75t_SL U23810 ( .A1(mult_x_1196_n784), .A2(mult_x_1196_n405), 
        .B(mult_x_1196_n396), .Y(mult_x_1196_n394) );
  XNOR2x2_ASAP7_75t_SL U23811 ( .A(mult_x_1196_n1767), .B(n22536), .Y(
        mult_x_1196_n1732) );
  XOR2x2_ASAP7_75t_SL U23812 ( .A(n24063), .B(n23397), .Y(n23421) );
  BUFx2_ASAP7_75t_SL U23813 ( .A(n24215), .Y(n18410) );
  XNOR2x1_ASAP7_75t_SL U23814 ( .A(n18411), .B(n23930), .Y(n23862) );
  XNOR2x1_ASAP7_75t_SL U23815 ( .A(n18412), .B(n23863), .Y(n18411) );
  INVx2_ASAP7_75t_SL U23816 ( .A(mult_x_1196_n1812), .Y(n18412) );
  XNOR2xp5_ASAP7_75t_SL U23817 ( .A(n24256), .B(mult_x_1196_n1834), .Y(n22888)
         );
  XOR2xp5_ASAP7_75t_SL U23818 ( .A(n18413), .B(n23590), .Y(mult_x_1196_n1834)
         );
  INVx1_ASAP7_75t_SL U23819 ( .A(n23591), .Y(n18413) );
  XNOR2x1_ASAP7_75t_SL U23820 ( .A(mult_x_1196_n1092), .B(n18562), .Y(
        mult_x_1196_n1094) );
  NOR2x1p5_ASAP7_75t_SL U23821 ( .A(n22792), .B(mult_x_1196_n3056), .Y(n23357)
         );
  INVx2_ASAP7_75t_SL U23822 ( .A(mult_x_1196_n3097), .Y(n23126) );
  BUFx5_ASAP7_75t_SL U23823 ( .A(n23959), .Y(n18414) );
  INVx2_ASAP7_75t_SL U23824 ( .A(n23373), .Y(n23113) );
  NOR3xp33_ASAP7_75t_SL U23825 ( .A(n24151), .B(n23374), .C(mult_x_1196_n3151), 
        .Y(n24166) );
  NOR2x1p5_ASAP7_75t_SL U23826 ( .A(n18611), .B(n23189), .Y(n23188) );
  XNOR2x1_ASAP7_75t_SL U23827 ( .A(mult_x_1196_n2436), .B(n23188), .Y(n23187)
         );
  INVx1_ASAP7_75t_SL U23828 ( .A(n23005), .Y(n23003) );
  BUFx6f_ASAP7_75t_SL U23829 ( .A(n24021), .Y(n22781) );
  XOR2x2_ASAP7_75t_SL U23830 ( .A(n23540), .B(n23539), .Y(mult_x_1196_n1091)
         );
  XOR2x1_ASAP7_75t_SL U23831 ( .A(mult_x_1196_n1091), .B(mult_x_1196_n1094), 
        .Y(n22972) );
  BUFx5_ASAP7_75t_SL U23832 ( .A(mult_x_1196_n787), .Y(n18416) );
  AND2x4_ASAP7_75t_SL U23833 ( .A(mult_x_1196_n2699), .B(mult_x_1196_n2635), 
        .Y(mult_x_1196_n2086) );
  OAI22x1_ASAP7_75t_SL U23834 ( .A1(mult_x_1196_n3211), .A2(n23989), .B1(
        mult_x_1196_n3210), .B2(n22248), .Y(mult_x_1196_n2635) );
  OAI21xp5_ASAP7_75t_SL U23835 ( .A1(mult_x_1196_n418), .A2(n22258), .B(n23134), .Y(n18417) );
  INVx1_ASAP7_75t_SL U23836 ( .A(mult_x_1196_n236), .Y(n18418) );
  XNOR2x1_ASAP7_75t_SL U23837 ( .A(n18419), .B(n22442), .Y(mult_x_1196_n2784)
         );
  INVx1_ASAP7_75t_SL U23838 ( .A(n23479), .Y(n18419) );
  HB1xp67_ASAP7_75t_SL U23839 ( .A(n25087), .Y(n18420) );
  XOR2x2_ASAP7_75t_SL U23840 ( .A(n18675), .B(n24190), .Y(mult_x_1196_n1730)
         );
  XOR2x2_ASAP7_75t_SL U23841 ( .A(n23397), .B(n24062), .Y(mult_x_1196_n3163)
         );
  NAND2x2_ASAP7_75t_SL U23842 ( .A(n25199), .B(n23640), .Y(mult_x_1196_n39) );
  INVx2_ASAP7_75t_SL U23843 ( .A(n18421), .Y(n23640) );
  NOR2x1_ASAP7_75t_SL U23844 ( .A(n27110), .B(n24686), .Y(n18421) );
  OAI22x1_ASAP7_75t_SL U23845 ( .A1(mult_x_1196_n2902), .A2(n24026), .B1(
        mult_x_1196_n2901), .B2(n24025), .Y(mult_x_1196_n2330) );
  NAND2x1p5_ASAP7_75t_SL U23846 ( .A(n18778), .B(n18777), .Y(mult_x_1196_n794)
         );
  OAI22x1_ASAP7_75t_SL U23847 ( .A1(n27257), .A2(n23559), .B1(n24689), .B2(
        n23551), .Y(u0_0_leon3x0_p0_muli[25]) );
  NOR2x1p5_ASAP7_75t_SL U23848 ( .A(mult_x_1196_n2985), .B(n23311), .Y(n18489)
         );
  NOR2x1p5_ASAP7_75t_SL U23849 ( .A(n30594), .B(n23559), .Y(n23621) );
  INVx2_ASAP7_75t_SL U23850 ( .A(n23621), .Y(n23620) );
  BUFx5_ASAP7_75t_SL U23851 ( .A(mult_x_1196_n489), .Y(n18422) );
  MAJIxp5_ASAP7_75t_SL U23852 ( .A(mult_x_1196_n1271), .B(mult_x_1196_n1274), 
        .C(mult_x_1196_n1264), .Y(mult_x_1196_n1265) );
  XNOR2xp5_ASAP7_75t_SL U23853 ( .A(mult_x_1196_n1269), .B(n22736), .Y(
        mult_x_1196_n1271) );
  BUFx5_ASAP7_75t_SL U23854 ( .A(n23968), .Y(n18423) );
  NAND2x1_ASAP7_75t_SL U23855 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__11_), .B(
        n23903), .Y(n25137) );
  XOR2x2_ASAP7_75t_SL U23856 ( .A(mult_x_1196_n2554), .B(n23135), .Y(
        mult_x_1196_n1836) );
  NAND2x1_ASAP7_75t_SL U23857 ( .A(n18737), .B(n18735), .Y(n24200) );
  INVx3_ASAP7_75t_SL U23858 ( .A(n22533), .Y(n23230) );
  NOR2x1p5_ASAP7_75t_SL U23859 ( .A(n23224), .B(n23230), .Y(n23222) );
  INVx1_ASAP7_75t_SL U23860 ( .A(mult_x_1196_n2256), .Y(n23654) );
  MAJIxp5_ASAP7_75t_SL U23861 ( .A(mult_x_1196_n2180), .B(mult_x_1196_n2241), 
        .C(mult_x_1196_n900), .Y(mult_x_1196_n885) );
  XOR2xp5_ASAP7_75t_SL U23862 ( .A(mult_x_1196_n886), .B(mult_x_1196_n898), 
        .Y(n22701) );
  XNOR2xp5_ASAP7_75t_SL U23863 ( .A(mult_x_1196_n2180), .B(n18424), .Y(
        mult_x_1196_n886) );
  XOR2xp5_ASAP7_75t_SL U23864 ( .A(mult_x_1196_n900), .B(mult_x_1196_n2241), 
        .Y(n18424) );
  NOR2x1p5_ASAP7_75t_SL U23865 ( .A(n18425), .B(n18436), .Y(n24422) );
  INVx2_ASAP7_75t_SL U23866 ( .A(n18426), .Y(n18425) );
  NAND2x1_ASAP7_75t_SL U23867 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__15_), .B(
        n22434), .Y(n18426) );
  XNOR2xp5_ASAP7_75t_SL U23868 ( .A(mult_x_1196_n1279), .B(mult_x_1196_n1283), 
        .Y(n22832) );
  OAI22x1_ASAP7_75t_SL U23869 ( .A1(n23394), .A2(n22464), .B1(
        mult_x_1196_n2882), .B2(n18305), .Y(mult_x_1196_n2313) );
  MAJIxp5_ASAP7_75t_SL U23870 ( .A(n18427), .B(mult_x_1196_n991), .C(
        mult_x_1196_n993), .Y(mult_x_1196_n969) );
  INVx1_ASAP7_75t_SL U23871 ( .A(n18429), .Y(n18427) );
  XNOR2xp5_ASAP7_75t_SL U23872 ( .A(mult_x_1196_n991), .B(n18428), .Y(
        mult_x_1196_n970) );
  XNOR2xp5_ASAP7_75t_SL U23873 ( .A(mult_x_1196_n993), .B(n18429), .Y(n18428)
         );
  XNOR2xp5_ASAP7_75t_SL U23874 ( .A(n23148), .B(n23145), .Y(n18429) );
  OAI21x1_ASAP7_75t_SL U23875 ( .A1(mult_x_1196_n678), .A2(mult_x_1196_n684), 
        .B(n24200), .Y(mult_x_1196_n677) );
  NOR2x1p5_ASAP7_75t_SL U23876 ( .A(n18737), .B(n18735), .Y(mult_x_1196_n678)
         );
  BUFx2_ASAP7_75t_SL U23877 ( .A(n23577), .Y(n22929) );
  XNOR2xp5_ASAP7_75t_SL U23878 ( .A(mult_x_1196_n230), .B(n18430), .Y(n18581)
         );
  OAI21xp5_ASAP7_75t_SL U23879 ( .A1(mult_x_1196_n350), .A2(n22533), .B(n18431), .Y(n18430) );
  INVx1_ASAP7_75t_SL U23880 ( .A(n18432), .Y(n18431) );
  NAND2xp5_ASAP7_75t_SL U23881 ( .A(n23670), .B(n23673), .Y(n18432) );
  NAND2x1p5_ASAP7_75t_SL U23882 ( .A(n18483), .B(n18482), .Y(n18591) );
  OAI21xp5_ASAP7_75t_SL U23883 ( .A1(n18434), .A2(n18433), .B(n22130), .Y(
        n4237) );
  XNOR2xp5_ASAP7_75t_SL U23884 ( .A(mult_x_1196_n251), .B(mult_x_1196_n566), 
        .Y(n18433) );
  INVx1_ASAP7_75t_SL U23885 ( .A(n22421), .Y(n18434) );
  AOI21x1_ASAP7_75t_SL U23886 ( .A1(n23577), .A2(mult_x_1196_n513), .B(
        mult_x_1196_n514), .Y(mult_x_1196_n223) );
  OAI21x1_ASAP7_75t_SL U23887 ( .A1(mult_x_1196_n582), .A2(n23745), .B(n23743), 
        .Y(n23577) );
  BUFx5_ASAP7_75t_SL U23888 ( .A(n24003), .Y(n18435) );
  BUFx10_ASAP7_75t_SL U23889 ( .A(u0_0_leon3x0_p0_muli[35]), .Y(n24047) );
  NOR2x1p5_ASAP7_75t_SL U23890 ( .A(n24686), .B(n26562), .Y(n18436) );
  INVx11_ASAP7_75t_SL U23891 ( .A(n24682), .Y(n24646) );
  BUFx3_ASAP7_75t_SL U23892 ( .A(mult_x_1196_n223), .Y(n22258) );
  OAI21x1_ASAP7_75t_SL U23893 ( .A1(mult_x_1196_n2787), .A2(n22412), .B(n23409), .Y(n23408) );
  BUFx5_ASAP7_75t_SL U23894 ( .A(mult_x_1196_n343), .Y(n18437) );
  AND2x4_ASAP7_75t_SL U23895 ( .A(n28380), .B(n23620), .Y(n23619) );
  OAI22x1_ASAP7_75t_SL U23896 ( .A1(mult_x_1196_n2878), .A2(n24026), .B1(
        n24025), .B2(mult_x_1196_n2877), .Y(mult_x_1196_n995) );
  XNOR2x1_ASAP7_75t_SL U23897 ( .A(n23089), .B(n24048), .Y(mult_x_1196_n2877)
         );
  BUFx6f_ASAP7_75t_SL U23898 ( .A(mult_x_1196_n126), .Y(n24034) );
  NAND2x1_ASAP7_75t_SL U23899 ( .A(n24147), .B(n24145), .Y(n24294) );
  XNOR2x1_ASAP7_75t_SL U23900 ( .A(n18612), .B(n24294), .Y(n18480) );
  OAI21xp5_ASAP7_75t_SL U23901 ( .A1(n18441), .A2(n18439), .B(n18438), .Y(
        n4239) );
  INVx1_ASAP7_75t_SL U23902 ( .A(n25277), .Y(n18438) );
  XNOR2xp5_ASAP7_75t_SL U23903 ( .A(n18440), .B(mult_x_1196_n577), .Y(n18439)
         );
  INVx1_ASAP7_75t_SL U23904 ( .A(n23908), .Y(n18440) );
  INVx1_ASAP7_75t_SL U23905 ( .A(n23229), .Y(n18441) );
  BUFx3_ASAP7_75t_SL U23906 ( .A(n24014), .Y(n18442) );
  OAI21xp5_ASAP7_75t_SL U23907 ( .A1(n18444), .A2(n18443), .B(n21677), .Y(
        n4233) );
  XNOR2xp5_ASAP7_75t_SL U23908 ( .A(mult_x_1196_n249), .B(mult_x_1196_n548), 
        .Y(n18443) );
  INVx1_ASAP7_75t_SL U23909 ( .A(n23229), .Y(n18444) );
  BUFx2_ASAP7_75t_SL U23910 ( .A(mult_x_1196_n1061), .Y(n18445) );
  OAI22x1_ASAP7_75t_SL U23911 ( .A1(mult_x_1196_n2855), .A2(n24031), .B1(
        n22743), .B2(mult_x_1196_n2854), .Y(mult_x_1196_n2289) );
  BUFx5_ASAP7_75t_SL U23912 ( .A(n23576), .Y(n18446) );
  INVx5_ASAP7_75t_SL U23913 ( .A(n18526), .Y(n22533) );
  XNOR2x1_ASAP7_75t_SL U23914 ( .A(n22511), .B(mult_x_1196_n1086), .Y(n22927)
         );
  OAI22x1_ASAP7_75t_SL U23915 ( .A1(mult_x_1196_n2970), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2969), .Y(mult_x_1196_n2398) );
  BUFx5_ASAP7_75t_SL U23916 ( .A(n18375), .Y(n18447) );
  XNOR2xp5_ASAP7_75t_SL U23917 ( .A(mult_x_1196_n246), .B(n18448), .Y(n18524)
         );
  XOR2xp5_ASAP7_75t_SL U23918 ( .A(n18449), .B(n18574), .Y(mult_x_1196_n1122)
         );
  INVx1_ASAP7_75t_SL U23919 ( .A(n23074), .Y(n18449) );
  OR2x2_ASAP7_75t_SL U23920 ( .A(mult_x_1196_n2983), .B(n23311), .Y(n18482) );
  AOI21x1_ASAP7_75t_SL U23921 ( .A1(n24310), .A2(mult_x_1196_n704), .B(
        mult_x_1196_n699), .Y(mult_x_1196_n697) );
  NAND2x1_ASAP7_75t_SL U23922 ( .A(n18555), .B(n18554), .Y(n24310) );
  BUFx5_ASAP7_75t_SL U23923 ( .A(mult_x_1196_n3227), .Y(n18450) );
  XNOR2x1_ASAP7_75t_SL U23924 ( .A(n18451), .B(n24238), .Y(n24259) );
  XNOR2x1_ASAP7_75t_SL U23925 ( .A(n18452), .B(mult_x_1196_n1240), .Y(n18451)
         );
  INVx2_ASAP7_75t_SL U23926 ( .A(mult_x_1196_n1270), .Y(n18452) );
  XNOR2x2_ASAP7_75t_SL U23927 ( .A(n24062), .B(n23089), .Y(mult_x_1196_n2891)
         );
  MAJIxp5_ASAP7_75t_SL U23928 ( .A(n22312), .B(mult_x_1196_n913), .C(
        mult_x_1196_n915), .Y(mult_x_1196_n907) );
  MAJIxp5_ASAP7_75t_SL U23929 ( .A(mult_x_1196_n921), .B(mult_x_1196_n911), 
        .C(n18454), .Y(mult_x_1196_n904) );
  XNOR2xp5_ASAP7_75t_SL U23930 ( .A(mult_x_1196_n921), .B(n18453), .Y(
        mult_x_1196_n905) );
  XOR2xp5_ASAP7_75t_SL U23931 ( .A(n18454), .B(mult_x_1196_n911), .Y(n18453)
         );
  XNOR2xp5_ASAP7_75t_SL U23932 ( .A(n18455), .B(n22312), .Y(n18454) );
  XNOR2xp5_ASAP7_75t_SL U23933 ( .A(n18456), .B(mult_x_1196_n913), .Y(n18455)
         );
  INVx1_ASAP7_75t_SL U23934 ( .A(mult_x_1196_n915), .Y(n18456) );
  OAI22xp5_ASAP7_75t_SL U23935 ( .A1(n23846), .A2(n23831), .B1(n24689), .B2(
        n26160), .Y(u0_0_leon3x0_p0_muli[23]) );
  XNOR2xp5_ASAP7_75t_SL U23936 ( .A(n18363), .B(n23178), .Y(mult_x_1196_n2009)
         );
  INVx8_ASAP7_75t_SL U23937 ( .A(n22424), .Y(n22395) );
  NAND2x1_ASAP7_75t_SL U23938 ( .A(mult_x_1196_n1093), .B(mult_x_1196_n1067), 
        .Y(n23693) );
  OAI22x1_ASAP7_75t_SL U23939 ( .A1(mult_x_1196_n2981), .A2(n24012), .B1(
        n23311), .B2(mult_x_1196_n2982), .Y(mult_x_1196_n2410) );
  INVx2_ASAP7_75t_SL U23940 ( .A(mult_x_1196_n2410), .Y(n23265) );
  OAI22x1_ASAP7_75t_SL U23941 ( .A1(n18537), .A2(mult_x_1196_n3005), .B1(
        mult_x_1196_n3004), .B2(n24011), .Y(mult_x_1196_n2433) );
  OAI22x1_ASAP7_75t_SL U23942 ( .A1(n18457), .A2(n24020), .B1(
        mult_x_1196_n2938), .B2(n24021), .Y(n23136) );
  OAI22xp5_ASAP7_75t_SL U23943 ( .A1(n18457), .A2(n24021), .B1(n24020), .B2(
        mult_x_1196_n2936), .Y(mult_x_1196_n2365) );
  XOR2x1_ASAP7_75t_SL U23944 ( .A(n18458), .B(n24074), .Y(n18457) );
  INVx3_ASAP7_75t_SL U23945 ( .A(n23969), .Y(n18458) );
  OAI22x1_ASAP7_75t_SL U23946 ( .A1(n23981), .A2(mult_x_1196_n3272), .B1(
        mult_x_1196_n3271), .B2(n23980), .Y(n18460) );
  INVx13_ASAP7_75t_SL U23947 ( .A(n18459), .Y(mult_x_1196_n2065) );
  XOR2xp5_ASAP7_75t_SL U23948 ( .A(mult_x_1196_n2632), .B(n18460), .Y(n23047)
         );
  MAJx2_ASAP7_75t_SL U23949 ( .A(mult_x_1196_n2632), .B(n18460), .C(n22331), 
        .Y(n18459) );
  MAJIxp5_ASAP7_75t_SL U23950 ( .A(n18461), .B(mult_x_1196_n1386), .C(
        mult_x_1196_n1380), .Y(mult_x_1196_n1368) );
  INVx1_ASAP7_75t_SL U23951 ( .A(n23852), .Y(n18461) );
  MAJx2_ASAP7_75t_SL U23952 ( .A(n23419), .B(mult_x_1196_n2231), .C(
        mult_x_1196_n2637), .Y(n23852) );
  XNOR2x1_ASAP7_75t_SL U23953 ( .A(n18462), .B(n22660), .Y(mult_x_1196_n982)
         );
  XOR2xp5_ASAP7_75t_SL U23954 ( .A(mult_x_1196_n1005), .B(mult_x_1196_n987), 
        .Y(n18462) );
  MAJIxp5_ASAP7_75t_SL U23955 ( .A(n22351), .B(mult_x_1196_n1353), .C(n22684), 
        .Y(n18463) );
  XNOR2xp5_ASAP7_75t_SL U23956 ( .A(mult_x_1196_n1310), .B(n18463), .Y(n22836)
         );
  MAJIxp5_ASAP7_75t_SL U23957 ( .A(mult_x_1196_n1308), .B(mult_x_1196_n1310), 
        .C(n18463), .Y(mult_x_1196_n1299) );
  NOR2x2_ASAP7_75t_SL U23958 ( .A(n18465), .B(n18464), .Y(n18466) );
  NOR2x1p5_ASAP7_75t_SL U23959 ( .A(n26680), .B(n23829), .Y(n18464) );
  NOR2x1p5_ASAP7_75t_SL U23960 ( .A(n23841), .B(n18997), .Y(n18465) );
  INVx13_ASAP7_75t_SL U23961 ( .A(n18467), .Y(n18469) );
  NOR2x1p5_ASAP7_75t_SL U23962 ( .A(n18469), .B(n18468), .Y(
        u0_0_leon3x0_p0_divi[15]) );
  INVxp67_ASAP7_75t_SL U23963 ( .A(n26681), .Y(n18468) );
  OR2x2_ASAP7_75t_SL U23964 ( .A(n24060), .B(n28769), .Y(n18467) );
  AOI22xp5_ASAP7_75t_SL U23965 ( .A1(n28631), .A2(n24060), .B1(n28835), .B2(
        n30333), .Y(n26673) );
  OAI21xp5_ASAP7_75t_SL U23966 ( .A1(n23536), .A2(n18470), .B(
        mult_x_1196_n1341), .Y(n22654) );
  INVx1_ASAP7_75t_SL U23967 ( .A(n18470), .Y(mult_x_1196_n1321) );
  BUFx6f_ASAP7_75t_SL U23968 ( .A(n24020), .Y(n18471) );
  OAI22xp5_ASAP7_75t_SL U23969 ( .A1(mult_x_1196_n2911), .A2(n22781), .B1(
        n18471), .B2(mult_x_1196_n2910), .Y(mult_x_1196_n2339) );
  OAI22xp5_ASAP7_75t_SL U23970 ( .A1(mult_x_1196_n2909), .A2(n22781), .B1(
        n18471), .B2(mult_x_1196_n2908), .Y(mult_x_1196_n2337) );
  OAI22xp5_ASAP7_75t_SL U23971 ( .A1(mult_x_1196_n2912), .A2(n22487), .B1(
        n24020), .B2(mult_x_1196_n2911), .Y(mult_x_1196_n2340) );
  AO21x1_ASAP7_75t_SL U23972 ( .A1(n18471), .A2(n22487), .B(mult_x_1196_n2907), 
        .Y(mult_x_1196_n2335) );
  OAI21xp5_ASAP7_75t_SL U23973 ( .A1(mult_x_1196_n1921), .A2(mult_x_1196_n1902), .B(n18472), .Y(n23204) );
  NAND2xp5_ASAP7_75t_SL U23974 ( .A(n18473), .B(mult_x_1196_n1918), .Y(n18472)
         );
  MAJIxp5_ASAP7_75t_SL U23975 ( .A(mult_x_1196_n1924), .B(mult_x_1196_n1943), 
        .C(n23761), .Y(mult_x_1196_n1918) );
  XNOR2xp5_ASAP7_75t_SL U23976 ( .A(n24148), .B(n23762), .Y(n23761) );
  MAJIxp5_ASAP7_75t_SL U23977 ( .A(n23578), .B(mult_x_1196_n2559), .C(n23199), 
        .Y(mult_x_1196_n1943) );
  XNOR2xp5_ASAP7_75t_SL U23978 ( .A(n23566), .B(n18621), .Y(mult_x_1196_n1924)
         );
  NAND2xp5_ASAP7_75t_SL U23979 ( .A(mult_x_1196_n1921), .B(mult_x_1196_n1902), 
        .Y(n18473) );
  INVx1_ASAP7_75t_SL U23980 ( .A(n22691), .Y(n18474) );
  OR2x2_ASAP7_75t_SL U23981 ( .A(n18474), .B(mult_x_1196_n2062), .Y(
        mult_x_1196_n829) );
  XNOR2xp5_ASAP7_75t_SL U23982 ( .A(mult_x_1196_n2064), .B(n18475), .Y(
        mult_x_1196_n2062) );
  XNOR2xp5_ASAP7_75t_SL U23983 ( .A(mult_x_1196_n2071), .B(n23046), .Y(n18475)
         );
  XOR2xp5_ASAP7_75t_SL U23984 ( .A(n18476), .B(n18965), .Y(mult_x_1196_n2064)
         );
  INVx1_ASAP7_75t_SL U23985 ( .A(n18967), .Y(n18476) );
  NAND2xp5_ASAP7_75t_SL U23986 ( .A(n18477), .B(mult_x_1196_n1844), .Y(n22242)
         );
  NAND2xp5_ASAP7_75t_SL U23987 ( .A(mult_x_1196_n788), .B(n23573), .Y(n23499)
         );
  OR2x2_ASAP7_75t_SL U23988 ( .A(mult_x_1196_n1036), .B(mult_x_1196_n1017), 
        .Y(n23573) );
  XOR2xp5_ASAP7_75t_SL U23989 ( .A(n18478), .B(n18479), .Y(mult_x_1196_n1017)
         );
  INVx1_ASAP7_75t_SL U23990 ( .A(mult_x_1196_n1020), .Y(n18478) );
  OR2x2_ASAP7_75t_SL U23991 ( .A(mult_x_1196_n1016), .B(mult_x_1196_n998), .Y(
        mult_x_1196_n788) );
  XNOR2xp5_ASAP7_75t_SL U23992 ( .A(n18613), .B(n18480), .Y(mult_x_1196_n998)
         );
  XNOR2xp5_ASAP7_75t_SL U23993 ( .A(n22499), .B(mult_x_1196_n1039), .Y(n18479)
         );
  XNOR2xp5_ASAP7_75t_SL U23994 ( .A(mult_x_1196_n1022), .B(n23687), .Y(n18613)
         );
  NOR2x1_ASAP7_75t_SL U23995 ( .A(n18977), .B(n18481), .Y(n18976) );
  AOI21xp5_ASAP7_75t_SL U23996 ( .A1(n18481), .A2(n18980), .B(n18979), .Y(
        n18973) );
  OAI21xp5_ASAP7_75t_SL U23997 ( .A1(mult_x_1196_n294), .A2(mult_x_1196_n298), 
        .B(mult_x_1196_n295), .Y(n18481) );
  INVxp67_ASAP7_75t_SL U23998 ( .A(n23828), .Y(n18483) );
  XNOR2xp5_ASAP7_75t_SL U23999 ( .A(n18484), .B(n18591), .Y(n23827) );
  INVx1_ASAP7_75t_SL U24000 ( .A(mult_x_1196_n2347), .Y(n18484) );
  NOR2x1_ASAP7_75t_SL U24001 ( .A(n18485), .B(n24034), .Y(n18768) );
  OAI22x1_ASAP7_75t_SL U24002 ( .A1(n24035), .A2(mult_x_1196_n2828), .B1(
        n22251), .B2(n18485), .Y(mult_x_1196_n2262) );
  XNOR2x1_ASAP7_75t_SL U24003 ( .A(n22395), .B(n24066), .Y(n18485) );
  MAJIxp5_ASAP7_75t_SL U24004 ( .A(n18486), .B(mult_x_1196_n2445), .C(
        mult_x_1196_n2381), .Y(mult_x_1196_n1281) );
  INVx1_ASAP7_75t_SL U24005 ( .A(n18488), .Y(n18486) );
  XNOR2xp5_ASAP7_75t_SL U24006 ( .A(n18488), .B(n18487), .Y(mult_x_1196_n1282)
         );
  XNOR2xp5_ASAP7_75t_SL U24007 ( .A(mult_x_1196_n2381), .B(mult_x_1196_n2445), 
        .Y(n18487) );
  NOR2x1_ASAP7_75t_SL U24008 ( .A(n18490), .B(n18489), .Y(n18488) );
  NOR2x1_ASAP7_75t_SL U24009 ( .A(mult_x_1196_n2984), .B(n24011), .Y(n18490)
         );
  BUFx6f_ASAP7_75t_SL U24010 ( .A(n22395), .Y(n18491) );
  XNOR2xp5_ASAP7_75t_SL U24011 ( .A(n18491), .B(n24054), .Y(mult_x_1196_n2815)
         );
  XNOR2xp5_ASAP7_75t_SL U24012 ( .A(n22395), .B(n24053), .Y(mult_x_1196_n2814)
         );
  XNOR2xp5_ASAP7_75t_SL U24013 ( .A(n22395), .B(n24058), .Y(mult_x_1196_n2819)
         );
  XNOR2xp5_ASAP7_75t_SL U24014 ( .A(n18491), .B(n18615), .Y(mult_x_1196_n2810)
         );
  XNOR2xp5_ASAP7_75t_SL U24015 ( .A(n22395), .B(n18534), .Y(mult_x_1196_n2820)
         );
  NAND2xp5_ASAP7_75t_SL U24016 ( .A(n18491), .B(u0_0_leon3x0_p0_divi[26]), .Y(
        add_x_735_n75) );
  NOR2x1_ASAP7_75t_SL U24017 ( .A(n18491), .B(u0_0_leon3x0_p0_divi[26]), .Y(
        add_x_735_n74) );
  XNOR2xp5_ASAP7_75t_SL U24018 ( .A(n18491), .B(n18541), .Y(mult_x_1196_n2805)
         );
  NAND2xp5_ASAP7_75t_SL U24019 ( .A(n18491), .B(n24577), .Y(n25466) );
  AOI22xp5_ASAP7_75t_SL U24020 ( .A1(n23091), .A2(n24578), .B1(n18491), .B2(
        n28982), .Y(n28871) );
  NAND2xp5_ASAP7_75t_SL U24021 ( .A(n18492), .B(n26891), .Y(n26892) );
  OAI22xp5_ASAP7_75t_SL U24022 ( .A1(n24572), .A2(n18493), .B1(n18491), .B2(
        n29148), .Y(n18492) );
  INVx1_ASAP7_75t_SL U24023 ( .A(n29150), .Y(n18493) );
  INVx1_ASAP7_75t_SL U24024 ( .A(n18491), .Y(n24572) );
  NAND2xp5_ASAP7_75t_SL U24025 ( .A(n18491), .B(n28402), .Y(n26340) );
  AOI22xp5_ASAP7_75t_SL U24026 ( .A1(n18491), .A2(n29583), .B1(n26950), .B2(
        n29598), .Y(n26900) );
  NOR2x1_ASAP7_75t_SL U24027 ( .A(n18494), .B(n21135), .Y(n3005) );
  INVx1_ASAP7_75t_SL U24028 ( .A(n18495), .Y(n18494) );
  XNOR2x2_ASAP7_75t_SL U24029 ( .A(n24158), .B(n18496), .Y(mult_x_1196_n1159)
         );
  XNOR2xp5_ASAP7_75t_SL U24030 ( .A(mult_x_1196_n2162), .B(n23913), .Y(n18496)
         );
  XNOR2x1_ASAP7_75t_SL U24031 ( .A(n18499), .B(n18497), .Y(mult_x_1196_n1148)
         );
  XNOR2xp5_ASAP7_75t_SL U24032 ( .A(mult_x_1196_n1159), .B(n22984), .Y(n18497)
         );
  XOR2xp5_ASAP7_75t_SL U24033 ( .A(n18498), .B(n18501), .Y(n22984) );
  INVx1_ASAP7_75t_SL U24034 ( .A(n23716), .Y(n18498) );
  INVx1_ASAP7_75t_SL U24035 ( .A(n22337), .Y(n18499) );
  XNOR2xp5_ASAP7_75t_SL U24036 ( .A(n18500), .B(mult_x_1196_n2345), .Y(n18501)
         );
  INVx1_ASAP7_75t_SL U24037 ( .A(mult_x_1196_n2223), .Y(n18500) );
  AOI31xp67_ASAP7_75t_SL U24038 ( .A1(mult_x_1196_n328), .A2(n23230), .A3(
        n18505), .B(n18503), .Y(n18502) );
  INVx1_ASAP7_75t_SL U24039 ( .A(n25316), .Y(n18503) );
  NAND2xp5_ASAP7_75t_SL U24040 ( .A(n18505), .B(n18508), .Y(n18504) );
  NOR2x1_ASAP7_75t_SL U24041 ( .A(n22427), .B(n18617), .Y(n18505) );
  NAND2xp5_ASAP7_75t_SL U24042 ( .A(n18507), .B(n18617), .Y(n18506) );
  INVx1_ASAP7_75t_SL U24043 ( .A(n22427), .Y(n18507) );
  NAND3xp33_ASAP7_75t_SL U24044 ( .A(n23682), .B(mult_x_1196_n331), .C(n23681), 
        .Y(n18508) );
  NAND2xp5_ASAP7_75t_SL U24045 ( .A(n18350), .B(n18509), .Y(mult_x_1196_n494)
         );
  NAND2xp5_ASAP7_75t_SL U24046 ( .A(n18510), .B(n18526), .Y(n18509) );
  INVx1_ASAP7_75t_SL U24047 ( .A(mult_x_1196_n495), .Y(n18510) );
  NAND2xp5_ASAP7_75t_SL U24048 ( .A(mult_x_1196_n485), .B(n18511), .Y(
        mult_x_1196_n483) );
  NAND2xp5_ASAP7_75t_SL U24049 ( .A(n18512), .B(n18526), .Y(n18511) );
  INVx1_ASAP7_75t_SL U24050 ( .A(mult_x_1196_n484), .Y(n18512) );
  NAND2xp5_ASAP7_75t_SL U24051 ( .A(mult_x_1196_n507), .B(n18513), .Y(
        mult_x_1196_n505) );
  NAND2xp5_ASAP7_75t_SL U24052 ( .A(n18514), .B(n18526), .Y(n18513) );
  INVx1_ASAP7_75t_SL U24053 ( .A(mult_x_1196_n506), .Y(n18514) );
  XNOR2xp5_ASAP7_75t_SL U24054 ( .A(n22342), .B(mult_x_1196_n1753), .Y(n23293)
         );
  XOR2xp5_ASAP7_75t_SL U24055 ( .A(mult_x_1196_n1760), .B(n24104), .Y(
        mult_x_1196_n1753) );
  MAJIxp5_ASAP7_75t_SL U24056 ( .A(mult_x_1196_n1425), .B(mult_x_1196_n1459), 
        .C(mult_x_1196_n1423), .Y(mult_x_1196_n1409) );
  XNOR2xp5_ASAP7_75t_SL U24057 ( .A(n23406), .B(n23404), .Y(mult_x_1196_n1423)
         );
  INVx8_ASAP7_75t_SL U24058 ( .A(n24681), .Y(n22428) );
  OAI21x1_ASAP7_75t_SL U24059 ( .A1(mult_x_1196_n648), .A2(n23455), .B(n18515), 
        .Y(n23700) );
  AOI21x1_ASAP7_75t_SL U24060 ( .A1(mult_x_1196_n639), .A2(n24304), .B(n23450), 
        .Y(n18515) );
  HB1xp67_ASAP7_75t_SL U24061 ( .A(n24201), .Y(n18516) );
  OAI21xp5_ASAP7_75t_SL U24062 ( .A1(mult_x_1196_n1520), .A2(n22329), .B(
        n23266), .Y(n22728) );
  OR2x2_ASAP7_75t_SL U24063 ( .A(mult_x_1196_n1525), .B(mult_x_1196_n1556), 
        .Y(n23266) );
  OAI22xp5_ASAP7_75t_SL U24064 ( .A1(n24005), .A2(mult_x_1196_n3045), .B1(
        mult_x_1196_n3046), .B2(n23637), .Y(mult_x_1196_n2474) );
  XNOR2xp5_ASAP7_75t_SL U24065 ( .A(n24046), .B(n24081), .Y(mult_x_1196_n3045)
         );
  INVx5_ASAP7_75t_SL U24066 ( .A(add_x_735_A_26_), .Y(n23970) );
  INVx13_ASAP7_75t_SL U24067 ( .A(n23970), .Y(n23971) );
  NAND2x1p5_ASAP7_75t_SL U24068 ( .A(n22294), .B(n22293), .Y(n23710) );
  INVx2_ASAP7_75t_SL U24069 ( .A(n23710), .Y(n23711) );
  AO21x2_ASAP7_75t_SL U24070 ( .A1(n23371), .A2(mult_x_1196_n1563), .B(n23370), 
        .Y(mult_x_1196_n1522) );
  BUFx2_ASAP7_75t_SL U24071 ( .A(n22792), .Y(n18561) );
  XNOR2xp5_ASAP7_75t_SL U24072 ( .A(n18518), .B(n18517), .Y(mult_x_1196_n1328)
         );
  XNOR2xp5_ASAP7_75t_SL U24073 ( .A(n24260), .B(mult_x_1196_n1362), .Y(n18517)
         );
  INVx1_ASAP7_75t_SL U24074 ( .A(n22905), .Y(n18518) );
  XNOR2xp5_ASAP7_75t_SL U24075 ( .A(mult_x_1196_n2266), .B(n18519), .Y(
        mult_x_1196_n1537) );
  XOR2xp5_ASAP7_75t_SL U24076 ( .A(mult_x_1196_n2324), .B(n23056), .Y(n18519)
         );
  MAJIxp5_ASAP7_75t_SL U24077 ( .A(mult_x_1196_n2166), .B(n18521), .C(
        mult_x_1196_n2508), .Y(mult_x_1196_n1285) );
  XOR2xp5_ASAP7_75t_SL U24078 ( .A(n18520), .B(mult_x_1196_n2508), .Y(
        mult_x_1196_n1286) );
  XNOR2xp5_ASAP7_75t_SL U24079 ( .A(n18521), .B(mult_x_1196_n2166), .Y(n18520)
         );
  OAI22xp5_ASAP7_75t_SL U24080 ( .A1(mult_x_1196_n2857), .A2(n24031), .B1(
        n24029), .B2(mult_x_1196_n2856), .Y(n18521) );
  AOI21x1_ASAP7_75t_SL U24081 ( .A1(mult_x_1196_n584), .A2(mult_x_1196_n597), 
        .B(n23744), .Y(n23743) );
  INVx2_ASAP7_75t_SL U24082 ( .A(n24259), .Y(n24184) );
  OAI22xp5_ASAP7_75t_SL U24083 ( .A1(n24230), .A2(mult_x_1196_n3153), .B1(
        n23992), .B2(mult_x_1196_n3152), .Y(mult_x_1196_n2577) );
  XOR2xp5_ASAP7_75t_SL U24084 ( .A(n18522), .B(n22760), .Y(mult_x_1196_n1963)
         );
  INVx1_ASAP7_75t_SL U24085 ( .A(n23793), .Y(n18522) );
  XNOR2x1_ASAP7_75t_SL U24086 ( .A(n23488), .B(mult_x_1196_n1387), .Y(n18700)
         );
  XOR2xp5_ASAP7_75t_SL U24087 ( .A(mult_x_1196_n1328), .B(n18523), .Y(n23338)
         );
  XNOR2xp5_ASAP7_75t_SL U24088 ( .A(n23636), .B(mult_x_1196_n1359), .Y(n18523)
         );
  OAI21xp5_ASAP7_75t_SL U24089 ( .A1(n18525), .A2(n18524), .B(n21188), .Y(
        n4227) );
  INVx1_ASAP7_75t_SL U24090 ( .A(n22421), .Y(n18525) );
  INVx2_ASAP7_75t_SL U24091 ( .A(mult_x_1196_n223), .Y(n18526) );
  INVx11_ASAP7_75t_SL U24092 ( .A(n24682), .Y(n22378) );
  XNOR2x1_ASAP7_75t_SL U24093 ( .A(n22566), .B(n18527), .Y(mult_x_1196_n1791)
         );
  XOR2x2_ASAP7_75t_SL U24094 ( .A(mult_x_1196_n2492), .B(n22243), .Y(n18527)
         );
  MAJIxp5_ASAP7_75t_SL U24095 ( .A(n22974), .B(mult_x_1196_n1408), .C(
        mult_x_1196_n1405), .Y(mult_x_1196_n1397) );
  INVx5_ASAP7_75t_SL U24096 ( .A(n23073), .Y(n24040) );
  XNOR2x2_ASAP7_75t_SL U24097 ( .A(n22285), .B(n25644), .Y(n23073) );
  INVx4_ASAP7_75t_SL U24098 ( .A(n24002), .Y(n22582) );
  OAI22x1_ASAP7_75t_SL U24099 ( .A1(mult_x_1196_n2893), .A2(n24026), .B1(
        mult_x_1196_n2892), .B2(n24025), .Y(n23585) );
  XNOR2xp5_ASAP7_75t_SL U24100 ( .A(mult_x_1196_n1516), .B(n23268), .Y(n23267)
         );
  XNOR2x2_ASAP7_75t_SL U24101 ( .A(n23269), .B(n23267), .Y(mult_x_1196_n1475)
         );
  NOR2x1_ASAP7_75t_SL U24102 ( .A(mult_x_1196_n2067), .B(mult_x_1196_n2070), 
        .Y(n18529) );
  BUFx5_ASAP7_75t_SL U24103 ( .A(add_x_735_A_32_), .Y(n18530) );
  INVx11_ASAP7_75t_SL U24104 ( .A(n24682), .Y(n22427) );
  INVx5_ASAP7_75t_SL U24105 ( .A(n18910), .Y(n24687) );
  NAND2x1p5_ASAP7_75t_SL U24106 ( .A(n18657), .B(n23112), .Y(n23368) );
  OAI22x1_ASAP7_75t_SL U24107 ( .A1(n22647), .A2(mult_x_1196_n3242), .B1(
        mult_x_1196_n3241), .B2(n23984), .Y(mult_x_1196_n2666) );
  INVx2_ASAP7_75t_SL U24108 ( .A(mult_x_1196_n2666), .Y(n23009) );
  BUFx5_ASAP7_75t_SL U24109 ( .A(n23920), .Y(n18531) );
  NOR2x1p5_ASAP7_75t_SL U24110 ( .A(n24005), .B(mult_x_1196_n3055), .Y(n23356)
         );
  NOR2x1p5_ASAP7_75t_SL U24111 ( .A(n23357), .B(n23356), .Y(n23355) );
  XOR2x2_ASAP7_75t_SL U24112 ( .A(mult_x_1196_n1421), .B(n24174), .Y(
        mult_x_1196_n1408) );
  XNOR2x1_ASAP7_75t_SL U24113 ( .A(n22395), .B(n24064), .Y(n18676) );
  BUFx5_ASAP7_75t_SL U24114 ( .A(n23829), .Y(n18532) );
  XNOR2x1_ASAP7_75t_SL U24115 ( .A(n22346), .B(mult_x_1196_n1229), .Y(n22773)
         );
  XNOR2xp5_ASAP7_75t_SL U24116 ( .A(mult_x_1196_n2170), .B(n23405), .Y(n23404)
         );
  BUFx5_ASAP7_75t_SL U24117 ( .A(n23573), .Y(n18533) );
  BUFx3_ASAP7_75t_SL U24118 ( .A(n24059), .Y(n18534) );
  HB1xp67_ASAP7_75t_SL U24119 ( .A(mult_x_1196_n617), .Y(n18535) );
  HB1xp67_ASAP7_75t_SL U24120 ( .A(n24023), .Y(n18536) );
  BUFx3_ASAP7_75t_SL U24121 ( .A(n24013), .Y(n18537) );
  HB1xp67_ASAP7_75t_SL U24122 ( .A(mult_x_1196_n1819), .Y(n18538) );
  HB1xp67_ASAP7_75t_SL U24123 ( .A(mult_x_1196_n810), .Y(n18539) );
  XOR2xp5_ASAP7_75t_SL U24124 ( .A(n23049), .B(n18540), .Y(mult_x_1196_n1809)
         );
  XNOR2xp5_ASAP7_75t_SL U24125 ( .A(mult_x_1196_n1835), .B(mult_x_1196_n1837), 
        .Y(n18540) );
  BUFx5_ASAP7_75t_SL U24126 ( .A(n24044), .Y(n18541) );
  MAJIxp5_ASAP7_75t_SL U24127 ( .A(mult_x_1196_n1080), .B(mult_x_1196_n2284), 
        .C(mult_x_1196_n2220), .Y(mult_x_1196_n1075) );
  NOR2x1_ASAP7_75t_SL U24128 ( .A(n24091), .B(n24092), .Y(mult_x_1196_n1080)
         );
  XNOR2xp5_ASAP7_75t_SL U24129 ( .A(mult_x_1196_n1671), .B(mult_x_1196_n1675), 
        .Y(n23440) );
  MAJIxp5_ASAP7_75t_SL U24130 ( .A(mult_x_1196_n2644), .B(mult_x_1196_n2328), 
        .C(mult_x_1196_n2238), .Y(mult_x_1196_n1675) );
  XNOR2x2_ASAP7_75t_SL U24131 ( .A(n23287), .B(n23285), .Y(mult_x_1196_n1127)
         );
  INVx2_ASAP7_75t_SL U24132 ( .A(mult_x_1196_n1127), .Y(n23864) );
  INVx1_ASAP7_75t_SL U24133 ( .A(n18542), .Y(n22281) );
  NOR2x1_ASAP7_75t_SL U24134 ( .A(n24040), .B(mult_x_1196_n2754), .Y(n18542)
         );
  XNOR2xp5_ASAP7_75t_SL U24135 ( .A(n24061), .B(n23975), .Y(mult_x_1196_n2754)
         );
  XNOR2x1_ASAP7_75t_SL U24136 ( .A(n18690), .B(n23407), .Y(mult_x_1196_n1098)
         );
  INVx1_ASAP7_75t_SL U24137 ( .A(n18543), .Y(n24268) );
  MAJIxp5_ASAP7_75t_SL U24138 ( .A(n23321), .B(n23127), .C(mult_x_1196_n1882), 
        .Y(n18543) );
  NAND3xp33_ASAP7_75t_SL U24139 ( .A(n23746), .B(n23640), .C(n25199), .Y(
        n23747) );
  INVx1_ASAP7_75t_SL U24140 ( .A(n25108), .Y(n18545) );
  OAI21x1_ASAP7_75t_SL U24141 ( .A1(mult_x_1196_n2864), .A2(n23449), .B(n18608), .Y(mult_x_1196_n2298) );
  OAI22x1_ASAP7_75t_SL U24142 ( .A1(n24106), .A2(mult_x_1196_n3184), .B1(
        n23522), .B2(mult_x_1196_n3185), .Y(mult_x_1196_n2609) );
  XOR2x2_ASAP7_75t_SL U24143 ( .A(mult_x_1196_n2609), .B(n23384), .Y(n23383)
         );
  XNOR2x1_ASAP7_75t_SL U24144 ( .A(mult_x_1196_n1340), .B(n22207), .Y(n18751)
         );
  XNOR2x1_ASAP7_75t_SL U24145 ( .A(n23718), .B(n18546), .Y(mult_x_1196_n1251)
         );
  XOR2x2_ASAP7_75t_SL U24146 ( .A(mult_x_1196_n2476), .B(mult_x_1196_n1255), 
        .Y(n18546) );
  BUFx3_ASAP7_75t_SL U24147 ( .A(mult_x_1196_n1694), .Y(n18913) );
  INVx1_ASAP7_75t_SL U24148 ( .A(mult_x_1196_n1350), .Y(n22709) );
  A2O1A1Ixp33_ASAP7_75t_SL U24149 ( .A1(n23778), .A2(mult_x_1196_n2319), .B(
        mult_x_1196_n2571), .C(n23776), .Y(mult_x_1196_n1350) );
  MAJIxp5_ASAP7_75t_SL U24150 ( .A(mult_x_1196_n1528), .B(n24255), .C(n23799), 
        .Y(mult_x_1196_n1490) );
  MAJIxp5_ASAP7_75t_SL U24151 ( .A(mult_x_1196_n2388), .B(mult_x_1196_n2356), 
        .C(mult_x_1196_n2452), .Y(mult_x_1196_n1528) );
  BUFx5_ASAP7_75t_SL U24152 ( .A(mult_x_1196_n1314), .Y(n18547) );
  XOR2x2_ASAP7_75t_SL U24153 ( .A(n23401), .B(n23399), .Y(mult_x_1196_n2058)
         );
  XNOR2x1_ASAP7_75t_SL U24154 ( .A(mult_x_1196_n2065), .B(mult_x_1196_n2058), 
        .Y(n22947) );
  XNOR2x1_ASAP7_75t_SL U24155 ( .A(n18548), .B(mult_x_1196_n2024), .Y(n22679)
         );
  INVx1_ASAP7_75t_SL U24156 ( .A(n22819), .Y(n18548) );
  INVx1_ASAP7_75t_SL U24157 ( .A(n18549), .Y(n22329) );
  NAND2xp5_ASAP7_75t_SL U24158 ( .A(mult_x_1196_n1556), .B(mult_x_1196_n1525), 
        .Y(n18549) );
  BUFx3_ASAP7_75t_SL U24159 ( .A(n24005), .Y(n18550) );
  INVx2_ASAP7_75t_SL U24160 ( .A(mult_x_1196_n1526), .Y(n22597) );
  MAJIxp5_ASAP7_75t_SL U24161 ( .A(n24078), .B(mult_x_1196_n1172), .C(
        mult_x_1196_n1169), .Y(mult_x_1196_n1139) );
  XNOR2xp5_ASAP7_75t_SL U24162 ( .A(n18551), .B(n23101), .Y(mult_x_1196_n1134)
         );
  INVx1_ASAP7_75t_SL U24163 ( .A(mult_x_1196_n1140), .Y(n18551) );
  XNOR2xp5_ASAP7_75t_SL U24164 ( .A(n24078), .B(n18552), .Y(mult_x_1196_n1140)
         );
  XNOR2xp5_ASAP7_75t_SL U24165 ( .A(n18553), .B(mult_x_1196_n1169), .Y(n18552)
         );
  INVx1_ASAP7_75t_SL U24166 ( .A(mult_x_1196_n1172), .Y(n18553) );
  NAND2x1p5_ASAP7_75t_SL U24167 ( .A(n25106), .B(n25105), .Y(
        u0_0_leon3x0_p0_muli[46]) );
  INVx1_ASAP7_75t_SL U24168 ( .A(mult_x_1196_n1968), .Y(n18554) );
  INVx2_ASAP7_75t_SL U24169 ( .A(mult_x_1196_n1969), .Y(n18555) );
  BUFx2_ASAP7_75t_SL U24170 ( .A(n24052), .Y(n18556) );
  BUFx12f_ASAP7_75t_SL U24171 ( .A(n24031), .Y(n23449) );
  XOR2x2_ASAP7_75t_SL U24172 ( .A(n22547), .B(n22546), .Y(n22208) );
  NAND2xp5_ASAP7_75t_SL U24173 ( .A(mult_x_1196_n1931), .B(mult_x_1196_n1911), 
        .Y(mult_x_1196_n684) );
  MAJIxp5_ASAP7_75t_SL U24174 ( .A(mult_x_1196_n1397), .B(mult_x_1196_n1367), 
        .C(mult_x_1196_n1365), .Y(mult_x_1196_n1359) );
  OAI22x1_ASAP7_75t_SL U24175 ( .A1(mult_x_1196_n2830), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2829), .Y(mult_x_1196_n2264) );
  XOR2x2_ASAP7_75t_SL U24176 ( .A(n23185), .B(mult_x_1196_n2264), .Y(n18626)
         );
  AND2x2_ASAP7_75t_SL U24177 ( .A(n18911), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__3_), .Y(n18601) );
  MAJIxp5_ASAP7_75t_SL U24178 ( .A(n18557), .B(mult_x_1196_n1606), .C(
        mult_x_1196_n1602), .Y(mult_x_1196_n1591) );
  INVx1_ASAP7_75t_SL U24179 ( .A(n22688), .Y(n18557) );
  MAJIxp5_ASAP7_75t_SL U24180 ( .A(n23439), .B(mult_x_1196_n1671), .C(
        mult_x_1196_n1675), .Y(n22688) );
  XNOR2x1_ASAP7_75t_SL U24181 ( .A(mult_x_1196_n2318), .B(n18656), .Y(n23789)
         );
  OAI21x1_ASAP7_75t_SL U24182 ( .A1(n23487), .A2(n22806), .B(n23485), .Y(
        n23484) );
  NOR2x1p5_ASAP7_75t_SL U24183 ( .A(n18945), .B(n18944), .Y(n23379) );
  INVx1_ASAP7_75t_SL U24184 ( .A(n23297), .Y(n23298) );
  XNOR2xp5_ASAP7_75t_SL U24185 ( .A(n23299), .B(n24108), .Y(n23297) );
  OAI22x1_ASAP7_75t_SL U24186 ( .A1(mult_x_1196_n3117), .A2(n23999), .B1(
        mult_x_1196_n3116), .B2(n23997), .Y(n23405) );
  BUFx5_ASAP7_75t_SL U24187 ( .A(n22351), .Y(n18558) );
  XNOR2xp5_ASAP7_75t_SL U24188 ( .A(n22699), .B(n24296), .Y(mult_x_1196_n2044)
         );
  XNOR2xp5_ASAP7_75t_SL U24189 ( .A(mult_x_1196_n2049), .B(n24116), .Y(n24296)
         );
  NOR2x2_ASAP7_75t_SL U24190 ( .A(n23423), .B(n23422), .Y(n23424) );
  OAI22x1_ASAP7_75t_SL U24191 ( .A1(n22647), .A2(mult_x_1196_n3241), .B1(
        mult_x_1196_n3240), .B2(n23984), .Y(mult_x_1196_n2665) );
  XNOR2x1_ASAP7_75t_SL U24192 ( .A(n23564), .B(mult_x_1196_n2665), .Y(n23563)
         );
  OAI22x1_ASAP7_75t_SL U24193 ( .A1(mult_x_1196_n3249), .A2(n23981), .B1(
        n22389), .B2(mult_x_1196_n3248), .Y(mult_x_1196_n2673) );
  XNOR2x1_ASAP7_75t_SL U24194 ( .A(n24046), .B(n18927), .Y(mult_x_1196_n3249)
         );
  BUFx3_ASAP7_75t_SL U24195 ( .A(n24006), .Y(n22792) );
  XOR2xp5_ASAP7_75t_SL U24196 ( .A(n18560), .B(n18559), .Y(mult_x_1196_n1956)
         );
  XNOR2xp5_ASAP7_75t_SL U24197 ( .A(mult_x_1196_n1975), .B(n22677), .Y(n18559)
         );
  INVx1_ASAP7_75t_SL U24198 ( .A(mult_x_1196_n1961), .Y(n18560) );
  XOR2xp5_ASAP7_75t_SL U24199 ( .A(n23240), .B(n18915), .Y(n23239) );
  XOR2xp5_ASAP7_75t_SL U24200 ( .A(n24224), .B(n22703), .Y(n23240) );
  XNOR2x1_ASAP7_75t_SL U24201 ( .A(n23094), .B(mult_x_1196_n1509), .Y(
        mult_x_1196_n1504) );
  NOR2x1p5_ASAP7_75t_SL U24202 ( .A(n22345), .B(mult_x_1196_n1504), .Y(
        mult_x_1196_n591) );
  INVx5_ASAP7_75t_SL U24203 ( .A(n18792), .Y(n24062) );
  XOR2xp5_ASAP7_75t_SL U24204 ( .A(mult_x_1196_n1100), .B(mult_x_1196_n1104), 
        .Y(n18562) );
  XNOR2x1_ASAP7_75t_SL U24205 ( .A(n18927), .B(n24054), .Y(mult_x_1196_n3257)
         );
  INVx2_ASAP7_75t_SL U24206 ( .A(mult_x_1196_n3257), .Y(n23290) );
  BUFx3_ASAP7_75t_SL U24207 ( .A(mult_x_1196_n2646), .Y(n18570) );
  BUFx5_ASAP7_75t_SL U24208 ( .A(n24019), .Y(n18563) );
  BUFx10_ASAP7_75t_SL U24209 ( .A(u0_0_leon3x0_p0_muli[33]), .Y(n24051) );
  NAND2x1_ASAP7_75t_SL U24210 ( .A(n18565), .B(n18564), .Y(mult_x_1196_n1383)
         );
  INVx1_ASAP7_75t_SL U24211 ( .A(n22938), .Y(n18564) );
  NAND2xp5_ASAP7_75t_SL U24212 ( .A(n22941), .B(n22940), .Y(n18565) );
  XNOR2x1_ASAP7_75t_SL U24213 ( .A(n23352), .B(n22709), .Y(n23351) );
  XNOR2x1_ASAP7_75t_SL U24214 ( .A(n23873), .B(n18566), .Y(n23352) );
  INVx2_ASAP7_75t_SL U24215 ( .A(mult_x_1196_n1323), .Y(n18566) );
  XNOR2xp5_ASAP7_75t_SL U24216 ( .A(mult_x_1196_n2468), .B(n23792), .Y(n22760)
         );
  XNOR2xp5_ASAP7_75t_SL U24217 ( .A(mult_x_1196_n1899), .B(n18721), .Y(
        mult_x_1196_n1877) );
  BUFx5_ASAP7_75t_SL U24218 ( .A(n22986), .Y(n18567) );
  NAND2x1p5_ASAP7_75t_SL U24219 ( .A(n25193), .B(n25192), .Y(
        u0_0_leon3x0_p0_muli[42]) );
  NOR2x1p5_ASAP7_75t_SL U24220 ( .A(mult_x_1196_n2996), .B(n23311), .Y(n23871)
         );
  BUFx5_ASAP7_75t_SL U24221 ( .A(n22220), .Y(n18568) );
  BUFx5_ASAP7_75t_SL U24222 ( .A(n30605), .Y(n18569) );
  XNOR2x1_ASAP7_75t_SL U24223 ( .A(n24217), .B(n24218), .Y(mult_x_1196_n1928)
         );
  OAI22x1_ASAP7_75t_SL U24224 ( .A1(mult_x_1196_n2866), .A2(n23449), .B1(
        n24030), .B2(mult_x_1196_n2865), .Y(mult_x_1196_n2300) );
  OAI22xp5_ASAP7_75t_SL U24225 ( .A1(n23992), .A2(mult_x_1196_n3146), .B1(
        mult_x_1196_n3147), .B2(n24287), .Y(mult_x_1196_n2571) );
  NAND3xp33_ASAP7_75t_SL U24226 ( .A(n18573), .B(n23227), .C(n18571), .Y(n4205) );
  NOR2x1_ASAP7_75t_SL U24227 ( .A(n23219), .B(n18572), .Y(n18571) );
  INVx1_ASAP7_75t_SL U24228 ( .A(n23218), .Y(n18572) );
  OAI21xp5_ASAP7_75t_SL U24229 ( .A1(n23223), .A2(n23222), .B(n23221), .Y(
        n18573) );
  XNOR2xp5_ASAP7_75t_SL U24230 ( .A(mult_x_1196_n1154), .B(mult_x_1196_n1156), 
        .Y(n18574) );
  NAND2x1_ASAP7_75t_SL U24231 ( .A(n18928), .B(mult_x_1196_n1745), .Y(
        mult_x_1196_n641) );
  NAND2x1p5_ASAP7_75t_SL U24232 ( .A(mult_x_1196_n555), .B(n18730), .Y(
        mult_x_1196_n549) );
  XNOR2xp5_ASAP7_75t_SL U24233 ( .A(n18575), .B(n22807), .Y(mult_x_1196_n1237)
         );
  INVx1_ASAP7_75t_SL U24234 ( .A(mult_x_1196_n1235), .Y(n18575) );
  OAI22x1_ASAP7_75t_SL U24235 ( .A1(n22953), .A2(mult_x_1196_n3238), .B1(
        mult_x_1196_n3237), .B2(n23984), .Y(mult_x_1196_n2662) );
  XNOR2x1_ASAP7_75t_SL U24236 ( .A(mult_x_1196_n2534), .B(mult_x_1196_n2662), 
        .Y(n22955) );
  BUFx5_ASAP7_75t_SL U24237 ( .A(n18399), .Y(n18576) );
  XNOR2xp5_ASAP7_75t_SL U24238 ( .A(n23965), .B(n24060), .Y(mult_x_1196_n2991)
         );
  XNOR2xp5_ASAP7_75t_SL U24239 ( .A(n22227), .B(n22449), .Y(mult_x_1196_n3245)
         );
  NAND2x1_ASAP7_75t_SL U24240 ( .A(n18577), .B(n22654), .Y(mult_x_1196_n1305)
         );
  INVx1_ASAP7_75t_SL U24241 ( .A(mult_x_1196_n2570), .Y(n18578) );
  INVx1_ASAP7_75t_SL U24242 ( .A(mult_x_1196_n1315), .Y(n18579) );
  INVx2_ASAP7_75t_SL U24243 ( .A(n22258), .Y(n22584) );
  XNOR2x1_ASAP7_75t_SL U24244 ( .A(n22903), .B(n24090), .Y(mult_x_1196_n1084)
         );
  OAI22x1_ASAP7_75t_SL U24245 ( .A1(n22251), .A2(mult_x_1196_n2838), .B1(
        n22918), .B2(n24034), .Y(mult_x_1196_n2130) );
  NAND2x1p5_ASAP7_75t_SL U24246 ( .A(n23104), .B(n23113), .Y(n24233) );
  NAND2x1p5_ASAP7_75t_SL U24247 ( .A(n18628), .B(n23435), .Y(n23434) );
  NAND2x1_ASAP7_75t_SL U24248 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__25_), .B(
        n24687), .Y(n23623) );
  XNOR2x1_ASAP7_75t_SL U24249 ( .A(n24073), .B(n23089), .Y(mult_x_1196_n2902)
         );
  BUFx5_ASAP7_75t_SL U24250 ( .A(mult_x_1196_n596), .Y(n18580) );
  OAI22x1_ASAP7_75t_SL U24251 ( .A1(mult_x_1196_n2973), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2972), .Y(mult_x_1196_n2401) );
  INVx2_ASAP7_75t_SL U24252 ( .A(mult_x_1196_n2401), .Y(n18650) );
  MAJIxp5_ASAP7_75t_SL U24253 ( .A(n24228), .B(n23330), .C(mult_x_1196_n2268), 
        .Y(n23350) );
  NAND2xp5_ASAP7_75t_SL U24254 ( .A(n24264), .B(n22286), .Y(n24228) );
  XNOR2x1_ASAP7_75t_SL U24255 ( .A(n22447), .B(mult_x_1196_n2295), .Y(n22588)
         );
  NOR2x1p5_ASAP7_75t_SL U24256 ( .A(n18780), .B(n18779), .Y(n18644) );
  OAI21xp5_ASAP7_75t_SL U24257 ( .A1(n18582), .A2(n18581), .B(n21919), .Y(
        n4195) );
  INVx1_ASAP7_75t_SL U24258 ( .A(n21918), .Y(n18582) );
  XNOR2xp5_ASAP7_75t_SL U24259 ( .A(n18584), .B(n18583), .Y(n23735) );
  OAI21xp5_ASAP7_75t_SL U24260 ( .A1(n23737), .A2(n22258), .B(n23736), .Y(
        n18583) );
  INVx1_ASAP7_75t_SL U24261 ( .A(mult_x_1196_n226), .Y(n18584) );
  NAND2x1_ASAP7_75t_SL U24262 ( .A(n23328), .B(n18644), .Y(n18643) );
  NAND2x1_ASAP7_75t_SL U24263 ( .A(n22848), .B(n22847), .Y(mult_x_1196_n1135)
         );
  MAJIxp5_ASAP7_75t_SL U24264 ( .A(n18585), .B(mult_x_1196_n2181), .C(
        mult_x_1196_n901), .Y(mult_x_1196_n896) );
  INVx1_ASAP7_75t_SL U24265 ( .A(n18587), .Y(n18585) );
  XNOR2xp5_ASAP7_75t_SL U24266 ( .A(n18587), .B(n18586), .Y(mult_x_1196_n897)
         );
  XNOR2xp5_ASAP7_75t_SL U24267 ( .A(mult_x_1196_n2181), .B(mult_x_1196_n901), 
        .Y(n18586) );
  MAJIxp5_ASAP7_75t_SL U24268 ( .A(mult_x_1196_n2182), .B(mult_x_1196_n929), 
        .C(n22682), .Y(n18587) );
  BUFx5_ASAP7_75t_SL U24269 ( .A(n18394), .Y(n18588) );
  NOR2x1_ASAP7_75t_SL U24270 ( .A(n24035), .B(n18589), .Y(n23494) );
  XNOR2xp5_ASAP7_75t_SL U24271 ( .A(n22395), .B(n22227), .Y(n18589) );
  INVx3_ASAP7_75t_SL U24272 ( .A(n24685), .Y(n22434) );
  NAND2x1p5_ASAP7_75t_SL U24273 ( .A(mult_x_1196_n1796), .B(mult_x_1196_n1772), 
        .Y(mult_x_1196_n646) );
  BUFx5_ASAP7_75t_SL U24274 ( .A(mult_x_1196_n1475), .Y(n18590) );
  BUFx2_ASAP7_75t_SL U24275 ( .A(mult_x_1196_n1578), .Y(n22644) );
  NAND2xp5_ASAP7_75t_SL U24276 ( .A(n24688), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__29_), .Y(n25709) );
  NAND2x1_ASAP7_75t_SL U24277 ( .A(n23558), .B(n25709), .Y(
        u0_0_leon3x0_p0_muli[35]) );
  MAJIxp5_ASAP7_75t_SL U24278 ( .A(n18591), .B(mult_x_1196_n2347), .C(
        mult_x_1196_n2443), .Y(mult_x_1196_n1216) );
  NAND2x1_ASAP7_75t_SL U24279 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__21_), .B(
        n22434), .Y(n18592) );
  BUFx5_ASAP7_75t_SL U24280 ( .A(n18388), .Y(n18593) );
  XOR2xp5_ASAP7_75t_SL U24281 ( .A(n18330), .B(n18594), .Y(mult_x_1196_n1112)
         );
  XNOR2xp5_ASAP7_75t_SL U24282 ( .A(n22710), .B(mult_x_1196_n1117), .Y(n18594)
         );
  XOR2xp5_ASAP7_75t_SL U24283 ( .A(mult_x_1196_n2426), .B(n22452), .Y(n22451)
         );
  OAI21xp5_ASAP7_75t_SL U24284 ( .A1(mult_x_1196_n2998), .A2(n24014), .B(
        n18595), .Y(mult_x_1196_n2426) );
  INVx1_ASAP7_75t_SL U24285 ( .A(n18596), .Y(n18595) );
  NOR2x1_ASAP7_75t_SL U24286 ( .A(mult_x_1196_n2997), .B(n24012), .Y(n18596)
         );
  BUFx5_ASAP7_75t_SL U24287 ( .A(n24121), .Y(n18597) );
  NOR2x1_ASAP7_75t_SL U24288 ( .A(n22248), .B(mult_x_1196_n3193), .Y(n22734)
         );
  NOR2x1p5_ASAP7_75t_SL U24289 ( .A(n22734), .B(n22733), .Y(n22732) );
  XNOR2xp5_ASAP7_75t_SL U24290 ( .A(n22314), .B(n22766), .Y(mult_x_1196_n1117)
         );
  XNOR2xp5_ASAP7_75t_SL U24291 ( .A(n18927), .B(n24060), .Y(mult_x_1196_n3263)
         );
  XNOR2x1_ASAP7_75t_SL U24292 ( .A(n23341), .B(n23604), .Y(mult_x_1196_n1766)
         );
  XNOR2x1_ASAP7_75t_SL U24293 ( .A(mult_x_1196_n1365), .B(n18598), .Y(n23344)
         );
  INVx2_ASAP7_75t_SL U24294 ( .A(mult_x_1196_n1367), .Y(n18598) );
  XNOR2x1_ASAP7_75t_SL U24295 ( .A(n18599), .B(n23424), .Y(n23986) );
  INVx2_ASAP7_75t_SL U24296 ( .A(n24551), .Y(n18599) );
  NOR2x2_ASAP7_75t_SL U24297 ( .A(n18601), .B(n18600), .Y(n24551) );
  INVx2_ASAP7_75t_SL U24298 ( .A(n24552), .Y(n18600) );
  OAI22x1_ASAP7_75t_SL U24299 ( .A1(mult_x_1196_n2967), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2966), .Y(mult_x_1196_n2395) );
  OAI22xp5_ASAP7_75t_SL U24300 ( .A1(mult_x_1196_n3001), .A2(n24014), .B1(
        mult_x_1196_n3000), .B2(n24012), .Y(mult_x_1196_n2429) );
  MAJIxp5_ASAP7_75t_SL U24301 ( .A(mult_x_1196_n1239), .B(mult_x_1196_n1202), 
        .C(mult_x_1196_n1212), .Y(mult_x_1196_n1203) );
  XNOR2xp5_ASAP7_75t_SL U24302 ( .A(n18603), .B(mult_x_1196_n1204), .Y(n22474)
         );
  XNOR2xp5_ASAP7_75t_SL U24303 ( .A(mult_x_1196_n1212), .B(n18602), .Y(
        mult_x_1196_n1204) );
  XOR2xp5_ASAP7_75t_SL U24304 ( .A(mult_x_1196_n1239), .B(mult_x_1196_n1202), 
        .Y(n18602) );
  INVx1_ASAP7_75t_SL U24305 ( .A(mult_x_1196_n1196), .Y(n18603) );
  HB1xp67_ASAP7_75t_SL U24306 ( .A(n24692), .Y(n18604) );
  INVx2_ASAP7_75t_SL U24307 ( .A(mult_x_1196_n2606), .Y(n23749) );
  MAJIxp5_ASAP7_75t_SL U24308 ( .A(mult_x_1196_n1501), .B(mult_x_1196_n1497), 
        .C(mult_x_1196_n1493), .Y(mult_x_1196_n1483) );
  INVx2_ASAP7_75t_SL U24309 ( .A(n22411), .Y(n18605) );
  XNOR2x1_ASAP7_75t_SL U24310 ( .A(mult_x_1196_n1173), .B(n22849), .Y(
        mult_x_1196_n1168) );
  XNOR2x1_ASAP7_75t_SL U24311 ( .A(mult_x_1196_n1669), .B(n24156), .Y(n18950)
         );
  OAI22x1_ASAP7_75t_SL U24312 ( .A1(mult_x_1196_n2865), .A2(n23449), .B1(
        n24030), .B2(mult_x_1196_n2864), .Y(mult_x_1196_n2299) );
  BUFx5_ASAP7_75t_SL U24313 ( .A(n22897), .Y(n18606) );
  NAND3xp33_ASAP7_75t_SL U24314 ( .A(n18607), .B(n23214), .C(n22368), .Y(n4193) );
  NAND2xp5_ASAP7_75t_SL U24315 ( .A(n23209), .B(n23208), .Y(n18607) );
  XNOR2x1_ASAP7_75t_SL U24316 ( .A(n22211), .B(mult_x_1196_n1913), .Y(n18732)
         );
  NAND2x1_ASAP7_75t_SL U24317 ( .A(n22764), .B(n23024), .Y(mult_x_1196_n1913)
         );
  OAI22x1_ASAP7_75t_SL U24318 ( .A1(mult_x_1196_n3261), .A2(n23982), .B1(
        n22389), .B2(mult_x_1196_n3260), .Y(n23112) );
  XNOR2x1_ASAP7_75t_SL U24319 ( .A(n18927), .B(n24058), .Y(mult_x_1196_n3261)
         );
  OAI22x1_ASAP7_75t_SL U24320 ( .A1(n24000), .A2(mult_x_1196_n3132), .B1(
        mult_x_1196_n3131), .B2(n23996), .Y(n23095) );
  OAI21x1_ASAP7_75t_SL U24321 ( .A1(mult_x_1196_n357), .A2(n22533), .B(
        mult_x_1196_n358), .Y(mult_x_1196_n356) );
  OAI22x1_ASAP7_75t_SL U24322 ( .A1(n24003), .A2(mult_x_1196_n3085), .B1(
        n18919), .B2(mult_x_1196_n3086), .Y(n24211) );
  NOR2x1p5_ASAP7_75t_SL U24323 ( .A(n23462), .B(n23463), .Y(n23461) );
  MAJIxp5_ASAP7_75t_SL U24324 ( .A(mult_x_1196_n2576), .B(n24212), .C(
        mult_x_1196_n2298), .Y(n23458) );
  INVx1_ASAP7_75t_SL U24325 ( .A(n18609), .Y(n18608) );
  NOR2x1_ASAP7_75t_SL U24326 ( .A(n24030), .B(mult_x_1196_n2863), .Y(n18609)
         );
  XNOR2xp5_ASAP7_75t_SL U24327 ( .A(n24067), .B(n23091), .Y(mult_x_1196_n3100)
         );
  XOR2xp5_ASAP7_75t_SL U24328 ( .A(n23851), .B(n22774), .Y(n23016) );
  INVx13_ASAP7_75t_SL U24329 ( .A(n23935), .Y(n24231) );
  XNOR2xp5_ASAP7_75t_SL U24330 ( .A(n24069), .B(n23089), .Y(mult_x_1196_n2898)
         );
  BUFx5_ASAP7_75t_SL U24331 ( .A(add_x_735_A_15_), .Y(n18610) );
  OAI22x1_ASAP7_75t_SL U24332 ( .A1(mult_x_1196_n3093), .A2(n23100), .B1(
        mult_x_1196_n3092), .B2(n18435), .Y(n23518) );
  NOR2x1_ASAP7_75t_SL U24333 ( .A(n23984), .B(mult_x_1196_n3231), .Y(n18611)
         );
  MAJIxp5_ASAP7_75t_SL U24334 ( .A(n24294), .B(mult_x_1196_n1004), .C(n18613), 
        .Y(mult_x_1196_n997) );
  INVx1_ASAP7_75t_SL U24335 ( .A(mult_x_1196_n1004), .Y(n18612) );
  NAND2x1p5_ASAP7_75t_SL U24336 ( .A(n24086), .B(mult_x_1196_n810), .Y(
        mult_x_1196_n616) );
  INVx1_ASAP7_75t_SL U24337 ( .A(mult_x_1196_n1314), .Y(n23794) );
  MAJIxp5_ASAP7_75t_SL U24338 ( .A(mult_x_1196_n2350), .B(mult_x_1196_n2167), 
        .C(n18962), .Y(mult_x_1196_n1314) );
  XNOR2xp5_ASAP7_75t_SL U24339 ( .A(n22870), .B(mult_x_1196_n1789), .Y(n22869)
         );
  XNOR2xp5_ASAP7_75t_SL U24340 ( .A(n22824), .B(n23560), .Y(mult_x_1196_n1789)
         );
  BUFx5_ASAP7_75t_SL U24341 ( .A(n22933), .Y(n18614) );
  INVx4_ASAP7_75t_SL U24342 ( .A(n24685), .Y(n23903) );
  NAND2x1_ASAP7_75t_SL U24343 ( .A(n23484), .B(n23486), .Y(mult_x_1196_n1744)
         );
  BUFx6f_ASAP7_75t_SL U24344 ( .A(n23639), .Y(n22448) );
  BUFx10_ASAP7_75t_SL U24345 ( .A(n24049), .Y(n18615) );
  BUFx5_ASAP7_75t_SL U24346 ( .A(mult_x_1196_n1167), .Y(n18616) );
  MAJIxp5_ASAP7_75t_SL U24347 ( .A(mult_x_1196_n2439), .B(mult_x_1196_n2407), 
        .C(mult_x_1196_n2375), .Y(mult_x_1196_n1099) );
  OAI22xp5_ASAP7_75t_SL U24348 ( .A1(mult_x_1196_n2947), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2946), .Y(mult_x_1196_n2375) );
  INVx1_ASAP7_75t_SL U24349 ( .A(mult_x_1196_n228), .Y(n18617) );
  OAI22x1_ASAP7_75t_SL U24350 ( .A1(n18919), .A2(mult_x_1196_n3082), .B1(
        mult_x_1196_n3081), .B2(n24003), .Y(mult_x_1196_n1322) );
  NAND2x1_ASAP7_75t_SL U24351 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__8_), .B(n18862), .Y(n25098) );
  XNOR2x1_ASAP7_75t_SL U24352 ( .A(n18618), .B(n24085), .Y(n24188) );
  MAJIxp5_ASAP7_75t_SL U24353 ( .A(n18618), .B(n18925), .C(mult_x_1196_n1719), 
        .Y(n18619) );
  XOR2x2_ASAP7_75t_SL U24354 ( .A(n24308), .B(n22803), .Y(n18618) );
  INVx1_ASAP7_75t_SL U24355 ( .A(n18619), .Y(n24270) );
  XNOR2xp5_ASAP7_75t_SL U24356 ( .A(n18952), .B(n18620), .Y(n23026) );
  XOR2xp5_ASAP7_75t_SL U24357 ( .A(mult_x_1196_n1924), .B(mult_x_1196_n1943), 
        .Y(n18620) );
  OAI22xp33_ASAP7_75t_SL U24358 ( .A1(mult_x_1196_n3135), .A2(n23999), .B1(
        n23996), .B2(mult_x_1196_n3134), .Y(mult_x_1196_n2559) );
  XOR2xp5_ASAP7_75t_SL U24359 ( .A(n23853), .B(mult_x_1196_n2498), .Y(n18621)
         );
  NOR2x1_ASAP7_75t_SL U24360 ( .A(n24031), .B(n18622), .Y(n23462) );
  OAI22x1_ASAP7_75t_SL U24361 ( .A1(n24007), .A2(mult_x_1196_n3067), .B1(
        n24005), .B2(mult_x_1196_n3066), .Y(mult_x_1196_n2495) );
  XOR2x1_ASAP7_75t_SL U24362 ( .A(mult_x_1196_n1860), .B(mult_x_1196_n1864), 
        .Y(n18651) );
  XNOR2x2_ASAP7_75t_SL U24363 ( .A(n18624), .B(n18623), .Y(mult_x_1196_n1864)
         );
  XNOR2xp5_ASAP7_75t_SL U24364 ( .A(mult_x_1196_n2651), .B(mult_x_1196_n2495), 
        .Y(n18623) );
  OAI22xp5_ASAP7_75t_SL U24365 ( .A1(mult_x_1196_n3226), .A2(n23984), .B1(
        mult_x_1196_n3227), .B2(n24121), .Y(mult_x_1196_n2651) );
  INVxp67_ASAP7_75t_SL U24366 ( .A(mult_x_1196_n2619), .Y(n18624) );
  OAI22xp33_ASAP7_75t_SL U24367 ( .A1(mult_x_1196_n3195), .A2(n23989), .B1(
        mult_x_1196_n3194), .B2(n23987), .Y(mult_x_1196_n2619) );
  XNOR2x1_ASAP7_75t_SL U24368 ( .A(n23129), .B(n18625), .Y(mult_x_1196_n1860)
         );
  XNOR2x1_ASAP7_75t_SL U24369 ( .A(mult_x_1196_n2399), .B(mult_x_1196_n2367), 
        .Y(n18625) );
  OAI22x1_ASAP7_75t_SL U24370 ( .A1(n23141), .A2(mult_x_1196_n2971), .B1(
        mult_x_1196_n2970), .B2(n24017), .Y(mult_x_1196_n2399) );
  NOR2xp67_ASAP7_75t_SL U24371 ( .A(n23131), .B(n23130), .Y(n23129) );
  XOR2xp5_ASAP7_75t_SL U24372 ( .A(mult_x_1196_n1490), .B(mult_x_1196_n1441), 
        .Y(n23336) );
  XNOR2xp5_ASAP7_75t_SL U24373 ( .A(n18627), .B(n18626), .Y(mult_x_1196_n1441)
         );
  INVx1_ASAP7_75t_SL U24374 ( .A(mult_x_1196_n2638), .Y(n18627) );
  OAI22xp5_ASAP7_75t_SL U24375 ( .A1(mult_x_1196_n3214), .A2(n24082), .B1(
        n22538), .B2(mult_x_1196_n3213), .Y(mult_x_1196_n2638) );
  XNOR2xp5_ASAP7_75t_SL U24376 ( .A(n24084), .B(n23800), .Y(n23799) );
  INVx2_ASAP7_75t_SL U24377 ( .A(n18629), .Y(n18628) );
  NOR2x1_ASAP7_75t_SL U24378 ( .A(mult_x_1196_n3060), .B(n24007), .Y(n18629)
         );
  MAJIxp5_ASAP7_75t_SL U24379 ( .A(n18630), .B(mult_x_1196_n1669), .C(
        mult_x_1196_n1677), .Y(n23809) );
  INVx1_ASAP7_75t_SL U24380 ( .A(n24156), .Y(n18630) );
  INVx1_ASAP7_75t_SL U24381 ( .A(n23809), .Y(n22477) );
  MAJx2_ASAP7_75t_SL U24382 ( .A(n23332), .B(n23931), .C(mult_x_1196_n2302), 
        .Y(n24156) );
  MAJIxp5_ASAP7_75t_SL U24383 ( .A(n23434), .B(mult_x_1196_n2392), .C(
        mult_x_1196_n2360), .Y(mult_x_1196_n1669) );
  OAI22xp5_ASAP7_75t_SL U24384 ( .A1(mult_x_1196_n2932), .A2(n24022), .B1(
        mult_x_1196_n2931), .B2(n24020), .Y(mult_x_1196_n2360) );
  MAJIxp5_ASAP7_75t_SL U24385 ( .A(mult_x_1196_n2516), .B(n23117), .C(
        mult_x_1196_n1711), .Y(mult_x_1196_n1677) );
  NOR2x1_ASAP7_75t_SL U24386 ( .A(n18632), .B(n18631), .Y(mult_x_1196_n1711)
         );
  INVx1_ASAP7_75t_SL U24387 ( .A(n23518), .Y(n18631) );
  INVx1_ASAP7_75t_SL U24388 ( .A(mult_x_1196_n2677), .Y(n18632) );
  MAJIxp5_ASAP7_75t_SL U24389 ( .A(n22782), .B(mult_x_1196_n1662), .C(n24301), 
        .Y(n18633) );
  MAJIxp5_ASAP7_75t_SL U24390 ( .A(n18633), .B(n22336), .C(n23583), .Y(
        mult_x_1196_n1583) );
  XNOR2xp5_ASAP7_75t_SL U24391 ( .A(n23250), .B(n18376), .Y(n23093) );
  INVx2_ASAP7_75t_SL U24392 ( .A(mult_x_1196_n1946), .Y(n23807) );
  XNOR2xp5_ASAP7_75t_SL U24393 ( .A(n23646), .B(n18634), .Y(mult_x_1196_n1946)
         );
  XOR2xp5_ASAP7_75t_SL U24394 ( .A(mult_x_1196_n2655), .B(mult_x_1196_n2623), 
        .Y(n18634) );
  OAI22x1_ASAP7_75t_SL U24395 ( .A1(mult_x_1196_n3199), .A2(n23072), .B1(
        mult_x_1196_n3198), .B2(n23987), .Y(mult_x_1196_n2623) );
  OAI22xp5_ASAP7_75t_SL U24396 ( .A1(mult_x_1196_n3167), .A2(n24230), .B1(
        n23992), .B2(mult_x_1196_n3166), .Y(n23646) );
  OAI22xp5_ASAP7_75t_SL U24397 ( .A1(n24040), .A2(mult_x_1196_n2770), .B1(
        n24041), .B2(n23974), .Y(mult_x_1196_n2128) );
  OAI22xp5_ASAP7_75t_SL U24398 ( .A1(n24017), .A2(mult_x_1196_n2960), .B1(
        n23142), .B2(mult_x_1196_n2961), .Y(mult_x_1196_n2389) );
  MAJIxp5_ASAP7_75t_SL U24399 ( .A(mult_x_1196_n2235), .B(mult_x_1196_n2545), 
        .C(mult_x_1196_n2389), .Y(mult_x_1196_n1567) );
  MAJIxp5_ASAP7_75t_SL U24400 ( .A(mult_x_1196_n2128), .B(mult_x_1196_n2357), 
        .C(mult_x_1196_n2453), .Y(mult_x_1196_n1565) );
  OAI22xp5_ASAP7_75t_SL U24401 ( .A1(mult_x_1196_n3025), .A2(n24009), .B1(
        n23442), .B2(mult_x_1196_n3024), .Y(mult_x_1196_n2453) );
  OAI22xp5_ASAP7_75t_SL U24402 ( .A1(mult_x_1196_n2929), .A2(n24021), .B1(
        n24020), .B2(mult_x_1196_n2928), .Y(mult_x_1196_n2357) );
  XNOR2x1_ASAP7_75t_SL U24403 ( .A(n18635), .B(n22754), .Y(mult_x_1196_n1527)
         );
  XNOR2xp5_ASAP7_75t_SL U24404 ( .A(mult_x_1196_n1567), .B(mult_x_1196_n1565), 
        .Y(n18635) );
  OAI22xp5_ASAP7_75t_SL U24405 ( .A1(mult_x_1196_n3121), .A2(n23999), .B1(
        n23996), .B2(mult_x_1196_n3120), .Y(mult_x_1196_n2545) );
  OAI22xp5_ASAP7_75t_SL U24406 ( .A1(mult_x_1196_n2801), .A2(n24038), .B1(
        mult_x_1196_n2800), .B2(n22391), .Y(mult_x_1196_n2235) );
  MAJx3_ASAP7_75t_SL U24407 ( .A(mult_x_1196_n1703), .B(mult_x_1196_n1705), 
        .C(mult_x_1196_n1676), .Y(n22344) );
  XNOR2xp5_ASAP7_75t_SL U24408 ( .A(mult_x_1196_n2644), .B(n18636), .Y(
        mult_x_1196_n1676) );
  XNOR2x1_ASAP7_75t_SL U24409 ( .A(mult_x_1196_n2328), .B(n22665), .Y(n18636)
         );
  OAI22x1_ASAP7_75t_SL U24410 ( .A1(mult_x_1196_n2900), .A2(n24026), .B1(
        mult_x_1196_n2899), .B2(n24025), .Y(mult_x_1196_n2328) );
  OAI21x1_ASAP7_75t_SL U24411 ( .A1(n24014), .A2(mult_x_1196_n3006), .B(n22304), .Y(n23853) );
  XNOR2x1_ASAP7_75t_SL U24412 ( .A(n18637), .B(mult_x_1196_n1927), .Y(
        mult_x_1196_n1900) );
  XNOR2xp5_ASAP7_75t_SL U24413 ( .A(n18638), .B(n23857), .Y(n18637) );
  MAJIxp5_ASAP7_75t_SL U24414 ( .A(mult_x_1196_n2498), .B(n23853), .C(n23566), 
        .Y(n23857) );
  OAI22xp5_ASAP7_75t_SL U24415 ( .A1(mult_x_1196_n3166), .A2(n23994), .B1(
        n23992), .B2(mult_x_1196_n3165), .Y(n23566) );
  OAI22xp5_ASAP7_75t_SL U24416 ( .A1(mult_x_1196_n3070), .A2(n23637), .B1(
        n24005), .B2(mult_x_1196_n3069), .Y(mult_x_1196_n2498) );
  INVx1_ASAP7_75t_SL U24417 ( .A(n24293), .Y(n18638) );
  XNOR2xp5_ASAP7_75t_SL U24418 ( .A(n23112), .B(n18657), .Y(n24293) );
  OAI211xp5_ASAP7_75t_SL U24419 ( .A1(n18644), .A2(n18787), .B(n18643), .C(
        n18639), .Y(n4203) );
  O2A1O1Ixp5_ASAP7_75t_SL U24420 ( .A1(n23225), .A2(n23226), .B(n18640), .C(
        n23327), .Y(n18639) );
  NOR2x1_ASAP7_75t_SL U24421 ( .A(n18642), .B(n18641), .Y(n18640) );
  INVx1_ASAP7_75t_SL U24422 ( .A(n22366), .Y(n18641) );
  NAND2xp5_ASAP7_75t_SL U24423 ( .A(n22421), .B(n18576), .Y(n18642) );
  XOR2xp5_ASAP7_75t_SL U24424 ( .A(mult_x_1196_n1904), .B(n23502), .Y(n18646)
         );
  XNOR2xp5_ASAP7_75t_SL U24425 ( .A(n23169), .B(n18645), .Y(mult_x_1196_n1904)
         );
  XOR2xp5_ASAP7_75t_SL U24426 ( .A(mult_x_1196_n2589), .B(mult_x_1196_n2433), 
        .Y(n18645) );
  XNOR2xp5_ASAP7_75t_SL U24427 ( .A(n18647), .B(n18646), .Y(n23027) );
  INVx1_ASAP7_75t_SL U24428 ( .A(mult_x_1196_n1906), .Y(n18647) );
  XNOR2xp5_ASAP7_75t_SL U24429 ( .A(n18649), .B(n18648), .Y(mult_x_1196_n1906)
         );
  XOR2x2_ASAP7_75t_SL U24430 ( .A(n18650), .B(n22814), .Y(n18648) );
  INVx2_ASAP7_75t_SL U24431 ( .A(mult_x_1196_n2653), .Y(n18649) );
  MAJIxp5_ASAP7_75t_SL U24432 ( .A(n22623), .B(n22620), .C(mult_x_1196_n1876), 
        .Y(mult_x_1196_n1846) );
  XNOR2xp5_ASAP7_75t_SL U24433 ( .A(n18651), .B(n23542), .Y(n22623) );
  AO21x1_ASAP7_75t_SL U24434 ( .A1(n22811), .A2(mult_x_1196_n1899), .B(n22812), 
        .Y(mult_x_1196_n1876) );
  MAJIxp5_ASAP7_75t_SL U24435 ( .A(n18998), .B(n24293), .C(mult_x_1196_n1927), 
        .Y(mult_x_1196_n1899) );
  XNOR2x1_ASAP7_75t_SL U24436 ( .A(mult_x_1196_n2650), .B(n22731), .Y(
        mult_x_1196_n1840) );
  MAJIxp5_ASAP7_75t_SL U24437 ( .A(n23366), .B(mult_x_1196_n2684), .C(n22244), 
        .Y(n23321) );
  NAND2x1_ASAP7_75t_SL U24438 ( .A(n22296), .B(n24236), .Y(n23049) );
  MAJIxp5_ASAP7_75t_SL U24439 ( .A(mult_x_1196_n1828), .B(mult_x_1196_n1809), 
        .C(mult_x_1196_n1830), .Y(mult_x_1196_n1801) );
  MAJIxp5_ASAP7_75t_SL U24440 ( .A(mult_x_1196_n1838), .B(mult_x_1196_n1840), 
        .C(mult_x_1196_n1859), .Y(mult_x_1196_n1830) );
  MAJIxp5_ASAP7_75t_SL U24441 ( .A(n23128), .B(mult_x_1196_n2399), .C(
        mult_x_1196_n2367), .Y(mult_x_1196_n1859) );
  XOR2xp5_ASAP7_75t_SL U24442 ( .A(n22450), .B(n23464), .Y(mult_x_1196_n1838)
         );
  MAJIxp5_ASAP7_75t_SL U24443 ( .A(n24268), .B(mult_x_1196_n1836), .C(n24306), 
        .Y(mult_x_1196_n1828) );
  XNOR2xp5_ASAP7_75t_SL U24444 ( .A(n24233), .B(n24234), .Y(n24306) );
  MAJIxp5_ASAP7_75t_SL U24445 ( .A(n23760), .B(mult_x_1196_n2588), .C(
        mult_x_1196_n2400), .Y(mult_x_1196_n1882) );
  MAJIxp5_ASAP7_75t_SL U24446 ( .A(mult_x_1196_n2496), .B(n24100), .C(n23095), 
        .Y(n23127) );
  XOR2xp5_ASAP7_75t_SL U24447 ( .A(n18653), .B(n18652), .Y(mult_x_1196_n1612)
         );
  XNOR2xp5_ASAP7_75t_SL U24448 ( .A(mult_x_1196_n2674), .B(mult_x_1196_n2514), 
        .Y(n18652) );
  OAI22xp5_ASAP7_75t_SL U24449 ( .A1(n22389), .A2(mult_x_1196_n3249), .B1(
        mult_x_1196_n3250), .B2(n23981), .Y(mult_x_1196_n2674) );
  INVx1_ASAP7_75t_SL U24450 ( .A(n24189), .Y(n18653) );
  BUFx6f_ASAP7_75t_SL U24451 ( .A(n18919), .Y(n18654) );
  OAI21xp5_ASAP7_75t_SL U24452 ( .A1(mult_x_1196_n3090), .A2(n18654), .B(
        n18655), .Y(mult_x_1196_n2514) );
  NAND2xp5_ASAP7_75t_SL U24453 ( .A(n23099), .B(n24246), .Y(n18655) );
  NAND2xp5_ASAP7_75t_SL U24454 ( .A(n18656), .B(n18712), .Y(n23296) );
  OAI21xp33_ASAP7_75t_SL U24455 ( .A1(n18712), .A2(n18656), .B(n23295), .Y(
        n23294) );
  NOR2x1p5_ASAP7_75t_SL U24456 ( .A(n23791), .B(n23790), .Y(n18656) );
  OAI22x1_ASAP7_75t_SL U24457 ( .A1(n24002), .A2(mult_x_1196_n3100), .B1(
        n18920), .B2(mult_x_1196_n3101), .Y(n18657) );
  INVx1_ASAP7_75t_SL U24458 ( .A(n18658), .Y(mult_x_1196_n3110) );
  NOR2x1_ASAP7_75t_SL U24459 ( .A(n18662), .B(n22227), .Y(n18658) );
  XNOR2xp5_ASAP7_75t_SL U24460 ( .A(n22394), .B(n24057), .Y(mult_x_1196_n3090)
         );
  XNOR2x1_ASAP7_75t_SL U24461 ( .A(n22394), .B(n24058), .Y(mult_x_1196_n3091)
         );
  NOR2x1_ASAP7_75t_SL U24462 ( .A(n18662), .B(n18920), .Y(n22696) );
  NAND2xp5_ASAP7_75t_SL U24463 ( .A(n22394), .B(n18659), .Y(n28683) );
  NAND2xp5_ASAP7_75t_SL U24464 ( .A(n28830), .B(u0_0_leon3x0_p0_divi[10]), .Y(
        n18659) );
  NAND2xp5_ASAP7_75t_SL U24465 ( .A(n18660), .B(n19792), .Y(n28668) );
  NAND2xp5_ASAP7_75t_SL U24466 ( .A(n22394), .B(n18661), .Y(n18660) );
  A2O1A1Ixp33_ASAP7_75t_SL U24467 ( .A1(n28827), .A2(u0_0_leon3x0_p0_divi[10]), 
        .B(n28678), .C(n18662), .Y(n28682) );
  INVx1_ASAP7_75t_SL U24468 ( .A(n22394), .Y(n18662) );
  XNOR2xp5_ASAP7_75t_SL U24469 ( .A(n18663), .B(mult_x_1196_n2430), .Y(n23464)
         );
  MAJIxp5_ASAP7_75t_SL U24470 ( .A(n23465), .B(mult_x_1196_n2430), .C(n18663), 
        .Y(mult_x_1196_n1837) );
  XNOR2x1_ASAP7_75t_SL U24471 ( .A(mult_x_1196_n1636), .B(n22985), .Y(n22840)
         );
  XNOR2x1_ASAP7_75t_SL U24472 ( .A(n24228), .B(n24229), .Y(n22985) );
  OAI22xp5_ASAP7_75t_SL U24473 ( .A1(mult_x_1196_n3097), .A2(n18920), .B1(
        n24002), .B2(n18664), .Y(mult_x_1196_n2521) );
  OAI21xp5_ASAP7_75t_SL U24474 ( .A1(n18654), .A2(n18664), .B(n23097), .Y(
        mult_x_1196_n2520) );
  XNOR2xp5_ASAP7_75t_SL U24475 ( .A(n22394), .B(n24063), .Y(n18664) );
  NAND2xp5_ASAP7_75t_SL U24476 ( .A(n18666), .B(n18665), .Y(mult_x_1196_n1463)
         );
  INVx1_ASAP7_75t_SL U24477 ( .A(n18668), .Y(n18665) );
  NAND2xp5_ASAP7_75t_SL U24478 ( .A(n18669), .B(n18667), .Y(n18666) );
  OAI21xp5_ASAP7_75t_SL U24479 ( .A1(n18669), .A2(n18668), .B(n18667), .Y(
        n18672) );
  NAND2xp5_ASAP7_75t_SL U24480 ( .A(n23185), .B(mult_x_1196_n2638), .Y(n18667)
         );
  NOR2xp67_ASAP7_75t_SL U24481 ( .A(n23185), .B(mult_x_1196_n2638), .Y(n18668)
         );
  INVx1_ASAP7_75t_SL U24482 ( .A(mult_x_1196_n2264), .Y(n18669) );
  MAJx2_ASAP7_75t_SL U24483 ( .A(mult_x_1196_n1411), .B(n22308), .C(n18670), 
        .Y(mult_x_1196_n1371) );
  INVx1_ASAP7_75t_SL U24484 ( .A(mult_x_1196_n1378), .Y(n18670) );
  NAND2xp5_ASAP7_75t_SL U24485 ( .A(n18673), .B(n18671), .Y(mult_x_1196_n1411)
         );
  OAI21xp5_ASAP7_75t_SL U24486 ( .A1(n18674), .A2(n23748), .B(n18672), .Y(
        n18671) );
  NAND2xp5_ASAP7_75t_SL U24487 ( .A(n23748), .B(n18674), .Y(n18673) );
  INVx1_ASAP7_75t_SL U24488 ( .A(mult_x_1196_n1454), .Y(n18674) );
  MAJIxp5_ASAP7_75t_SL U24489 ( .A(mult_x_1196_n2354), .B(mult_x_1196_n2171), 
        .C(mult_x_1196_n2386), .Y(mult_x_1196_n1454) );
  XNOR2xp5_ASAP7_75t_SL U24490 ( .A(mult_x_1196_n2540), .B(n23476), .Y(
        mult_x_1196_n1378) );
  MAJIxp5_ASAP7_75t_SL U24491 ( .A(mult_x_1196_n1738), .B(mult_x_1196_n1765), 
        .C(n18675), .Y(n24226) );
  XOR2xp5_ASAP7_75t_SL U24492 ( .A(n18570), .B(n22778), .Y(n18675) );
  NOR2x1_ASAP7_75t_SL U24493 ( .A(n18676), .B(n24035), .Y(n23312) );
  XNOR2xp5_ASAP7_75t_SL U24494 ( .A(mult_x_1196_n1718), .B(mult_x_1196_n1689), 
        .Y(n18770) );
  XNOR2xp5_ASAP7_75t_SL U24495 ( .A(n23238), .B(n18677), .Y(mult_x_1196_n1689)
         );
  XOR2xp5_ASAP7_75t_SL U24496 ( .A(mult_x_1196_n1699), .B(mult_x_1196_n1697), 
        .Y(n18677) );
  XOR2xp5_ASAP7_75t_SL U24497 ( .A(n18678), .B(n23689), .Y(mult_x_1196_n1699)
         );
  INVx1_ASAP7_75t_SL U24498 ( .A(n23691), .Y(n18678) );
  MAJIxp5_ASAP7_75t_SL U24499 ( .A(mult_x_1196_n1749), .B(n22213), .C(n22750), 
        .Y(mult_x_1196_n1718) );
  XNOR2xp5_ASAP7_75t_SL U24500 ( .A(mult_x_1196_n1756), .B(n18679), .Y(n22750)
         );
  XNOR2xp5_ASAP7_75t_SL U24501 ( .A(n23512), .B(mult_x_1196_n1754), .Y(n18679)
         );
  XNOR2xp5_ASAP7_75t_SL U24502 ( .A(n18681), .B(n18680), .Y(n22213) );
  XOR2xp5_ASAP7_75t_SL U24503 ( .A(mult_x_1196_n1734), .B(mult_x_1196_n1736), 
        .Y(n18680) );
  INVx1_ASAP7_75t_SL U24504 ( .A(n23105), .Y(n18681) );
  MAJIxp5_ASAP7_75t_SL U24505 ( .A(mult_x_1196_n1755), .B(mult_x_1196_n1781), 
        .C(mult_x_1196_n1757), .Y(mult_x_1196_n1749) );
  XNOR2xp5_ASAP7_75t_SL U24506 ( .A(n23017), .B(n23018), .Y(mult_x_1196_n1757)
         );
  XNOR2xp5_ASAP7_75t_SL U24507 ( .A(mult_x_1196_n1762), .B(n22485), .Y(
        mult_x_1196_n1755) );
  XNOR2x1_ASAP7_75t_SL U24508 ( .A(n22966), .B(n22693), .Y(n18682) );
  XOR2xp5_ASAP7_75t_SL U24509 ( .A(n23819), .B(n18682), .Y(mult_x_1196_n1426)
         );
  NAND2xp5_ASAP7_75t_SL U24510 ( .A(n22724), .B(n18682), .Y(n22723) );
  XNOR2x1_ASAP7_75t_SL U24511 ( .A(n18683), .B(n22840), .Y(n23251) );
  INVx2_ASAP7_75t_SL U24512 ( .A(n22841), .Y(n18683) );
  MAJIxp5_ASAP7_75t_SL U24513 ( .A(n23251), .B(n18685), .C(n18684), .Y(n24288)
         );
  INVx1_ASAP7_75t_SL U24514 ( .A(mult_x_1196_n1599), .Y(n18684) );
  INVx1_ASAP7_75t_SL U24515 ( .A(mult_x_1196_n1630), .Y(n18685) );
  MAJIxp5_ASAP7_75t_SL U24516 ( .A(mult_x_1196_n1069), .B(mult_x_1196_n1072), 
        .C(mult_x_1196_n1090), .Y(mult_x_1196_n1063) );
  MAJIxp5_ASAP7_75t_SL U24517 ( .A(mult_x_1196_n1124), .B(mult_x_1196_n1102), 
        .C(mult_x_1196_n1098), .Y(mult_x_1196_n1090) );
  AO21x1_ASAP7_75t_SL U24518 ( .A1(n18687), .A2(mult_x_1196_n1160), .B(n18686), 
        .Y(mult_x_1196_n1124) );
  NOR2x1_ASAP7_75t_SL U24519 ( .A(mult_x_1196_n2161), .B(mult_x_1196_n2440), 
        .Y(n18686) );
  NAND2xp5_ASAP7_75t_SL U24520 ( .A(n18689), .B(n18688), .Y(n18687) );
  INVx1_ASAP7_75t_SL U24521 ( .A(n24119), .Y(n18688) );
  INVx1_ASAP7_75t_SL U24522 ( .A(n24117), .Y(n18689) );
  XNOR2xp5_ASAP7_75t_SL U24523 ( .A(n18692), .B(n18691), .Y(mult_x_1196_n1072)
         );
  XOR2xp5_ASAP7_75t_SL U24524 ( .A(n23478), .B(mult_x_1196_n1101), .Y(n18691)
         );
  INVx1_ASAP7_75t_SL U24525 ( .A(mult_x_1196_n1103), .Y(n18692) );
  MAJIxp5_ASAP7_75t_SL U24526 ( .A(n18701), .B(mult_x_1196_n2253), .C(n23201), 
        .Y(mult_x_1196_n1103) );
  XNOR2xp5_ASAP7_75t_SL U24527 ( .A(n18693), .B(mult_x_1196_n1076), .Y(
        mult_x_1196_n1069) );
  XNOR2xp5_ASAP7_75t_SL U24528 ( .A(n18694), .B(mult_x_1196_n1097), .Y(n18693)
         );
  MAJIxp5_ASAP7_75t_SL U24529 ( .A(mult_x_1196_n2343), .B(mult_x_1196_n2471), 
        .C(n23408), .Y(mult_x_1196_n1097) );
  INVx1_ASAP7_75t_SL U24530 ( .A(mult_x_1196_n1099), .Y(n18694) );
  NAND2xp5_ASAP7_75t_SL U24531 ( .A(n18696), .B(n18695), .Y(n23542) );
  OAI21xp5_ASAP7_75t_SL U24532 ( .A1(mult_x_1196_n1901), .A2(mult_x_1196_n1903), .B(mult_x_1196_n1905), .Y(n18695) );
  MAJIxp5_ASAP7_75t_SL U24533 ( .A(n22814), .B(mult_x_1196_n2401), .C(
        mult_x_1196_n2653), .Y(mult_x_1196_n1905) );
  OAI21xp5_ASAP7_75t_SL U24534 ( .A1(n23984), .A2(mult_x_1196_n3228), .B(
        n24170), .Y(mult_x_1196_n2653) );
  NAND2xp5_ASAP7_75t_SL U24535 ( .A(mult_x_1196_n1903), .B(mult_x_1196_n1901), 
        .Y(n18696) );
  MAJIxp5_ASAP7_75t_SL U24536 ( .A(mult_x_1196_n2134), .B(mult_x_1196_n2465), 
        .C(n23519), .Y(mult_x_1196_n1901) );
  MAJIxp5_ASAP7_75t_SL U24537 ( .A(mult_x_1196_n2589), .B(n23169), .C(
        mult_x_1196_n2433), .Y(mult_x_1196_n1903) );
  NOR2x1_ASAP7_75t_SL U24538 ( .A(n18697), .B(n24008), .Y(n23629) );
  OAI22xp5_ASAP7_75t_SL U24539 ( .A1(n24008), .A2(mult_x_1196_n3039), .B1(
        n18697), .B2(n24009), .Y(mult_x_1196_n2468) );
  XNOR2xp5_ASAP7_75t_SL U24540 ( .A(n18698), .B(n24075), .Y(n18697) );
  INVx1_ASAP7_75t_SL U24541 ( .A(n23963), .Y(n18698) );
  OAI22x1_ASAP7_75t_SL U24542 ( .A1(mult_x_1196_n2767), .A2(n24040), .B1(
        mult_x_1196_n2768), .B2(n24041), .Y(n18699) );
  MAJIxp5_ASAP7_75t_SL U24543 ( .A(n23354), .B(n18699), .C(n23851), .Y(
        mult_x_1196_n1532) );
  XNOR2xp5_ASAP7_75t_SL U24544 ( .A(n18699), .B(n23355), .Y(n22774) );
  INVx1_ASAP7_75t_SL U24545 ( .A(mult_x_1196_n1387), .Y(n23107) );
  MAJIxp5_ASAP7_75t_SL U24546 ( .A(n22916), .B(mult_x_1196_n1420), .C(n22482), 
        .Y(mult_x_1196_n1373) );
  XNOR2xp5_ASAP7_75t_SL U24547 ( .A(n23782), .B(n18700), .Y(n22916) );
  OAI22xp5_ASAP7_75t_SL U24548 ( .A1(n24287), .A2(mult_x_1196_n3148), .B1(
        mult_x_1196_n3147), .B2(n23992), .Y(n23488) );
  XNOR2x2_ASAP7_75t_SL U24549 ( .A(mult_x_1196_n1133), .B(n23201), .Y(n23200)
         );
  INVx1_ASAP7_75t_SL U24550 ( .A(mult_x_1196_n1133), .Y(n18701) );
  NOR2x1p5_ASAP7_75t_SL U24551 ( .A(n22983), .B(n23394), .Y(n18702) );
  XNOR2xp5_ASAP7_75t_SL U24552 ( .A(mult_x_1196_n1591), .B(n18703), .Y(n23753)
         );
  XNOR2xp5_ASAP7_75t_SL U24553 ( .A(n18710), .B(n18704), .Y(mult_x_1196_n1561)
         );
  XNOR2xp5_ASAP7_75t_SL U24554 ( .A(n18711), .B(mult_x_1196_n2578), .Y(
        mult_x_1196_n1606) );
  XNOR2xp5_ASAP7_75t_SL U24555 ( .A(n18705), .B(n18706), .Y(mult_x_1196_n1602)
         );
  XOR2xp5_ASAP7_75t_SL U24556 ( .A(mult_x_1196_n1603), .B(mult_x_1196_n1605), 
        .Y(n18704) );
  AO21x1_ASAP7_75t_SL U24557 ( .A1(n18708), .A2(n18707), .B(n18709), .Y(n23632) );
  XNOR2x1_ASAP7_75t_SL U24558 ( .A(mult_x_1196_n2358), .B(n23633), .Y(n18705)
         );
  OAI21x1_ASAP7_75t_SL U24559 ( .A1(n18709), .A2(n18708), .B(n18707), .Y(
        n18706) );
  NAND2x1_ASAP7_75t_SL U24560 ( .A(mult_x_1196_n2269), .B(mult_x_1196_n2327), 
        .Y(n18707) );
  INVx2_ASAP7_75t_SL U24561 ( .A(n24130), .Y(n18708) );
  NOR2xp67_ASAP7_75t_SL U24562 ( .A(mult_x_1196_n2269), .B(mult_x_1196_n2327), 
        .Y(n18709) );
  INVx1_ASAP7_75t_SL U24563 ( .A(n24105), .Y(n18710) );
  XOR2xp5_ASAP7_75t_SL U24564 ( .A(mult_x_1196_n2422), .B(n22708), .Y(n18711)
         );
  INVx2_ASAP7_75t_SL U24565 ( .A(n18712), .Y(mult_x_1196_n2570) );
  NOR2x1p5_ASAP7_75t_SL U24566 ( .A(n18713), .B(n23430), .Y(n18712) );
  NOR2x1p5_ASAP7_75t_SL U24567 ( .A(n24287), .B(mult_x_1196_n3146), .Y(n18713)
         );
  MAJx2_ASAP7_75t_SL U24568 ( .A(n18714), .B(mult_x_1196_n2419), .C(n24180), 
        .Y(n24300) );
  INVx1_ASAP7_75t_SL U24569 ( .A(n22932), .Y(n18714) );
  NOR2x1_ASAP7_75t_SL U24570 ( .A(n18720), .B(n24040), .Y(n18716) );
  XNOR2x1_ASAP7_75t_SL U24571 ( .A(n18718), .B(n18717), .Y(n22653) );
  XNOR2x1_ASAP7_75t_SL U24572 ( .A(mult_x_1196_n2368), .B(n23244), .Y(n18717)
         );
  OAI22x1_ASAP7_75t_SL U24573 ( .A1(n23989), .A2(mult_x_1196_n3196), .B1(
        n24106), .B2(mult_x_1196_n3195), .Y(n23244) );
  INVx2_ASAP7_75t_SL U24574 ( .A(mult_x_1196_n2652), .Y(n18718) );
  OAI21x1_ASAP7_75t_SL U24575 ( .A1(n23984), .A2(n18450), .B(n18719), .Y(
        mult_x_1196_n2652) );
  NAND3x1_ASAP7_75t_SL U24576 ( .A(n23309), .B(n22791), .C(n22538), .Y(n18719)
         );
  OAI22xp5_ASAP7_75t_SL U24577 ( .A1(mult_x_1196_n2765), .A2(n24040), .B1(
        n24041), .B2(n18720), .Y(n23912) );
  XOR2xp5_ASAP7_75t_SL U24578 ( .A(n23204), .B(n18722), .Y(n22758) );
  XOR2xp5_ASAP7_75t_SL U24579 ( .A(n18941), .B(n18723), .Y(mult_x_1196_n1879)
         );
  XNOR2xp5_ASAP7_75t_SL U24580 ( .A(mult_x_1196_n1903), .B(mult_x_1196_n1905), 
        .Y(n18723) );
  XNOR2x1_ASAP7_75t_SL U24581 ( .A(n24048), .B(n18927), .Y(mult_x_1196_n3251)
         );
  NOR2x2_ASAP7_75t_SL U24582 ( .A(n23832), .B(n18724), .Y(n26917) );
  NOR2x1p5_ASAP7_75t_SL U24583 ( .A(n26916), .B(n23830), .Y(n18724) );
  OAI21x1_ASAP7_75t_SL U24584 ( .A1(n18725), .A2(n22467), .B(mult_x_1196_n460), 
        .Y(n18727) );
  AOI21x1_ASAP7_75t_SL U24585 ( .A1(mult_x_1196_n491), .A2(mult_x_1196_n472), 
        .B(mult_x_1196_n473), .Y(n22467) );
  INVx2_ASAP7_75t_SL U24586 ( .A(n23732), .Y(n18725) );
  OAI21x1_ASAP7_75t_SL U24587 ( .A1(n18350), .A2(n18728), .B(n18726), .Y(
        mult_x_1196_n456) );
  INVx2_ASAP7_75t_SL U24588 ( .A(n18727), .Y(n18726) );
  NAND2x1_ASAP7_75t_SL U24589 ( .A(n23732), .B(n18729), .Y(n18728) );
  INVx2_ASAP7_75t_SL U24590 ( .A(mult_x_1196_n470), .Y(n18729) );
  NOR2x2_ASAP7_75t_SL U24591 ( .A(n23731), .B(n23730), .Y(mult_x_1196_n496) );
  NAND2x1_ASAP7_75t_SL U24592 ( .A(mult_x_1196_n472), .B(mult_x_1196_n793), 
        .Y(mult_x_1196_n470) );
  OAI21x1_ASAP7_75t_SL U24593 ( .A1(mult_x_1196_n470), .A2(mult_x_1196_n496), 
        .B(n22467), .Y(mult_x_1196_n465) );
  NOR2x1_ASAP7_75t_SL U24594 ( .A(mult_x_1196_n578), .B(mult_x_1196_n575), .Y(
        n18730) );
  NAND2xp5_ASAP7_75t_SL U24595 ( .A(n18730), .B(mult_x_1196_n801), .Y(
        mult_x_1196_n560) );
  XNOR2x1_ASAP7_75t_SL U24596 ( .A(n18731), .B(n24220), .Y(mult_x_1196_n1358)
         );
  XOR2x2_ASAP7_75t_SL U24597 ( .A(mult_x_1196_n1394), .B(mult_x_1196_n1363), 
        .Y(n18731) );
  XNOR2x1_ASAP7_75t_SL U24598 ( .A(mult_x_1196_n1934), .B(n22325), .Y(n18734)
         );
  MAJx2_ASAP7_75t_SL U24599 ( .A(n18740), .B(n18739), .C(n18738), .Y(n18737)
         );
  XOR2xp5_ASAP7_75t_SL U24600 ( .A(n23025), .B(n22543), .Y(n18740) );
  MAJIxp5_ASAP7_75t_SL U24601 ( .A(n22324), .B(n18935), .C(n18733), .Y(
        mult_x_1196_n1931) );
  INVx1_ASAP7_75t_SL U24602 ( .A(n23020), .Y(n18733) );
  XNOR2xp5_ASAP7_75t_SL U24603 ( .A(n18734), .B(n18740), .Y(mult_x_1196_n1911)
         );
  INVx1_ASAP7_75t_SL U24604 ( .A(n22979), .Y(n18736) );
  INVx1_ASAP7_75t_SL U24605 ( .A(n22325), .Y(n18738) );
  INVx1_ASAP7_75t_SL U24606 ( .A(mult_x_1196_n1934), .Y(n18739) );
  XNOR2x1_ASAP7_75t_SL U24607 ( .A(n23340), .B(n18741), .Y(n22253) );
  XNOR2x1_ASAP7_75t_SL U24608 ( .A(n18742), .B(n23878), .Y(n18741) );
  INVx2_ASAP7_75t_SL U24609 ( .A(mult_x_1196_n2395), .Y(n18742) );
  XNOR2xp5_ASAP7_75t_SL U24610 ( .A(n18743), .B(mult_x_1196_n1376), .Y(n18746)
         );
  INVx1_ASAP7_75t_SL U24611 ( .A(mult_x_1196_n1409), .Y(n18743) );
  XNOR2x2_ASAP7_75t_SL U24612 ( .A(mult_x_1196_n1369), .B(n18744), .Y(
        mult_x_1196_n1365) );
  XNOR2xp5_ASAP7_75t_SL U24613 ( .A(mult_x_1196_n1404), .B(n18745), .Y(n18744)
         );
  INVx1_ASAP7_75t_SL U24614 ( .A(mult_x_1196_n1407), .Y(n18745) );
  MAJIxp5_ASAP7_75t_SL U24615 ( .A(mult_x_1196_n1452), .B(mult_x_1196_n1419), 
        .C(mult_x_1196_n1415), .Y(mult_x_1196_n1404) );
  XNOR2x2_ASAP7_75t_SL U24616 ( .A(mult_x_1196_n1374), .B(n18746), .Y(
        mult_x_1196_n1367) );
  XNOR2x1_ASAP7_75t_SL U24617 ( .A(n18747), .B(n23920), .Y(n18992) );
  MAJIxp5_ASAP7_75t_SL U24618 ( .A(mult_x_1196_n1395), .B(n18531), .C(n18401), 
        .Y(mult_x_1196_n1391) );
  MAJx2_ASAP7_75t_SL U24619 ( .A(n24095), .B(mult_x_1196_n1440), .C(n24089), 
        .Y(n18747) );
  XNOR2xp5_ASAP7_75t_SL U24620 ( .A(n18748), .B(n22758), .Y(mult_x_1196_n1869)
         );
  XNOR2xp5_ASAP7_75t_SL U24621 ( .A(n22326), .B(mult_x_1196_n1891), .Y(n18748)
         );
  MAJIxp5_ASAP7_75t_SL U24622 ( .A(n23027), .B(mult_x_1196_n1900), .C(
        mult_x_1196_n1916), .Y(mult_x_1196_n1891) );
  XNOR2x1_ASAP7_75t_SL U24623 ( .A(n22867), .B(n22866), .Y(mult_x_1196_n1665)
         );
  XNOR2xp5_ASAP7_75t_SL U24624 ( .A(n18750), .B(mult_x_1196_n1658), .Y(n22546)
         );
  XNOR2xp5_ASAP7_75t_SL U24625 ( .A(mult_x_1196_n1665), .B(n18749), .Y(
        mult_x_1196_n1658) );
  XOR2xp5_ASAP7_75t_SL U24626 ( .A(mult_x_1196_n1696), .B(mult_x_1196_n1668), 
        .Y(n18749) );
  INVx1_ASAP7_75t_SL U24627 ( .A(mult_x_1196_n1691), .Y(n18750) );
  MAJIxp5_ASAP7_75t_SL U24628 ( .A(mult_x_1196_n1727), .B(mult_x_1196_n1690), 
        .C(n18366), .Y(mult_x_1196_n1691) );
  MAJIxp5_ASAP7_75t_SL U24629 ( .A(n23105), .B(mult_x_1196_n1736), .C(
        mult_x_1196_n1734), .Y(mult_x_1196_n1727) );
  XNOR2xp5_ASAP7_75t_SL U24630 ( .A(n22973), .B(n23594), .Y(mult_x_1196_n1734)
         );
  XNOR2xp5_ASAP7_75t_SL U24631 ( .A(mult_x_1196_n2550), .B(n22451), .Y(
        mult_x_1196_n1736) );
  NOR2x1_ASAP7_75t_SL U24632 ( .A(n22323), .B(n23096), .Y(n23105) );
  XOR2xp5_ASAP7_75t_SL U24633 ( .A(n22833), .B(n24141), .Y(mult_x_1196_n1668)
         );
  MAJIxp5_ASAP7_75t_SL U24634 ( .A(n23446), .B(mult_x_1196_n1708), .C(
        mult_x_1196_n1735), .Y(mult_x_1196_n1696) );
  XNOR2xp5_ASAP7_75t_SL U24635 ( .A(mult_x_1196_n1415), .B(n23472), .Y(
        mult_x_1196_n1405) );
  XNOR2xp5_ASAP7_75t_SL U24636 ( .A(n23320), .B(n18987), .Y(n22974) );
  XNOR2xp5_ASAP7_75t_SL U24637 ( .A(n18752), .B(n18751), .Y(n23636) );
  INVx1_ASAP7_75t_SL U24638 ( .A(mult_x_1196_n1364), .Y(n18752) );
  MAJIxp5_ASAP7_75t_SL U24639 ( .A(mult_x_1196_n1369), .B(mult_x_1196_n1404), 
        .C(n22581), .Y(mult_x_1196_n1364) );
  NAND2x2_ASAP7_75t_SL U24640 ( .A(n18753), .B(n23289), .Y(n23288) );
  XNOR2x1_ASAP7_75t_SL U24641 ( .A(n18927), .B(n24055), .Y(n18754) );
  NOR2x1_ASAP7_75t_SL U24642 ( .A(n22389), .B(n18754), .Y(n23115) );
  XNOR2xp5_ASAP7_75t_SL U24643 ( .A(mult_x_1196_n2306), .B(n18755), .Y(n22835)
         );
  MAJIxp5_ASAP7_75t_SL U24644 ( .A(n18755), .B(mult_x_1196_n2306), .C(n22834), 
        .Y(mult_x_1196_n1792) );
  OAI22xp5_ASAP7_75t_SL U24645 ( .A1(n24025), .A2(mult_x_1196_n2903), .B1(
        mult_x_1196_n2904), .B2(n23116), .Y(n18755) );
  XNOR2x2_ASAP7_75t_SL U24646 ( .A(n18757), .B(n22469), .Y(n22471) );
  XNOR2x1_ASAP7_75t_SL U24647 ( .A(mult_x_1196_n2515), .B(n18756), .Y(n22469)
         );
  INVx2_ASAP7_75t_SL U24648 ( .A(mult_x_1196_n2675), .Y(n18756) );
  INVx2_ASAP7_75t_SL U24649 ( .A(mult_x_1196_n2129), .Y(n18757) );
  INVx8_ASAP7_75t_SL U24650 ( .A(n18758), .Y(n24069) );
  INVx13_ASAP7_75t_SL U24651 ( .A(n18759), .Y(n18760) );
  NOR2x1p5_ASAP7_75t_SL U24652 ( .A(n18760), .B(n18761), .Y(
        u0_0_leon3x0_p0_divi[6]) );
  OR2x2_ASAP7_75t_SL U24653 ( .A(n24069), .B(n28769), .Y(n18759) );
  OA22x2_ASAP7_75t_SL U24654 ( .A1(n28767), .A2(n24689), .B1(n23848), .B2(
        n23831), .Y(n18758) );
  INVxp67_ASAP7_75t_SL U24655 ( .A(n28768), .Y(n18761) );
  MAJIxp5_ASAP7_75t_SL U24656 ( .A(n18763), .B(mult_x_1196_n2352), .C(
        mult_x_1196_n2169), .Y(mult_x_1196_n1379) );
  XOR2xp5_ASAP7_75t_SL U24657 ( .A(n18762), .B(mult_x_1196_n2352), .Y(
        mult_x_1196_n1380) );
  XNOR2xp5_ASAP7_75t_SL U24658 ( .A(n18763), .B(mult_x_1196_n2169), .Y(n18762)
         );
  OAI22xp5_ASAP7_75t_SL U24659 ( .A1(mult_x_1196_n2955), .A2(n24016), .B1(
        mult_x_1196_n2956), .B2(n23142), .Y(n18763) );
  MAJIxp5_ASAP7_75t_SL U24660 ( .A(mult_x_1196_n1387), .B(n18764), .C(n18767), 
        .Y(n22925) );
  INVx1_ASAP7_75t_SL U24661 ( .A(n23616), .Y(n18764) );
  NOR2x1_ASAP7_75t_SL U24662 ( .A(n18766), .B(n18765), .Y(n23616) );
  NOR2x1_ASAP7_75t_SL U24663 ( .A(mult_x_1196_n2762), .B(n24040), .Y(n18765)
         );
  NOR2x1_ASAP7_75t_SL U24664 ( .A(n24041), .B(mult_x_1196_n2763), .Y(n18766)
         );
  INVx1_ASAP7_75t_SL U24665 ( .A(n23618), .Y(n18767) );
  NOR2x1_ASAP7_75t_SL U24666 ( .A(n18769), .B(n18768), .Y(n23618) );
  NOR2x1_ASAP7_75t_SL U24667 ( .A(mult_x_1196_n2826), .B(n22251), .Y(n18769)
         );
  XNOR2x1_ASAP7_75t_SL U24668 ( .A(n18770), .B(n23448), .Y(n18918) );
  INVx3_ASAP7_75t_SL U24669 ( .A(n23971), .Y(n18771) );
  XNOR2xp5_ASAP7_75t_SL U24670 ( .A(n18772), .B(mult_x_1196_n2614), .Y(n22564)
         );
  MAJIxp5_ASAP7_75t_SL U24671 ( .A(mult_x_1196_n2614), .B(mult_x_1196_n2490), 
        .C(n18772), .Y(mult_x_1196_n1737) );
  XNOR2xp5_ASAP7_75t_SL U24672 ( .A(n18934), .B(n23054), .Y(mult_x_1196_n1268)
         );
  XNOR2xp5_ASAP7_75t_SL U24673 ( .A(mult_x_1196_n1286), .B(n23703), .Y(n18934)
         );
  XNOR2xp5_ASAP7_75t_SL U24674 ( .A(n18776), .B(n18773), .Y(mult_x_1196_n1425)
         );
  XOR2xp5_ASAP7_75t_SL U24675 ( .A(n24211), .B(n24210), .Y(n18773) );
  NOR2x1_ASAP7_75t_SL U24676 ( .A(n18774), .B(n18775), .Y(n24210) );
  NOR2x1_ASAP7_75t_SL U24677 ( .A(mult_x_1196_n2829), .B(n24035), .Y(n18774)
         );
  NOR2x1_ASAP7_75t_SL U24678 ( .A(mult_x_1196_n2828), .B(n22251), .Y(n18775)
         );
  INVx1_ASAP7_75t_SL U24679 ( .A(n23322), .Y(n18776) );
  NOR2x1p5_ASAP7_75t_SL U24680 ( .A(mult_x_1196_n474), .B(mult_x_1196_n481), 
        .Y(mult_x_1196_n472) );
  NOR2x1_ASAP7_75t_SL U24681 ( .A(mult_x_1196_n1084), .B(mult_x_1196_n1081), 
        .Y(mult_x_1196_n481) );
  NOR2x1_ASAP7_75t_SL U24682 ( .A(mult_x_1196_n1059), .B(mult_x_1196_n1083), 
        .Y(mult_x_1196_n474) );
  INVx2_ASAP7_75t_SL U24683 ( .A(mult_x_1196_n794), .Y(n22894) );
  INVx2_ASAP7_75t_SL U24684 ( .A(mult_x_1196_n1135), .Y(n18777) );
  INVx2_ASAP7_75t_SL U24685 ( .A(mult_x_1196_n1134), .Y(n18778) );
  INVx1_ASAP7_75t_SL U24686 ( .A(n22491), .Y(n23263) );
  INVx2_ASAP7_75t_SL U24687 ( .A(n22584), .Y(n18779) );
  NAND2x1_ASAP7_75t_SL U24688 ( .A(n18781), .B(n22517), .Y(n18780) );
  INVx1_ASAP7_75t_SL U24689 ( .A(n18782), .Y(n18781) );
  NAND2xp5_ASAP7_75t_SL U24690 ( .A(n18399), .B(n18446), .Y(n18782) );
  NOR2x1_ASAP7_75t_SL U24691 ( .A(n22404), .B(n23134), .Y(n23226) );
  OAI21xp5_ASAP7_75t_SL U24692 ( .A1(n18784), .A2(n23134), .B(n18783), .Y(
        n18787) );
  AOI21xp5_ASAP7_75t_SL U24693 ( .A1(n23225), .A2(n18576), .B(n23329), .Y(
        n18783) );
  INVx1_ASAP7_75t_SL U24694 ( .A(n18785), .Y(n18784) );
  NOR2x1_ASAP7_75t_SL U24695 ( .A(n18786), .B(n22404), .Y(n18785) );
  INVx1_ASAP7_75t_SL U24696 ( .A(n18576), .Y(n18786) );
  BUFx6f_ASAP7_75t_SL U24697 ( .A(n24050), .Y(n18788) );
  NOR2x1p5_ASAP7_75t_SL U24698 ( .A(n18791), .B(n18790), .Y(
        u0_0_leon3x0_p0_divi[25]) );
  INVxp67_ASAP7_75t_SL U24699 ( .A(n25487), .Y(n18790) );
  NOR2x1_ASAP7_75t_SL U24700 ( .A(n18788), .B(n28769), .Y(n18791) );
  NAND2xp5_ASAP7_75t_SL U24701 ( .A(n18788), .B(n28631), .Y(n25484) );
  OA21x2_ASAP7_75t_SL U24702 ( .A1(n26236), .A2(n23849), .B(n25483), .Y(n18789) );
  NOR2xp33_ASAP7_75t_SL U24703 ( .A(n24062), .B(n28769), .Y(n27193) );
  AND2x2_ASAP7_75t_SL U24704 ( .A(n27192), .B(n23554), .Y(n18792) );
  OAI21x1_ASAP7_75t_SL U24705 ( .A1(n31997), .A2(n22415), .B(n25253), .Y(
        n32879) );
  INVx2_ASAP7_75t_SL U24706 ( .A(n32879), .Y(n32801) );
  NOR2x1_ASAP7_75t_SL U24707 ( .A(n32879), .B(n31737), .Y(n32723) );
  NOR2x1_ASAP7_75t_SL U24708 ( .A(n32728), .B(n31704), .Y(n31730) );
  NOR2x1_ASAP7_75t_SL U24709 ( .A(add_x_735_n183), .B(add_x_735_n149), .Y(
        add_x_735_n147) );
  NAND2x1_ASAP7_75t_SL U24710 ( .A(add_x_735_n167), .B(add_x_735_n151), .Y(
        add_x_735_n149) );
  HB1xp67_ASAP7_75t_SL U24711 ( .A(n31435), .Y(n18793) );
  OAI21xp5_ASAP7_75t_SL U24712 ( .A1(n30514), .A2(n22415), .B(n30513), .Y(
        n33011) );
  AOI21x1_ASAP7_75t_SL U24713 ( .A1(n32785), .A2(n32784), .B(n32783), .Y(
        n32816) );
  NAND3x2_ASAP7_75t_SL U24714 ( .A(n26352), .B(n26757), .C(n30115), .Y(n32153)
         );
  NOR2x1p5_ASAP7_75t_SL U24715 ( .A(n24679), .B(n31813), .Y(n32068) );
  NAND2x1p5_ASAP7_75t_SL U24716 ( .A(n24736), .B(n32153), .Y(n31813) );
  NAND2x1_ASAP7_75t_SL U24717 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_), 
        .B(n31262), .Y(n32443) );
  NAND2x1p5_ASAP7_75t_SL U24718 ( .A(n13499), .B(n32443), .Y(n31582) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24719 ( .A1(n31544), .A2(n31543), .B(n31542), 
        .C(n31541), .Y(n4348) );
  NOR2x1_ASAP7_75t_SL U24720 ( .A(n26157), .B(n24470), .Y(n27210) );
  NOR2x1p5_ASAP7_75t_SL U24721 ( .A(n28448), .B(n28447), .Y(n29789) );
  INVx1_ASAP7_75t_SL U24722 ( .A(n28446), .Y(n28447) );
  OAI21xp5_ASAP7_75t_SL U24723 ( .A1(n26937), .A2(n28987), .B(n25119), .Y(
        n29608) );
  NOR2x1_ASAP7_75t_SL U24724 ( .A(n25044), .B(n25022), .Y(n24573) );
  AND2x4_ASAP7_75t_SL U24725 ( .A(n18857), .B(n31890), .Y(n31830) );
  NOR2x1_ASAP7_75t_SL U24726 ( .A(n31702), .B(n31743), .Y(n32695) );
  NAND2x1_ASAP7_75t_SL U24727 ( .A(n32707), .B(n31707), .Y(n31742) );
  OAI21x1_ASAP7_75t_SL U24728 ( .A1(n32707), .A2(n31708), .B(n31742), .Y(
        n11260) );
  NAND2x1_ASAP7_75t_SL U24729 ( .A(n32716), .B(n31755), .Y(n32707) );
  NOR2x1_ASAP7_75t_SL U24730 ( .A(n31695), .B(n32786), .Y(n31705) );
  NAND2xp5_ASAP7_75t_SL U24731 ( .A(n31706), .B(n31705), .Y(n31731) );
  NOR2x1p5_ASAP7_75t_SL U24732 ( .A(n22378), .B(n30793), .Y(n30794) );
  AOI21x1_ASAP7_75t_SL U24733 ( .A1(n29626), .A2(n22432), .B(n28864), .Y(
        n30793) );
  NOR2x1p5_ASAP7_75t_SL U24734 ( .A(n22378), .B(n31012), .Y(n31013) );
  AOI21x1_ASAP7_75t_SL U24735 ( .A1(n30473), .A2(n22432), .B(n28955), .Y(
        n31012) );
  NOR2x2_ASAP7_75t_SL U24736 ( .A(n25033), .B(n25032), .Y(n30130) );
  INVx2_ASAP7_75t_SL U24737 ( .A(n25044), .Y(n25032) );
  XOR2xp5_ASAP7_75t_SL U24738 ( .A(n18795), .B(DP_OP_5187J1_124_3275_n160), 
        .Y(u0_0_leon3x0_p0_div0_addout_20_) );
  AND2x2_ASAP7_75t_SL U24739 ( .A(DP_OP_5187J1_124_3275_n159), .B(
        DP_OP_5187J1_124_3275_n319), .Y(n18795) );
  NAND2x1_ASAP7_75t_SL U24740 ( .A(n24978), .B(n32705), .Y(n31306) );
  NAND2x1p5_ASAP7_75t_SL U24741 ( .A(n25570), .B(n32705), .Y(n32662) );
  INVx3_ASAP7_75t_SL U24742 ( .A(n32705), .Y(n22393) );
  NOR2x1_ASAP7_75t_SL U24743 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_STPEND_), 
        .B(n31306), .Y(n25014) );
  NAND2x1_ASAP7_75t_SL U24744 ( .A(n31001), .B(n30013), .Y(n31488) );
  INVx4_ASAP7_75t_SL U24745 ( .A(n28869), .Y(n28847) );
  AOI21xp5_ASAP7_75t_SL U24746 ( .A1(u0_0_leon3x0_p0_dci[36]), .A2(n22398), 
        .B(n25206), .Y(n29815) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24747 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__31_), .B(n31343), .C(n30949), .Y(n30950)
         );
  NAND2x1_ASAP7_75t_SL U24748 ( .A(n25509), .B(n25508), .Y(n29800) );
  XOR2xp5_ASAP7_75t_SL U24749 ( .A(n18796), .B(DP_OP_5187J1_124_3275_n95), .Y(
        u0_0_leon3x0_p0_div0_addout_27_) );
  AND2x2_ASAP7_75t_SL U24750 ( .A(DP_OP_5187J1_124_3275_n94), .B(
        DP_OP_5187J1_124_3275_n312), .Y(n18796) );
  INVx1_ASAP7_75t_SL U24751 ( .A(n25883), .Y(n18797) );
  INVx2_ASAP7_75t_SL U24752 ( .A(n18797), .Y(n18798) );
  NAND2x1p5_ASAP7_75t_SL U24753 ( .A(n24733), .B(n24734), .Y(n25883) );
  BUFx2_ASAP7_75t_SL U24754 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__0_), .Y(
        n18799) );
  BUFx2_ASAP7_75t_SL U24755 ( .A(n4081), .Y(n18800) );
  HB1xp67_ASAP7_75t_SL U24756 ( .A(n31629), .Y(n18801) );
  XOR2xp5_ASAP7_75t_SL U24757 ( .A(n18802), .B(DP_OP_5187J1_124_3275_n122), 
        .Y(u0_0_leon3x0_p0_div0_addout_24_) );
  AND2x2_ASAP7_75t_SL U24758 ( .A(DP_OP_5187J1_124_3275_n121), .B(
        DP_OP_5187J1_124_3275_n315), .Y(n18802) );
  XOR2xp5_ASAP7_75t_SL U24759 ( .A(n18803), .B(DP_OP_5187J1_124_3275_n142), 
        .Y(u0_0_leon3x0_p0_div0_addout_22_) );
  AND2x2_ASAP7_75t_SL U24760 ( .A(DP_OP_5187J1_124_3275_n141), .B(
        DP_OP_5187J1_124_3275_n317), .Y(n18803) );
  INVx3_ASAP7_75t_SL U24761 ( .A(n28977), .Y(n28975) );
  OAI21xp5_ASAP7_75t_SL U24762 ( .A1(n30007), .A2(n27218), .B(n27217), .Y(
        n30495) );
  XOR2xp5_ASAP7_75t_SL U24763 ( .A(n18804), .B(DP_OP_5187J1_124_3275_n178), 
        .Y(u0_0_leon3x0_p0_div0_addout_18_) );
  AND2x2_ASAP7_75t_SL U24764 ( .A(DP_OP_5187J1_124_3275_n177), .B(
        DP_OP_5187J1_124_3275_n321), .Y(n18804) );
  BUFx6f_ASAP7_75t_SL U24765 ( .A(n29010), .Y(n18805) );
  BUFx3_ASAP7_75t_SL U24766 ( .A(n29010), .Y(n18806) );
  NOR2x1_ASAP7_75t_SL U24767 ( .A(n25366), .B(n25171), .Y(n29010) );
  NOR2x1_ASAP7_75t_SL U24768 ( .A(n24646), .B(n30646), .Y(n31874) );
  XOR2xp5_ASAP7_75t_SL U24769 ( .A(n18807), .B(DP_OP_5187J1_124_3275_n189), 
        .Y(u0_0_leon3x0_p0_div0_addout_17_) );
  AND2x2_ASAP7_75t_SL U24770 ( .A(DP_OP_5187J1_124_3275_n188), .B(
        DP_OP_5187J1_124_3275_n322), .Y(n18807) );
  NAND2xp5_ASAP7_75t_SL U24771 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), 
        .B(n25379), .Y(n25171) );
  XOR2xp5_ASAP7_75t_SL U24772 ( .A(n18808), .B(DP_OP_5187J1_124_3275_n133), 
        .Y(u0_0_leon3x0_p0_div0_addout_23_) );
  AND2x2_ASAP7_75t_SL U24773 ( .A(DP_OP_5187J1_124_3275_n132), .B(
        DP_OP_5187J1_124_3275_n316), .Y(n18808) );
  XOR2xp5_ASAP7_75t_SL U24774 ( .A(n18809), .B(DP_OP_5187J1_124_3275_n153), 
        .Y(u0_0_leon3x0_p0_div0_addout_21_) );
  AND2x2_ASAP7_75t_SL U24775 ( .A(DP_OP_5187J1_124_3275_n152), .B(
        DP_OP_5187J1_124_3275_n318), .Y(n18809) );
  XOR2xp5_ASAP7_75t_SL U24776 ( .A(n18810), .B(DP_OP_5187J1_124_3275_n171), 
        .Y(u0_0_leon3x0_p0_div0_addout_19_) );
  AND2x2_ASAP7_75t_SL U24777 ( .A(DP_OP_5187J1_124_3275_n170), .B(
        DP_OP_5187J1_124_3275_n320), .Y(n18810) );
  XNOR2xp5_ASAP7_75t_SRAM U24778 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__7_), 
        .B(n32171), .Y(n26862) );
  INVx2_ASAP7_75t_SL U24779 ( .A(n25783), .Y(n18811) );
  INVx2_ASAP7_75t_SL U24780 ( .A(n18811), .Y(n18812) );
  INVx3_ASAP7_75t_SL U24781 ( .A(n18811), .Y(n18813) );
  INVx2_ASAP7_75t_SL U24782 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__30_), .Y(
        n18814) );
  NOR2x1_ASAP7_75t_SL U24783 ( .A(n18814), .B(n32051), .Y(n18815) );
  INVx3_ASAP7_75t_SL U24784 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__30_), .Y(
        n30909) );
  INVx4_ASAP7_75t_SL U24785 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__31_), .Y(
        n32051) );
  XOR2xp5_ASAP7_75t_SL U24786 ( .A(n18816), .B(DP_OP_5187J1_124_3275_n75), .Y(
        u0_0_leon3x0_p0_div0_addout_29_) );
  AND2x2_ASAP7_75t_SL U24787 ( .A(DP_OP_5187J1_124_3275_n74), .B(
        DP_OP_5187J1_124_3275_n310), .Y(n18816) );
  XOR2xp5_ASAP7_75t_SL U24788 ( .A(n18817), .B(DP_OP_5187J1_124_3275_n64), .Y(
        u0_0_leon3x0_p0_div0_addout_30_) );
  AND2x2_ASAP7_75t_SL U24789 ( .A(DP_OP_5187J1_124_3275_n63), .B(
        DP_OP_5187J1_124_3275_n60), .Y(n18817) );
  BUFx3_ASAP7_75t_SL U24790 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__22_), .Y(
        n18818) );
  BUFx2_ASAP7_75t_SL U24791 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__22_), .Y(
        n18819) );
  OAI21xp5_ASAP7_75t_SL U24792 ( .A1(n31857), .A2(n26815), .B(n24880), .Y(
        n25216) );
  OAI21xp5_ASAP7_75t_SL U24793 ( .A1(n24740), .A2(n31857), .B(n24745), .Y(
        n24741) );
  NOR2x1p5_ASAP7_75t_SL U24794 ( .A(n28096), .B(n31238), .Y(n27496) );
  NAND2x1p5_ASAP7_75t_SL U24795 ( .A(n31325), .B(n27473), .Y(n31238) );
  HB1xp67_ASAP7_75t_SL U24796 ( .A(n24877), .Y(n18820) );
  NAND2xp5_ASAP7_75t_SL U24797 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(
        DP_OP_1196_128_7433_n456), .Y(n18821) );
  OAI21xp33_ASAP7_75t_SRAM U24798 ( .A1(n32083), .A2(n30909), .B(n30908), .Y(
        DP_OP_1196_128_7433_n475) );
  OAI21xp33_ASAP7_75t_SRAM U24799 ( .A1(n30907), .A2(n30909), .B(n30908), .Y(
        DP_OP_1196_128_7433_n477) );
  NAND2x1_ASAP7_75t_SL U24800 ( .A(n24745), .B(n18815), .Y(n24746) );
  AND2x2_ASAP7_75t_SL U24801 ( .A(n25884), .B(n25883), .Y(n29059) );
  NAND2x1p5_ASAP7_75t_SL U24802 ( .A(n25882), .B(n25883), .Y(n31885) );
  XOR2xp5_ASAP7_75t_SL U24803 ( .A(n18822), .B(mult_x_1196_n707), .Y(n23883)
         );
  NAND2xp5_ASAP7_75t_SL U24804 ( .A(mult_x_1196_n706), .B(n24273), .Y(n18822)
         );
  INVx2_ASAP7_75t_SL U24805 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), .Y(
        n18823) );
  INVx1_ASAP7_75t_SL U24806 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), .Y(
        n24745) );
  INVx2_ASAP7_75t_SL U24807 ( .A(n26298), .Y(n28845) );
  INVxp33_ASAP7_75t_SRAM U24808 ( .A(n26850), .Y(n18824) );
  INVxp33_ASAP7_75t_SRAM U24809 ( .A(n18824), .Y(n18825) );
  NAND2x2_ASAP7_75t_SL U24810 ( .A(n31627), .B(n31629), .Y(n32719) );
  NOR2x1_ASAP7_75t_SL U24811 ( .A(n32709), .B(n32695), .Y(n31755) );
  NAND2x1_ASAP7_75t_SL U24812 ( .A(n30639), .B(n30638), .Y(n31350) );
  NAND2xp5_ASAP7_75t_SL U24813 ( .A(n32187), .B(n30940), .Y(n24865) );
  NAND2xp5_ASAP7_75t_SL U24814 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__4_), .B(
        n32164), .Y(n24826) );
  INVx1_ASAP7_75t_SL U24815 ( .A(n30714), .Y(n18826) );
  INVx2_ASAP7_75t_SL U24816 ( .A(n18826), .Y(n18827) );
  BUFx3_ASAP7_75t_SL U24817 ( .A(n24635), .Y(n18828) );
  BUFx12f_ASAP7_75t_SL U24818 ( .A(n24635), .Y(n18829) );
  BUFx12f_ASAP7_75t_SL U24819 ( .A(n24635), .Y(n18830) );
  INVx4_ASAP7_75t_SL U24820 ( .A(n30714), .Y(n24635) );
  INVxp33_ASAP7_75t_SRAM U24821 ( .A(n32188), .Y(n18831) );
  INVx1_ASAP7_75t_SL U24822 ( .A(n18831), .Y(n18832) );
  NOR2x1_ASAP7_75t_SL U24823 ( .A(n22379), .B(n30017), .Y(n30208) );
  NOR2x1p5_ASAP7_75t_SL U24824 ( .A(n25016), .B(n25015), .Y(n30017) );
  AOI21xp5_ASAP7_75t_SL U24825 ( .A1(DP_OP_5187J1_124_3275_n193), .A2(
        DP_OP_5187J1_124_3275_n261), .B(DP_OP_5187J1_124_3275_n194), .Y(
        DP_OP_5187J1_124_3275_n2) );
  NOR2x1_ASAP7_75t_SL U24826 ( .A(n24778), .B(n18850), .Y(n30934) );
  NOR2x1p5_ASAP7_75t_SL U24827 ( .A(n32689), .B(n18827), .Y(n32060) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24828 ( .A1(n18832), .A2(n30943), .B(n32192), 
        .C(n30942), .Y(n4350) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24829 ( .A1(n18832), .A2(n32190), .B(n32192), 
        .C(n32107), .Y(n32108) );
  OAI21xp33_ASAP7_75t_SRAM U24830 ( .A1(n18819), .A2(n22377), .B(n24917), .Y(
        n4177) );
  INVx1_ASAP7_75t_SL U24831 ( .A(n30934), .Y(n24806) );
  NAND2xp33_ASAP7_75t_SRAM U24832 ( .A(n18819), .B(n24999), .Y(n24854) );
  NOR2x1_ASAP7_75t_SL U24833 ( .A(DP_OP_5187J1_124_3275_n237), .B(
        DP_OP_5187J1_124_3275_n244), .Y(DP_OP_5187J1_124_3275_n235) );
  NAND2x1_ASAP7_75t_SL U24834 ( .A(DP_OP_5187J1_124_3275_n249), .B(
        DP_OP_5187J1_124_3275_n235), .Y(DP_OP_5187J1_124_3275_n229) );
  HB1xp67_ASAP7_75t_SL U24835 ( .A(DP_OP_5187J1_124_3275_n250), .Y(n18833) );
  NOR2x2_ASAP7_75t_SL U24836 ( .A(n18814), .B(n32051), .Y(n32086) );
  NOR2x1_ASAP7_75t_SL U24837 ( .A(n25045), .B(n25044), .Y(n31473) );
  AND2x2_ASAP7_75t_SL U24838 ( .A(n18846), .B(n26854), .Y(n32164) );
  AOI22xp5_ASAP7_75t_SL U24839 ( .A1(n26853), .A2(n26852), .B1(
        u0_0_leon3x0_p0_iu_v_X__CTRL__RD__5_), .B2(n26851), .Y(n26866) );
  INVx1_ASAP7_75t_SL U24840 ( .A(n26853), .Y(n32166) );
  NAND2x2_ASAP7_75t_SL U24841 ( .A(n24681), .B(n31890), .Y(n30714) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24842 ( .A1(n24893), .A2(n24892), .B(n31890), 
        .C(n24891), .Y(n25219) );
  NAND2x2_ASAP7_75t_SL U24843 ( .A(n30503), .B(n30504), .Y(n31890) );
  NOR2x1p5_ASAP7_75t_SL U24844 ( .A(n30505), .B(n30504), .Y(n32123) );
  NAND2x1p5_ASAP7_75t_SL U24845 ( .A(n24888), .B(n25214), .Y(n30504) );
  INVx1_ASAP7_75t_SL U24846 ( .A(DP_OP_5187J1_124_3275_n206), .Y(n20560) );
  NOR2x1_ASAP7_75t_SL U24847 ( .A(u0_0_leon3x0_p0_div0_vaddin1[14]), .B(
        u0_0_leon3x0_p0_div0_b[14]), .Y(DP_OP_5187J1_124_3275_n206) );
  INVx2_ASAP7_75t_SL U24848 ( .A(n24775), .Y(n24796) );
  HB1xp67_ASAP7_75t_SL U24849 ( .A(DP_OP_5187J1_124_3275_n288), .Y(n18834) );
  HB1xp67_ASAP7_75t_SL U24850 ( .A(DP_OP_5187J1_124_3275_n277), .Y(n18835) );
  BUFx2_ASAP7_75t_SL U24851 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__21_), .Y(
        n18841) );
  NOR2x2_ASAP7_75t_SL U24852 ( .A(n24479), .B(n31627), .Y(n31877) );
  INVx2_ASAP7_75t_SL U24853 ( .A(n30191), .Y(n32120) );
  HB1xp67_ASAP7_75t_SL U24854 ( .A(DP_OP_5187J1_124_3275_n297), .Y(n18836) );
  NOR2x1_ASAP7_75t_SL U24855 ( .A(n25044), .B(n25022), .Y(n29991) );
  INVx1_ASAP7_75t_SL U24856 ( .A(n23831), .Y(n18837) );
  BUFx2_ASAP7_75t_SL U24857 ( .A(n24796), .Y(n18838) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24858 ( .A1(n26298), .A2(n18813), .B(n26390), 
        .C(n25111), .Y(n25460) );
  AOI21xp33_ASAP7_75t_SRAM U24859 ( .A1(n22416), .A2(n23365), .B(n18813), .Y(
        n25116) );
  AOI21xp33_ASAP7_75t_SRAM U24860 ( .A1(n22416), .A2(n23969), .B(n18813), .Y(
        n25194) );
  INVx2_ASAP7_75t_SL U24861 ( .A(n18812), .Y(n25476) );
  NAND2x1p5_ASAP7_75t_SL U24862 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), .Y(n24877) );
  INVx4_ASAP7_75t_SL U24863 ( .A(n18818), .Y(n32079) );
  NOR2x1_ASAP7_75t_SL U24864 ( .A(n31585), .B(n18852), .Y(n32272) );
  NOR2x1p5_ASAP7_75t_SL U24865 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .Y(n25226) );
  NOR2x1_ASAP7_75t_SL U24866 ( .A(u0_0_leon3x0_p0_ici[49]), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .Y(DP_OP_1196_128_7433_n147)
         );
  NAND2xp5_ASAP7_75t_SL U24867 ( .A(u0_0_leon3x0_p0_ici[49]), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .Y(DP_OP_1196_128_7433_n148)
         );
  INVx1_ASAP7_75t_SL U24868 ( .A(n25226), .Y(n32078) );
  NOR2x2_ASAP7_75t_SL U24869 ( .A(n31380), .B(n24796), .Y(n24786) );
  BUFx6f_ASAP7_75t_SL U24870 ( .A(DP_OP_5187J1_124_3275_n2), .Y(n22225) );
  INVxp33_ASAP7_75t_SRAM U24871 ( .A(n32171), .Y(n26849) );
  INVxp33_ASAP7_75t_SRAM U24872 ( .A(n24998), .Y(n24744) );
  INVxp33_ASAP7_75t_SRAM U24873 ( .A(n26855), .Y(n18846) );
  AOI22xp5_ASAP7_75t_SL U24874 ( .A1(n22416), .A2(n24231), .B1(n22449), .B2(
        n25200), .Y(n25907) );
  INVx6_ASAP7_75t_SL U24875 ( .A(n24469), .Y(n22416) );
  NAND2xp5_ASAP7_75t_SL U24876 ( .A(n23091), .B(n22416), .Y(n25478) );
  NAND2xp5_ASAP7_75t_SL U24877 ( .A(n23958), .B(n22416), .Y(n25784) );
  AOI211x1_ASAP7_75t_SL U24878 ( .A1(n27098), .A2(n25794), .B(n25793), .C(
        n25792), .Y(n28503) );
  O2A1O1Ixp5_ASAP7_75t_SL U24879 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__7_), 
        .A2(n32186), .B(n19208), .C(n19209), .Y(n19210) );
  NOR2x1_ASAP7_75t_SL U24880 ( .A(n28110), .B(n26470), .Y(n28111) );
  INVxp33_ASAP7_75t_SRAM U24881 ( .A(n31862), .Y(n18843) );
  NAND2xp5_ASAP7_75t_SL U24882 ( .A(DP_OP_5187J1_124_3275_n256), .B(
        DP_OP_5187J1_124_3275_n330), .Y(DP_OP_5187J1_124_3275_n30) );
  XNOR2x2_ASAP7_75t_SL U24883 ( .A(u0_0_leon3x0_p0_iu_de_icc_1_), .B(
        u0_0_leon3x0_p0_iu_de_icc_3_), .Y(n24873) );
  NAND2xp5_ASAP7_75t_SL U24884 ( .A(u0_0_leon3x0_p0_div0_vaddin1[14]), .B(
        u0_0_leon3x0_p0_div0_b[14]), .Y(DP_OP_5187J1_124_3275_n209) );
  NOR2x1_ASAP7_75t_SL U24885 ( .A(n24776), .B(n23899), .Y(n24783) );
  NAND3x1_ASAP7_75t_SL U24886 ( .A(n30016), .B(n30015), .C(n31474), .Y(n31483)
         );
  NOR2x1_ASAP7_75t_SL U24887 ( .A(n25438), .B(n25445), .Y(n30016) );
  INVxp33_ASAP7_75t_SRAM U24888 ( .A(n30909), .Y(n18839) );
  XOR2xp5_ASAP7_75t_SL U24889 ( .A(n18840), .B(n30938), .Y(n24798) );
  INVx13_ASAP7_75t_SL U24890 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__1_), .Y(
        n18840) );
  NAND2x1_ASAP7_75t_SL U24891 ( .A(n27085), .B(n27084), .Y(n31545) );
  NAND2x1_ASAP7_75t_SL U24892 ( .A(n26945), .B(n26944), .Y(n28275) );
  BUFx6f_ASAP7_75t_SL U24893 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__21_), 
        .Y(n18842) );
  NAND2x2_ASAP7_75t_SL U24894 ( .A(n18841), .B(n32079), .Y(n31857) );
  AO21x2_ASAP7_75t_SL U24895 ( .A1(n23997), .A2(n18397), .B(mult_x_1196_n3111), 
        .Y(mult_x_1196_n2535) );
  OAI22xp33_ASAP7_75t_SRAM U24896 ( .A1(mult_x_1196_n3138), .A2(n24000), .B1(
        n23996), .B2(mult_x_1196_n3137), .Y(mult_x_1196_n2562) );
  NOR2x1_ASAP7_75t_SL U24897 ( .A(n24000), .B(n18958), .Y(n18957) );
  OAI21xp5_ASAP7_75t_SL U24898 ( .A1(mult_x_1196_n3239), .A2(n22953), .B(
        n22705), .Y(mult_x_1196_n2663) );
  XNOR2xp5_ASAP7_75t_SL U24899 ( .A(n24069), .B(n22926), .Y(mult_x_1196_n2762)
         );
  OAI21x1_ASAP7_75t_SL U24900 ( .A1(timer0_vtimers_1__LOAD_), .A2(n28111), .B(
        n31841), .Y(n31847) );
  BUFx12f_ASAP7_75t_SL U24901 ( .A(n31847), .Y(n22399) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24902 ( .A1(n31857), .A2(n25601), .B(n24876), 
        .C(n24859), .Y(n24860) );
  NAND2x1_ASAP7_75t_SL U24903 ( .A(n31584), .B(n32272), .Y(n31599) );
  NOR2x1_ASAP7_75t_SL U24904 ( .A(n25039), .B(n25038), .Y(n25440) );
  INVx1_ASAP7_75t_SL U24905 ( .A(n25440), .Y(n30018) );
  NAND2xp5_ASAP7_75t_SL U24906 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), 
        .B(n24882), .Y(n24753) );
  INVx1_ASAP7_75t_SL U24907 ( .A(n26817), .Y(n25217) );
  NAND2x1p5_ASAP7_75t_SL U24908 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__0_), 
        .B(n18823), .Y(n26817) );
  INVx2_ASAP7_75t_SL U24909 ( .A(n18843), .Y(n18844) );
  NOR2x1_ASAP7_75t_SL U24910 ( .A(n24746), .B(n31862), .Y(n18867) );
  NOR2xp33_ASAP7_75t_SL U24911 ( .A(n29638), .B(n30706), .Y(n18845) );
  NAND2x1_ASAP7_75t_SL U24912 ( .A(n31960), .B(n30212), .Y(n29638) );
  AND2x6_ASAP7_75t_SL U24913 ( .A(n26471), .B(n26470), .Y(n31845) );
  NAND2x1p5_ASAP7_75t_SL U24914 ( .A(n28847), .B(n28982), .Y(n28970) );
  AOI21xp5_ASAP7_75t_SL U24915 ( .A1(n28873), .A2(n28975), .B(n28872), .Y(
        n28971) );
  INVx2_ASAP7_75t_SL U24916 ( .A(n24363), .Y(n24419) );
  NOR2x1_ASAP7_75t_SL U24917 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_), 
        .B(n23899), .Y(n24808) );
  XNOR2x2_ASAP7_75t_SL U24918 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__1_), .B(
        n30938), .Y(n30921) );
  NOR2x1p5_ASAP7_75t_SL U24919 ( .A(n24418), .B(n24419), .Y(n24365) );
  INVx1_ASAP7_75t_SL U24920 ( .A(n18852), .Y(n18859) );
  INVxp33_ASAP7_75t_SRAM U24921 ( .A(n32524), .Y(n18847) );
  INVx1_ASAP7_75t_SL U24922 ( .A(n18847), .Y(n18848) );
  NAND2xp5_ASAP7_75t_SL U24923 ( .A(n24353), .B(n24396), .Y(n24354) );
  AND2x4_ASAP7_75t_SL U24924 ( .A(n24417), .B(n24365), .Y(n24420) );
  NOR2x1_ASAP7_75t_SL U24925 ( .A(n26777), .B(n18821), .Y(n24765) );
  NOR2x1p5_ASAP7_75t_SL U24926 ( .A(n24786), .B(n24783), .Y(n32186) );
  OAI21x1_ASAP7_75t_SL U24927 ( .A1(n32169), .A2(n24764), .B(n32167), .Y(
        n32170) );
  OR2x2_ASAP7_75t_SL U24928 ( .A(n24807), .B(n24774), .Y(n18849) );
  NOR2x1_ASAP7_75t_SL U24929 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_), 
        .B(n24796), .Y(n24807) );
  NOR2x1_ASAP7_75t_SL U24930 ( .A(n31586), .B(n31462), .Y(n31262) );
  NOR2x1p5_ASAP7_75t_SL U24931 ( .A(n31001), .B(n30014), .Y(n31486) );
  OAI21x1_ASAP7_75t_SL U24932 ( .A1(n29914), .A2(n29913), .B(n31474), .Y(
        n30014) );
  NOR2xp33_ASAP7_75t_SL U24933 ( .A(n24780), .B(n24779), .Y(n18850) );
  BUFx3_ASAP7_75t_SL U24934 ( .A(n31547), .Y(n18851) );
  NAND2xp5_ASAP7_75t_SL U24935 ( .A(n32030), .B(n29997), .Y(n31547) );
  INVx1_ASAP7_75t_SL U24936 ( .A(n24549), .Y(n31620) );
  NOR2x1_ASAP7_75t_SL U24937 ( .A(n32038), .B(n24696), .Y(ahb0_v_HREADY_) );
  NOR2x1p5_ASAP7_75t_SL U24938 ( .A(ahb0_r_DEFSLV_), .B(n32037), .Y(n24696) );
  AOI21xp33_ASAP7_75t_SRAM U24939 ( .A1(n30652), .A2(
        u0_0_leon3x0_p0_iu_de_icc_2_), .B(n24679), .Y(n29131) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24940 ( .A1(u0_0_leon3x0_p0_iu_r_D__ANNUL_), 
        .A2(n25882), .B(n18798), .C(n30681), .Y(n24893) );
  INVxp33_ASAP7_75t_SRAM U24941 ( .A(u0_0_leon3x0_p0_iu_de_icc_2_), .Y(n29173)
         );
  AOI22xp5_ASAP7_75t_SL U24942 ( .A1(n24807), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__28_), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_), .B2(n24808), .Y(n24777) );
  NOR2x1_ASAP7_75t_SL U24943 ( .A(n25572), .B(n18830), .Y(n18900) );
  NOR2x1_ASAP7_75t_SL U24944 ( .A(n25572), .B(n18829), .Y(n18901) );
  NAND2x1p5_ASAP7_75t_SL U24945 ( .A(n32197), .B(n24978), .Y(n31697) );
  NOR2x1_ASAP7_75t_SL U24946 ( .A(n18800), .B(n31602), .Y(n24978) );
  OR3x1_ASAP7_75t_SL U24947 ( .A(n31257), .B(n24530), .C(n32198), .Y(n18852)
         );
  INVx3_ASAP7_75t_SL U24948 ( .A(n31574), .Y(n32198) );
  NOR2x1_ASAP7_75t_SL U24949 ( .A(n28869), .B(n28868), .Y(n28980) );
  OAI22xp33_ASAP7_75t_SRAM U24950 ( .A1(n27144), .A2(n25110), .B1(n18380), 
        .B2(n25190), .Y(n25111) );
  OAI21xp5_ASAP7_75t_SL U24951 ( .A1(n24691), .A2(n25190), .B(n25476), .Y(
        n25191) );
  NAND2xp5_ASAP7_75t_SL U24952 ( .A(n28845), .B(n22416), .Y(n25190) );
  NAND2xp5_ASAP7_75t_SL U24953 ( .A(n24681), .B(n26735), .Y(n26452) );
  BUFx6f_ASAP7_75t_SL U24954 ( .A(n28961), .Y(n22410) );
  NAND2x1p5_ASAP7_75t_SL U24955 ( .A(n28975), .B(n28845), .Y(n28850) );
  INVx3_ASAP7_75t_SL U24956 ( .A(n28850), .Y(n27098) );
  NOR2x1_ASAP7_75t_SL U24957 ( .A(n24766), .B(n24764), .Y(n26853) );
  NOR2x1_ASAP7_75t_SL U24958 ( .A(n24747), .B(n26854), .Y(n24764) );
  NOR2x1p5_ASAP7_75t_SL U24959 ( .A(n18876), .B(n31890), .Y(n26204) );
  INVx3_ASAP7_75t_SL U24960 ( .A(n28835), .Y(n29595) );
  NOR2x1p5_ASAP7_75t_SL U24961 ( .A(n24427), .B(n26176), .Y(n28835) );
  OAI21xp5_ASAP7_75t_SL U24962 ( .A1(n30282), .A2(n29595), .B(n27070), .Y(
        n27071) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24963 ( .A1(n18799), .A2(n25214), .B(n24914), 
        .C(n24913), .Y(n24916) );
  INVxp33_ASAP7_75t_SRAM U24964 ( .A(n25214), .Y(n31818) );
  INVxp33_ASAP7_75t_SRAM U24965 ( .A(n24319), .Y(n18853) );
  INVxp33_ASAP7_75t_SRAM U24966 ( .A(n18853), .Y(n18854) );
  INVxp33_ASAP7_75t_SRAM U24967 ( .A(n24333), .Y(n18855) );
  INVxp33_ASAP7_75t_SRAM U24968 ( .A(n18855), .Y(n18856) );
  NOR2x1p5_ASAP7_75t_SL U24969 ( .A(n5061), .B(n2846), .Y(timer0_N91) );
  NOR2x1_ASAP7_75t_SL U24970 ( .A(n24831), .B(n24830), .Y(n26850) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U24971 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__7_), .A2(n32171), .B(n24752), .C(n24751), .Y(n24758) );
  NOR2x1_ASAP7_75t_SL U24972 ( .A(DP_OP_5187J1_124_3275_n151), .B(
        DP_OP_5187J1_124_3275_n158), .Y(DP_OP_5187J1_124_3275_n145) );
  NOR2x1_ASAP7_75t_SL U24973 ( .A(u0_0_leon3x0_p0_div0_vaddin1[21]), .B(
        u0_0_leon3x0_p0_div0_b[21]), .Y(DP_OP_5187J1_124_3275_n151) );
  NAND2x1_ASAP7_75t_SL U24974 ( .A(DP_OP_5187J1_124_3275_n129), .B(
        DP_OP_5187J1_124_3275_n145), .Y(DP_OP_5187J1_124_3275_n127) );
  NOR2x1_ASAP7_75t_SL U24975 ( .A(DP_OP_5187J1_124_3275_n131), .B(
        DP_OP_5187J1_124_3275_n138), .Y(DP_OP_5187J1_124_3275_n129) );
  NOR2x1_ASAP7_75t_SL U24976 ( .A(n29206), .B(n31809), .Y(n31426) );
  INVx2_ASAP7_75t_SL U24977 ( .A(n31426), .Y(n26807) );
  NAND2x1p5_ASAP7_75t_SL U24978 ( .A(n24872), .B(n30683), .Y(n31809) );
  NAND2x1_ASAP7_75t_SL U24979 ( .A(n26775), .B(n26807), .Y(n31435) );
  AND2x2_ASAP7_75t_SL U24980 ( .A(n26202), .B(n26203), .Y(n18857) );
  HB1xp67_ASAP7_75t_SL U24981 ( .A(n32667), .Y(n18858) );
  NOR2x1_ASAP7_75t_SL U24982 ( .A(n29009), .B(n29008), .Y(n32119) );
  AOI22xp33_ASAP7_75t_SRAM U24983 ( .A1(u0_0_leon3x0_p0_dci[8]), .A2(n31828), 
        .B1(n31830), .B2(u0_0_leon3x0_p0_iu_N5467), .Y(n30910) );
  INVxp33_ASAP7_75t_SRAM U24984 ( .A(n31830), .Y(n19219) );
  AND2x4_ASAP7_75t_SL U24985 ( .A(n22379), .B(n31830), .Y(n31994) );
  AOI21xp5_ASAP7_75t_SL U24986 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_4_), .A2(n31833), .B(n29479), .Y(n32692) );
  NOR3xp33_ASAP7_75t_SL U24987 ( .A(n31257), .B(n24530), .C(n32198), .Y(n32281) );
  NAND2x2_ASAP7_75t_SL U24988 ( .A(n3065), .B(n31563), .Y(n32545) );
  AO21x2_ASAP7_75t_SL U24989 ( .A1(n31549), .A2(n32281), .B(n31548), .Y(n31563) );
  HB1xp67_ASAP7_75t_SL U24990 ( .A(n5061), .Y(n18860) );
  HB1xp67_ASAP7_75t_SL U24991 ( .A(n24349), .Y(n18861) );
  XNOR2xp5_ASAP7_75t_SL U24992 ( .A(n24064), .B(n23955), .Y(mult_x_1196_n3233)
         );
  INVx6_ASAP7_75t_SL U24993 ( .A(n32719), .Y(n24583) );
  INVx1_ASAP7_75t_SL U24994 ( .A(n23834), .Y(n18897) );
  INVxp33_ASAP7_75t_SRAM U24995 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__0_), .Y(
        n23834) );
  NAND2x1p5_ASAP7_75t_SL U24996 ( .A(n18568), .B(n26739), .Y(
        u0_0_leon3x0_p0_divi[0]) );
  OAI22xp5_ASAP7_75t_SL U24997 ( .A1(mult_x_1196_n3206), .A2(n22802), .B1(
        mult_x_1196_n3205), .B2(n22248), .Y(n18863) );
  XNOR2xp5_ASAP7_75t_SL U24998 ( .A(n23168), .B(mult_x_1196_n2630), .Y(n23167)
         );
  OAI22xp5_ASAP7_75t_SL U24999 ( .A1(mult_x_1196_n3206), .A2(n22802), .B1(
        mult_x_1196_n3205), .B2(n22248), .Y(mult_x_1196_n2630) );
  INVx2_ASAP7_75t_SL U25000 ( .A(n32086), .Y(n26818) );
  NOR2x1_ASAP7_75t_SL U25001 ( .A(n24871), .B(n24870), .Y(n30683) );
  HB1xp67_ASAP7_75t_SL U25002 ( .A(n18860), .Y(n18864) );
  INVxp33_ASAP7_75t_SRAM U25003 ( .A(n24414), .Y(n18865) );
  NOR2x1p5_ASAP7_75t_SL U25004 ( .A(n24746), .B(n31862), .Y(n18866) );
  NOR2x1_ASAP7_75t_SL U25005 ( .A(n24746), .B(n31862), .Y(n32095) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25006 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__4_), .A2(n32164), .B(n26864), .C(n26863), .Y(n26865) );
  NAND2x1p5_ASAP7_75t_SL U25007 ( .A(n25128), .B(n25127), .Y(n29150) );
  INVx1_ASAP7_75t_SL U25008 ( .A(n25901), .Y(n25128) );
  NAND2x1_ASAP7_75t_SL U25009 ( .A(n26583), .B(n26582), .Y(n28578) );
  NAND2x1_ASAP7_75t_SL U25010 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__3_), .B(n23903), .Y(n24552) );
  BUFx2_ASAP7_75t_SL U25011 ( .A(mult_x_1196_n667), .Y(n23902) );
  NAND3x1_ASAP7_75t_SL U25012 ( .A(n24769), .B(n24768), .C(n24767), .Y(n30810)
         );
  NAND2xp5_ASAP7_75t_SL U25013 ( .A(n30810), .B(n30809), .Y(n32172) );
  INVx3_ASAP7_75t_SL U25014 ( .A(n28967), .Y(n28986) );
  NOR2x1p5_ASAP7_75t_SL U25015 ( .A(n26298), .B(n28975), .Y(n28967) );
  AOI22xp33_ASAP7_75t_SRAM U25016 ( .A1(n28980), .A2(add_x_735_A_2_), .B1(
        n28967), .B2(n28966), .Y(n28969) );
  NOR3xp33_ASAP7_75t_SL U25017 ( .A(n18856), .B(timer0_N77), .C(timer0_N78), 
        .Y(n18868) );
  NAND2x1_ASAP7_75t_SL U25018 ( .A(n24331), .B(n24405), .Y(n24333) );
  XOR2xp5_ASAP7_75t_SL U25019 ( .A(n18869), .B(mult_x_1196_n629), .Y(n23897)
         );
  AND2x2_ASAP7_75t_SL U25020 ( .A(n18539), .B(n23925), .Y(n18869) );
  INVx1_ASAP7_75t_SL U25021 ( .A(n24806), .Y(n18870) );
  BUFx16f_ASAP7_75t_SL U25022 ( .A(n29128), .Y(n22373) );
  NAND2x1p5_ASAP7_75t_SL U25023 ( .A(n25362), .B(n18805), .Y(n29128) );
  NOR2x2_ASAP7_75t_SL U25024 ( .A(n3878), .B(n18866), .Y(
        DP_OP_1196_128_7433_n456) );
  NOR2x1_ASAP7_75t_SL U25025 ( .A(n4927), .B(n32095), .Y(
        DP_OP_1196_128_7433_n452) );
  NOR2x1_ASAP7_75t_SL U25026 ( .A(u0_0_leon3x0_p0_ici[34]), .B(
        DP_OP_1196_128_7433_n456), .Y(DP_OP_1196_128_7433_n338) );
  NOR3xp33_ASAP7_75t_SL U25027 ( .A(n18854), .B(timer0_N83), .C(timer0_N84), 
        .Y(n18871) );
  NAND2x1_ASAP7_75t_SL U25028 ( .A(n24381), .B(n24411), .Y(n24319) );
  OAI21x1_ASAP7_75t_SL U25029 ( .A1(u0_0_leon3x0_p0_iu_v_A__CWP__2_), .A2(
        n24811), .B(n24810), .Y(n32185) );
  HB1xp67_ASAP7_75t_SL U25030 ( .A(n5061), .Y(n18872) );
  INVxp33_ASAP7_75t_SRAM U25031 ( .A(n24331), .Y(n18873) );
  INVx1_ASAP7_75t_SL U25032 ( .A(n18873), .Y(n18874) );
  NOR3xp33_ASAP7_75t_SL U25033 ( .A(n24325), .B(timer0_N80), .C(timer0_N81), 
        .Y(n24331) );
  NOR2x1p5_ASAP7_75t_SL U25034 ( .A(n24813), .B(n24812), .Y(n32188) );
  INVxp33_ASAP7_75t_SRAM U25035 ( .A(n18864), .Y(n24683) );
  NOR2xp67_ASAP7_75t_SRAM U25036 ( .A(n18872), .B(n4456), .Y(timer0_N81) );
  NOR2x1p5_ASAP7_75t_SL U25037 ( .A(n22380), .B(n31587), .Y(n31596) );
  NOR2x2_ASAP7_75t_SL U25038 ( .A(n4930), .B(n18866), .Y(
        DP_OP_1196_128_7433_n455) );
  XNOR2xp5_ASAP7_75t_SRAM U25039 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__6_), 
        .B(n32170), .Y(n26867) );
  XNOR2x2_ASAP7_75t_SL U25040 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__6_), .B(
        n32185), .Y(n24812) );
  AOI21x1_ASAP7_75t_SL U25041 ( .A1(n26204), .A2(n31884), .B(n26198), .Y(
        n31826) );
  OAI22xp33_ASAP7_75t_SRAM U25042 ( .A1(n18842), .A2(n24495), .B1(n23229), 
        .B2(u0_0_leon3x0_p0_iu_r_A__IMM__31_), .Y(n26370) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25043 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__5_), .A2(n30934), .B(n30933), .C(n30932), .Y(n30937) );
  OAI22xp33_ASAP7_75t_SRAM U25044 ( .A1(n18819), .A2(n24858), .B1(n18842), 
        .B2(n32083), .Y(n24743) );
  INVxp33_ASAP7_75t_SRAM U25045 ( .A(n18842), .Y(n32087) );
  NOR2x1_ASAP7_75t_SL U25046 ( .A(n32180), .B(n32181), .Y(n32183) );
  NOR2x1_ASAP7_75t_SL U25047 ( .A(n24788), .B(n24787), .Y(n32181) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25048 ( .A1(n22415), .A2(n31936), .B(
        u0_0_leon3x0_p0_c0mmu_mcii[0]), .C(n31935), .Y(n31938) );
  AOI22xp33_ASAP7_75t_SRAM U25049 ( .A1(u0_0_leon3x0_p0_c0mmu_mcii[9]), .A2(
        n31877), .B1(u0_0_leon3x0_p0_c0mmu_mcdi[45]), .B2(n24583), .Y(n33004)
         );
  NAND2xp33_ASAP7_75t_SRAM U25050 ( .A(n25334), .B(n31877), .Y(n25335) );
  NAND2xp33_ASAP7_75t_SRAM U25051 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[4]), .B(
        n31877), .Y(n25261) );
  NAND2xp33_ASAP7_75t_SRAM U25052 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[3]), .B(
        n31877), .Y(n25263) );
  OAI21xp33_ASAP7_75t_SRAM U25053 ( .A1(n30530), .A2(n22415), .B(n30529), .Y(
        n33008) );
  OAI21xp33_ASAP7_75t_SRAM U25054 ( .A1(n25250), .A2(n22415), .B(n25249), .Y(
        n32776) );
  OAI21xp33_ASAP7_75t_SRAM U25055 ( .A1(n31782), .A2(n22415), .B(n25248), .Y(
        n33046) );
  OAI21xp33_ASAP7_75t_SRAM U25056 ( .A1(n30832), .A2(n22415), .B(n30831), .Y(
        n33026) );
  OAI21xp33_ASAP7_75t_SRAM U25057 ( .A1(n25257), .A2(n22415), .B(n25256), .Y(
        n33052) );
  OAI21xp33_ASAP7_75t_SRAM U25058 ( .A1(n31792), .A2(n22415), .B(n31791), .Y(
        n33023) );
  OAI21xp33_ASAP7_75t_SRAM U25059 ( .A1(n30537), .A2(n22415), .B(n30536), .Y(
        n33017) );
  AO21x2_ASAP7_75t_SL U25060 ( .A1(n32732), .A2(n24583), .B(n31877), .Y(n32728) );
  OAI21xp33_ASAP7_75t_SRAM U25061 ( .A1(n30521), .A2(n22415), .B(n30520), .Y(
        n33014) );
  OAI21xp33_ASAP7_75t_SRAM U25062 ( .A1(n30544), .A2(n22415), .B(n30543), .Y(
        n33020) );
  NOR2x1p5_ASAP7_75t_SL U25063 ( .A(n25251), .B(n22415), .Y(n25252) );
  INVx4_ASAP7_75t_SL U25064 ( .A(n31877), .Y(n22415) );
  XNOR2xp5_ASAP7_75t_SL U25065 ( .A(n18875), .B(mult_x_1196_n622), .Y(n23900)
         );
  AND2x2_ASAP7_75t_SL U25066 ( .A(n24083), .B(n24087), .Y(n18875) );
  BUFx6f_ASAP7_75t_SL U25067 ( .A(n31885), .Y(n18876) );
  BUFx6f_ASAP7_75t_SL U25068 ( .A(n32736), .Y(n24645) );
  BUFx6f_ASAP7_75t_SL U25069 ( .A(n31042), .Y(n22400) );
  OAI22xp33_ASAP7_75t_SRAM U25070 ( .A1(n32361), .A2(n24637), .B1(n32365), 
        .B2(n22383), .Y(n27248) );
  NAND2x1p5_ASAP7_75t_SL U25071 ( .A(n3055), .B(n30189), .Y(n30166) );
  NOR2x2_ASAP7_75t_SL U25072 ( .A(ahb0_v_HREADY_), .B(n24699), .Y(n32705) );
  AOI21xp5_ASAP7_75t_SL U25073 ( .A1(u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__1_), 
        .A2(n30017), .B(n25017), .Y(n25439) );
  NOR2x1_ASAP7_75t_SL U25074 ( .A(mult_x_1196_n651), .B(mult_x_1196_n654), .Y(
        n23451) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25075 ( .A1(n31585), .A2(n31263), .B(n31574), 
        .C(n31568), .Y(n31613) );
  OAI21x1_ASAP7_75t_SL U25076 ( .A1(n25073), .A2(n25072), .B(n25447), .Y(
        n30578) );
  OAI21x1_ASAP7_75t_SL U25077 ( .A1(n25071), .A2(n29912), .B(n25070), .Y(
        n25447) );
  INVx3_ASAP7_75t_SL U25078 ( .A(n23894), .Y(n18877) );
  INVx3_ASAP7_75t_SL U25079 ( .A(n23894), .Y(n31633) );
  AND2x2_ASAP7_75t_SL U25080 ( .A(n25592), .B(n18878), .Y(n32731) );
  AND2x2_ASAP7_75t_SL U25081 ( .A(n32022), .B(n18879), .Y(n18878) );
  INVxp33_ASAP7_75t_SRAM U25082 ( .A(n30507), .Y(n18879) );
  BUFx3_ASAP7_75t_SL U25083 ( .A(add_x_746_n1), .Y(n18880) );
  HB1xp67_ASAP7_75t_SL U25084 ( .A(n24347), .Y(n18881) );
  HB1xp67_ASAP7_75t_SL U25085 ( .A(timer0_res_31_), .Y(n18882) );
  NOR2x1p5_ASAP7_75t_SL U25086 ( .A(n22380), .B(n30166), .Y(n30182) );
  NAND2x1_ASAP7_75t_SL U25087 ( .A(n25592), .B(n32022), .Y(n18883) );
  XNOR2x2_ASAP7_75t_SL U25088 ( .A(add_x_746_n78), .B(n18880), .Y(
        u0_0_leon3x0_p0_iu_fe_npc_18_) );
  NOR2x1p5_ASAP7_75t_SL U25089 ( .A(n32079), .B(n24877), .Y(n24998) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25090 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), .A2(n24878), .B(n31858), .C(
        n24998), .Y(n24771) );
  AND3x1_ASAP7_75t_SL U25091 ( .A(n24999), .B(n24998), .C(n25226), .Y(n25000)
         );
  NOR2x1_ASAP7_75t_SL U25092 ( .A(n24766), .B(n32168), .Y(n32165) );
  INVx1_ASAP7_75t_SL U25093 ( .A(n23830), .Y(n18884) );
  NOR4xp75_ASAP7_75t_SL U25094 ( .A(u0_0_leon3x0_p0_dci[29]), .B(
        u0_0_leon3x0_p0_dci[28]), .C(u0_0_leon3x0_p0_dci[27]), .D(
        u0_0_leon3x0_p0_dci[30]), .Y(n25355) );
  NAND2x1_ASAP7_75t_SL U25095 ( .A(n26466), .B(timer0_res_31_), .Y(n26470) );
  INVx8_ASAP7_75t_SL U25096 ( .A(n18911), .Y(n24686) );
  AOI22xp33_ASAP7_75t_SRAM U25097 ( .A1(n31824), .A2(n29729), .B1(n31828), 
        .B2(u0_0_leon3x0_p0_dci[14]), .Y(n26200) );
  NOR2x1p5_ASAP7_75t_SL U25098 ( .A(u0_0_leon3x0_p0_dci[15]), .B(
        u0_0_leon3x0_p0_dci[14]), .Y(n25345) );
  AOI21xp5_ASAP7_75t_SL U25099 ( .A1(n18886), .A2(add_x_735_n230), .B(
        add_x_735_n231), .Y(add_x_735_n229) );
  AOI21x1_ASAP7_75t_SL U25100 ( .A1(add_x_735_n223), .A2(n18886), .B(
        add_x_735_n224), .Y(add_x_735_n222) );
  INVxp33_ASAP7_75t_SRAM U25101 ( .A(add_x_735_n247), .Y(add_x_735_n298) );
  XOR2x1_ASAP7_75t_SL U25102 ( .A(add_x_735_n26), .B(add_x_735_n229), .Y(
        u0_0_leon3x0_p0_dci[14]) );
  INVxp33_ASAP7_75t_SRAM U25103 ( .A(add_x_735_n299), .Y(n18885) );
  OAI21xp5_ASAP7_75t_SL U25104 ( .A1(n18997), .A2(n23229), .B(n31871), .Y(
        n2818) );
  NAND2x1_ASAP7_75t_SL U25105 ( .A(n18997), .B(n25081), .Y(n26351) );
  OAI21x1_ASAP7_75t_SL U25106 ( .A1(n22228), .A2(add_x_735_n39), .B(
        add_x_735_n40), .Y(add_x_735_n38) );
  XNOR2x1_ASAP7_75t_SL U25107 ( .A(add_x_735_n4), .B(add_x_735_n38), .Y(
        u0_0_leon3x0_p0_dci[36]) );
  AO21x2_ASAP7_75t_SL U25108 ( .A1(add_x_735_n253), .A2(add_x_735_n245), .B(
        add_x_735_n246), .Y(n18886) );
  BUFx16f_ASAP7_75t_SL U25109 ( .A(n32731), .Y(n22381) );
  INVx1_ASAP7_75t_SL U25110 ( .A(u0_0_leon3x0_p0_dci[10]), .Y(n25342) );
  INVxp33_ASAP7_75t_SRAM U25111 ( .A(u0_0_leon3x0_p0_dci[35]), .Y(n31991) );
  NOR4xp75_ASAP7_75t_SL U25112 ( .A(u0_0_leon3x0_p0_dci[25]), .B(
        u0_0_leon3x0_p0_dci[34]), .C(u0_0_leon3x0_p0_dci[35]), .D(
        u0_0_leon3x0_p0_dci[31]), .Y(n25354) );
  AOI21xp5_ASAP7_75t_SL U25113 ( .A1(add_x_735_n2), .A2(add_x_735_n61), .B(
        add_x_735_n62), .Y(add_x_735_n60) );
  HB1xp67_ASAP7_75t_SL U25114 ( .A(u0_0_leon3x0_p0_dci[13]), .Y(n18887) );
  XOR2xp5_ASAP7_75t_SL U25115 ( .A(add_x_735_n27), .B(add_x_735_n238), .Y(
        u0_0_leon3x0_p0_dci[13]) );
  NOR2xp33_ASAP7_75t_SL U25116 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[9]), .Y(
        n27139) );
  NOR2x1_ASAP7_75t_SL U25117 ( .A(n22837), .B(u0_0_leon3x0_p0_divi[9]), .Y(
        add_x_735_n220) );
  INVx1_ASAP7_75t_SL U25118 ( .A(n25516), .Y(n25517) );
  NOR2x1p5_ASAP7_75t_SL U25119 ( .A(n24462), .B(n27138), .Y(
        u0_0_leon3x0_p0_divi[9]) );
  OAI21xp5_ASAP7_75t_SL U25120 ( .A1(add_x_735_n81), .A2(add_x_735_n116), .B(
        add_x_735_n82), .Y(add_x_735_n2) );
  NOR2x1_ASAP7_75t_SL U25121 ( .A(add_x_735_n209), .B(add_x_735_n212), .Y(
        add_x_735_n203) );
  NOR2x1_ASAP7_75t_SL U25122 ( .A(n22721), .B(u0_0_leon3x0_p0_divi[11]), .Y(
        add_x_735_n209) );
  NOR2x1_ASAP7_75t_SL U25123 ( .A(add_x_735_n198), .B(add_x_735_n191), .Y(
        add_x_735_n189) );
  NAND2xp5_ASAP7_75t_SL U25124 ( .A(add_x_735_n99), .B(add_x_735_n117), .Y(
        add_x_735_n97) );
  NOR2x1_ASAP7_75t_SL U25125 ( .A(add_x_735_n112), .B(add_x_735_n105), .Y(
        add_x_735_n99) );
  NAND2xp5_ASAP7_75t_SL U25126 ( .A(add_x_735_n90), .B(add_x_735_n117), .Y(
        add_x_735_n88) );
  NOR2x1p5_ASAP7_75t_SL U25127 ( .A(n24467), .B(n25891), .Y(
        u0_0_leon3x0_p0_divi[28]) );
  NAND2xp5_ASAP7_75t_SL U25128 ( .A(n18588), .B(u0_0_leon3x0_p0_divi[6]), .Y(
        add_x_735_n242) );
  NOR2x1p5_ASAP7_75t_SL U25129 ( .A(n24465), .B(n26416), .Y(
        u0_0_leon3x0_p0_divi[22]) );
  INVx1_ASAP7_75t_SL U25130 ( .A(add_x_735_n287), .Y(n18888) );
  INVx1_ASAP7_75t_SL U25131 ( .A(add_x_735_n160), .Y(add_x_735_n287) );
  OAI21x1_ASAP7_75t_SL U25132 ( .A1(n18895), .A2(add_x_735_n236), .B(
        add_x_735_n237), .Y(add_x_735_n231) );
  AOI21xp5_ASAP7_75t_SL U25133 ( .A1(add_x_735_n231), .A2(add_x_735_n218), .B(
        add_x_735_n219), .Y(add_x_735_n217) );
  NOR2x1_ASAP7_75t_SL U25134 ( .A(n23964), .B(u0_0_leon3x0_p0_divi[14]), .Y(
        add_x_735_n180) );
  INVx1_ASAP7_75t_SL U25135 ( .A(add_x_735_n180), .Y(add_x_735_n289) );
  AOI22xp33_ASAP7_75t_SRAM U25136 ( .A1(u0_0_leon3x0_p0_divi[14]), .A2(n27200), 
        .B1(n28830), .B2(n26567), .Y(n26568) );
  INVxp33_ASAP7_75t_SRAM U25137 ( .A(u0_0_leon3x0_p0_divi[14]), .Y(n26565) );
  HB1xp67_ASAP7_75t_SL U25138 ( .A(add_x_735_n145), .Y(n18889) );
  BUFx3_ASAP7_75t_SL U25139 ( .A(u0_0_leon3x0_p0_divi[8]), .Y(n18890) );
  NOR2xp33_ASAP7_75t_SL U25140 ( .A(n27112), .B(n27111), .Y(
        u0_0_leon3x0_p0_divi[8]) );
  NOR2x1p5_ASAP7_75t_SL U25141 ( .A(n24461), .B(n26703), .Y(
        u0_0_leon3x0_p0_divi[16]) );
  NOR2x1_ASAP7_75t_SL U25142 ( .A(n23154), .B(u0_0_leon3x0_p0_divi[13]), .Y(
        add_x_735_n191) );
  NOR2x1p5_ASAP7_75t_SL U25143 ( .A(n24459), .B(n27193), .Y(
        u0_0_leon3x0_p0_divi[13]) );
  OAI21xp5_ASAP7_75t_SL U25144 ( .A1(n18889), .A2(add_x_735_n141), .B(
        add_x_735_n142), .Y(add_x_735_n136) );
  NOR4xp75_ASAP7_75t_SL U25145 ( .A(u0_0_leon3x0_p0_dci[33]), .B(
        u0_0_leon3x0_p0_dci[36]), .C(u0_0_leon3x0_p0_dci[24]), .D(
        u0_0_leon3x0_p0_dci[21]), .Y(n25353) );
  NAND2xp5_ASAP7_75t_SL U25146 ( .A(n23396), .B(u0_0_leon3x0_p0_divi[12]), .Y(
        add_x_735_n199) );
  OR2x2_ASAP7_75t_SL U25147 ( .A(n23548), .B(n24689), .Y(n18891) );
  INVx8_ASAP7_75t_SL U25148 ( .A(n18891), .Y(n28769) );
  NOR4xp75_ASAP7_75t_SL U25149 ( .A(n32438), .B(u0_0_leon3x0_p0_dci[9]), .C(
        u0_0_leon3x0_p0_dci[6]), .D(u0_0_leon3x0_p0_dci[7]), .Y(n25341) );
  NAND2xp5_ASAP7_75t_SL U25150 ( .A(n18884), .B(n25088), .Y(n28820) );
  XNOR2x2_ASAP7_75t_SL U25151 ( .A(add_x_735_n28), .B(n18886), .Y(
        u0_0_leon3x0_p0_dci[12]) );
  NAND2xp5_ASAP7_75t_SL U25152 ( .A(u0_0_leon3x0_p0_iu_fe_pc_18_), .B(n18880), 
        .Y(add_x_746_n76) );
  NAND2xp5_ASAP7_75t_SL U25153 ( .A(add_x_746_n58), .B(n18880), .Y(
        add_x_746_n57) );
  NOR2x1_ASAP7_75t_SL U25154 ( .A(n24468), .B(n28381), .Y(
        u0_0_leon3x0_p0_divi[29]) );
  HB1xp67_ASAP7_75t_SL U25155 ( .A(add_x_735_n268), .Y(n18892) );
  NOR3x1_ASAP7_75t_SL U25156 ( .A(n24349), .B(timer0_N71), .C(timer0_N72), .Y(
        n24353) );
  XNOR2x1_ASAP7_75t_SL U25157 ( .A(n2307), .B(n31419), .Y(n29114) );
  INVx1_ASAP7_75t_SL U25158 ( .A(n31419), .Y(n21549) );
  HB1xp67_ASAP7_75t_SL U25159 ( .A(add_x_735_n256), .Y(n18893) );
  AOI21xp5_ASAP7_75t_SL U25160 ( .A1(add_x_735_n253), .A2(add_x_735_n245), .B(
        add_x_735_n246), .Y(n18894) );
  NAND2xp5_ASAP7_75t_SL U25161 ( .A(u0_0_leon3x0_p0_div0_vaddin1[9]), .B(
        u0_0_leon3x0_p0_div0_b[9]), .Y(DP_OP_5187J1_124_3275_n256) );
  INVx1_ASAP7_75t_SL U25162 ( .A(DP_OP_5187J1_124_3275_n230), .Y(
        DP_OP_5187J1_124_3275_n232) );
  NAND2x1p5_ASAP7_75t_SL U25163 ( .A(n28977), .B(n26298), .Y(n28869) );
  NOR2x1_ASAP7_75t_SL U25164 ( .A(n22378), .B(n29013), .Y(n30489) );
  INVx1_ASAP7_75t_SL U25165 ( .A(u0_0_leon3x0_p0_dci[8]), .Y(n25340) );
  INVx3_ASAP7_75t_SL U25166 ( .A(add_x_735_n215), .Y(add_x_735_n214) );
  BUFx6f_ASAP7_75t_SL U25167 ( .A(n31039), .Y(n22383) );
  OAI21x1_ASAP7_75t_SL U25168 ( .A1(n31460), .A2(n32274), .B(n25410), .Y(
        n31039) );
  NAND3x1_ASAP7_75t_SL U25169 ( .A(n25342), .B(n25340), .C(n25341), .Y(n25343)
         );
  NOR2x1_ASAP7_75t_SL U25170 ( .A(add_x_735_n81), .B(add_x_735_n115), .Y(
        add_x_735_n3) );
  NAND2xp5_ASAP7_75t_SL U25171 ( .A(add_x_735_n52), .B(add_x_735_n3), .Y(
        add_x_735_n50) );
  NAND2xp5_ASAP7_75t_SL U25172 ( .A(add_x_735_n61), .B(add_x_735_n3), .Y(
        add_x_735_n59) );
  NAND2xp5_ASAP7_75t_SL U25173 ( .A(add_x_735_n72), .B(add_x_735_n3), .Y(
        add_x_735_n70) );
  NOR2x1p5_ASAP7_75t_SL U25174 ( .A(n26564), .B(n26563), .Y(
        u0_0_leon3x0_p0_divi[14]) );
  BUFx2_ASAP7_75t_SL U25175 ( .A(add_x_735_n242), .Y(n18895) );
  OA21x2_ASAP7_75t_SL U25176 ( .A1(n18895), .A2(add_x_735_n236), .B(
        add_x_735_n237), .Y(n18896) );
  NOR2x1_ASAP7_75t_SL U25177 ( .A(n24479), .B(n25245), .Y(n31629) );
  NAND2x1p5_ASAP7_75t_SL U25178 ( .A(n32705), .B(n31734), .Y(n32786) );
  AOI21x1_ASAP7_75t_SL U25179 ( .A1(n24583), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[63]), .B(n25252), .Y(n31734) );
  NOR2x1_ASAP7_75t_SL U25180 ( .A(n25439), .B(n31364), .Y(n28411) );
  OR2x6_ASAP7_75t_SL U25181 ( .A(n30208), .B(n25018), .Y(n31364) );
  AO21x2_ASAP7_75t_SL U25182 ( .A1(n22607), .A2(n23325), .B(n22606), .Y(
        mult_x_1196_n2024) );
  NAND2x1p5_ASAP7_75t_SL U25183 ( .A(n24271), .B(n22319), .Y(n23183) );
  NAND2xp5_ASAP7_75t_SL U25184 ( .A(n18897), .B(n24689), .Y(n22220) );
  BUFx2_ASAP7_75t_SL U25185 ( .A(n24688), .Y(n18997) );
  INVx1_ASAP7_75t_SL U25186 ( .A(n18882), .Y(n20910) );
  BUFx12f_ASAP7_75t_SL U25187 ( .A(n32684), .Y(n22405) );
  NAND2x1_ASAP7_75t_SL U25188 ( .A(n24684), .B(n31934), .Y(n32684) );
  AOI22xp33_ASAP7_75t_SRAM U25189 ( .A1(n31824), .A2(n29731), .B1(n31828), 
        .B2(u0_0_leon3x0_p0_dci[16]), .Y(n28659) );
  NOR2x1p5_ASAP7_75t_SL U25190 ( .A(n31461), .B(n25516), .Y(n30509) );
  NOR2x1_ASAP7_75t_SL U25191 ( .A(u0_0_leon3x0_p0_div0_vaddin1[6]), .B(
        u0_0_leon3x0_p0_div0_b[6]), .Y(DP_OP_5187J1_124_3275_n271) );
  NAND2x1p5_ASAP7_75t_SL U25192 ( .A(u0_0_leon3x0_p0_divi[30]), .B(n22919), 
        .Y(n31419) );
  NAND2xp5_ASAP7_75t_SL U25193 ( .A(u0_0_leon3x0_p0_div0_vaddin1[6]), .B(
        u0_0_leon3x0_p0_div0_b[6]), .Y(DP_OP_5187J1_124_3275_n274) );
  NOR2x1_ASAP7_75t_SL U25194 ( .A(n23858), .B(n26920), .Y(
        u0_0_leon3x0_p0_divi[27]) );
  NOR2xp33_ASAP7_75t_SL U25195 ( .A(n24048), .B(n28769), .Y(n23858) );
  NOR2x1_ASAP7_75t_SL U25196 ( .A(add_x_735_n74), .B(add_x_735_n67), .Y(
        add_x_735_n61) );
  NOR2x1_ASAP7_75t_SL U25197 ( .A(add_x_735_A_29_), .B(
        u0_0_leon3x0_p0_divi[27]), .Y(add_x_735_n67) );
  OR2x2_ASAP7_75t_SL U25198 ( .A(add_x_735_n180), .B(add_x_735_n173), .Y(
        n18898) );
  INVx6_ASAP7_75t_SL U25199 ( .A(n18898), .Y(add_x_735_n167) );
  NAND3x2_ASAP7_75t_SL U25200 ( .A(n24998), .B(n18842), .C(n25226), .Y(n31862)
         );
  NOR2x1p5_ASAP7_75t_SL U25201 ( .A(n4928), .B(n18867), .Y(
        DP_OP_1196_128_7433_n453) );
  HB1xp67_ASAP7_75t_SL U25202 ( .A(n23929), .Y(n18899) );
  AOI21xp5_ASAP7_75t_SL U25203 ( .A1(n18886), .A2(add_x_735_n297), .B(
        add_x_735_n240), .Y(add_x_735_n238) );
  INVx1_ASAP7_75t_SL U25204 ( .A(add_x_735_n262), .Y(n21259) );
  NOR2x1_ASAP7_75t_SL U25205 ( .A(u0_0_leon3x0_p0_divi[1]), .B(n22939), .Y(
        add_x_735_n262) );
  OAI21xp5_ASAP7_75t_SL U25206 ( .A1(n30913), .A2(n22405), .B(n30912), .Y(
        u0_0_leon3x0_p0_c0mmu_icache0_v_WADDRESS__2_) );
  INVx13_ASAP7_75t_SL U25207 ( .A(n22405), .Y(n22385) );
  BUFx6f_ASAP7_75t_SL U25208 ( .A(n29019), .Y(n24630) );
  NOR2x1_ASAP7_75t_SL U25209 ( .A(u0_0_leon3x0_p0_divi[2]), .B(n18393), .Y(
        add_x_735_n259) );
  NOR2x2_ASAP7_75t_SL U25210 ( .A(n24432), .B(n28677), .Y(
        u0_0_leon3x0_p0_divi[10]) );
  NOR2x1_ASAP7_75t_SL U25211 ( .A(n23091), .B(u0_0_leon3x0_p0_divi[10]), .Y(
        add_x_735_n212) );
  INVx5_ASAP7_75t_SL U25212 ( .A(n22403), .Y(n22384) );
  OAI21x1_ASAP7_75t_SL U25213 ( .A1(add_x_735_n266), .A2(add_x_735_n268), .B(
        add_x_735_n267), .Y(add_x_735_n265) );
  INVx4_ASAP7_75t_SL U25214 ( .A(n32059), .Y(n22403) );
  NOR4xp75_ASAP7_75t_SL U25215 ( .A(u0_0_leon3x0_p0_dci[13]), .B(n25343), .C(
        u0_0_leon3x0_p0_dci[11]), .D(u0_0_leon3x0_p0_dci[12]), .Y(n25346) );
  AOI22xp33_ASAP7_75t_SRAM U25216 ( .A1(n31824), .A2(n30709), .B1(n31828), 
        .B2(n18887), .Y(n30710) );
  NOR2x1_ASAP7_75t_SL U25217 ( .A(DP_OP_5187J1_124_3275_n219), .B(
        DP_OP_5187J1_124_3275_n226), .Y(DP_OP_5187J1_124_3275_n213) );
  NOR2x1_ASAP7_75t_SL U25218 ( .A(u0_0_leon3x0_p0_div0_vaddin1[13]), .B(
        u0_0_leon3x0_p0_div0_b[13]), .Y(DP_OP_5187J1_124_3275_n219) );
  NAND4xp75_ASAP7_75t_SL U25219 ( .A(n25935), .B(n25934), .C(n25933), .D(
        n25932), .Y(n28377) );
  NOR3x1_ASAP7_75t_SL U25220 ( .A(n25931), .B(u0_0_leon3x0_p0_div0_addout_31_), 
        .C(n25930), .Y(n25935) );
  NOR2x1_ASAP7_75t_SL U25221 ( .A(u0_0_leon3x0_p0_div0_vaddin1[5]), .B(
        u0_0_leon3x0_p0_div0_b[5]), .Y(DP_OP_5187J1_124_3275_n282) );
  HB1xp67_ASAP7_75t_SL U25222 ( .A(n23504), .Y(n22775) );
  NOR2x2_ASAP7_75t_SL U25223 ( .A(n26205), .B(n26204), .Y(n31833) );
  AOI21x1_ASAP7_75t_SL U25224 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_5_), .A2(n31833), 
        .B(n29679), .Y(n32568) );
  NOR2x1_ASAP7_75t_SL U25225 ( .A(n5061), .B(n2842), .Y(timer0_N89) );
  INVxp33_ASAP7_75t_SRAM U25226 ( .A(n32030), .Y(n18902) );
  INVxp33_ASAP7_75t_SRAM U25227 ( .A(n18902), .Y(n18903) );
  XOR2x2_ASAP7_75t_SL U25228 ( .A(add_x_735_n25), .B(add_x_735_n222), .Y(
        u0_0_leon3x0_p0_dci[15]) );
  BUFx2_ASAP7_75t_SL U25229 ( .A(u0_0_leon3x0_p0_divi[7]), .Y(n18904) );
  BUFx12f_ASAP7_75t_SL U25230 ( .A(u0_0_leon3x0_p0_muli[26]), .Y(n24058) );
  XNOR2xp5_ASAP7_75t_SL U25231 ( .A(n24058), .B(n23967), .Y(mult_x_1196_n2955)
         );
  XNOR2xp5_ASAP7_75t_SL U25232 ( .A(n24058), .B(n23955), .Y(mult_x_1196_n3227)
         );
  XNOR2xp5_ASAP7_75t_SL U25233 ( .A(n23969), .B(n24058), .Y(mult_x_1196_n2921)
         );
  BUFx16f_ASAP7_75t_SL U25234 ( .A(n32062), .Y(n22402) );
  NAND2x1p5_ASAP7_75t_SL U25235 ( .A(n32689), .B(n22403), .Y(n32062) );
  NAND2x1_ASAP7_75t_SL U25236 ( .A(u0_0_leon3x0_p0_div0_vaddin1[8]), .B(
        u0_0_leon3x0_p0_div0_b[8]), .Y(DP_OP_5187J1_124_3275_n259) );
  OAI21x1_ASAP7_75t_SL U25237 ( .A1(DP_OP_5187J1_124_3275_n259), .A2(
        DP_OP_5187J1_124_3275_n255), .B(DP_OP_5187J1_124_3275_n256), .Y(
        DP_OP_5187J1_124_3275_n250) );
  OR2x2_ASAP7_75t_SL U25238 ( .A(mult_x_1196_n1580), .B(mult_x_1196_n1544), 
        .Y(mult_x_1196_n603) );
  AOI22xp33_ASAP7_75t_SRAM U25239 ( .A1(n31824), .A2(n29739), .B1(
        u0_0_leon3x0_p0_dci[15]), .B2(n31828), .Y(n28702) );
  AOI21xp33_ASAP7_75t_SRAM U25240 ( .A1(n18904), .A2(n24580), .B(n28722), .Y(
        n28723) );
  NOR2x1_ASAP7_75t_SL U25241 ( .A(DP_OP_5187J1_124_3275_n266), .B(
        DP_OP_5187J1_124_3275_n271), .Y(DP_OP_5187J1_124_3275_n264) );
  NOR2x1_ASAP7_75t_SL U25242 ( .A(n24002), .B(mult_x_1196_n3108), .Y(n23599)
         );
  INVx1_ASAP7_75t_SL U25243 ( .A(mult_x_1196_n1268), .Y(n24191) );
  BUFx6f_ASAP7_75t_SL U25244 ( .A(n31040), .Y(n24637) );
  NOR2x1_ASAP7_75t_SL U25245 ( .A(n4929), .B(n32095), .Y(
        DP_OP_1196_128_7433_n454) );
  NOR2x2_ASAP7_75t_SL U25246 ( .A(n25572), .B(n18828), .Y(n32059) );
  INVx1_ASAP7_75t_SL U25247 ( .A(mult_x_1196_n1053), .Y(n18905) );
  INVx2_ASAP7_75t_SL U25248 ( .A(n18905), .Y(n18906) );
  HB1xp67_ASAP7_75t_SL U25249 ( .A(mult_x_1196_n1046), .Y(n18907) );
  NAND2xp5_ASAP7_75t_SL U25250 ( .A(add_x_735_n251), .B(add_x_735_n299), .Y(
        add_x_735_n30) );
  NAND2xp5_ASAP7_75t_SL U25251 ( .A(n23958), .B(u0_0_leon3x0_p0_divi[4]), .Y(
        add_x_735_n251) );
  XNOR2x2_ASAP7_75t_SL U25252 ( .A(mult_x_1196_n1794), .B(n23532), .Y(
        mult_x_1196_n1760) );
  NAND2xp5_ASAP7_75t_SL U25253 ( .A(n18569), .B(n26351), .Y(n18908) );
  NAND2xp5_ASAP7_75t_SL U25254 ( .A(n18569), .B(n26351), .Y(n18909) );
  BUFx6f_ASAP7_75t_SL U25255 ( .A(u0_0_leon3x0_p0_iu_r_E__LDBP1_), .Y(n18910)
         );
  BUFx6f_ASAP7_75t_SL U25256 ( .A(u0_0_leon3x0_p0_iu_r_E__LDBP1_), .Y(n18911)
         );
  XNOR2xp5_ASAP7_75t_SL U25257 ( .A(mult_x_1196_n1627), .B(mult_x_1196_n1597), 
        .Y(n22857) );
  OAI22xp5_ASAP7_75t_SL U25258 ( .A1(mult_x_1196_n3278), .A2(n18319), .B1(
        n23980), .B2(mult_x_1196_n3277), .Y(mult_x_1196_n2702) );
  HB1xp67_ASAP7_75t_SL U25259 ( .A(mult_x_1196_n1696), .Y(n18912) );
  INVx3_ASAP7_75t_SL U25260 ( .A(n24550), .Y(n23375) );
  XOR2x2_ASAP7_75t_SL U25261 ( .A(n23264), .B(mult_x_1196_n1918), .Y(n22211)
         );
  AOI22xp33_ASAP7_75t_SRAM U25262 ( .A1(n30622), .A2(n18908), .B1(
        u0_0_leon3x0_p0_iu_r_E__CWP__1_), .B2(n30621), .Y(n30623) );
  INVx1_ASAP7_75t_SL U25263 ( .A(n21758), .Y(n18914) );
  OAI21xp5_ASAP7_75t_SL U25264 ( .A1(mult_x_1196_n547), .A2(mult_x_1196_n539), 
        .B(mult_x_1196_n540), .Y(mult_x_1196_n534) );
  BUFx2_ASAP7_75t_SL U25265 ( .A(mult_x_1196_n1494), .Y(n18915) );
  BUFx2_ASAP7_75t_SL U25266 ( .A(mult_x_1196_n1806), .Y(n18916) );
  OAI22xp5_ASAP7_75t_SL U25267 ( .A1(n23997), .A2(mult_x_1196_n3144), .B1(
        n22578), .B2(n23999), .Y(mult_x_1196_n2139) );
  XOR2xp5_ASAP7_75t_SL U25268 ( .A(mult_x_1196_n1727), .B(n18917), .Y(n24295)
         );
  XNOR2xp5_ASAP7_75t_SL U25269 ( .A(n24226), .B(mult_x_1196_n1690), .Y(n18917)
         );
  INVx2_ASAP7_75t_SL U25270 ( .A(mult_x_1196_n1686), .Y(n23448) );
  OR2x6_ASAP7_75t_SL U25271 ( .A(n18993), .B(n22965), .Y(n18919) );
  OR2x6_ASAP7_75t_SL U25272 ( .A(n22965), .B(n18993), .Y(n18920) );
  HB1xp67_ASAP7_75t_SL U25273 ( .A(mult_x_1196_n550), .Y(n18921) );
  NAND2x1p5_ASAP7_75t_SL U25274 ( .A(n23808), .B(n23754), .Y(mult_x_1196_n1596) );
  INVxp33_ASAP7_75t_SRAM U25275 ( .A(mult_x_1196_n677), .Y(n18922) );
  INVx1_ASAP7_75t_SL U25276 ( .A(n18922), .Y(n18923) );
  XOR2x2_ASAP7_75t_SL U25277 ( .A(mult_x_1196_n1944), .B(n23806), .Y(n22324)
         );
  XNOR2xp5_ASAP7_75t_SL U25278 ( .A(mult_x_1196_n1955), .B(n22324), .Y(n23019)
         );
  MAJIxp5_ASAP7_75t_SL U25279 ( .A(n23860), .B(n18916), .C(n23859), .Y(n18924)
         );
  HB1xp67_ASAP7_75t_SL U25280 ( .A(mult_x_1196_n1747), .Y(n18925) );
  INVx2_ASAP7_75t_SL U25281 ( .A(n23862), .Y(n23859) );
  HB1xp67_ASAP7_75t_SL U25282 ( .A(mult_x_1196_n1991), .Y(n23934) );
  BUFx3_ASAP7_75t_SL U25283 ( .A(n23953), .Y(n18926) );
  BUFx16f_ASAP7_75t_SL U25284 ( .A(n23953), .Y(n18927) );
  INVx2_ASAP7_75t_SL U25285 ( .A(n23951), .Y(n23953) );
  BUFx2_ASAP7_75t_SL U25286 ( .A(mult_x_1196_n1771), .Y(n18928) );
  NAND2xp33_ASAP7_75t_SRAM U25287 ( .A(n18928), .B(mult_x_1196_n1745), .Y(
        n18929) );
  HB1xp67_ASAP7_75t_SL U25288 ( .A(mult_x_1196_n1976), .Y(n18930) );
  HB1xp67_ASAP7_75t_SL U25289 ( .A(mult_x_1196_n1203), .Y(n18931) );
  OAI21x1_ASAP7_75t_SL U25290 ( .A1(mult_x_1196_n470), .A2(mult_x_1196_n496), 
        .B(n22467), .Y(n18932) );
  MAJIxp5_ASAP7_75t_SL U25291 ( .A(mult_x_1196_n1570), .B(mult_x_1196_n1572), 
        .C(n24284), .Y(n18933) );
  HB1xp67_ASAP7_75t_SL U25292 ( .A(mult_x_1196_n1955), .Y(n18935) );
  XNOR2x2_ASAP7_75t_SL U25293 ( .A(n18933), .B(mult_x_1196_n1525), .Y(n18968)
         );
  BUFx2_ASAP7_75t_SL U25294 ( .A(mult_x_1196_n1813), .Y(n18936) );
  XNOR2x1_ASAP7_75t_SL U25295 ( .A(n22423), .B(n22424), .Y(mult_x_1196_n3317)
         );
  OAI22x1_ASAP7_75t_SL U25296 ( .A1(n24007), .A2(mult_x_1196_n3071), .B1(
        n24005), .B2(mult_x_1196_n3070), .Y(n23199) );
  INVx5_ASAP7_75t_SL U25297 ( .A(n22206), .Y(n23959) );
  INVx2_ASAP7_75t_SL U25298 ( .A(n23779), .Y(n23778) );
  HB1xp67_ASAP7_75t_SL U25299 ( .A(n22335), .Y(n18937) );
  XOR2xp5_ASAP7_75t_SL U25300 ( .A(n23868), .B(n23869), .Y(mult_x_1196_n1672)
         );
  XNOR2x1_ASAP7_75t_SL U25301 ( .A(n23861), .B(n22772), .Y(mult_x_1196_n1777)
         );
  XNOR2x1_ASAP7_75t_SL U25302 ( .A(n23012), .B(n18938), .Y(n18939) );
  INVx2_ASAP7_75t_SL U25303 ( .A(n23011), .Y(n18938) );
  MAJIxp5_ASAP7_75t_SL U25304 ( .A(n18939), .B(n22885), .C(n22697), .Y(
        mult_x_1196_n1820) );
  NOR2xp33_ASAP7_75t_SL U25305 ( .A(n18940), .B(mult_x_1196_n1790), .Y(n22323)
         );
  INVxp67_ASAP7_75t_SL U25306 ( .A(n23533), .Y(n18940) );
  XNOR2xp5_ASAP7_75t_SL U25307 ( .A(n23533), .B(mult_x_1196_n1790), .Y(n23532)
         );
  INVx1_ASAP7_75t_SL U25308 ( .A(n22758), .Y(n22842) );
  INVx1_ASAP7_75t_SL U25309 ( .A(DP_OP_5187J1_124_3275_n229), .Y(
        DP_OP_5187J1_124_3275_n231) );
  NOR2x1_ASAP7_75t_SL U25310 ( .A(DP_OP_5187J1_124_3275_n255), .B(
        DP_OP_5187J1_124_3275_n258), .Y(DP_OP_5187J1_124_3275_n249) );
  NOR2x1_ASAP7_75t_SL U25311 ( .A(u0_0_leon3x0_p0_div0_vaddin1[8]), .B(
        u0_0_leon3x0_p0_div0_b[8]), .Y(DP_OP_5187J1_124_3275_n258) );
  NOR2x1_ASAP7_75t_SL U25312 ( .A(u0_0_leon3x0_p0_div0_vaddin1[9]), .B(
        u0_0_leon3x0_p0_div0_b[9]), .Y(DP_OP_5187J1_124_3275_n255) );
  INVx1_ASAP7_75t_SL U25313 ( .A(n24214), .Y(n18941) );
  NAND2xp5_ASAP7_75t_SL U25314 ( .A(n18946), .B(n18942), .Y(n22537) );
  OAI21xp5_ASAP7_75t_SL U25315 ( .A1(mult_x_1196_n2363), .A2(n23380), .B(
        n18943), .Y(n18942) );
  INVx1_ASAP7_75t_SL U25316 ( .A(n23379), .Y(n18943) );
  NOR2x1_ASAP7_75t_SL U25317 ( .A(n24008), .B(mult_x_1196_n3030), .Y(n18944)
         );
  NOR2x1_ASAP7_75t_SL U25318 ( .A(mult_x_1196_n3031), .B(n24009), .Y(n18945)
         );
  NAND2xp5_ASAP7_75t_SL U25319 ( .A(mult_x_1196_n2363), .B(n23380), .Y(n18946)
         );
  XOR2xp5_ASAP7_75t_SL U25320 ( .A(n18948), .B(mult_x_1196_n2009), .Y(n22478)
         );
  NAND2xp5_ASAP7_75t_SL U25321 ( .A(n18949), .B(n18947), .Y(n22332) );
  OAI21xp5_ASAP7_75t_SL U25322 ( .A1(n22635), .A2(mult_x_1196_n2006), .B(
        n18948), .Y(n18947) );
  MAJIxp5_ASAP7_75t_SL U25323 ( .A(mult_x_1196_n2029), .B(mult_x_1196_n2027), 
        .C(n22821), .Y(n18948) );
  NAND2xp5_ASAP7_75t_SL U25324 ( .A(n22635), .B(mult_x_1196_n2006), .Y(n18949)
         );
  INVx1_ASAP7_75t_SL U25325 ( .A(n22671), .Y(n22669) );
  XNOR2xp5_ASAP7_75t_SL U25326 ( .A(n18951), .B(n18950), .Y(n22671) );
  INVx1_ASAP7_75t_SL U25327 ( .A(mult_x_1196_n1677), .Y(n18951) );
  NAND2xp5_ASAP7_75t_SL U25328 ( .A(n18953), .B(n23026), .Y(n23024) );
  INVx1_ASAP7_75t_SL U25329 ( .A(n23761), .Y(n18952) );
  NAND2xp5_ASAP7_75t_SL U25330 ( .A(mult_x_1196_n1912), .B(mult_x_1196_n1937), 
        .Y(n18953) );
  MAJIxp5_ASAP7_75t_SL U25331 ( .A(mult_x_1196_n1936), .B(mult_x_1196_n1946), 
        .C(mult_x_1196_n1944), .Y(mult_x_1196_n1937) );
  XOR2xp5_ASAP7_75t_SL U25332 ( .A(n18954), .B(n23579), .Y(mult_x_1196_n1944)
         );
  INVx1_ASAP7_75t_SL U25333 ( .A(mult_x_1196_n2559), .Y(n18954) );
  MAJx2_ASAP7_75t_SL U25334 ( .A(mult_x_1196_n1982), .B(mult_x_1196_n1959), 
        .C(n23052), .Y(mult_x_1196_n1936) );
  NAND2xp5_ASAP7_75t_SL U25335 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__18_), .B(
        n23903), .Y(n25105) );
  NAND2xp5_ASAP7_75t_SL U25336 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__18_), .B(
        n18910), .Y(n25106) );
  INVx2_ASAP7_75t_SL U25337 ( .A(n24016), .Y(n24015) );
  XNOR2x1_ASAP7_75t_SL U25338 ( .A(n18955), .B(u0_0_leon3x0_p0_muli[46]), .Y(
        n24016) );
  NAND2xp5_ASAP7_75t_SL U25339 ( .A(n23770), .B(n22266), .Y(n18955) );
  OR2x2_ASAP7_75t_SL U25340 ( .A(n23771), .B(n18910), .Y(n22266) );
  NAND2xp5_ASAP7_75t_SL U25341 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__17_), .B(
        n18911), .Y(n23770) );
  INVx2_ASAP7_75t_SL U25342 ( .A(n18957), .Y(n18956) );
  XNOR2x1_ASAP7_75t_SL U25343 ( .A(n24062), .B(n23658), .Y(n18958) );
  INVxp33_ASAP7_75t_SL U25344 ( .A(mult_x_1196_n549), .Y(n23914) );
  XNOR2xp5_ASAP7_75t_SL U25345 ( .A(n18960), .B(n18959), .Y(n22819) );
  MAJIxp5_ASAP7_75t_SL U25346 ( .A(n23183), .B(mult_x_1196_n2629), .C(n24243), 
        .Y(n23325) );
  XOR2xp5_ASAP7_75t_SL U25347 ( .A(mult_x_1196_n2137), .B(mult_x_1196_n2563), 
        .Y(n18959) );
  INVx1_ASAP7_75t_SL U25348 ( .A(mult_x_1196_n2503), .Y(n18960) );
  OAI22xp5_ASAP7_75t_SL U25349 ( .A1(mult_x_1196_n3075), .A2(n24007), .B1(
        n24005), .B2(mult_x_1196_n3074), .Y(mult_x_1196_n2503) );
  XNOR2xp5_ASAP7_75t_SL U25350 ( .A(n18961), .B(mult_x_1196_n1185), .Y(n22930)
         );
  MAJIxp5_ASAP7_75t_SL U25351 ( .A(mult_x_1196_n1185), .B(mult_x_1196_n1183), 
        .C(n18961), .Y(mult_x_1196_n1152) );
  AOI21xp5_ASAP7_75t_SL U25352 ( .A1(n18920), .A2(n18435), .B(
        mult_x_1196_n3077), .Y(n18961) );
  INVx1_ASAP7_75t_SL U25353 ( .A(n18962), .Y(n18964) );
  OAI22xp5_ASAP7_75t_SL U25354 ( .A1(mult_x_1196_n2954), .A2(n23142), .B1(
        mult_x_1196_n2953), .B2(n24017), .Y(n18962) );
  XNOR2xp5_ASAP7_75t_SL U25355 ( .A(n18964), .B(n18963), .Y(mult_x_1196_n1315)
         );
  XNOR2xp5_ASAP7_75t_SL U25356 ( .A(mult_x_1196_n2167), .B(mult_x_1196_n2350), 
        .Y(n18963) );
  MAJIxp5_ASAP7_75t_SL U25357 ( .A(mult_x_1196_n2664), .B(mult_x_1196_n2568), 
        .C(n18966), .Y(mult_x_1196_n2063) );
  XNOR2xp5_ASAP7_75t_SL U25358 ( .A(mult_x_1196_n2568), .B(n18966), .Y(n18965)
         );
  OAI22xp5_ASAP7_75t_SL U25359 ( .A1(mult_x_1196_n3176), .A2(n24230), .B1(
        n23992), .B2(mult_x_1196_n3175), .Y(n18966) );
  INVx1_ASAP7_75t_SL U25360 ( .A(mult_x_1196_n2664), .Y(n18967) );
  MAJIxp5_ASAP7_75t_SL U25361 ( .A(mult_x_1196_n1570), .B(mult_x_1196_n1572), 
        .C(n24284), .Y(mult_x_1196_n1556) );
  XNOR2xp5_ASAP7_75t_SL U25362 ( .A(n18969), .B(n18968), .Y(n23471) );
  INVx1_ASAP7_75t_SL U25363 ( .A(mult_x_1196_n1520), .Y(n18969) );
  XNOR2xp5_ASAP7_75t_SL U25364 ( .A(n18971), .B(mult_x_1196_n1537), .Y(n18970)
         );
  NAND2xp5_ASAP7_75t_SL U25365 ( .A(n18976), .B(n18975), .Y(n18974) );
  INVx1_ASAP7_75t_SL U25366 ( .A(n18978), .Y(n18977) );
  NOR2x1_ASAP7_75t_SL U25367 ( .A(n23589), .B(mult_x_1196_n224), .Y(n18978) );
  INVx1_ASAP7_75t_SL U25368 ( .A(n26372), .Y(n18979) );
  AND2x2_ASAP7_75t_SL U25369 ( .A(n18981), .B(mult_x_1196_n224), .Y(n18980) );
  INVx1_ASAP7_75t_SL U25370 ( .A(n23589), .Y(n18981) );
  XOR2xp5_ASAP7_75t_SL U25371 ( .A(mult_x_1196_n1810), .B(mult_x_1196_n1791), 
        .Y(n23075) );
  XOR2x2_ASAP7_75t_SL U25372 ( .A(n23759), .B(n23758), .Y(mult_x_1196_n1883)
         );
  OAI21x1_ASAP7_75t_SL U25373 ( .A1(n22621), .A2(mult_x_1196_n1872), .B(n22321), .Y(n22620) );
  XNOR2x1_ASAP7_75t_SL U25374 ( .A(n23964), .B(n22227), .Y(mult_x_1196_n3041)
         );
  HB1xp67_ASAP7_75t_SL U25375 ( .A(mult_x_1196_n1882), .Y(n18982) );
  INVxp33_ASAP7_75t_SRAM U25376 ( .A(mult_x_1196_n611), .Y(n23702) );
  XNOR2x1_ASAP7_75t_SL U25377 ( .A(n22901), .B(n22900), .Y(mult_x_1196_n1797)
         );
  OAI22x1_ASAP7_75t_SL U25378 ( .A1(mult_x_1196_n3208), .A2(n23072), .B1(
        mult_x_1196_n3207), .B2(n23987), .Y(mult_x_1196_n2632) );
  BUFx2_ASAP7_75t_SL U25379 ( .A(mult_x_1196_n1271), .Y(n22928) );
  HB1xp67_ASAP7_75t_SL U25380 ( .A(n24200), .Y(n18983) );
  HB1xp67_ASAP7_75t_SL U25381 ( .A(n22227), .Y(n18984) );
  OAI21x1_ASAP7_75t_SL U25382 ( .A1(mult_x_1196_n3177), .A2(n23994), .B(n22318), .Y(n23564) );
  XNOR2x1_ASAP7_75t_SL U25383 ( .A(n23272), .B(mult_x_1196_n1463), .Y(n23319)
         );
  OAI21xp33_ASAP7_75t_SRAM U25384 ( .A1(mult_x_1196_n579), .A2(
        mult_x_1196_n575), .B(n18516), .Y(n18985) );
  XOR2xp5_ASAP7_75t_SL U25385 ( .A(n24180), .B(n23648), .Y(n18986) );
  OAI21xp5_ASAP7_75t_SL U25386 ( .A1(n25104), .A2(n24686), .B(n25103), .Y(
        u0_0_leon3x0_p0_muli[40]) );
  OAI22xp5_ASAP7_75t_SL U25387 ( .A1(mult_x_1196_n2988), .A2(n24014), .B1(
        n24012), .B2(mult_x_1196_n2987), .Y(n23782) );
  NOR2x1_ASAP7_75t_SL U25388 ( .A(mult_x_1196_n3007), .B(n24014), .Y(n23581)
         );
  XOR2xp5_ASAP7_75t_SL U25389 ( .A(n23319), .B(n22370), .Y(n18987) );
  HB1xp67_ASAP7_75t_SL U25390 ( .A(mult_x_1196_n529), .Y(n18988) );
  INVx2_ASAP7_75t_SL U25391 ( .A(mult_x_1196_n1395), .Y(n23772) );
  NAND2x1_ASAP7_75t_SL U25392 ( .A(mult_x_1196_n596), .B(mult_x_1196_n584), 
        .Y(mult_x_1196_n582) );
  NOR2x1_ASAP7_75t_SL U25393 ( .A(mult_x_1196_n602), .B(mult_x_1196_n607), .Y(
        mult_x_1196_n596) );
  HB1xp67_ASAP7_75t_SL U25394 ( .A(mult_x_1196_n1229), .Y(n18989) );
  XNOR2x1_ASAP7_75t_SL U25395 ( .A(n22845), .B(n23612), .Y(n23613) );
  XNOR2x1_ASAP7_75t_SL U25396 ( .A(n22865), .B(n23752), .Y(n22845) );
  INVxp33_ASAP7_75t_SRAM U25397 ( .A(mult_x_1196_n639), .Y(n18990) );
  INVx1_ASAP7_75t_SL U25398 ( .A(n18990), .Y(n18991) );
  OAI22x1_ASAP7_75t_SL U25399 ( .A1(mult_x_1196_n3001), .A2(n24012), .B1(
        n18537), .B2(mult_x_1196_n3002), .Y(mult_x_1196_n2430) );
  XOR2x2_ASAP7_75t_SL U25400 ( .A(mult_x_1196_n1830), .B(mult_x_1196_n1828), 
        .Y(n22853) );
  NAND2x1_ASAP7_75t_SL U25401 ( .A(n25187), .B(n25188), .Y(
        u0_0_leon3x0_p0_muli[39]) );
  BUFx2_ASAP7_75t_SL U25402 ( .A(u0_0_leon3x0_p0_muli[39]), .Y(n22864) );
  INVx2_ASAP7_75t_SL U25403 ( .A(u0_0_leon3x0_p0_muli[39]), .Y(n23951) );
  XNOR2x1_ASAP7_75t_SL U25404 ( .A(n22787), .B(n22786), .Y(mult_x_1196_n1234)
         );
  XNOR2x1_ASAP7_75t_SL U25405 ( .A(n18992), .B(n23772), .Y(mult_x_1196_n1392)
         );
  AND2x2_ASAP7_75t_SL U25406 ( .A(n23961), .B(n24109), .Y(n18993) );
  INVxp33_ASAP7_75t_SRAM U25407 ( .A(mult_x_1196_n638), .Y(n18994) );
  INVxp33_ASAP7_75t_SRAM U25408 ( .A(n18994), .Y(n18995) );
  HB1xp67_ASAP7_75t_SL U25409 ( .A(mult_x_1196_n533), .Y(n18996) );
  OAI22x1_ASAP7_75t_SL U25410 ( .A1(mult_x_1196_n2976), .A2(n24012), .B1(
        n24014), .B2(mult_x_1196_n2977), .Y(mult_x_1196_n2405) );
  NAND2x1p5_ASAP7_75t_SL U25411 ( .A(n24681), .B(n24585), .Y(n31988) );
  BUFx6f_ASAP7_75t_SL U25412 ( .A(n31826), .Y(n24585) );
  NOR2x2_ASAP7_75t_SL U25413 ( .A(DP_OP_1196_128_7433_n456), .B(
        DP_OP_1196_128_7433_n455), .Y(n32171) );
  XNOR2x2_ASAP7_75t_SL U25414 ( .A(n18326), .B(n22829), .Y(mult_x_1196_n1417)
         );
  XNOR2x1_ASAP7_75t_SL U25415 ( .A(n23118), .B(mult_x_1196_n1711), .Y(
        mult_x_1196_n1678) );
  XNOR2x1_ASAP7_75t_SL U25416 ( .A(n22597), .B(mult_x_1196_n1480), .Y(n22596)
         );
  XNOR2x1_ASAP7_75t_SL U25417 ( .A(n23304), .B(n22596), .Y(n23268) );
  HB1xp67_ASAP7_75t_SL U25418 ( .A(n23857), .Y(n18998) );
  HB1xp67_ASAP7_75t_SL U25419 ( .A(mult_x_1196_n1394), .Y(n18999) );
  NOR2x1_ASAP7_75t_SL U25420 ( .A(add_x_735_n241), .B(add_x_735_n236), .Y(
        add_x_735_n230) );
  NOR2x1_ASAP7_75t_SL U25421 ( .A(add_x_735_A_9_), .B(u0_0_leon3x0_p0_divi[7]), 
        .Y(add_x_735_n236) );
  INVx2_ASAP7_75t_SL U25422 ( .A(mult_x_1196_n1780), .Y(n22610) );
  NAND2xp5_ASAP7_75t_SL U25423 ( .A(n23809), .B(n23335), .Y(n23808) );
  NAND2x1_ASAP7_75t_SL U25424 ( .A(n23775), .B(n23774), .Y(n23773) );
  INVx1_ASAP7_75t_SL U25425 ( .A(mult_x_1196_n2862), .Y(n23774) );
  NOR2x1_ASAP7_75t_SL U25426 ( .A(n23115), .B(n23114), .Y(n23373) );
  AND3x1_ASAP7_75t_SL U25427 ( .A(n23574), .B(n23573), .C(mult_x_1196_n788), 
        .Y(n23669) );
  NOR2x1_ASAP7_75t_SL U25428 ( .A(n22404), .B(mult_x_1196_n393), .Y(
        mult_x_1196_n391) );
  NOR2x1_ASAP7_75t_SL U25429 ( .A(mult_x_1196_n613), .B(mult_x_1196_n616), .Y(
        mult_x_1196_n611) );
  AND2x2_ASAP7_75t_SL U25430 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__14_), .B(n24687), .Y(n22273) );
  OAI22xp5_ASAP7_75t_SL U25431 ( .A1(mult_x_1196_n2821), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2820), .Y(mult_x_1196_n2255) );
  NOR2xp33_ASAP7_75t_SL U25432 ( .A(mult_x_1196_n2885), .B(n24026), .Y(n23734)
         );
  XNOR2xp5_ASAP7_75t_SL U25433 ( .A(n23261), .B(mult_x_1196_n1129), .Y(n23511)
         );
  HB1xp67_ASAP7_75t_SL U25434 ( .A(mult_x_1196_n1139), .Y(n22810) );
  BUFx3_ASAP7_75t_SL U25435 ( .A(n22391), .Y(n22481) );
  XOR2xp5_ASAP7_75t_SL U25436 ( .A(mult_x_1196_n1178), .B(n22501), .Y(n22341)
         );
  HB1xp67_ASAP7_75t_SL U25437 ( .A(n22339), .Y(n22521) );
  HB1xp67_ASAP7_75t_SL U25438 ( .A(mult_x_1196_n1089), .Y(n22528) );
  NOR2xp33_ASAP7_75t_SL U25439 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[28]), .Y(
        n26988) );
  XNOR2xp5_ASAP7_75t_SL U25440 ( .A(n23441), .B(mult_x_1196_n882), .Y(n22313)
         );
  XNOR2xp5_ASAP7_75t_SL U25441 ( .A(mult_x_1196_n2050), .B(n23376), .Y(
        mult_x_1196_n2035) );
  HB1xp67_ASAP7_75t_SL U25442 ( .A(mult_x_1196_n2046), .Y(n22490) );
  NOR2xp33_ASAP7_75t_SL U25443 ( .A(mult_x_1196_n2982), .B(n24012), .Y(n23828)
         );
  NOR2xp33_ASAP7_75t_SL U25444 ( .A(mult_x_1196_n387), .B(mult_x_1196_n312), 
        .Y(n23393) );
  AOI21xp5_ASAP7_75t_SL U25445 ( .A1(mult_x_1196_n465), .A2(mult_x_1196_n420), 
        .B(mult_x_1196_n421), .Y(n23134) );
  AND4x1_ASAP7_75t_SL U25446 ( .A(n18514), .B(n23263), .C(mult_x_1196_n793), 
        .D(n23732), .Y(mult_x_1196_n455) );
  HB1xp67_ASAP7_75t_SL U25447 ( .A(mult_x_1196_n526), .Y(n22468) );
  BUFx2_ASAP7_75t_SL U25448 ( .A(n18423), .Y(n23061) );
  HB1xp67_ASAP7_75t_SL U25449 ( .A(n18406), .Y(n23666) );
  INVx2_ASAP7_75t_SL U25450 ( .A(n23746), .Y(u0_0_leon3x0_p0_muli[44]) );
  BUFx3_ASAP7_75t_SL U25451 ( .A(n33058), .Y(n24682) );
  HB1xp67_ASAP7_75t_SL U25452 ( .A(mult_x_1196_n1619), .Y(n22652) );
  NOR2x1_ASAP7_75t_SL U25453 ( .A(n22247), .B(n25236), .Y(n23979) );
  INVx3_ASAP7_75t_SL U25454 ( .A(n24422), .Y(add_x_735_A_16_) );
  BUFx3_ASAP7_75t_SL U25455 ( .A(add_x_735_A_25_), .Y(n23002) );
  BUFx3_ASAP7_75t_SL U25456 ( .A(u0_0_leon3x0_p0_muli[45]), .Y(n22721) );
  OAI21xp5_ASAP7_75t_SL U25457 ( .A1(n23702), .A2(mult_x_1196_n629), .B(n23701), .Y(n23929) );
  HB1xp67_ASAP7_75t_SL U25458 ( .A(mult_x_1196_n753), .Y(n22664) );
  HB1xp67_ASAP7_75t_SL U25459 ( .A(n24262), .Y(n22624) );
  NOR4xp25_ASAP7_75t_SL U25460 ( .A(add_x_735_A_10_), .B(n22449), .C(n18325), 
        .D(n22556), .Y(n31669) );
  BUFx3_ASAP7_75t_SL U25461 ( .A(u0_0_leon3x0_p0_muli[44]), .Y(n22837) );
  OAI22xp5_ASAP7_75t_SL U25462 ( .A1(mult_x_1196_n2760), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2759), .Y(mult_x_1196_n2197) );
  XNOR2xp5_ASAP7_75t_SL U25463 ( .A(n23481), .B(n23480), .Y(n22209) );
  NAND2xp5_ASAP7_75t_SL U25464 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__2_), .B(
        n24687), .Y(n25103) );
  NOR2x1_ASAP7_75t_SL U25465 ( .A(n24686), .B(n25115), .Y(n23153) );
  BUFx3_ASAP7_75t_SL U25466 ( .A(n24009), .Y(n22563) );
  BUFx2_ASAP7_75t_SL U25467 ( .A(n23972), .Y(n23076) );
  BUFx2_ASAP7_75t_SL U25468 ( .A(n24120), .Y(n22538) );
  BUFx6f_ASAP7_75t_SL U25469 ( .A(n24057), .Y(n22442) );
  BUFx3_ASAP7_75t_SL U25470 ( .A(n23962), .Y(n22961) );
  BUFx12f_ASAP7_75t_SL U25471 ( .A(u0_0_leon3x0_p0_muli[15]), .Y(n24072) );
  BUFx6f_ASAP7_75t_SL U25472 ( .A(u0_0_leon3x0_p0_muli[22]), .Y(n24064) );
  INVx6_ASAP7_75t_SL U25473 ( .A(n23588), .Y(n24041) );
  XNOR2xp5_ASAP7_75t_SL U25474 ( .A(n25644), .B(n23415), .Y(n23587) );
  XNOR2xp5_ASAP7_75t_SL U25475 ( .A(n24045), .B(n18926), .Y(mult_x_1196_n3248)
         );
  XNOR2xp5_ASAP7_75t_SL U25476 ( .A(n24061), .B(n23964), .Y(mult_x_1196_n3026)
         );
  AO21x1_ASAP7_75t_SL U25477 ( .A1(n25237), .A2(n18911), .B(n32012), .Y(n22247) );
  OAI22xp5_ASAP7_75t_SL U25478 ( .A1(mult_x_1196_n2858), .A2(n24031), .B1(
        n24030), .B2(mult_x_1196_n2857), .Y(mult_x_1196_n2292) );
  XNOR2xp5_ASAP7_75t_SL U25479 ( .A(n24066), .B(n23960), .Y(mult_x_1196_n3167)
         );
  XNOR2xp5_ASAP7_75t_SL U25480 ( .A(n24056), .B(n23396), .Y(mult_x_1196_n3055)
         );
  XOR2xp5_ASAP7_75t_SL U25481 ( .A(n24205), .B(n24074), .Y(mult_x_1196_n3209)
         );
  INVx1_ASAP7_75t_SL U25482 ( .A(n24031), .Y(n22446) );
  XOR2xp5_ASAP7_75t_SL U25483 ( .A(n24205), .B(n24066), .Y(mult_x_1196_n3201)
         );
  INVx1_ASAP7_75t_SL U25484 ( .A(n24005), .Y(n22460) );
  XNOR2xp5_ASAP7_75t_SL U25485 ( .A(n24054), .B(n23964), .Y(mult_x_1196_n3019)
         );
  XNOR2xp5_ASAP7_75t_SL U25486 ( .A(n24067), .B(add_x_735_A_10_), .Y(
        mult_x_1196_n3134) );
  OAI22xp5_ASAP7_75t_SL U25487 ( .A1(n24021), .A2(mult_x_1196_n2935), .B1(
        mult_x_1196_n2934), .B2(n24020), .Y(mult_x_1196_n2363) );
  XNOR2xp5_ASAP7_75t_SL U25488 ( .A(n24068), .B(n23971), .Y(mult_x_1196_n2863)
         );
  XNOR2xp5_ASAP7_75t_SL U25489 ( .A(n24057), .B(n23967), .Y(mult_x_1196_n2954)
         );
  NOR2xp33_ASAP7_75t_SL U25490 ( .A(n23358), .B(mult_x_1196_n3229), .Y(n22636)
         );
  OAI22xp5_ASAP7_75t_SL U25491 ( .A1(n22647), .A2(mult_x_1196_n3221), .B1(
        mult_x_1196_n3220), .B2(n22538), .Y(mult_x_1196_n2645) );
  OAI22xp5_ASAP7_75t_SL U25492 ( .A1(n23081), .A2(n23421), .B1(n23992), .B2(
        mult_x_1196_n3163), .Y(mult_x_1196_n2588) );
  OAI22xp5_ASAP7_75t_SL U25493 ( .A1(mult_x_1196_n2824), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2823), .Y(mult_x_1196_n2258) );
  BUFx2_ASAP7_75t_SL U25494 ( .A(mult_x_1196_n1748), .Y(n22806) );
  OAI21xp5_ASAP7_75t_SL U25495 ( .A1(mult_x_1196_n3202), .A2(n23522), .B(
        n22315), .Y(n24244) );
  XNOR2xp5_ASAP7_75t_SL U25496 ( .A(n24057), .B(n18926), .Y(mult_x_1196_n3260)
         );
  XNOR2xp5_ASAP7_75t_SL U25497 ( .A(n24067), .B(n23971), .Y(mult_x_1196_n2862)
         );
  OAI22xp5_ASAP7_75t_SL U25498 ( .A1(mult_x_1196_n3223), .A2(n22647), .B1(
        mult_x_1196_n3222), .B2(n22538), .Y(mult_x_1196_n2647) );
  XNOR2xp5_ASAP7_75t_SL U25499 ( .A(n24057), .B(n23964), .Y(mult_x_1196_n3022)
         );
  XNOR2xp5_ASAP7_75t_SL U25500 ( .A(n24072), .B(add_x_735_A_10_), .Y(
        mult_x_1196_n3139) );
  OAI22xp5_ASAP7_75t_SL U25501 ( .A1(mult_x_1196_n3126), .A2(n18397), .B1(
        n23996), .B2(mult_x_1196_n3125), .Y(mult_x_1196_n2550) );
  NOR2xp33_ASAP7_75t_SL U25502 ( .A(mult_x_1196_n3173), .B(n23992), .Y(n22958)
         );
  NOR2xp33_ASAP7_75t_SL U25503 ( .A(mult_x_1196_n2728), .B(n24043), .Y(
        mult_x_1196_n2166) );
  OAI22xp5_ASAP7_75t_SL U25504 ( .A1(mult_x_1196_n3265), .A2(n23982), .B1(
        n22389), .B2(mult_x_1196_n3264), .Y(mult_x_1196_n2689) );
  OAI22xp5_ASAP7_75t_SL U25505 ( .A1(mult_x_1196_n2798), .A2(n24039), .B1(
        mult_x_1196_n2797), .B2(n22391), .Y(mult_x_1196_n2232) );
  NOR2xp33_ASAP7_75t_SL U25506 ( .A(n22756), .B(mult_x_1196_n3093), .Y(n23110)
         );
  NOR2xp33_ASAP7_75t_SL U25507 ( .A(mult_x_1196_n3252), .B(n23982), .Y(n23120)
         );
  NOR2xp33_ASAP7_75t_SL U25508 ( .A(mult_x_1196_n3267), .B(n23982), .Y(n23206)
         );
  NOR2xp33_ASAP7_75t_SL U25509 ( .A(n22389), .B(mult_x_1196_n3266), .Y(n23207)
         );
  XNOR2xp5_ASAP7_75t_SL U25510 ( .A(n24056), .B(n23964), .Y(mult_x_1196_n3021)
         );
  XNOR2xp5_ASAP7_75t_SL U25511 ( .A(n24055), .B(n23964), .Y(mult_x_1196_n3020)
         );
  OAI22xp5_ASAP7_75t_SL U25512 ( .A1(n18528), .A2(mult_x_1196_n3200), .B1(
        mult_x_1196_n3199), .B2(n23987), .Y(mult_x_1196_n2624) );
  NOR2xp33_ASAP7_75t_SL U25513 ( .A(mult_x_1196_n3006), .B(n24012), .Y(n23582)
         );
  NOR2xp33_ASAP7_75t_SL U25514 ( .A(mult_x_1196_n2889), .B(n24026), .Y(n23788)
         );
  NOR2xp33_ASAP7_75t_SL U25515 ( .A(mult_x_1196_n2760), .B(n24040), .Y(n23855)
         );
  XNOR2xp5_ASAP7_75t_SL U25516 ( .A(n24180), .B(n23648), .Y(n23647) );
  XOR2x2_ASAP7_75t_SL U25517 ( .A(n23535), .B(n23060), .Y(n22354) );
  NOR2x1p5_ASAP7_75t_SL U25518 ( .A(n23599), .B(n23598), .Y(n23597) );
  XNOR2xp5_ASAP7_75t_SL U25519 ( .A(mult_x_1196_n2356), .B(mult_x_1196_n2452), 
        .Y(n22843) );
  NOR2xp33_ASAP7_75t_SL U25520 ( .A(mult_x_1196_n2008), .B(n22320), .Y(n23437)
         );
  XOR2xp5_ASAP7_75t_SL U25521 ( .A(n23088), .B(n22690), .Y(n22335) );
  INVx1_ASAP7_75t_SL U25522 ( .A(n23368), .Y(n23366) );
  XNOR2xp5_ASAP7_75t_SL U25523 ( .A(mult_x_1196_n1972), .B(n23567), .Y(
        mult_x_1196_n1974) );
  XOR2xp5_ASAP7_75t_SL U25524 ( .A(n23520), .B(n23519), .Y(n22625) );
  XNOR2xp5_ASAP7_75t_SL U25525 ( .A(n23179), .B(n24265), .Y(n23178) );
  NOR2xp33_ASAP7_75t_SL U25526 ( .A(n24312), .B(mult_x_1196_n1531), .Y(n23370)
         );
  XOR2xp5_ASAP7_75t_SL U25527 ( .A(mult_x_1196_n1327), .B(mult_x_1196_n1298), 
        .Y(n22539) );
  XNOR2xp5_ASAP7_75t_SL U25528 ( .A(mult_x_1196_n1811), .B(n23133), .Y(
        mult_x_1196_n1805) );
  NOR2xp33_ASAP7_75t_SL U25529 ( .A(n23116), .B(mult_x_1196_n2901), .Y(n24160)
         );
  HB1xp67_ASAP7_75t_SL U25530 ( .A(mult_x_1196_n1569), .Y(n22651) );
  NAND2xp5_ASAP7_75t_SL U25531 ( .A(mult_x_1196_n2628), .B(mult_x_1196_n2504), 
        .Y(n23181) );
  HB1xp67_ASAP7_75t_SL U25532 ( .A(n24288), .Y(n22571) );
  NAND2xp5_ASAP7_75t_SL U25533 ( .A(n23775), .B(n23697), .Y(n23696) );
  NOR2xp33_ASAP7_75t_SL U25534 ( .A(mult_x_1196_n3174), .B(n23081), .Y(n22957)
         );
  HB1xp67_ASAP7_75t_SL U25535 ( .A(n23937), .Y(n22935) );
  HB1xp67_ASAP7_75t_SL U25536 ( .A(mult_x_1196_n1422), .Y(n22482) );
  HB1xp67_ASAP7_75t_SL U25537 ( .A(n23005), .Y(n22595) );
  HB1xp67_ASAP7_75t_SL U25538 ( .A(mult_x_1196_n1351), .Y(n22655) );
  NOR2xp33_ASAP7_75t_SL U25539 ( .A(mult_x_1196_n2010), .B(mult_x_1196_n2012), 
        .Y(n22456) );
  HB1xp67_ASAP7_75t_SL U25540 ( .A(n22944), .Y(n22529) );
  HB1xp67_ASAP7_75t_SL U25541 ( .A(mult_x_1196_n1512), .Y(n22761) );
  OAI22xp5_ASAP7_75t_SL U25542 ( .A1(mult_x_1196_n3139), .A2(n24000), .B1(
        n23996), .B2(mult_x_1196_n3138), .Y(mult_x_1196_n2563) );
  NOR2xp33_ASAP7_75t_SL U25543 ( .A(mult_x_1196_n3033), .B(n24008), .Y(n22950)
         );
  HB1xp67_ASAP7_75t_SL U25544 ( .A(mult_x_1196_n3329), .Y(n22791) );
  HB1xp67_ASAP7_75t_SL U25545 ( .A(mult_x_1196_n1822), .Y(n22550) );
  NOR2xp33_ASAP7_75t_SL U25546 ( .A(mult_x_1196_n2564), .B(mult_x_1196_n2596), 
        .Y(n22606) );
  BUFx2_ASAP7_75t_SL U25547 ( .A(n22424), .Y(n22918) );
  HB1xp67_ASAP7_75t_SL U25548 ( .A(mult_x_1196_n1846), .Y(n22697) );
  HB1xp67_ASAP7_75t_SL U25549 ( .A(mult_x_1196_n2009), .Y(n22635) );
  HB1xp67_ASAP7_75t_SL U25550 ( .A(n22688), .Y(n22638) );
  NAND2xp5_ASAP7_75t_SL U25551 ( .A(n23103), .B(n23977), .Y(n23102) );
  HAxp5_ASAP7_75t_SL U25552 ( .A(n19194), .B(n19197), .CON(), .SN(n19000) );
  O2A1O1Ixp33_ASAP7_75t_SL U25553 ( .A1(n19199), .A2(n19198), .B(n19000), .C(
        n19001), .Y(mult_x_1196_n874) );
  INVxp33_ASAP7_75t_SRAM U25554 ( .A(n23947), .Y(n19008) );
  INVxp33_ASAP7_75t_SRAM U25555 ( .A(DP_OP_1196_128_7433_n347), .Y(n19015) );
  AND2x2_ASAP7_75t_SL U25556 ( .A(n19016), .B(DP_OP_1196_128_7433_n351), .Y(
        n19017) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25557 ( .A1(DP_OP_1196_128_7433_n352), .A2(
        DP_OP_1196_128_7433_n350), .B(DP_OP_1196_128_7433_n351), .C(n19016), 
        .Y(n19018) );
  O2A1O1Ixp33_ASAP7_75t_SL U25558 ( .A1(DP_OP_1196_128_7433_n352), .A2(
        DP_OP_1196_128_7433_n350), .B(n19017), .C(n19018), .Y(
        u0_0_leon3x0_p0_iu_N5469) );
  INVxp33_ASAP7_75t_SRAM U25559 ( .A(ahbso_0__HRDATA__8_), .Y(n19020) );
  NAND3xp33_ASAP7_75t_SL U25560 ( .A(DP_OP_1196_128_7433_n374), .B(
        DP_OP_1196_128_7433_n222), .C(n19031), .Y(n19032) );
  A2O1A1Ixp33_ASAP7_75t_SL U25561 ( .A1(DP_OP_1196_128_7433_n222), .A2(
        DP_OP_1196_128_7433_n374), .B(n19031), .C(n19032), .Y(
        u0_0_leon3x0_p0_iu_N5479) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25562 ( .A1(n19037), .A2(n19038), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_), .C(n19039), .Y(n19040) );
  INVxp33_ASAP7_75t_SRAM U25563 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__27_), 
        .Y(n19041) );
  A2O1A1Ixp33_ASAP7_75t_SL U25564 ( .A1(n19043), .A2(n19044), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__27_), .C(n32102), .Y(n19045) );
  INVxp33_ASAP7_75t_SRAM U25565 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_), 
        .Y(n19047) );
  O2A1O1Ixp5_ASAP7_75t_SL U25566 ( .A1(n19042), .A2(n19045), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__28_), .C(n19051), .Y(n29177) );
  INVx1_ASAP7_75t_SL U25567 ( .A(add_x_735_n266), .Y(n19054) );
  A2O1A1Ixp33_ASAP7_75t_SL U25568 ( .A1(add_x_735_n267), .A2(n19054), .B(
        n18892), .C(n19055), .Y(u0_0_leon3x0_p0_dci[7]) );
  INVx1_ASAP7_75t_SL U25569 ( .A(n19065), .Y(n19066) );
  INVx1_ASAP7_75t_SL U25570 ( .A(n32319), .Y(n19068) );
  INVx1_ASAP7_75t_SL U25571 ( .A(n32542), .Y(n19072) );
  A2O1A1Ixp33_ASAP7_75t_SL U25572 ( .A1(n29109), .A2(n29110), .B(
        u0_0_leon3x0_p0_div0_r_NEG_), .C(n19076), .Y(n19077) );
  O2A1O1Ixp33_ASAP7_75t_SL U25573 ( .A1(n30595), .A2(n19084), .B(n19085), .C(
        n19086), .Y(n2588) );
  INVxp33_ASAP7_75t_SRAM U25574 ( .A(n22433), .Y(n19087) );
  A2O1A1Ixp33_ASAP7_75t_SL U25575 ( .A1(sr1_r_WS__2_), .A2(n31714), .B(n31717), 
        .C(n31718), .Y(n19092) );
  INVx1_ASAP7_75t_SL U25576 ( .A(n29350), .Y(n19097) );
  OAI21xp5_ASAP7_75t_SL U25577 ( .A1(uart1_r_IRQCNT__4_), .A2(n19097), .B(
        n29344), .Y(n19098) );
  A2O1A1Ixp33_ASAP7_75t_SL U25578 ( .A1(n29350), .A2(uart1_r_IRQCNT__4_), .B(
        n29344), .C(n19098), .Y(n1760) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25579 ( .A1(n27313), .A2(n27394), .B(n27393), 
        .C(n27317), .Y(n19101) );
  INVx1_ASAP7_75t_SL U25580 ( .A(n19102), .Y(n19103) );
  INVxp33_ASAP7_75t_SRAM U25581 ( .A(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__4_), .Y(n19106) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25582 ( .A1(n32564), .A2(n19106), .B(n32512), 
        .C(n19107), .Y(n19108) );
  A2O1A1Ixp33_ASAP7_75t_SL U25583 ( .A1(n22396), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_READ_), .B(n19114), .C(n24684), .Y(
        n3076) );
  INVxp33_ASAP7_75t_SRAM U25584 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__10_), 
        .Y(n19116) );
  INVxp33_ASAP7_75t_SRAM U25585 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__3_), 
        .Y(n19118) );
  INVxp33_ASAP7_75t_SRAM U25586 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__25_), 
        .Y(n19124) );
  INVxp33_ASAP7_75t_SRAM U25587 ( .A(n18844), .Y(n19126) );
  A2O1A1Ixp33_ASAP7_75t_SL U25588 ( .A1(n24648), .A2(
        u0_0_leon3x0_p0_iu_r_A__WUNF_), .B(n19127), .C(n31439), .Y(n3524) );
  INVxp33_ASAP7_75t_SRAM U25589 ( .A(n27020), .Y(n19128) );
  A2O1A1Ixp33_ASAP7_75t_SL U25590 ( .A1(n32069), .A2(n19128), .B(n24680), .C(
        n19129), .Y(n3576) );
  INVxp33_ASAP7_75t_SRAM U25591 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__29_), 
        .Y(n19133) );
  INVxp33_ASAP7_75t_SRAM U25592 ( .A(u0_0_dbgo_OPTYPE__5_), .Y(n19139) );
  INVx1_ASAP7_75t_SL U25593 ( .A(n24197), .Y(n19143) );
  NAND3xp33_ASAP7_75t_SL U25594 ( .A(mult_x_1196_n829), .B(n19143), .C(n19142), 
        .Y(n19144) );
  A2O1A1Ixp33_ASAP7_75t_SL U25595 ( .A1(n19143), .A2(mult_x_1196_n829), .B(
        n19142), .C(n19144), .Y(n19145) );
  O2A1O1Ixp5_ASAP7_75t_SL U25596 ( .A1(n19151), .A2(n19152), .B(n24684), .C(
        n19153), .Y(n4317) );
  INVxp33_ASAP7_75t_SRAM U25597 ( .A(timer0_r_RELOAD__0_), .Y(n19154) );
  A2O1A1Ixp33_ASAP7_75t_SL U25598 ( .A1(n30266), .A2(n31415), .B(n19163), .C(
        n19164), .Y(n4421) );
  INVxp33_ASAP7_75t_SRAM U25599 ( .A(n31249), .Y(n19169) );
  INVxp33_ASAP7_75t_SRAM U25600 ( .A(n1752), .Y(n19176) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25601 ( .A1(uart1_r_DPAR_), .A2(n19185), .B(
        n27539), .C(n24695), .Y(n19186) );
  INVxp33_ASAP7_75t_SRAM U25602 ( .A(n24043), .Y(n19195) );
  OAI21xp33_ASAP7_75t_SRAM U25603 ( .A1(n24043), .A2(n24050), .B(n22642), .Y(
        n19196) );
  A2O1A1Ixp33_ASAP7_75t_SL U25604 ( .A1(n24050), .A2(n19195), .B(n22642), .C(
        n19196), .Y(n19197) );
  NAND2xp33_ASAP7_75t_SRAM U25605 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__7_), 
        .B(n32186), .Y(n19208) );
  XOR2xp5_ASAP7_75t_SL U25606 ( .A(n26819), .B(n30939), .Y(n19209) );
  INVx1_ASAP7_75t_SL U25607 ( .A(n19210), .Y(n24838) );
  INVxp33_ASAP7_75t_SRAM U25608 ( .A(add_x_735_n99), .Y(n19211) );
  INVxp33_ASAP7_75t_SRAM U25609 ( .A(n24585), .Y(n19218) );
  INVx1_ASAP7_75t_SL U25610 ( .A(n28491), .Y(n19226) );
  A2O1A1Ixp33_ASAP7_75t_SL U25611 ( .A1(u0_0_leon3x0_p0_divi[21]), .A2(n28827), 
        .B(n19229), .C(n28490), .Y(n19230) );
  A2O1A1Ixp33_ASAP7_75t_SL U25612 ( .A1(u0_0_leon3x0_p0_divi[21]), .A2(n28680), 
        .B(n19225), .C(n19231), .Y(n30276) );
  INVxp33_ASAP7_75t_SRAM U25613 ( .A(n30209), .Y(n19233) );
  INVx1_ASAP7_75t_SL U25614 ( .A(n24907), .Y(n19241) );
  O2A1O1Ixp33_ASAP7_75t_SL U25615 ( .A1(n19244), .A2(n19249), .B(n19254), .C(
        n19255), .Y(u0_0_leon3x0_p0_iu_N5495) );
  INVxp33_ASAP7_75t_SRAM U25616 ( .A(DP_OP_5187J1_124_3275_n258), .Y(n19256)
         );
  NAND3xp33_ASAP7_75t_SL U25617 ( .A(DP_OP_5187J1_124_3275_n259), .B(n19256), 
        .C(n23887), .Y(n19257) );
  A2O1A1Ixp33_ASAP7_75t_SL U25618 ( .A1(n19256), .A2(
        DP_OP_5187J1_124_3275_n259), .B(n23887), .C(n19257), .Y(
        u0_0_leon3x0_p0_div0_addout_8_) );
  INVxp33_ASAP7_75t_SRAM U25619 ( .A(n22427), .Y(n19265) );
  INVx1_ASAP7_75t_SL U25620 ( .A(n19268), .Y(n19269) );
  INVx1_ASAP7_75t_SL U25621 ( .A(n32542), .Y(n19282) );
  INVxp33_ASAP7_75t_SRAM U25622 ( .A(n22433), .Y(n19287) );
  INVx1_ASAP7_75t_SL U25623 ( .A(n29342), .Y(n19290) );
  A2O1A1Ixp33_ASAP7_75t_SL U25624 ( .A1(uart1_r_IRQCNT__1_), .A2(n19290), .B(
        n29338), .C(n19291), .Y(n1763) );
  INVx1_ASAP7_75t_SL U25625 ( .A(n19294), .Y(uart1_v_TXCLK__2_) );
  INVxp33_ASAP7_75t_SRAM U25626 ( .A(n32743), .Y(n19295) );
  INVxp33_ASAP7_75t_SRAM U25627 ( .A(u0_0_leon3x0_p0_iu_v_E__CWP__1_), .Y(
        n19302) );
  OAI21xp33_ASAP7_75t_SRAM U25628 ( .A1(u0_0_leon3x0_p0_div0_addout_32_), .A2(
        n31417), .B(n19304), .Y(n19306) );
  A2O1A1Ixp33_ASAP7_75t_SL U25629 ( .A1(n31417), .A2(
        u0_0_leon3x0_p0_div0_addout_32_), .B(n19306), .C(n19305), .Y(n18172)
         );
  INVxp33_ASAP7_75t_SRAM U25630 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__10_), 
        .Y(n19308) );
  INVxp33_ASAP7_75t_SRAM U25631 ( .A(u0_0_leon3x0_p0_ici[20]), .Y(n19310) );
  INVxp33_ASAP7_75t_SRAM U25632 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__8_), 
        .Y(n19312) );
  INVxp33_ASAP7_75t_SRAM U25633 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__8_), 
        .Y(n19315) );
  INVxp33_ASAP7_75t_SRAM U25634 ( .A(n24291), .Y(n19330) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25635 ( .A1(mult_x_1196_n744), .A2(n19330), .B(
        mult_x_1196_n747), .C(n22427), .Y(n19331) );
  A2O1A1Ixp33_ASAP7_75t_SL U25636 ( .A1(n28809), .A2(n19342), .B(n19343), .C(
        n19344), .Y(n4376) );
  INVxp33_ASAP7_75t_SRAM U25637 ( .A(n30386), .Y(n19349) );
  INVxp33_ASAP7_75t_SRAM U25638 ( .A(n31404), .Y(n19352) );
  A2O1A1Ixp33_ASAP7_75t_SL U25639 ( .A1(n31415), .A2(n19349), .B(n19356), .C(
        n19357), .Y(n4445) );
  A2O1A1Ixp33_ASAP7_75t_SL U25640 ( .A1(n4082), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_BMEXC_), .B(n19428), .C(n32201), .Y(
        n19429) );
  INVx1_ASAP7_75t_SL U25641 ( .A(add_x_735_n254), .Y(n19430) );
  NAND3xp33_ASAP7_75t_SL U25642 ( .A(add_x_735_n255), .B(n19430), .C(
        add_x_735_n256), .Y(n19431) );
  A2O1A1Ixp33_ASAP7_75t_SL U25643 ( .A1(n19430), .A2(add_x_735_n255), .B(
        n18893), .C(n19431), .Y(u0_0_leon3x0_p0_dci[9]) );
  INVxp33_ASAP7_75t_SRAM U25644 ( .A(u0_0_leon3x0_p0_iu_fe_pc_2_), .Y(n19437)
         );
  INVxp33_ASAP7_75t_SRAM U25645 ( .A(DP_OP_5187J1_124_3275_n296), .Y(n19444)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U25646 ( .A1(n18836), .A2(n19444), .B(
        DP_OP_5187J1_124_3275_n298), .C(n19445), .Y(
        u0_0_leon3x0_p0_div0_addout_2_) );
  INVxp33_ASAP7_75t_SRAM U25647 ( .A(DP_OP_1196_128_7433_n50), .Y(n19453) );
  INVxp33_ASAP7_75t_SRAM U25648 ( .A(n29422), .Y(n19469) );
  INVx1_ASAP7_75t_SL U25649 ( .A(n32542), .Y(n19481) );
  INVx1_ASAP7_75t_SL U25650 ( .A(n31939), .Y(n19483) );
  INVx1_ASAP7_75t_SL U25651 ( .A(address[13]), .Y(n19484) );
  INVxp33_ASAP7_75t_SRAM U25652 ( .A(n22433), .Y(n19486) );
  INVx1_ASAP7_75t_SL U25653 ( .A(n26776), .Y(n19501) );
  INVxp33_ASAP7_75t_SRAM U25654 ( .A(n31417), .Y(n19502) );
  A2O1A1Ixp33_ASAP7_75t_SL U25655 ( .A1(n31419), .A2(n19502), .B(n19503), .C(
        n31662), .Y(n19504) );
  INVxp33_ASAP7_75t_SRAM U25656 ( .A(irqctrl0_r_ILEVEL__4_), .Y(n19505) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25657 ( .A1(n32562), .A2(n32583), .B(n19507), 
        .C(n31563), .Y(n19508) );
  INVxp33_ASAP7_75t_SRAM U25658 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__PC__2_), 
        .Y(n19509) );
  INVxp33_ASAP7_75t_SRAM U25659 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__23_), 
        .Y(n19511) );
  INVxp33_ASAP7_75t_SRAM U25660 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__29_), 
        .Y(n19513) );
  INVxp33_ASAP7_75t_SRAM U25661 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__27_), 
        .Y(n19517) );
  A2O1A1Ixp33_ASAP7_75t_SL U25662 ( .A1(n30819), .A2(n19521), .B(n30818), .C(
        n19522), .Y(n3562) );
  INVxp33_ASAP7_75t_SRAM U25663 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__22_), .Y(
        n19524) );
  INVxp33_ASAP7_75t_SRAM U25664 ( .A(u0_0_leon3x0_p0_iu_r_D__DIVRDY_), .Y(
        n19526) );
  INVxp33_ASAP7_75t_SRAM U25665 ( .A(n3897), .Y(n19529) );
  A2O1A1Ixp33_ASAP7_75t_SL U25666 ( .A1(n19540), .A2(n28802), .B(n19541), .C(
        n19542), .Y(n4402) );
  INVxp33_ASAP7_75t_SRAM U25667 ( .A(n30789), .Y(n19554) );
  INVxp33_ASAP7_75t_SRAM U25668 ( .A(u0_0_leon3x0_p0_divi[28]), .Y(n19636) );
  O2A1O1Ixp33_ASAP7_75t_SL U25669 ( .A1(n24541), .A2(n30966), .B(n19648), .C(
        n24659), .Y(n30818) );
  INVxp33_ASAP7_75t_SRAM U25670 ( .A(DP_OP_5187J1_124_3275_n274), .Y(n19649)
         );
  INVxp33_ASAP7_75t_SRAM U25671 ( .A(n26456), .Y(n19653) );
  INVxp33_ASAP7_75t_SRAM U25672 ( .A(n22433), .Y(n19682) );
  INVx1_ASAP7_75t_SL U25673 ( .A(uart1_r_TXCLK__1_), .Y(n19686) );
  INVxp33_ASAP7_75t_SRAM U25674 ( .A(n31731), .Y(n19689) );
  INVxp33_ASAP7_75t_SRAM U25675 ( .A(irqctrl0_r_ILEVEL__2_), .Y(n19694) );
  INVxp33_ASAP7_75t_SRAM U25676 ( .A(n31549), .Y(n19698) );
  INVxp33_ASAP7_75t_SRAM U25677 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__2_), 
        .Y(n19703) );
  INVxp33_ASAP7_75t_SRAM U25678 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__7_), 
        .Y(n19705) );
  INVxp33_ASAP7_75t_SRAM U25679 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__4_), 
        .Y(n19707) );
  INVxp33_ASAP7_75t_SRAM U25680 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__14_), 
        .Y(n19715) );
  INVxp33_ASAP7_75t_SRAM U25681 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__15_), .Y(
        n19717) );
  A2O1A1Ixp33_ASAP7_75t_SL U25682 ( .A1(n24647), .A2(n19717), .B(n30114), .C(
        n28701), .Y(n19718) );
  A2O1A1Ixp33_ASAP7_75t_SL U25683 ( .A1(n24909), .A2(n24900), .B(n24908), .C(
        n19719), .Y(n3723) );
  INVx1_ASAP7_75t_SL U25684 ( .A(n30706), .Y(n19720) );
  INVxp33_ASAP7_75t_SRAM U25685 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__26_), 
        .Y(n19722) );
  INVxp33_ASAP7_75t_SRAM U25686 ( .A(u0_0_leon3x0_p0_dci[6]), .Y(n19734) );
  INVxp33_ASAP7_75t_SRAM U25687 ( .A(u0_0_leon3x0_p0_dci[7]), .Y(n19735) );
  INVx1_ASAP7_75t_SL U25688 ( .A(n22664), .Y(n19738) );
  INVxp33_ASAP7_75t_SRAM U25689 ( .A(u0_0_leon3x0_p0_divi[40]), .Y(n19745) );
  INVxp33_ASAP7_75t_SRAM U25690 ( .A(n31664), .Y(n19757) );
  A2O1A1Ixp33_ASAP7_75t_SL U25691 ( .A1(n19770), .A2(n19777), .B(n31673), .C(
        n31677), .Y(n19778) );
  O2A1O1Ixp33_ASAP7_75t_SL U25692 ( .A1(n19779), .A2(n4517), .B(n29952), .C(
        n24695), .Y(n17445) );
  HAxp5_ASAP7_75t_SL U25693 ( .A(n24053), .B(n22642), .CON(), .SN(n19780) );
  INVx1_ASAP7_75t_SL U25694 ( .A(n32356), .Y(n19788) );
  INVx1_ASAP7_75t_SL U25695 ( .A(n31352), .Y(n19791) );
  INVxp33_ASAP7_75t_SRAM U25696 ( .A(u0_0_leon3x0_p0_iu_fe_pc_28_), .Y(n19800)
         );
  INVxp33_ASAP7_75t_SRAM U25697 ( .A(n29433), .Y(n19821) );
  INVx1_ASAP7_75t_SL U25698 ( .A(n31963), .Y(n19840) );
  INVxp33_ASAP7_75t_SRAM U25699 ( .A(n22433), .Y(n19843) );
  INVxp33_ASAP7_75t_SRAM U25700 ( .A(n32705), .Y(n19846) );
  INVxp33_ASAP7_75t_SRAM U25701 ( .A(n27515), .Y(n19854) );
  A2O1A1Ixp33_ASAP7_75t_SL U25702 ( .A1(n24605), .A2(n19862), .B(n24604), .C(
        n19863), .Y(n19864) );
  A2O1A1Ixp33_ASAP7_75t_SL U25703 ( .A1(n28174), .A2(n19864), .B(n19868), .C(
        n28154), .Y(n2879) );
  INVxp33_ASAP7_75t_SRAM U25704 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__23_), 
        .Y(n19869) );
  INVxp33_ASAP7_75t_SRAM U25705 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__7_), 
        .Y(n19871) );
  INVxp33_ASAP7_75t_SRAM U25706 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__11_), .Y(
        n19873) );
  A2O1A1Ixp33_ASAP7_75t_SL U25707 ( .A1(n24647), .A2(n19873), .B(n29207), .C(
        n24495), .Y(n19874) );
  INVxp33_ASAP7_75t_SRAM U25708 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__10_), 
        .Y(n19876) );
  INVxp33_ASAP7_75t_SRAM U25709 ( .A(u0_0_dbgo_OPTYPE__4_), .Y(n19878) );
  INVxp33_ASAP7_75t_SRAM U25710 ( .A(n30809), .Y(n19882) );
  INVxp33_ASAP7_75t_SRAM U25711 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__1_), 
        .Y(n19889) );
  O2A1O1Ixp33_ASAP7_75t_SL U25712 ( .A1(n30595), .A2(n19897), .B(n19898), .C(
        n19899), .Y(n4346) );
  A2O1A1Ixp33_ASAP7_75t_SL U25713 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[22]), .B(n19900), .C(n31638), .Y(n4355) );
  A2O1A1Ixp33_ASAP7_75t_SL U25714 ( .A1(n22413), .A2(n19905), .B(n31488), .C(
        n19913), .Y(n19914) );
  A2O1A1Ixp33_ASAP7_75t_SL U25715 ( .A1(n29953), .A2(uart1_r_PAREN_), .B(
        n29952), .C(n19915), .Y(n19916) );
  INVxp33_ASAP7_75t_SRAM U25716 ( .A(n31706), .Y(n19974) );
  INVxp33_ASAP7_75t_SRAM U25717 ( .A(n31803), .Y(n19976) );
  A2O1A1Ixp33_ASAP7_75t_SL U25718 ( .A1(n32703), .A2(n19974), .B(n19975), .C(
        n19976), .Y(n4722) );
  HAxp5_ASAP7_75t_SL U25719 ( .A(n24061), .B(n22642), .CON(), .SN(n19977) );
  INVx1_ASAP7_75t_SL U25720 ( .A(n24043), .Y(n19978) );
  A2O1A1Ixp33_ASAP7_75t_SL U25721 ( .A1(n24047), .A2(n19978), .B(n22642), .C(
        n19979), .Y(n21252) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25722 ( .A1(n25198), .A2(n28621), .B(n19993), 
        .C(n28850), .Y(n19994) );
  INVx1_ASAP7_75t_SL U25723 ( .A(n27505), .Y(n20000) );
  INVxp33_ASAP7_75t_SRAM U25724 ( .A(n32186), .Y(n20008) );
  O2A1O1Ixp33_ASAP7_75t_SL U25725 ( .A1(n32178), .A2(n20008), .B(n22379), .C(
        n20009), .Y(n31333) );
  INVx1_ASAP7_75t_SL U25726 ( .A(DP_OP_1196_128_7433_n77), .Y(n20013) );
  NAND3xp33_ASAP7_75t_SL U25727 ( .A(DP_OP_1196_128_7433_n80), .B(n20013), .C(
        n20016), .Y(n20017) );
  A2O1A1Ixp33_ASAP7_75t_SL U25728 ( .A1(n20013), .A2(DP_OP_1196_128_7433_n80), 
        .B(n20016), .C(n20017), .Y(u0_0_leon3x0_p0_iu_N5491) );
  INVxp33_ASAP7_75t_SRAM U25729 ( .A(DP_OP_5187J1_124_3275_n237), .Y(n20024)
         );
  NAND3xp33_ASAP7_75t_SL U25730 ( .A(DP_OP_5187J1_124_3275_n238), .B(n20024), 
        .C(n20023), .Y(n20025) );
  A2O1A1Ixp33_ASAP7_75t_SL U25731 ( .A1(n20024), .A2(
        DP_OP_5187J1_124_3275_n238), .B(n20023), .C(n20025), .Y(
        u0_0_leon3x0_p0_div0_addout_11_) );
  A2O1A1Ixp33_ASAP7_75t_SL U25732 ( .A1(n24694), .A2(uart1_r_TWADDR__1_), .B(
        n29356), .C(n20055), .Y(n2269) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25733 ( .A1(u0_0_leon3x0_p0_divo[31]), .A2(
        n24423), .B(n31654), .C(n24659), .Y(n20056) );
  INVxp33_ASAP7_75t_SRAM U25734 ( .A(n29971), .Y(n20062) );
  INVxp33_ASAP7_75t_SRAM U25735 ( .A(n31892), .Y(n20065) );
  INVxp33_ASAP7_75t_SRAM U25736 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__2_), 
        .Y(n20071) );
  INVxp33_ASAP7_75t_SRAM U25737 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__28_), 
        .Y(n20073) );
  INVxp33_ASAP7_75t_SRAM U25738 ( .A(u0_0_leon3x0_p0_ici[2]), .Y(n20076) );
  INVxp33_ASAP7_75t_SRAM U25739 ( .A(u0_0_leon3x0_p0_iu_r_X__DCI__SIGNED_), 
        .Y(n20078) );
  A2O1A1Ixp33_ASAP7_75t_SL U25740 ( .A1(n24648), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__6_), .B(n20082), .C(n24495), .Y(n3678) );
  INVxp33_ASAP7_75t_SRAM U25741 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RETT_), .Y(
        n20083) );
  A2O1A1Ixp33_ASAP7_75t_SL U25742 ( .A1(u0_0_leon3x0_p0_iu_r_M__CTRL__RETT_), 
        .A2(n25604), .B(n22378), .C(n20084), .Y(n3694) );
  A2O1A1Ixp33_ASAP7_75t_SL U25743 ( .A1(n22421), .A2(n29695), .B(n20089), .C(
        n25610), .Y(n3731) );
  INVxp33_ASAP7_75t_SRAM U25744 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__6_), 
        .Y(n20093) );
  INVxp33_ASAP7_75t_SRAM U25745 ( .A(n31625), .Y(n20095) );
  INVxp33_ASAP7_75t_SRAM U25746 ( .A(n31897), .Y(n20096) );
  A2O1A1Ixp33_ASAP7_75t_SL U25747 ( .A1(n30679), .A2(n30678), .B(n30945), .C(
        n20102), .Y(n4338) );
  INVxp33_ASAP7_75t_SRAM U25748 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__27_), .Y(
        n20103) );
  O2A1O1Ixp33_ASAP7_75t_SL U25749 ( .A1(n30595), .A2(n20116), .B(n20117), .C(
        n20118), .Y(n4423) );
  A2O1A1Ixp33_ASAP7_75t_SL U25750 ( .A1(n20119), .A2(n20120), .B(n24549), .C(
        n20121), .Y(n20122) );
  A2O1A1Ixp33_ASAP7_75t_SL U25751 ( .A1(n18859), .A2(n30210), .B(n20122), .C(
        n20123), .Y(n4480) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25752 ( .A1(apbi[29]), .A2(n29652), .B(n29651), 
        .C(n29236), .Y(n20129) );
  INVxp33_ASAP7_75t_SRAM U25753 ( .A(n29238), .Y(n20130) );
  A2O1A1Ixp33_ASAP7_75t_SL U25754 ( .A1(irqctrl0_r_IFORCE__0__13_), .A2(n20128), .B(n20129), .C(n20130), .Y(n4664) );
  INVxp33_ASAP7_75t_SRAM U25755 ( .A(uart1_r_RCNT__3_), .Y(n20131) );
  INVx1_ASAP7_75t_SL U25756 ( .A(n32008), .Y(n20134) );
  O2A1O1Ixp5_ASAP7_75t_SL U25757 ( .A1(uart1_r_TPAR_), .A2(n20136), .B(n20138), 
        .C(n20139), .Y(n4700) );
  INVxp33_ASAP7_75t_SRAM U25758 ( .A(n32717), .Y(n20141) );
  INVxp33_ASAP7_75t_SRAM U25759 ( .A(n31728), .Y(n20143) );
  A2O1A1Ixp33_ASAP7_75t_SL U25760 ( .A1(sr1_r_MCFG2__RAMWWS__0_), .A2(n20143), 
        .B(n20146), .C(n31729), .Y(n20147) );
  A2O1A1Ixp33_ASAP7_75t_SL U25761 ( .A1(sr1_r_WS__0_), .A2(n31740), .B(n20142), 
        .C(n20147), .Y(n20148) );
  HAxp5_ASAP7_75t_SL U25762 ( .A(n18556), .B(n22642), .CON(), .SN(n20152) );
  XOR2xp5_ASAP7_75t_SL U25763 ( .A(n22573), .B(mult_x_1196_n2150), .Y(n22572)
         );
  INVxp33_ASAP7_75t_SRAM U25764 ( .A(DP_OP_5187J1_124_3275_n300), .Y(n20192)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U25765 ( .A1(DP_OP_5187J1_124_3275_n301), .A2(
        n20192), .B(n24317), .C(n20193), .Y(u0_0_leon3x0_p0_div0_addout_1_) );
  INVx1_ASAP7_75t_SL U25766 ( .A(n23887), .Y(n20197) );
  NAND3xp33_ASAP7_75t_SL U25767 ( .A(DP_OP_5187J1_124_3275_n329), .B(
        DP_OP_5187J1_124_3275_n245), .C(n20198), .Y(n20199) );
  A2O1A1Ixp33_ASAP7_75t_SL U25768 ( .A1(DP_OP_5187J1_124_3275_n245), .A2(
        DP_OP_5187J1_124_3275_n329), .B(n20198), .C(n20199), .Y(
        u0_0_leon3x0_p0_div0_addout_10_) );
  INVx1_ASAP7_75t_SL U25769 ( .A(n23941), .Y(n20200) );
  A2O1A1Ixp33_ASAP7_75t_SL U25770 ( .A1(DP_OP_1196_128_7433_n95), .A2(
        DP_OP_1196_128_7433_n98), .B(n20201), .C(n20202), .Y(
        u0_0_leon3x0_p0_iu_N5489) );
  INVxp33_ASAP7_75t_SRAM U25771 ( .A(n27986), .Y(n20220) );
  A2O1A1Ixp33_ASAP7_75t_SL U25772 ( .A1(uart1_r_TRADDR__0_), .A2(n20217), .B(
        n20229), .C(n20252), .Y(n30871) );
  INVxp33_ASAP7_75t_SRAM U25773 ( .A(n22433), .Y(n20276) );
  INVxp33_ASAP7_75t_SRAM U25774 ( .A(n22433), .Y(n20279) );
  INVxp33_ASAP7_75t_SRAM U25775 ( .A(n27308), .Y(n20282) );
  A2O1A1Ixp33_ASAP7_75t_SL U25776 ( .A1(n24694), .A2(n20282), .B(n27327), .C(
        n20284), .Y(n2266) );
  INVxp33_ASAP7_75t_SRAM U25777 ( .A(n30653), .Y(n20285) );
  INVx1_ASAP7_75t_SL U25778 ( .A(n29977), .Y(n20288) );
  A2O1A1Ixp33_ASAP7_75t_SL U25779 ( .A1(n29978), .A2(n29987), .B(n29985), .C(
        n20289), .Y(n2462) );
  A2O1A1Ixp33_ASAP7_75t_SL U25780 ( .A1(n27493), .A2(n29325), .B(n20291), .C(
        n20294), .Y(n2697) );
  A2O1A1Ixp33_ASAP7_75t_SL U25781 ( .A1(n24595), .A2(n24604), .B(n24603), .C(
        n20297), .Y(n20298) );
  A2O1A1Ixp33_ASAP7_75t_SL U25782 ( .A1(n28174), .A2(n20298), .B(n20302), .C(
        n28153), .Y(n2880) );
  INVxp33_ASAP7_75t_SRAM U25783 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__29_), .Y(
        n20303) );
  INVxp33_ASAP7_75t_SRAM U25784 ( .A(n22390), .Y(n20308) );
  INVxp33_ASAP7_75t_SRAM U25785 ( .A(u0_0_leon3x0_p0_iu_r_W__S__WIM__7_), .Y(
        n20314) );
  INVxp33_ASAP7_75t_SRAM U25786 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__1_), 
        .Y(n20316) );
  INVxp33_ASAP7_75t_SRAM U25787 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__5_), 
        .Y(n20318) );
  INVx1_ASAP7_75t_SL U25788 ( .A(n30580), .Y(n20324) );
  INVx1_ASAP7_75t_SL U25789 ( .A(n29207), .Y(n20325) );
  INVxp33_ASAP7_75t_SRAM U25790 ( .A(n31657), .Y(n20326) );
  A2O1A1Ixp33_ASAP7_75t_SL U25791 ( .A1(n31660), .A2(n20326), .B(n31659), .C(
        n20327), .Y(n18174) );
  INVxp33_ASAP7_75t_SRAM U25792 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__26_), 
        .Y(n20328) );
  INVxp33_ASAP7_75t_SRAM U25793 ( .A(n32038), .Y(n20330) );
  INVxp33_ASAP7_75t_SRAM U25794 ( .A(mult_x_1196_n760), .Y(n20332) );
  A2O1A1Ixp33_ASAP7_75t_SL U25795 ( .A1(mult_x_1196_n761), .A2(n20332), .B(
        n22624), .C(n20333), .Y(n20334) );
  A2O1A1Ixp33_ASAP7_75t_SL U25796 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[25]), .B(n20340), .C(n31638), .Y(n4386) );
  INVxp33_ASAP7_75t_SRAM U25797 ( .A(n22379), .Y(n20341) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25798 ( .A1(n29883), .A2(
        u0_0_leon3x0_p0_iu_r_M__CTRL__TT__5_), .B(n20356), .C(n20357), .Y(
        n4564) );
  A2O1A1Ixp33_ASAP7_75t_SL U25799 ( .A1(n30030), .A2(timer0_vtimers_1__IRQEN_), 
        .B(n20358), .C(n24694), .Y(n4690) );
  HAxp5_ASAP7_75t_SL U25800 ( .A(n24055), .B(n22642), .CON(), .SN(n20363) );
  HAxp5_ASAP7_75t_SL U25801 ( .A(n24060), .B(n22642), .CON(), .SN(n20364) );
  HAxp5_ASAP7_75t_SL U25802 ( .A(n24048), .B(n22642), .CON(), .SN(n20365) );
  INVx1_ASAP7_75t_SL U25803 ( .A(add_x_746_n135), .Y(n20372) );
  INVx1_ASAP7_75t_SL U25804 ( .A(n2388), .Y(n20373) );
  INVxp33_ASAP7_75t_SRAM U25805 ( .A(n31308), .Y(n20376) );
  INVxp33_ASAP7_75t_SRAM U25806 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUCIN_), .Y(
        n20384) );
  INVxp33_ASAP7_75t_SRAM U25807 ( .A(n30939), .Y(n20388) );
  INVx1_ASAP7_75t_SL U25808 ( .A(DP_OP_5187J1_124_3275_n213), .Y(n20391) );
  INVxp33_ASAP7_75t_SRAM U25809 ( .A(DP_OP_5187J1_124_3275_n206), .Y(n20395)
         );
  INVxp33_ASAP7_75t_SRAM U25810 ( .A(DP_OP_5187J1_124_3275_n199), .Y(n20399)
         );
  NAND3xp33_ASAP7_75t_SL U25811 ( .A(DP_OP_5187J1_124_3275_n200), .B(n20399), 
        .C(n20398), .Y(n20400) );
  A2O1A1Ixp33_ASAP7_75t_SL U25812 ( .A1(n20399), .A2(
        DP_OP_5187J1_124_3275_n200), .B(n20398), .C(n20400), .Y(
        u0_0_leon3x0_p0_div0_addout_15_) );
  INVx1_ASAP7_75t_SL U25813 ( .A(n32319), .Y(n20415) );
  INVx1_ASAP7_75t_SL U25814 ( .A(n32542), .Y(n20426) );
  A2O1A1Ixp33_ASAP7_75t_SL U25815 ( .A1(n31262), .A2(n31459), .B(n22380), .C(
        n20439), .Y(n20440) );
  INVxp33_ASAP7_75t_SRAM U25816 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__5_), 
        .Y(n20444) );
  INVxp33_ASAP7_75t_SRAM U25817 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__2_), 
        .Y(n20448) );
  INVxp33_ASAP7_75t_SRAM U25818 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__9_), 
        .Y(n20453) );
  INVxp33_ASAP7_75t_SRAM U25819 ( .A(u0_0_leon3x0_p0_iu_r_E__CTRL__RETT_), .Y(
        n20455) );
  A2O1A1Ixp33_ASAP7_75t_SL U25820 ( .A1(n31811), .A2(
        u0_0_leon3x0_p0_iu_r_A__CTRL__RETT_), .B(n24678), .C(n20456), .Y(n3698) );
  O2A1O1Ixp33_ASAP7_75t_SL U25821 ( .A1(n31672), .A2(n31662), .B(n31661), .C(
        n20457), .Y(n20458) );
  INVxp33_ASAP7_75t_SRAM U25822 ( .A(n3730), .Y(n20460) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25823 ( .A1(n32660), .A2(n32122), .B(n32676), 
        .C(n22380), .Y(n20464) );
  INVxp33_ASAP7_75t_SRAM U25824 ( .A(n26811), .Y(n20465) );
  A2O1A1Ixp33_ASAP7_75t_SL U25825 ( .A1(n26808), .A2(n20465), .B(n20468), .C(
        n20469), .Y(n20470) );
  INVx1_ASAP7_75t_SL U25826 ( .A(n20470), .Y(n4012) );
  INVxp33_ASAP7_75t_SRAM U25827 ( .A(u0_0_leon3x0_p0_iu_r_X__LADDR__1_), .Y(
        n20471) );
  A2O1A1Ixp33_ASAP7_75t_SL U25828 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[27]), .B(n20479), .C(n31638), .Y(n4415) );
  INVx1_ASAP7_75t_SL U25829 ( .A(n30393), .Y(n20480) );
  INVxp33_ASAP7_75t_SRAM U25830 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__8_), .Y(
        n20481) );
  O2A1O1Ixp33_ASAP7_75t_SL U25831 ( .A1(n30395), .A2(n20480), .B(n30394), .C(
        n20485), .Y(n20486) );
  INVxp33_ASAP7_75t_SRAM U25832 ( .A(n23229), .Y(n20488) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U25833 ( .A1(apbi[30]), .A2(n29652), .B(n29651), 
        .C(n30547), .Y(n20502) );
  O2A1O1Ixp33_ASAP7_75t_SL U25834 ( .A1(apbi[30]), .A2(n29650), .B(n29649), 
        .C(n29655), .Y(n20503) );
  INVxp33_ASAP7_75t_SRAM U25835 ( .A(n29656), .Y(n20504) );
  A2O1A1Ixp33_ASAP7_75t_SL U25836 ( .A1(n20506), .A2(n20507), .B(
        mult_x_1196_n849), .C(n20508), .Y(mult_x_1196_n843) );
  INVx1_ASAP7_75t_SL U25837 ( .A(n2387), .Y(n20527) );
  INVx1_ASAP7_75t_SL U25838 ( .A(n32256), .Y(n20529) );
  INVxp33_ASAP7_75t_SRAM U25839 ( .A(n23229), .Y(n20530) );
  INVx1_ASAP7_75t_SL U25840 ( .A(n26084), .Y(n20531) );
  INVxp33_ASAP7_75t_SRAM U25841 ( .A(u0_0_leon3x0_p0_iu_fe_pc_16_), .Y(n20535)
         );
  INVxp33_ASAP7_75t_SRAM U25842 ( .A(DP_OP_1196_128_7433_n90), .Y(n20536) );
  INVxp33_ASAP7_75t_SRAM U25843 ( .A(u0_0_leon3x0_p0_muli[10]), .Y(n20540) );
  INVx1_ASAP7_75t_SL U25844 ( .A(n31894), .Y(n20549) );
  INVxp33_ASAP7_75t_SRAM U25845 ( .A(u0_0_leon3x0_p0_iu_fe_pc_24_), .Y(n20555)
         );
  NAND3xp33_ASAP7_75t_SL U25846 ( .A(DP_OP_5187J1_124_3275_n209), .B(n20560), 
        .C(n20559), .Y(n20561) );
  A2O1A1Ixp33_ASAP7_75t_SL U25847 ( .A1(n20560), .A2(
        DP_OP_5187J1_124_3275_n209), .B(n20559), .C(n20561), .Y(
        u0_0_leon3x0_p0_div0_addout_14_) );
  INVx1_ASAP7_75t_SL U25848 ( .A(n32542), .Y(n20582) );
  INVxp33_ASAP7_75t_SRAM U25849 ( .A(n22433), .Y(n20586) );
  INVxp33_ASAP7_75t_SRAM U25850 ( .A(n22433), .Y(n20589) );
  INVxp33_ASAP7_75t_SRAM U25851 ( .A(n29356), .Y(n20592) );
  A2O1A1Ixp33_ASAP7_75t_SL U25852 ( .A1(n24694), .A2(n20592), .B(n27357), .C(
        n20594), .Y(n2270) );
  A2O1A1Ixp33_ASAP7_75t_SL U25853 ( .A1(n24583), .A2(n20599), .B(n32786), .C(
        n20600), .Y(n2362) );
  INVxp33_ASAP7_75t_SRAM U25854 ( .A(n30653), .Y(n20601) );
  INVxp33_ASAP7_75t_SRAM U25855 ( .A(n22390), .Y(n20606) );
  INVxp33_ASAP7_75t_SRAM U25856 ( .A(n26802), .Y(n20609) );
  INVxp33_ASAP7_75t_SRAM U25857 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__25_), 
        .Y(n20613) );
  INVxp33_ASAP7_75t_SRAM U25858 ( .A(n22390), .Y(n20615) );
  INVxp33_ASAP7_75t_SRAM U25859 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__29_), 
        .Y(n20621) );
  INVxp33_ASAP7_75t_SRAM U25860 ( .A(n30472), .Y(n20623) );
  INVxp33_ASAP7_75t_SRAM U25861 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__5_), 
        .Y(n20624) );
  INVxp33_ASAP7_75t_SRAM U25862 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__4_), 
        .Y(n20626) );
  INVx1_ASAP7_75t_SL U25863 ( .A(n31874), .Y(n20632) );
  INVxp33_ASAP7_75t_SRAM U25864 ( .A(n30980), .Y(n20642) );
  INVx1_ASAP7_75t_SL U25865 ( .A(mult_x_1196_n771), .Y(n20650) );
  O2A1O1Ixp33_ASAP7_75t_SL U25866 ( .A1(n30595), .A2(n20662), .B(n20663), .C(
        n20664), .Y(n4465) );
  INVxp33_ASAP7_75t_SRAM U25867 ( .A(n33023), .Y(n20683) );
  INVxp33_ASAP7_75t_SRAM U25868 ( .A(irqctrl0_r_IFORCE__0__13_), .Y(n20690) );
  A2O1A1Ixp33_ASAP7_75t_SL U25869 ( .A1(apbi[13]), .A2(n29657), .B(n20689), 
        .C(n20692), .Y(n4663) );
  INVx1_ASAP7_75t_SL U25870 ( .A(mult_x_1196_n870), .Y(n20697) );
  INVx1_ASAP7_75t_SL U25871 ( .A(n32802), .Y(n20704) );
  INVxp33_ASAP7_75t_SRAM U25872 ( .A(u0_0_leon3x0_p0_dci[40]), .Y(n20713) );
  INVx1_ASAP7_75t_SL U25873 ( .A(n20726), .Y(n30783) );
  INVx1_ASAP7_75t_SL U25874 ( .A(n32542), .Y(n20750) );
  INVx1_ASAP7_75t_SL U25875 ( .A(n25238), .Y(n20756) );
  INVxp33_ASAP7_75t_SRAM U25876 ( .A(n22433), .Y(n20757) );
  INVxp33_ASAP7_75t_SRAM U25877 ( .A(u0_0_leon3x0_p0_ici[19]), .Y(n20760) );
  A2O1A1Ixp33_ASAP7_75t_SL U25878 ( .A1(n30819), .A2(n20769), .B(n30489), .C(
        n20770), .Y(n2703) );
  INVxp33_ASAP7_75t_SRAM U25879 ( .A(n32167), .Y(n20773) );
  A2O1A1Ixp33_ASAP7_75t_SL U25880 ( .A1(n24594), .A2(n24603), .B(n24602), .C(
        n20778), .Y(n20779) );
  A2O1A1Ixp33_ASAP7_75t_SL U25881 ( .A1(n28174), .A2(n20779), .B(n20783), .C(
        n28152), .Y(n2881) );
  INVxp33_ASAP7_75t_SRAM U25882 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__14_), 
        .Y(n20792) );
  INVxp33_ASAP7_75t_SRAM U25883 ( .A(u0_0_leon3x0_p0_ici[8]), .Y(n20795) );
  INVxp33_ASAP7_75t_SRAM U25884 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__5_), 
        .Y(n20797) );
  INVxp33_ASAP7_75t_SRAM U25885 ( .A(u0_0_leon3x0_p0_iu_r_A__MULSTART_), .Y(
        n20801) );
  A2O1A1Ixp33_ASAP7_75t_SL U25886 ( .A1(n32049), .A2(n32048), .B(n24680), .C(
        n20802), .Y(n3867) );
  INVxp33_ASAP7_75t_SRAM U25887 ( .A(u0_0_leon3x0_p0_iu_r_X__LADDR__0_), .Y(
        n20810) );
  INVx1_ASAP7_75t_SL U25888 ( .A(n26812), .Y(n20813) );
  INVxp33_ASAP7_75t_SRAM U25889 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__31_), 
        .Y(n20815) );
  A2O1A1Ixp33_ASAP7_75t_SL U25890 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[24]), .B(n20818), .C(n31638), .Y(n4498) );
  INVxp33_ASAP7_75t_SRAM U25891 ( .A(n22379), .Y(n20820) );
  A2O1A1Ixp33_ASAP7_75t_SL U25892 ( .A1(n30246), .A2(n31415), .B(n20837), .C(
        n20838), .Y(n4607) );
  INVxp33_ASAP7_75t_SRAM U25893 ( .A(sr1_r_MCFG2__RAMRWS__1_), .Y(n20846) );
  INVxp33_ASAP7_75t_SRAM U25894 ( .A(sr1_r_MCFG2__RAMWWS__1_), .Y(n20848) );
  INVxp33_ASAP7_75t_SRAM U25895 ( .A(sr1_r_MCFG1__IOWS__1_), .Y(n20850) );
  O2A1O1Ixp33_ASAP7_75t_SL U25896 ( .A1(n4724), .A2(n31724), .B(n31723), .C(
        n31722), .Y(n20854) );
  O2A1O1Ixp5_ASAP7_75t_SL U25897 ( .A1(n20847), .A2(n20849), .B(n31729), .C(
        n20857), .Y(n20858) );
  INVxp33_ASAP7_75t_SRAM U25898 ( .A(n29443), .Y(n20859) );
  O2A1O1Ixp33_ASAP7_75t_SL U25899 ( .A1(n29665), .A2(n20859), .B(n20860), .C(
        n29407), .Y(n20861) );
  O2A1O1Ixp33_ASAP7_75t_SL U25900 ( .A1(n20861), .A2(n29414), .B(n29880), .C(
        n20862), .Y(n20863) );
  INVx1_ASAP7_75t_SL U25901 ( .A(n20867), .Y(n20868) );
  HAxp5_ASAP7_75t_SL U25902 ( .A(n24054), .B(n23978), .CON(), .SN(n20869) );
  INVx1_ASAP7_75t_SL U25903 ( .A(DP_OP_5187J1_124_3275_n289), .Y(n20885) );
  NAND3xp33_ASAP7_75t_SL U25904 ( .A(n20885), .B(DP_OP_5187J1_124_3275_n335), 
        .C(n18834), .Y(n20886) );
  A2O1A1Ixp33_ASAP7_75t_SL U25905 ( .A1(DP_OP_5187J1_124_3275_n335), .A2(
        n18834), .B(n20885), .C(n20886), .Y(u0_0_leon3x0_p0_div0_addout_4_) );
  INVxp33_ASAP7_75t_SRAM U25906 ( .A(DP_OP_1196_128_7433_n66), .Y(n20888) );
  INVxp33_ASAP7_75t_SRAM U25907 ( .A(DP_OP_1196_128_7433_n57), .Y(n20894) );
  NAND3xp33_ASAP7_75t_SL U25908 ( .A(DP_OP_1196_128_7433_n60), .B(n20894), .C(
        n20893), .Y(n20895) );
  A2O1A1Ixp33_ASAP7_75t_SL U25909 ( .A1(n20894), .A2(DP_OP_1196_128_7433_n60), 
        .B(n20893), .C(n20895), .Y(u0_0_leon3x0_p0_iu_N5493) );
  INVxp33_ASAP7_75t_SRAM U25910 ( .A(n18437), .Y(n20896) );
  INVxp33_ASAP7_75t_SRAM U25911 ( .A(mult_x_1196_n552), .Y(n20897) );
  INVxp33_ASAP7_75t_SRAM U25912 ( .A(add_x_746_n12), .Y(n20898) );
  INVx1_ASAP7_75t_SL U25913 ( .A(u0_0_leon3x0_p0_iu_r_A__TICC_), .Y(n20900) );
  INVx1_ASAP7_75t_SL U25914 ( .A(n4388), .Y(n20904) );
  INVxp33_ASAP7_75t_SRAM U25915 ( .A(n28115), .Y(n20909) );
  INVx1_ASAP7_75t_SL U25916 ( .A(n32542), .Y(n20916) );
  INVx1_ASAP7_75t_SL U25917 ( .A(n31199), .Y(n20922) );
  INVxp33_ASAP7_75t_SRAM U25918 ( .A(n22433), .Y(n20923) );
  INVxp33_ASAP7_75t_SRAM U25919 ( .A(n22390), .Y(n20928) );
  INVxp33_ASAP7_75t_SRAM U25920 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__22_), 
        .Y(n20933) );
  INVxp33_ASAP7_75t_SRAM U25921 ( .A(uart1_r_BRATE__11_), .Y(n20942) );
  INVxp33_ASAP7_75t_SRAM U25922 ( .A(n22390), .Y(n20948) );
  INVxp33_ASAP7_75t_SRAM U25923 ( .A(n22390), .Y(n20953) );
  INVxp33_ASAP7_75t_SRAM U25924 ( .A(u0_0_leon3x0_p0_ici[12]), .Y(n20958) );
  INVx1_ASAP7_75t_SL U25925 ( .A(n31946), .Y(n20960) );
  INVxp33_ASAP7_75t_SRAM U25926 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__3_), 
        .Y(n20968) );
  INVxp33_ASAP7_75t_SRAM U25927 ( .A(u0_0_leon3x0_p0_iu_r_E__ET_), .Y(n20970)
         );
  INVxp33_ASAP7_75t_SRAM U25928 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__25_), .Y(
        n20972) );
  INVxp33_ASAP7_75t_SRAM U25929 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__11_), 
        .Y(n20974) );
  INVxp33_ASAP7_75t_SRAM U25930 ( .A(u0_0_leon3x0_p0_ici[4]), .Y(n20977) );
  INVxp33_ASAP7_75t_SRAM U25931 ( .A(u0_0_leon3x0_p0_ici[1]), .Y(n20980) );
  INVxp33_ASAP7_75t_SRAM U25932 ( .A(u0_0_leon3x0_p0_iu_r_M__MUL_), .Y(n20984)
         );
  INVx1_ASAP7_75t_SL U25933 ( .A(n20990), .Y(n20991) );
  INVxp33_ASAP7_75t_SRAM U25934 ( .A(u0_0_leon3x0_p0_iu_r_E__CWP__2_), .Y(
        n20996) );
  INVx1_ASAP7_75t_SL U25935 ( .A(n32008), .Y(n20998) );
  O2A1O1Ixp33_ASAP7_75t_SL U25936 ( .A1(n31652), .A2(n31653), .B(n21003), .C(
        n31656), .Y(n21004) );
  A2O1A1Ixp33_ASAP7_75t_SL U25937 ( .A1(n31656), .A2(n21002), .B(n21004), .C(
        n31663), .Y(n18176) );
  A2O1A1Ixp33_ASAP7_75t_SL U25938 ( .A1(n21024), .A2(n28802), .B(n21025), .C(
        n21026), .Y(n4592) );
  INVxp33_ASAP7_75t_SRAM U25939 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__25_), .Y(
        n21027) );
  INVxp33_ASAP7_75t_SRAM U25940 ( .A(n32705), .Y(n21035) );
  O2A1O1Ixp33_ASAP7_75t_SL U25941 ( .A1(n4715), .A2(n25997), .B(n21041), .C(
        n24695), .Y(n17455) );
  A2O1A1Ixp33_ASAP7_75t_SL U25942 ( .A1(u0_0_leon3x0_p0_divi[30]), .A2(n22410), 
        .B(n21051), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[31]) );
  INVx1_ASAP7_75t_SL U25943 ( .A(mult_x_1196_n347), .Y(n21060) );
  INVxp33_ASAP7_75t_SRAM U25944 ( .A(n31578), .Y(n21073) );
  INVxp33_ASAP7_75t_SRAM U25945 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__WICC_), .Y(
        n21074) );
  INVx1_ASAP7_75t_SL U25946 ( .A(n29630), .Y(n21081) );
  INVxp33_ASAP7_75t_SRAM U25947 ( .A(timer0_N60), .Y(n21090) );
  INVx1_ASAP7_75t_SL U25948 ( .A(n33062), .Y(n21096) );
  INVxp33_ASAP7_75t_SRAM U25949 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__22_), 
        .Y(n21099) );
  INVxp33_ASAP7_75t_SRAM U25950 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__13_), .Y(
        n21107) );
  INVxp33_ASAP7_75t_SRAM U25951 ( .A(n22390), .Y(n21115) );
  INVxp33_ASAP7_75t_SRAM U25952 ( .A(irqctrl0_r_ILEVEL__1_), .Y(n21118) );
  A2O1A1Ixp33_ASAP7_75t_SL U25953 ( .A1(n24602), .A2(n21121), .B(n24601), .C(
        n21122), .Y(n21123) );
  A2O1A1Ixp33_ASAP7_75t_SL U25954 ( .A1(n28174), .A2(n21123), .B(n21127), .C(
        n28151), .Y(n2882) );
  INVx1_ASAP7_75t_SL U25955 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__4_), 
        .Y(n21129) );
  INVxp33_ASAP7_75t_SRAM U25956 ( .A(n32683), .Y(n21130) );
  AOI21xp33_ASAP7_75t_SRAM U25957 ( .A1(n21129), .A2(n32682), .B(n22405), .Y(
        n21131) );
  O2A1O1Ixp33_ASAP7_75t_SL U25958 ( .A1(n21129), .A2(n32682), .B(n21131), .C(
        n21130), .Y(n32685) );
  INVxp33_ASAP7_75t_SRAM U25959 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__12_), 
        .Y(n21138) );
  INVxp33_ASAP7_75t_SRAM U25960 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__15_), 
        .Y(n21146) );
  INVxp33_ASAP7_75t_SRAM U25961 ( .A(u0_0_leon3x0_p0_iu_r_W__S__WIM__6_), .Y(
        n21148) );
  INVxp33_ASAP7_75t_SRAM U25962 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__11_), 
        .Y(n21150) );
  INVxp33_ASAP7_75t_SRAM U25963 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__4_), 
        .Y(n21152) );
  INVxp33_ASAP7_75t_SRAM U25964 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__9_), 
        .Y(n21160) );
  A2O1A1Ixp33_ASAP7_75t_SL U25965 ( .A1(n24647), .A2(
        u0_0_leon3x0_p0_iu_r_A__IMM__9_), .B(n21161), .C(n24495), .Y(n3651) );
  INVxp33_ASAP7_75t_SRAM U25966 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__RETT_), .Y(
        n21162) );
  A2O1A1Ixp33_ASAP7_75t_SL U25967 ( .A1(u0_0_leon3x0_p0_iu_r_E__CTRL__RETT_), 
        .A2(n32069), .B(n24678), .C(n21163), .Y(n3696) );
  A2O1A1Ixp33_ASAP7_75t_SL U25968 ( .A1(n24905), .A2(
        u0_0_leon3x0_p0_div0_r_CNT__2_), .B(u0_0_leon3x0_p0_div0_r_CNT__3_), 
        .C(n21164), .Y(n3721) );
  INVxp33_ASAP7_75t_SRAM U25969 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__1_), 
        .Y(n21165) );
  INVxp33_ASAP7_75t_SRAM U25970 ( .A(u0_0_dbgo_OPTYPE__2_), .Y(n21184) );
  INVxp33_ASAP7_75t_SRAM U25971 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__18_), 
        .Y(n21186) );
  INVxp33_ASAP7_75t_SRAM U25972 ( .A(u0_0_leon3x0_p0_iu_r_X__ICC__1_), .Y(
        n21193) );
  INVx1_ASAP7_75t_SL U25973 ( .A(n32008), .Y(n21195) );
  O2A1O1Ixp33_ASAP7_75t_SL U25974 ( .A1(n31818), .A2(n21211), .B(n25219), .C(
        n21212), .Y(n4493) );
  INVx1_ASAP7_75t_SL U25975 ( .A(n28053), .Y(n21213) );
  O2A1O1Ixp5_ASAP7_75t_SL U25976 ( .A1(uart1_r_TCNT__4_), .A2(n28052), .B(
        uart1_r_TCNT__5_), .C(n21213), .Y(n5590) );
  INVxp33_ASAP7_75t_SRAM U25977 ( .A(n22378), .Y(n21224) );
  INVxp33_ASAP7_75t_SRAM U25978 ( .A(n33026), .Y(n21241) );
  A2O1A1Ixp33_ASAP7_75t_SL U25979 ( .A1(apbi[14]), .A2(n29657), .B(n21246), 
        .C(n21248), .Y(n4735) );
  FAx1_ASAP7_75t_SL U25980 ( .A(n21251), .B(mult_x_1196_n855), .CI(n21252), 
        .CON(), .SN(mult_x_1196_n850) );
  INVx1_ASAP7_75t_SL U25981 ( .A(mult_x_1196_n855), .Y(n21253) );
  INVx1_ASAP7_75t_SL U25982 ( .A(mult_x_1196_n881), .Y(n21256) );
  INVxp33_ASAP7_75t_SRAM U25983 ( .A(mult_x_1196_n874), .Y(n21257) );
  NAND3xp33_ASAP7_75t_SL U25984 ( .A(add_x_735_n263), .B(n21259), .C(
        add_x_735_n264), .Y(n21260) );
  A2O1A1Ixp33_ASAP7_75t_SL U25985 ( .A1(n21259), .A2(add_x_735_n263), .B(
        add_x_735_n264), .C(n21260), .Y(u0_0_leon3x0_p0_iu_ex_jump_address_2_)
         );
  INVxp33_ASAP7_75t_SRAM U25986 ( .A(DP_OP_5187J1_124_3275_n304), .Y(n21268)
         );
  INVxp33_ASAP7_75t_SRAM U25987 ( .A(u0_0_leon3x0_p0_div0_b[0]), .Y(n21269) );
  NAND3xp33_ASAP7_75t_SL U25988 ( .A(n21269), .B(DP_OP_5187J1_124_3275_n305), 
        .C(n21268), .Y(n21270) );
  A2O1A1Ixp33_ASAP7_75t_SL U25989 ( .A1(DP_OP_5187J1_124_3275_n305), .A2(
        n21268), .B(n21269), .C(n21270), .Y(u0_0_leon3x0_p0_div0_addout_0_) );
  A2O1A1Ixp33_ASAP7_75t_SL U25990 ( .A1(n28827), .A2(n18890), .B(n21281), .C(
        n22578), .Y(n21282) );
  INVxp33_ASAP7_75t_SRAM U25991 ( .A(n31335), .Y(n21291) );
  INVxp33_ASAP7_75t_SRAM U25992 ( .A(n24694), .Y(n21308) );
  INVxp33_ASAP7_75t_SRAM U25993 ( .A(n22433), .Y(n21309) );
  INVxp33_ASAP7_75t_SRAM U25994 ( .A(n22433), .Y(n21312) );
  INVxp33_ASAP7_75t_SRAM U25995 ( .A(n32829), .Y(n21316) );
  INVxp33_ASAP7_75t_SRAM U25996 ( .A(n27501), .Y(n21320) );
  INVx1_ASAP7_75t_SL U25997 ( .A(n27509), .Y(n21322) );
  INVxp33_ASAP7_75t_SRAM U25998 ( .A(n22390), .Y(n21340) );
  A2O1A1Ixp33_ASAP7_75t_SL U25999 ( .A1(n28042), .A2(n24694), .B(n29374), .C(
        n21348), .Y(n2895) );
  INVx1_ASAP7_75t_SL U26000 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__25_), .Y(n21349) );
  INVx1_ASAP7_75t_SL U26001 ( .A(n3054), .Y(n21354) );
  INVxp33_ASAP7_75t_SRAM U26002 ( .A(n30180), .Y(n21357) );
  INVxp33_ASAP7_75t_SRAM U26003 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__13_), 
        .Y(n21360) );
  A2O1A1Ixp33_ASAP7_75t_SL U26004 ( .A1(n31598), .A2(n24684), .B(n31587), .C(
        n31586), .Y(n21364) );
  INVxp33_ASAP7_75t_SRAM U26005 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__15_), 
        .Y(n21370) );
  INVxp33_ASAP7_75t_SRAM U26006 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__11_), 
        .Y(n21377) );
  INVxp33_ASAP7_75t_SRAM U26007 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__7_), 
        .Y(n21379) );
  INVx1_ASAP7_75t_SL U26008 ( .A(n32018), .Y(n21385) );
  INVxp33_ASAP7_75t_SRAM U26009 ( .A(n24904), .Y(n21389) );
  INVx1_ASAP7_75t_SL U26010 ( .A(n30387), .Y(n21397) );
  INVxp33_ASAP7_75t_SRAM U26011 ( .A(u0_0_leon3x0_p0_iu_v_E__CWP__2_), .Y(
        n21405) );
  INVxp33_ASAP7_75t_SRAM U26012 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__17_), 
        .Y(n21407) );
  OAI21xp5_ASAP7_75t_SL U26013 ( .A1(mult_x_1196_n530), .A2(mult_x_1196_n247), 
        .B(n23229), .Y(n21413) );
  A2O1A1Ixp33_ASAP7_75t_SL U26014 ( .A1(mult_x_1196_n247), .A2(
        mult_x_1196_n530), .B(n21413), .C(n21414), .Y(n4229) );
  INVx1_ASAP7_75t_SL U26015 ( .A(mult_x_1196_n764), .Y(n21415) );
  A2O1A1Ixp33_ASAP7_75t_SL U26016 ( .A1(mult_x_1196_n765), .A2(n21415), .B(
        mult_x_1196_n766), .C(n21416), .Y(n21417) );
  INVxp33_ASAP7_75t_SRAM U26017 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__31_), 
        .Y(n21419) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U26018 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), 
        .A2(n27018), .B(n21434), .C(n30667), .Y(n21435) );
  INVxp33_ASAP7_75t_SRAM U26019 ( .A(n30774), .Y(n21440) );
  INVxp33_ASAP7_75t_SRAM U26020 ( .A(n29803), .Y(n21446) );
  A2O1A1Ixp33_ASAP7_75t_SL U26021 ( .A1(n28809), .A2(n21457), .B(n21458), .C(
        n21459), .Y(n4629) );
  A2O1A1Ixp33_ASAP7_75t_SL U26022 ( .A1(sr1_r_WS__3_), .A2(n21467), .B(n21471), 
        .C(n24694), .Y(n4725) );
  INVxp33_ASAP7_75t_SRAM U26023 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[1]), .Y(n21472) );
  A2O1A1Ixp33_ASAP7_75t_SL U26024 ( .A1(n31697), .A2(n21472), .B(n32719), .C(
        n21473), .Y(n21474) );
  INVxp33_ASAP7_75t_SRAM U26025 ( .A(n24043), .Y(n21540) );
  OAI21xp33_ASAP7_75t_SRAM U26026 ( .A1(n24043), .A2(n24062), .B(n22642), .Y(
        n21541) );
  A2O1A1Ixp33_ASAP7_75t_SL U26027 ( .A1(n24062), .A2(n21540), .B(n22642), .C(
        n21541), .Y(n24251) );
  INVx1_ASAP7_75t_SL U26028 ( .A(n23739), .Y(n21543) );
  INVx1_ASAP7_75t_SL U26029 ( .A(mult_x_1196_n2749), .Y(n21545) );
  A2O1A1Ixp33_ASAP7_75t_SL U26030 ( .A1(u0_0_leon3x0_p0_divi[29]), .A2(n22410), 
        .B(n21547), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[30]) );
  INVx1_ASAP7_75t_SL U26031 ( .A(add_x_735_n61), .Y(n21548) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U26032 ( .A1(n22227), .A2(n22538), .B(n24082), 
        .C(n23954), .Y(mult_x_1196_n2142) );
  A2O1A1Ixp33_ASAP7_75t_SL U26033 ( .A1(n22410), .A2(n21549), .B(n21550), .C(
        n24629), .Y(u0_0_leon3x0_p0_div0_b[32]) );
  INVx1_ASAP7_75t_SL U26034 ( .A(n29653), .Y(n21565) );
  INVx1_ASAP7_75t_SL U26035 ( .A(n32319), .Y(n21569) );
  INVxp33_ASAP7_75t_SRAM U26036 ( .A(n22390), .Y(n21581) );
  INVx1_ASAP7_75t_SL U26037 ( .A(n4643), .Y(n21584) );
  INVxp33_ASAP7_75t_SRAM U26038 ( .A(n22390), .Y(n21586) );
  INVxp33_ASAP7_75t_SRAM U26039 ( .A(n22390), .Y(n21596) );
  INVxp33_ASAP7_75t_SRAM U26040 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__4_), .Y(
        n21599) );
  INVxp33_ASAP7_75t_SRAM U26041 ( .A(n22390), .Y(n21606) );
  INVxp33_ASAP7_75t_SRAM U26042 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__0_), .Y(
        n21609) );
  INVx1_ASAP7_75t_SL U26043 ( .A(n21615), .Y(n2778) );
  INVxp33_ASAP7_75t_SRAM U26044 ( .A(n28182), .Y(n21617) );
  INVxp33_ASAP7_75t_SRAM U26045 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__9_), 
        .Y(n21626) );
  INVxp33_ASAP7_75t_SRAM U26046 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__7_), 
        .Y(n21628) );
  INVxp33_ASAP7_75t_SRAM U26047 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__29_), 
        .Y(n21631) );
  INVxp33_ASAP7_75t_SRAM U26048 ( .A(n22390), .Y(n21633) );
  INVxp33_ASAP7_75t_SRAM U26049 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__15_), 
        .Y(n21636) );
  INVxp33_ASAP7_75t_SRAM U26050 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__29_), 
        .Y(n21638) );
  INVxp33_ASAP7_75t_SRAM U26051 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__4_), 
        .Y(n21640) );
  INVx1_ASAP7_75t_SL U26052 ( .A(n21643), .Y(n21644) );
  INVxp33_ASAP7_75t_SRAM U26053 ( .A(n30395), .Y(n21654) );
  INVxp33_ASAP7_75t_SRAM U26054 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__6_), .Y(
        n21667) );
  INVxp33_ASAP7_75t_SRAM U26055 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__4_), 
        .Y(n21669) );
  INVxp33_ASAP7_75t_SRAM U26056 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__0_), 
        .Y(n21672) );
  A2O1A1Ixp33_ASAP7_75t_SL U26057 ( .A1(mult_x_1196_n225), .A2(
        mult_x_1196_n296), .B(n21675), .C(n21676), .Y(n4185) );
  A2O1A1Ixp33_ASAP7_75t_SL U26058 ( .A1(n18984), .A2(n22999), .B(n24646), .C(
        n21678), .Y(n4309) );
  INVxp33_ASAP7_75t_SRAM U26059 ( .A(u0_0_leon3x0_p0_div0_r_ZERO2_), .Y(n21679) );
  INVxp33_ASAP7_75t_SRAM U26060 ( .A(n31456), .Y(n21685) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U26061 ( .A1(n31458), .A2(n21686), .B(n31574), 
        .C(n21687), .Y(n21688) );
  INVxp33_ASAP7_75t_SRAM U26062 ( .A(n31568), .Y(n21693) );
  INVxp33_ASAP7_75t_SRAM U26063 ( .A(apb0_r_STATE__0_), .Y(n21698) );
  INVxp33_ASAP7_75t_SRAM U26064 ( .A(n32041), .Y(n21699) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U26065 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PV_), 
        .A2(n30681), .B(n30684), .C(n25723), .Y(n21704) );
  INVxp33_ASAP7_75t_SRAM U26066 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__10_), 
        .Y(n21705) );
  INVxp33_ASAP7_75t_SRAM U26067 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__5_), 
        .Y(n21711) );
  A2O1A1Ixp33_ASAP7_75t_SL U26068 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[26]), .B(n21713), .C(n31638), .Y(n4574) );
  INVxp33_ASAP7_75t_SRAM U26069 ( .A(uart1_r_LOOPB_), .Y(n21728) );
  A2O1A1Ixp33_ASAP7_75t_SL U26070 ( .A1(n21731), .A2(n21732), .B(n32452), .C(
        n31937), .Y(n21733) );
  A2O1A1Ixp33_ASAP7_75t_SL U26071 ( .A1(n21734), .A2(u0_0_leon3x0_p0_ici[62]), 
        .B(n21735), .C(n21736), .Y(n21737) );
  A2O1A1Ixp33_ASAP7_75t_SL U26072 ( .A1(n32689), .A2(n21733), .B(n21737), .C(
        n24684), .Y(n4730) );
  INVx1_ASAP7_75t_SL U26073 ( .A(mult_x_1196_n844), .Y(n21750) );
  INVxp33_ASAP7_75t_SRAM U26074 ( .A(n24043), .Y(n21751) );
  OAI21xp33_ASAP7_75t_SRAM U26075 ( .A1(n24043), .A2(n24045), .B(n23978), .Y(
        n21752) );
  A2O1A1Ixp33_ASAP7_75t_SL U26076 ( .A1(n24045), .A2(n21751), .B(n23978), .C(
        n21752), .Y(n21753) );
  FAx1_ASAP7_75t_SL U26077 ( .A(n21749), .B(n21750), .CI(n21753), .CON(), .SN(
        mult_x_1196_n839) );
  A2O1A1Ixp33_ASAP7_75t_SL U26078 ( .A1(u0_0_leon3x0_p0_divi[28]), .A2(n22410), 
        .B(n21754), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[29]) );
  INVxp33_ASAP7_75t_SRAM U26079 ( .A(mult_x_1196_n316), .Y(n21755) );
  INVxp33_ASAP7_75t_SRAM U26080 ( .A(n31714), .Y(n21771) );
  INVxp33_ASAP7_75t_SRAM U26081 ( .A(n32170), .Y(n21774) );
  INVx1_ASAP7_75t_SL U26082 ( .A(n31939), .Y(n21798) );
  INVxp33_ASAP7_75t_SRAM U26083 ( .A(n22433), .Y(n21799) );
  INVxp33_ASAP7_75t_SRAM U26084 ( .A(n22433), .Y(n21802) );
  INVx1_ASAP7_75t_SL U26085 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__30_), .Y(n21808) );
  INVxp33_ASAP7_75t_SRAM U26086 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__24_), 
        .Y(n21811) );
  INVxp33_ASAP7_75t_SRAM U26087 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__22_), 
        .Y(n21814) );
  INVxp33_ASAP7_75t_SRAM U26088 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__13_), 
        .Y(n21825) );
  INVxp33_ASAP7_75t_SRAM U26089 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__3_), .Y(
        n21829) );
  INVxp33_ASAP7_75t_SRAM U26090 ( .A(n31411), .Y(n21836) );
  INVxp33_ASAP7_75t_SRAM U26091 ( .A(irqctrl0_r_ILEVEL__12_), .Y(n21837) );
  INVx1_ASAP7_75t_SL U26092 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__26_), .Y(n21839) );
  INVxp33_ASAP7_75t_SRAM U26093 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__14_), 
        .Y(n21853) );
  INVxp33_ASAP7_75t_SRAM U26094 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__15_), 
        .Y(n21855) );
  INVxp33_ASAP7_75t_SRAM U26095 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__16_), 
        .Y(n21857) );
  INVxp33_ASAP7_75t_SRAM U26096 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__28_), 
        .Y(n21861) );
  INVxp33_ASAP7_75t_SRAM U26097 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__9_), 
        .Y(n21878) );
  INVxp33_ASAP7_75t_SRAM U26098 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__7_), 
        .Y(n21880) );
  INVxp33_ASAP7_75t_SRAM U26099 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__6_), 
        .Y(n21882) );
  INVx1_ASAP7_75t_SL U26100 ( .A(u0_0_leon3x0_p0_div0_r_CNT__4_), .Y(n21886)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U26101 ( .A1(n24909), .A2(n31655), .B(n24908), .C(
        n21887), .Y(n3726) );
  INVxp33_ASAP7_75t_SRAM U26102 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__29_), 
        .Y(n21888) );
  INVxp33_ASAP7_75t_SRAM U26103 ( .A(n30957), .Y(n21890) );
  INVxp33_ASAP7_75t_SRAM U26104 ( .A(u0_0_leon3x0_p0_iu_v_M__MUL_), .Y(n21891)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U26105 ( .A1(n25231), .A2(n21890), .B(n24680), .C(
        n21892), .Y(n3780) );
  A2O1A1Ixp33_ASAP7_75t_SL U26106 ( .A1(n33054), .A2(n21902), .B(n24680), .C(
        n21903), .Y(n3914) );
  INVxp33_ASAP7_75t_SRAM U26107 ( .A(n22390), .Y(n21907) );
  INVxp33_ASAP7_75t_SRAM U26108 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__18_), 
        .Y(n21916) );
  INVxp33_ASAP7_75t_SRAM U26109 ( .A(n24646), .Y(n21918) );
  OAI21xp5_ASAP7_75t_SL U26110 ( .A1(mult_x_1196_n559), .A2(mult_x_1196_n250), 
        .B(n22421), .Y(n21920) );
  A2O1A1Ixp33_ASAP7_75t_SL U26111 ( .A1(mult_x_1196_n250), .A2(
        mult_x_1196_n559), .B(n21920), .C(n21921), .Y(n4235) );
  A2O1A1Ixp33_ASAP7_75t_SL U26112 ( .A1(n29818), .A2(n30679), .B(n30944), .C(
        n21923), .Y(n4326) );
  INVx1_ASAP7_75t_SL U26113 ( .A(n30203), .Y(n21935) );
  O2A1O1Ixp33_ASAP7_75t_SL U26114 ( .A1(n30595), .A2(n21944), .B(n21945), .C(
        n21946), .Y(n4551) );
  A2O1A1Ixp33_ASAP7_75t_SL U26115 ( .A1(n24648), .A2(
        u0_0_leon3x0_p0_iu_r_A__WOVF_), .B(n21947), .C(n31439), .Y(n4569) );
  INVx1_ASAP7_75t_SL U26116 ( .A(n29804), .Y(n21952) );
  INVxp33_ASAP7_75t_SRAM U26117 ( .A(n28186), .Y(n21966) );
  INVxp33_ASAP7_75t_SRAM U26118 ( .A(n29948), .Y(n21967) );
  INVxp33_ASAP7_75t_SRAM U26119 ( .A(n31838), .Y(n21968) );
  INVxp33_ASAP7_75t_SRAM U26120 ( .A(n32791), .Y(n21969) );
  A2O1A1Ixp33_ASAP7_75t_SL U26121 ( .A1(n32827), .A2(n21969), .B(n31752), .C(
        n32789), .Y(n21970) );
  INVxp33_ASAP7_75t_SRAM U26122 ( .A(n32824), .Y(n21971) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U26123 ( .A1(n32723), .A2(n32787), .B(n21970), 
        .C(n21971), .Y(n4727) );
  INVx1_ASAP7_75t_SL U26124 ( .A(n29881), .Y(n21976) );
  A2O1A1Ixp33_ASAP7_75t_SL U26125 ( .A1(timer0_vtimers_1__IRQEN_), .A2(n30739), 
        .B(timer0_vtimers_1__IRQPEN_), .C(n21978), .Y(n4769) );
  INVxp33_ASAP7_75t_SRAM U26126 ( .A(n31249), .Y(n21984) );
  INVxp33_ASAP7_75t_SRAM U26127 ( .A(n30873), .Y(n22036) );
  HAxp5_ASAP7_75t_SL U26128 ( .A(n24056), .B(n22642), .CON(), .SN(n22041) );
  XOR2xp5_ASAP7_75t_SL U26129 ( .A(mult_x_1196_n1054), .B(mult_x_1196_n1052), 
        .Y(n23283) );
  FAx1_ASAP7_75t_SL U26130 ( .A(mult_x_1196_n850), .B(n22042), .CI(
        mult_x_1196_n853), .CON(), .SN(mult_x_1196_n848) );
  INVx1_ASAP7_75t_SL U26131 ( .A(mult_x_1196_n853), .Y(n22043) );
  A2O1A1Ixp33_ASAP7_75t_SL U26132 ( .A1(n22481), .A2(n22412), .B(
        mult_x_1196_n2771), .C(n22043), .Y(n22044) );
  A2O1A1Ixp33_ASAP7_75t_SL U26133 ( .A1(n22042), .A2(mult_x_1196_n853), .B(
        mult_x_1196_n850), .C(n22044), .Y(mult_x_1196_n847) );
  A2O1A1Ixp33_ASAP7_75t_SL U26134 ( .A1(u0_0_leon3x0_p0_divi[20]), .A2(n22410), 
        .B(n22045), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL U26135 ( .A1(u0_0_leon3x0_p0_divi[26]), .A2(n22410), 
        .B(n22046), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[27]) );
  INVx1_ASAP7_75t_SL U26136 ( .A(mult_x_1196_n324), .Y(n22049) );
  INVx1_ASAP7_75t_SL U26137 ( .A(n27513), .Y(n22050) );
  INVx1_ASAP7_75t_SL U26138 ( .A(n29991), .Y(n22051) );
  INVx1_ASAP7_75t_SL U26139 ( .A(n31556), .Y(n22052) );
  INVx1_ASAP7_75t_SL U26140 ( .A(n22468), .Y(n22054) );
  INVx1_ASAP7_75t_SL U26141 ( .A(n29406), .Y(n22056) );
  INVx1_ASAP7_75t_SL U26142 ( .A(n32319), .Y(n22061) );
  INVx1_ASAP7_75t_SL U26143 ( .A(n32542), .Y(n22065) );
  INVx1_ASAP7_75t_SL U26144 ( .A(n2236), .Y(n22070) );
  INVx1_ASAP7_75t_SL U26145 ( .A(n25996), .Y(n22072) );
  INVx1_ASAP7_75t_SL U26146 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__12_), .Y(
        n22078) );
  INVx1_ASAP7_75t_SL U26147 ( .A(u0_0_leon3x0_p0_iu_r_A__RFA2__5_), .Y(n22082)
         );
  INVx1_ASAP7_75t_SL U26148 ( .A(n2851), .Y(n22084) );
  INVx1_ASAP7_75t_SL U26149 ( .A(n24694), .Y(n22086) );
  OAI21xp33_ASAP7_75t_SL U26150 ( .A1(n29356), .A2(n22086), .B(n29357), .Y(
        n22087) );
  A2O1A1Ixp33_ASAP7_75t_SL U26151 ( .A1(n24694), .A2(n29356), .B(n29357), .C(
        n22087), .Y(n2896) );
  INVx1_ASAP7_75t_SL U26152 ( .A(sr1_r_MCFG1__IOWIDTH__0_), .Y(n22088) );
  INVx1_ASAP7_75t_SL U26153 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__2_), 
        .Y(n22094) );
  A2O1A1Ixp33_ASAP7_75t_SL U26154 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__2_), .A2(n30166), .B(n22380), 
        .C(n22096), .Y(n22097) );
  INVx1_ASAP7_75t_SL U26155 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__17_), .Y(
        n22098) );
  INVx1_ASAP7_75t_SL U26156 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__18_), .Y(
        n22100) );
  INVx1_ASAP7_75t_SL U26157 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__19_), .Y(
        n22102) );
  INVx1_ASAP7_75t_SL U26158 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__21_), .Y(
        n22104) );
  INVx1_ASAP7_75t_SL U26159 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__24_), .Y(
        n22106) );
  INVx1_ASAP7_75t_SL U26160 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__26_), .Y(
        n22108) );
  INVx1_ASAP7_75t_SL U26161 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__27_), .Y(
        n22110) );
  INVx1_ASAP7_75t_SL U26162 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__30_), .Y(
        n22112) );
  INVx1_ASAP7_75t_SL U26163 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__31_), .Y(
        n22114) );
  INVx1_ASAP7_75t_SL U26164 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__3_), .Y(
        n22116) );
  INVx1_ASAP7_75t_SL U26165 ( .A(n30114), .Y(n22120) );
  OAI21xp33_ASAP7_75t_SL U26166 ( .A1(mult_x_1196_n245), .A2(n23230), .B(
        n23229), .Y(n22129) );
  A2O1A1Ixp33_ASAP7_75t_SL U26167 ( .A1(mult_x_1196_n245), .A2(n18403), .B(
        n22129), .C(n22128), .Y(n4225) );
  O2A1O1Ixp33_ASAP7_75t_SL U26168 ( .A1(n31818), .A2(n31817), .B(n22135), .C(
        n31816), .Y(n22136) );
  INVx1_ASAP7_75t_SL U26169 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__8_), .Y(
        n22137) );
  INVx1_ASAP7_75t_SL U26170 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__31_), .Y(
        n22147) );
  INVx1_ASAP7_75t_SL U26171 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__28_), .Y(n22154) );
  INVx1_ASAP7_75t_SL U26172 ( .A(n22379), .Y(n22171) );
  O2A1O1Ixp33_ASAP7_75t_SL U26173 ( .A1(n29744), .A2(n29743), .B(
        irqctrl0_r_IPEND__8_), .C(n29745), .Y(n22183) );
  A2O1A1Ixp33_ASAP7_75t_SL U26174 ( .A1(timer0_vtimers_1__IRQEN_), .A2(
        timer0_gpto_TICK__1_), .B(n22184), .C(n24694), .Y(n15075) );
  INVx1_ASAP7_75t_SL U26175 ( .A(n4741), .Y(n22187) );
  INVx1_ASAP7_75t_SL U26176 ( .A(timer0_r_SCALER__7_), .Y(n22200) );
  INVx1_ASAP7_75t_SL U26177 ( .A(timer0_r_RELOAD__7_), .Y(n22203) );
  NAND2x1p5_ASAP7_75t_SL U26178 ( .A(n25144), .B(n25143), .Y(n22206) );
  INVx11_ASAP7_75t_SL U26179 ( .A(n22698), .Y(n23964) );
  INVx6_ASAP7_75t_SL U26180 ( .A(n24042), .Y(n24043) );
  INVx5_ASAP7_75t_SL U26181 ( .A(n23995), .Y(n23997) );
  INVx3_ASAP7_75t_SL U26182 ( .A(n23516), .Y(n23995) );
  NOR2xp33_ASAP7_75t_SL U26183 ( .A(n23833), .B(n24688), .Y(n23832) );
  AND2x2_ASAP7_75t_SL U26184 ( .A(n23686), .B(n23685), .Y(n22207) );
  MAJIxp5_ASAP7_75t_SL U26185 ( .A(mult_x_1196_n1805), .B(n23709), .C(n18415), 
        .Y(n22210) );
  INVx2_ASAP7_75t_SL U26186 ( .A(n23757), .Y(n23988) );
  INVx4_ASAP7_75t_SL U26187 ( .A(n23757), .Y(n22248) );
  INVx3_ASAP7_75t_SL U26188 ( .A(n23757), .Y(n24106) );
  XOR2x2_ASAP7_75t_SL U26189 ( .A(n24301), .B(n22783), .Y(n22212) );
  OA21x2_ASAP7_75t_SL U26190 ( .A1(mult_x_1196_n347), .A2(mult_x_1196_n355), 
        .B(mult_x_1196_n348), .Y(n22214) );
  OR2x2_ASAP7_75t_SL U26191 ( .A(mult_x_1196_n2994), .B(n23644), .Y(n22215) );
  AND2x4_ASAP7_75t_SL U26192 ( .A(n22266), .B(n23770), .Y(n22216) );
  OA21x2_ASAP7_75t_SL U26193 ( .A1(n29861), .A2(n22402), .B(n29860), .Y(n22217) );
  NAND2xp5_ASAP7_75t_SL U26194 ( .A(mult_x_1196_n1298), .B(mult_x_1196_n1327), 
        .Y(n22218) );
  AO21x1_ASAP7_75t_SL U26195 ( .A1(n23926), .A2(n23393), .B(n23389), .Y(n22219) );
  INVx1_ASAP7_75t_SL U26196 ( .A(n22248), .Y(n23159) );
  XOR2x2_ASAP7_75t_SL U26197 ( .A(n22525), .B(n22524), .Y(n22221) );
  INVx2_ASAP7_75t_SL U26198 ( .A(mult_x_1196_n330), .Y(n23683) );
  XOR2xp5_ASAP7_75t_SL U26199 ( .A(n23077), .B(mult_x_1196_n2698), .Y(n22222)
         );
  OR2x4_ASAP7_75t_SL U26200 ( .A(n32198), .B(n31572), .Y(n32729) );
  INVx1_ASAP7_75t_SL U26201 ( .A(mult_x_1196_n457), .Y(n23732) );
  AND2x2_ASAP7_75t_SL U26202 ( .A(mult_x_1196_n368), .B(n24279), .Y(n22223) );
  INVx6_ASAP7_75t_SL U26203 ( .A(n33053), .Y(n22386) );
  INVx8_ASAP7_75t_SL U26204 ( .A(n24425), .Y(n22376) );
  OR2x2_ASAP7_75t_SL U26205 ( .A(n23835), .B(n18884), .Y(n22224) );
  BUFx3_ASAP7_75t_SL U26206 ( .A(n23953), .Y(add_x_735_A_2_) );
  BUFx3_ASAP7_75t_SL U26207 ( .A(n23951), .Y(n22933) );
  OR2x4_ASAP7_75t_SL U26208 ( .A(n25080), .B(n32141), .Y(n30007) );
  INVx11_ASAP7_75t_SL U26209 ( .A(n30007), .Y(n22375) );
  NOR2x1p5_ASAP7_75t_SL U26210 ( .A(n4316), .B(n4318), .Y(n33058) );
  BUFx10_ASAP7_75t_SL U26211 ( .A(n33058), .Y(n24681) );
  INVx8_ASAP7_75t_SL U26212 ( .A(n24646), .Y(n22421) );
  BUFx8_ASAP7_75t_SL U26213 ( .A(n33058), .Y(n22379) );
  BUFx6f_ASAP7_75t_SL U26214 ( .A(rstn), .Y(n24694) );
  INVx6_ASAP7_75t_SL U26215 ( .A(rstn), .Y(n24695) );
  INVx8_ASAP7_75t_SL U26216 ( .A(n24684), .Y(n22380) );
  INVx5_ASAP7_75t_SL U26217 ( .A(n4818), .Y(n24684) );
  INVx1_ASAP7_75t_SL U26218 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__19_), .Y(n23845)
         );
  INVx1_ASAP7_75t_SL U26219 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__16_), .Y(n23841)
         );
  INVx1_ASAP7_75t_SL U26220 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__13_), .Y(n23846)
         );
  INVx1_ASAP7_75t_SL U26221 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__24_), .Y(n23836)
         );
  INVx1_ASAP7_75t_SL U26222 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__15_), .Y(n23840)
         );
  INVx1_ASAP7_75t_SL U26223 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__6_), .Y(n23847)
         );
  INVx1_ASAP7_75t_SL U26224 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__7_), .Y(n23848)
         );
  INVx1_ASAP7_75t_SL U26225 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__25_), .Y(n23842)
         );
  INVx1_ASAP7_75t_SL U26226 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__27_), .Y(n23843)
         );
  INVx1_ASAP7_75t_SL U26227 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__9_), .Y(n23839)
         );
  NAND2x1p5_ASAP7_75t_SL U26228 ( .A(n23838), .B(n30603), .Y(
        u0_0_leon3x0_p0_muli[15]) );
  XNOR2x1_ASAP7_75t_SL U26229 ( .A(n23657), .B(n23643), .Y(mult_x_1196_n3117)
         );
  NOR2xp33_ASAP7_75t_SL U26230 ( .A(mult_x_1196_n2761), .B(n24041), .Y(n23854)
         );
  OAI22x1_ASAP7_75t_SL U26231 ( .A1(n24035), .A2(mult_x_1196_n2835), .B1(
        n22251), .B2(mult_x_1196_n2834), .Y(mult_x_1196_n2269) );
  XOR2x1_ASAP7_75t_SL U26232 ( .A(mult_x_1196_n2327), .B(mult_x_1196_n2269), 
        .Y(n24129) );
  XNOR2x2_ASAP7_75t_SL U26233 ( .A(n24073), .B(n23971), .Y(mult_x_1196_n2868)
         );
  HB1xp67_ASAP7_75t_SL U26234 ( .A(n23337), .Y(n22591) );
  OAI22xp5_ASAP7_75t_SL U26235 ( .A1(mult_x_1196_n2936), .A2(n24022), .B1(
        mult_x_1196_n2935), .B2(n24020), .Y(mult_x_1196_n2364) );
  NOR2xp33_ASAP7_75t_SL U26236 ( .A(n18532), .B(n25085), .Y(n28880) );
  NOR2xp33_ASAP7_75t_SL U26237 ( .A(n18532), .B(n25083), .Y(n28926) );
  INVxp33_ASAP7_75t_SRAM U26238 ( .A(mult_x_1196_n565), .Y(mult_x_1196_n563)
         );
  NAND4xp75_ASAP7_75t_SL U26239 ( .A(n25352), .B(n25354), .C(n25355), .D(
        n25353), .Y(n29869) );
  OAI22x1_ASAP7_75t_SL U26240 ( .A1(n24035), .A2(mult_x_1196_n2834), .B1(
        n22251), .B2(mult_x_1196_n2833), .Y(mult_x_1196_n2268) );
  NOR2x1_ASAP7_75t_SL U26241 ( .A(mult_x_1196_n3259), .B(n23982), .Y(n23114)
         );
  XNOR2xp5_ASAP7_75t_SL U26242 ( .A(n22285), .B(n25644), .Y(n22226) );
  XNOR2x2_ASAP7_75t_SL U26243 ( .A(n24056), .B(n23957), .Y(mult_x_1196_n3191)
         );
  XNOR2x1_ASAP7_75t_SL U26244 ( .A(n22591), .B(n23336), .Y(mult_x_1196_n1443)
         );
  XNOR2x2_ASAP7_75t_SL U26245 ( .A(n24073), .B(n23965), .Y(mult_x_1196_n3004)
         );
  XNOR2x2_ASAP7_75t_SL U26246 ( .A(n24050), .B(n22394), .Y(mult_x_1196_n3083)
         );
  XOR2x2_ASAP7_75t_SL U26247 ( .A(n18534), .B(n23479), .Y(mult_x_1196_n2786)
         );
  XNOR2x2_ASAP7_75t_SL U26248 ( .A(n24059), .B(n23975), .Y(mult_x_1196_n2752)
         );
  XNOR2x2_ASAP7_75t_SL U26249 ( .A(n24059), .B(add_x_735_A_10_), .Y(
        mult_x_1196_n3126) );
  XNOR2x2_ASAP7_75t_SL U26250 ( .A(n24059), .B(n23971), .Y(mult_x_1196_n2854)
         );
  XNOR2x2_ASAP7_75t_SL U26251 ( .A(n24059), .B(n22642), .Y(mult_x_1196_n2718)
         );
  XNOR2x2_ASAP7_75t_SL U26252 ( .A(n24059), .B(n23089), .Y(mult_x_1196_n2888)
         );
  XNOR2x2_ASAP7_75t_SL U26253 ( .A(n24059), .B(n23964), .Y(mult_x_1196_n3024)
         );
  XNOR2x2_ASAP7_75t_SL U26254 ( .A(n24059), .B(n23952), .Y(mult_x_1196_n3262)
         );
  XNOR2x2_ASAP7_75t_SL U26255 ( .A(n24059), .B(n22394), .Y(mult_x_1196_n3092)
         );
  XNOR2x2_ASAP7_75t_SL U26256 ( .A(n24059), .B(n23957), .Y(mult_x_1196_n3194)
         );
  XOR2x2_ASAP7_75t_SL U26257 ( .A(n24059), .B(n23397), .Y(mult_x_1196_n3160)
         );
  XOR2x2_ASAP7_75t_SL U26258 ( .A(n23972), .B(n24071), .Y(mult_x_1196_n2798)
         );
  BUFx6f_ASAP7_75t_SL U26259 ( .A(u0_0_leon3x0_p0_muli[16]), .Y(n24071) );
  NOR3x1_ASAP7_75t_SL U26260 ( .A(timer0_N90), .B(timer0_N89), .C(timer0_N91), 
        .Y(n24373) );
  NOR2x1_ASAP7_75t_SL U26261 ( .A(n5061), .B(n2844), .Y(timer0_N90) );
  BUFx10_ASAP7_75t_SL U26262 ( .A(u0_0_leon3x0_p0_muli[11]), .Y(n22227) );
  OAI22x1_ASAP7_75t_SL U26263 ( .A1(mult_x_1196_n3081), .A2(n18920), .B1(
        mult_x_1196_n3080), .B2(n18435), .Y(mult_x_1196_n2508) );
  XNOR2x1_ASAP7_75t_SL U26264 ( .A(n24048), .B(n22394), .Y(mult_x_1196_n3081)
         );
  BUFx6f_ASAP7_75t_SL U26265 ( .A(u0_0_leon3x0_p0_muli[36]), .Y(n24045) );
  NAND2x1p5_ASAP7_75t_SL U26266 ( .A(n23555), .B(n25124), .Y(
        u0_0_leon3x0_p0_muli[36]) );
  BUFx6f_ASAP7_75t_SL U26267 ( .A(u0_0_leon3x0_p0_muli[34]), .Y(n24049) );
  BUFx6f_ASAP7_75t_SL U26268 ( .A(u0_0_leon3x0_p0_muli[21]), .Y(n24065) );
  XNOR2x2_ASAP7_75t_SL U26269 ( .A(n24073), .B(n22395), .Y(mult_x_1196_n2834)
         );
  INVx2_ASAP7_75t_SL U26270 ( .A(mult_x_1196_n2323), .Y(n23800) );
  BUFx12f_ASAP7_75t_SL U26271 ( .A(u0_0_leon3x0_p0_muli[13]), .Y(n24074) );
  BUFx6f_ASAP7_75t_SL U26272 ( .A(u0_0_leon3x0_p0_muli[31]), .Y(n24053) );
  XOR2x1_ASAP7_75t_SL U26273 ( .A(n24069), .B(n22918), .Y(mult_x_1196_n2830)
         );
  XNOR2x1_ASAP7_75t_SL U26274 ( .A(n24060), .B(n23969), .Y(mult_x_1196_n2923)
         );
  XNOR2x1_ASAP7_75t_SL U26275 ( .A(n18927), .B(n24044), .Y(mult_x_1196_n3247)
         );
  BUFx6f_ASAP7_75t_SL U26276 ( .A(add_x_735_n1), .Y(n22228) );
  XNOR2xp5_ASAP7_75t_SL U26277 ( .A(n24061), .B(n23969), .Y(mult_x_1196_n2924)
         );
  XNOR2xp5_ASAP7_75t_SL U26278 ( .A(n24061), .B(n23957), .Y(mult_x_1196_n3196)
         );
  BUFx6f_ASAP7_75t_SL U26279 ( .A(u0_0_leon3x0_p0_muli[24]), .Y(n24061) );
  XNOR2xp5_ASAP7_75t_SL U26280 ( .A(n24059), .B(n23969), .Y(mult_x_1196_n2922)
         );
  BUFx6f_ASAP7_75t_SL U26281 ( .A(u0_0_leon3x0_p0_muli[20]), .Y(n24066) );
  OAI22x1_ASAP7_75t_SL U26282 ( .A1(n23830), .A2(n25768), .B1(n18997), .B2(
        n23845), .Y(u0_0_leon3x0_p0_muli[27]) );
  OAI21xp33_ASAP7_75t_SL U26283 ( .A1(n11260), .A2(n24695), .B(n24694), .Y(
        n22229) );
  INVx1_ASAP7_75t_SL U26284 ( .A(n22231), .Y(n22230) );
  INVx1_ASAP7_75t_SL U26285 ( .A(n22234), .Y(n22233) );
  NOR2xp33_ASAP7_75t_SL U26286 ( .A(n17271), .B(n17270), .Y(n22234) );
  TIEHIx1_ASAP7_75t_SL U26287 ( .H(rf_ce_w) );
  TIEHIx1_ASAP7_75t_SL U26288 ( .H(dt_ce) );
  TIEHIx1_ASAP7_75t_SL U26289 ( .H(dc_ce) );
  TIEHIx1_ASAP7_75t_SL U26290 ( .H(it_ce) );
  TIEHIx1_ASAP7_75t_SL U26291 ( .H(ic_ce) );
  TIEHIx1_ASAP7_75t_SL U26292 ( .H(ramsn[4]) );
  INVx1_ASAP7_75t_SL U26293 ( .A(n22242), .Y(mult_x_1196_n657) );
  OAI22x1_ASAP7_75t_SL U26294 ( .A1(mult_x_1196_n3192), .A2(n23989), .B1(
        n24106), .B2(mult_x_1196_n3191), .Y(n22243) );
  MAJIxp5_ASAP7_75t_SL U26295 ( .A(mult_x_1196_n2492), .B(n22243), .C(
        mult_x_1196_n2584), .Y(mult_x_1196_n1790) );
  XNOR2xp5_ASAP7_75t_SL U26296 ( .A(mult_x_1196_n2684), .B(n22244), .Y(n23367)
         );
  OAI22xp5_ASAP7_75t_SL U26297 ( .A1(mult_x_1196_n3100), .A2(n18919), .B1(
        n22756), .B2(mult_x_1196_n3099), .Y(n22244) );
  NAND2xp33_ASAP7_75t_SL U26298 ( .A(mult_x_1196_n1973), .B(n22245), .Y(n23795) );
  INVxp67_ASAP7_75t_SL U26299 ( .A(n23798), .Y(n22245) );
  XNOR2x2_ASAP7_75t_SL U26300 ( .A(n22457), .B(n18298), .Y(n23798) );
  INVx1_ASAP7_75t_SL U26301 ( .A(mult_x_1196_n2141), .Y(n23253) );
  NAND2xp5_ASAP7_75t_SL U26302 ( .A(mult_x_1196_n2083), .B(mult_x_1196_n2082), 
        .Y(mult_x_1196_n758) );
  XNOR2xp5_ASAP7_75t_SL U26303 ( .A(mult_x_1196_n2087), .B(n22246), .Y(
        mult_x_1196_n2082) );
  XOR2xp5_ASAP7_75t_SL U26304 ( .A(mult_x_1196_n2141), .B(n24135), .Y(n22246)
         );
  XNOR2x1_ASAP7_75t_SL U26305 ( .A(n23415), .B(n23979), .Y(n24042) );
  INVx2_ASAP7_75t_SL U26306 ( .A(n23979), .Y(n23977) );
  OA21x2_ASAP7_75t_SL U26307 ( .A1(mult_x_1196_n3202), .A2(n22802), .B(n22315), 
        .Y(n22249) );
  INVx6_ASAP7_75t_SL U26308 ( .A(n23645), .Y(n24011) );
  OAI22xp5_ASAP7_75t_SL U26309 ( .A1(mult_x_1196_n2798), .A2(n24038), .B1(
        mult_x_1196_n2797), .B2(n22391), .Y(n22250) );
  NOR2xp33_ASAP7_75t_SL U26310 ( .A(mult_x_1196_n3035), .B(n24009), .Y(n23130)
         );
  XOR2xp5_ASAP7_75t_SL U26311 ( .A(n23511), .B(n23509), .Y(n22338) );
  BUFx10_ASAP7_75t_SL U26312 ( .A(n24033), .Y(n22251) );
  INVxp33_ASAP7_75t_SRAM U26313 ( .A(n24033), .Y(n24032) );
  HB1xp67_ASAP7_75t_SL U26314 ( .A(n18991), .Y(n22252) );
  INVxp33_ASAP7_75t_SRAM U26315 ( .A(mult_x_1196_n648), .Y(n22254) );
  NAND2xp5_ASAP7_75t_SL U26316 ( .A(mult_x_1196_n6), .B(mult_x_1196_n3330), 
        .Y(n22255) );
  NAND2xp5_ASAP7_75t_SL U26317 ( .A(mult_x_1196_n6), .B(mult_x_1196_n3330), 
        .Y(mult_x_1196_n9) );
  XOR2x1_ASAP7_75t_SL U26318 ( .A(n22864), .B(u0_0_leon3x0_p0_muli[38]), .Y(
        mult_x_1196_n3330) );
  NAND2x2_ASAP7_75t_SL U26319 ( .A(n24208), .B(n24209), .Y(mult_x_1196_n784)
         );
  INVx2_ASAP7_75t_SL U26320 ( .A(mult_x_1196_n933), .Y(n24209) );
  OAI21x1_ASAP7_75t_SL U26321 ( .A1(mult_x_1196_n2781), .A2(n22412), .B(n22283), .Y(n23334) );
  XOR2x2_ASAP7_75t_SL U26322 ( .A(n23167), .B(mult_x_1196_n2059), .Y(
        mult_x_1196_n2051) );
  NOR2xp33_ASAP7_75t_SL U26323 ( .A(n28904), .B(n18884), .Y(n22256) );
  AO21x2_ASAP7_75t_SL U26324 ( .A1(n23992), .A2(n24287), .B(mult_x_1196_n3145), 
        .Y(mult_x_1196_n2569) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U26325 ( .A1(n31406), .A2(n18997), .B(n31405), 
        .C(n31404), .Y(n31409) );
  HB1xp67_ASAP7_75t_SL U26326 ( .A(n23166), .Y(n23165) );
  INVx1_ASAP7_75t_SL U26327 ( .A(n22499), .Y(n22257) );
  BUFx3_ASAP7_75t_SL U26328 ( .A(mult_x_1196_n432), .Y(n23926) );
  OAI21x1_ASAP7_75t_SL U26329 ( .A1(mult_x_1196_n2466), .A2(mult_x_1196_n2558), 
        .B(n23721), .Y(mult_x_1196_n1921) );
  HB1xp67_ASAP7_75t_SL U26330 ( .A(mult_x_1196_n1913), .Y(n22259) );
  XNOR2x1_ASAP7_75t_SL U26331 ( .A(mult_x_1196_n1383), .B(n22769), .Y(
        mult_x_1196_n1345) );
  BUFx3_ASAP7_75t_SL U26332 ( .A(n24422), .Y(n22698) );
  XNOR2x1_ASAP7_75t_SL U26333 ( .A(n22680), .B(n22679), .Y(mult_x_1196_n2006)
         );
  XOR2xp5_ASAP7_75t_SL U26334 ( .A(mult_x_1196_n1810), .B(mult_x_1196_n1791), 
        .Y(n22263) );
  XNOR2x1_ASAP7_75t_SL U26335 ( .A(mult_x_1196_n1317), .B(n23351), .Y(
        mult_x_1196_n1308) );
  HB1xp67_ASAP7_75t_SL U26336 ( .A(mult_x_1196_n1359), .Y(n22260) );
  OAI22xp5_ASAP7_75t_SL U26337 ( .A1(mult_x_1196_n2817), .A2(n24034), .B1(
        n18402), .B2(mult_x_1196_n2816), .Y(mult_x_1196_n2251) );
  HB1xp67_ASAP7_75t_SL U26338 ( .A(n24191), .Y(n22261) );
  INVx8_ASAP7_75t_SL U26339 ( .A(add_x_735_A_20_), .Y(n23935) );
  XNOR2xp5_ASAP7_75t_SL U26340 ( .A(n22610), .B(n22263), .Y(n22262) );
  XNOR2xp5_ASAP7_75t_SL U26341 ( .A(n22610), .B(n23075), .Y(n24110) );
  INVx1_ASAP7_75t_SL U26342 ( .A(mult_x_1196_n1372), .Y(n22463) );
  INVxp33_ASAP7_75t_SRAM U26343 ( .A(mult_x_1196_n612), .Y(n23701) );
  XNOR2x2_ASAP7_75t_SL U26344 ( .A(n24072), .B(n18393), .Y(mult_x_1196_n3241)
         );
  XNOR2x2_ASAP7_75t_SL U26345 ( .A(n24066), .B(n18393), .Y(mult_x_1196_n3235)
         );
  BUFx5_ASAP7_75t_SL U26346 ( .A(add_x_735_A_4_), .Y(n22449) );
  OAI21xp33_ASAP7_75t_SRAM U26347 ( .A1(mult_x_1196_n748), .A2(n24196), .B(
        n22504), .Y(n23889) );
  INVxp33_ASAP7_75t_SRAM U26348 ( .A(mult_x_1196_n748), .Y(mult_x_1196_n747)
         );
  OAI22xp5_ASAP7_75t_SL U26349 ( .A1(n24017), .A2(mult_x_1196_n2941), .B1(
        mult_x_1196_n2942), .B2(n22779), .Y(mult_x_1196_n2370) );
  OAI21x1_ASAP7_75t_SL U26350 ( .A1(mult_x_1196_n3210), .A2(n22802), .B(n23079), .Y(n23078) );
  NOR2x1_ASAP7_75t_SL U26351 ( .A(mult_x_1196_n3194), .B(n23522), .Y(n22733)
         );
  BUFx2_ASAP7_75t_SL U26352 ( .A(n23026), .Y(n22543) );
  NAND2x1_ASAP7_75t_SL U26353 ( .A(n22330), .B(mult_x_1196_n1949), .Y(
        mult_x_1196_n693) );
  INVx1_ASAP7_75t_SL U26354 ( .A(n24017), .Y(n22265) );
  BUFx2_ASAP7_75t_SL U26355 ( .A(n24017), .Y(n22694) );
  NOR2x1p5_ASAP7_75t_SL U26356 ( .A(mult_x_1196_n1392), .B(n22359), .Y(
        mult_x_1196_n575) );
  NAND2x1p5_ASAP7_75t_SL U26357 ( .A(n22359), .B(mult_x_1196_n1392), .Y(n24201) );
  INVxp33_ASAP7_75t_SRAM U26358 ( .A(n23046), .Y(n23045) );
  INVx1_ASAP7_75t_SL U26359 ( .A(mult_x_1196_n535), .Y(n22264) );
  INVx1_ASAP7_75t_SL U26360 ( .A(n18996), .Y(mult_x_1196_n535) );
  INVx4_ASAP7_75t_SL U26361 ( .A(n24015), .Y(n24017) );
  OAI22x1_ASAP7_75t_SL U26362 ( .A1(n23830), .A2(n26260), .B1(n23559), .B2(
        n23847), .Y(u0_0_leon3x0_p0_muli[17]) );
  INVx8_ASAP7_75t_SL U26363 ( .A(n22216), .Y(n23965) );
  NOR2xp33_ASAP7_75t_SL U26364 ( .A(n22227), .B(n18423), .Y(n22267) );
  OR2x2_ASAP7_75t_SL U26365 ( .A(n26514), .B(n24686), .Y(n22268) );
  INVx3_ASAP7_75t_SL U26366 ( .A(add_x_735_A_24_), .Y(n24692) );
  INVx11_ASAP7_75t_SL U26367 ( .A(n23954), .Y(n23955) );
  AND2x2_ASAP7_75t_SL U26368 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__30_), .B(n24687), .Y(n22269) );
  OAI21xp5_ASAP7_75t_SL U26369 ( .A1(n31475), .A2(n18567), .B(n18420), .Y(
        u0_0_leon3x0_p0_muli[41]) );
  OR2x2_ASAP7_75t_SL U26370 ( .A(mult_x_1196_n2904), .B(n24025), .Y(n22270) );
  OR2x2_ASAP7_75t_SL U26371 ( .A(n24186), .B(n23788), .Y(n22271) );
  AOI21xp33_ASAP7_75t_SRAM U26372 ( .A1(n24025), .A2(n22464), .B(
        mult_x_1196_n2873), .Y(n22272) );
  INVx4_ASAP7_75t_SL U26373 ( .A(n23155), .Y(add_x_735_A_15_) );
  INVx1_ASAP7_75t_SL U26374 ( .A(u0_0_leon3x0_p0_muli[38]), .Y(mult_x_1196_n6)
         );
  OR2x2_ASAP7_75t_SL U26375 ( .A(u0_0_leon3x0_p0_divi[0]), .B(n22999), .Y(
        n22274) );
  BUFx2_ASAP7_75t_SL U26376 ( .A(u0_0_leon3x0_p0_muli[38]), .Y(n22999) );
  BUFx3_ASAP7_75t_SL U26377 ( .A(mult_x_1196_n6), .Y(n23980) );
  OR2x2_ASAP7_75t_SL U26378 ( .A(mult_x_1196_n3060), .B(n24005), .Y(n22275) );
  OR2x2_ASAP7_75t_SL U26379 ( .A(n24005), .B(mult_x_1196_n3048), .Y(n22276) );
  OR2x2_ASAP7_75t_SL U26380 ( .A(mult_x_1196_n3071), .B(n24005), .Y(n22277) );
  INVx5_ASAP7_75t_SL U26381 ( .A(n23415), .Y(add_x_735_A_32_) );
  OR2x2_ASAP7_75t_SL U26382 ( .A(n29801), .B(n18911), .Y(n22278) );
  BUFx2_ASAP7_75t_SL U26383 ( .A(n24550), .Y(n22902) );
  XOR2xp5_ASAP7_75t_SL U26384 ( .A(n22442), .B(n22642), .Y(n22279) );
  OR2x2_ASAP7_75t_SL U26385 ( .A(mult_x_1196_n2753), .B(n24040), .Y(n22280) );
  OR2x2_ASAP7_75t_SL U26386 ( .A(mult_x_1196_n2764), .B(n24040), .Y(n22282) );
  OAI22xp33_ASAP7_75t_SRAM U26387 ( .A1(n24040), .A2(mult_x_1196_n2747), .B1(
        n24041), .B2(n23534), .Y(mult_x_1196_n2185) );
  OR2x2_ASAP7_75t_SL U26388 ( .A(mult_x_1196_n2780), .B(n22481), .Y(n22283) );
  OR2x2_ASAP7_75t_SL U26389 ( .A(n22391), .B(mult_x_1196_n2781), .Y(n22284) );
  OAI22xp5_ASAP7_75t_SL U26390 ( .A1(mult_x_1196_n2789), .A2(n24039), .B1(
        mult_x_1196_n2788), .B2(n22936), .Y(mult_x_1196_n2223) );
  NAND2x1p5_ASAP7_75t_SL U26391 ( .A(n24546), .B(n24545), .Y(n22285) );
  OR2x2_ASAP7_75t_SL U26392 ( .A(mult_x_1196_n3122), .B(n23999), .Y(n22286) );
  OR2x2_ASAP7_75t_SL U26393 ( .A(n23996), .B(mult_x_1196_n3142), .Y(n22287) );
  OR2x2_ASAP7_75t_SL U26394 ( .A(n23996), .B(mult_x_1196_n3139), .Y(n22288) );
  MAJx2_ASAP7_75t_SL U26395 ( .A(mult_x_1196_n2371), .B(mult_x_1196_n2156), 
        .C(n22531), .Y(n22289) );
  OR2x2_ASAP7_75t_SL U26396 ( .A(n24017), .B(n22579), .Y(n22290) );
  OR2x2_ASAP7_75t_SL U26397 ( .A(mult_x_1196_n3036), .B(n23442), .Y(n22291) );
  OA22x2_ASAP7_75t_SL U26398 ( .A1(mult_x_1196_n3032), .A2(n22815), .B1(
        mult_x_1196_n3031), .B2(n23442), .Y(n22292) );
  OR2x2_ASAP7_75t_SL U26399 ( .A(mult_x_1196_n3020), .B(n24009), .Y(n22293) );
  OR2x2_ASAP7_75t_SL U26400 ( .A(mult_x_1196_n3019), .B(n23442), .Y(n22294) );
  OR2x2_ASAP7_75t_SL U26401 ( .A(n22389), .B(mult_x_1196_n3254), .Y(n22295) );
  OAI22x1_ASAP7_75t_SL U26402 ( .A1(mult_x_1196_n3257), .A2(n23981), .B1(
        n22389), .B2(mult_x_1196_n3256), .Y(n23932) );
  OR2x2_ASAP7_75t_SL U26403 ( .A(n23288), .B(n23125), .Y(n22296) );
  AND2x2_ASAP7_75t_SL U26404 ( .A(n23205), .B(mult_x_1196_n2531), .Y(n22297)
         );
  OR2x2_ASAP7_75t_SL U26405 ( .A(mult_x_1196_n2686), .B(mult_x_1196_n2526), 
        .Y(n22298) );
  XOR2x2_ASAP7_75t_SL U26406 ( .A(n18447), .B(n23070), .Y(n22299) );
  INVx11_ASAP7_75t_SL U26407 ( .A(n23358), .Y(n23984) );
  OR2x2_ASAP7_75t_SL U26408 ( .A(mult_x_1196_n2990), .B(n24011), .Y(n22300) );
  OR2x2_ASAP7_75t_SL U26409 ( .A(mult_x_1196_n2986), .B(n24011), .Y(n22301) );
  OR2x2_ASAP7_75t_SL U26410 ( .A(mult_x_1196_n2999), .B(n24011), .Y(n22302) );
  OR2x2_ASAP7_75t_SL U26411 ( .A(mult_x_1196_n2983), .B(n24011), .Y(n22303) );
  OR2x2_ASAP7_75t_SL U26412 ( .A(mult_x_1196_n3005), .B(n24011), .Y(n22304) );
  OR2x2_ASAP7_75t_SL U26413 ( .A(mult_x_1196_n3003), .B(n24012), .Y(n22305) );
  XNOR2x2_ASAP7_75t_SL U26414 ( .A(n22593), .B(mult_x_1196_n2377), .Y(n22306)
         );
  XOR2xp5_ASAP7_75t_SL U26415 ( .A(n22494), .B(mult_x_1196_n1948), .Y(n22307)
         );
  XOR2xp5_ASAP7_75t_SL U26416 ( .A(n22545), .B(n22544), .Y(n22308) );
  OR2x2_ASAP7_75t_SL U26417 ( .A(mult_x_1196_n2830), .B(n22251), .Y(n22309) );
  MAJx2_ASAP7_75t_SL U26418 ( .A(mult_x_1196_n1243), .B(mult_x_1196_n1285), 
        .C(n23426), .Y(n22310) );
  XOR2xp5_ASAP7_75t_SL U26419 ( .A(n22925), .B(n22922), .Y(n22311) );
  XNOR2x2_ASAP7_75t_SL U26420 ( .A(mult_x_1196_n1034), .B(n22838), .Y(
        mult_x_1196_n1015) );
  MAJx2_ASAP7_75t_SL U26421 ( .A(mult_x_1196_n926), .B(mult_x_1196_n944), .C(
        n22495), .Y(n22312) );
  NOR2x1_ASAP7_75t_SL U26422 ( .A(mult_x_1196_n869), .B(mult_x_1196_n860), .Y(
        mult_x_1196_n323) );
  MAJx2_ASAP7_75t_SL U26423 ( .A(mult_x_1196_n1161), .B(mult_x_1196_n1187), 
        .C(n23174), .Y(n22314) );
  OR2x2_ASAP7_75t_SL U26424 ( .A(mult_x_1196_n3201), .B(n22248), .Y(n22315) );
  OR2x2_ASAP7_75t_SL U26425 ( .A(n22248), .B(mult_x_1196_n3212), .Y(n22316) );
  OR2x2_ASAP7_75t_SL U26426 ( .A(mult_x_1196_n3179), .B(n23988), .Y(n22317) );
  INVx6_ASAP7_75t_SL U26427 ( .A(n23956), .Y(n23957) );
  OR2x2_ASAP7_75t_SL U26428 ( .A(mult_x_1196_n3176), .B(n23992), .Y(n22318) );
  OR2x2_ASAP7_75t_SL U26429 ( .A(mult_x_1196_n3173), .B(n24230), .Y(n22319) );
  XOR2xp5_ASAP7_75t_SL U26430 ( .A(n23044), .B(n23042), .Y(n22320) );
  OR2x2_ASAP7_75t_SL U26431 ( .A(mult_x_1196_n1887), .B(mult_x_1196_n1883), 
        .Y(n22321) );
  AND2x2_ASAP7_75t_SL U26432 ( .A(mult_x_1196_n2418), .B(mult_x_1196_n2574), 
        .Y(n22322) );
  XOR2x2_ASAP7_75t_SL U26433 ( .A(mult_x_1196_n1872), .B(n22618), .Y(n22326)
         );
  AND2x2_ASAP7_75t_SL U26434 ( .A(n23796), .B(n23798), .Y(n22327) );
  AND2x2_ASAP7_75t_SL U26435 ( .A(n23795), .B(mult_x_1196_n1956), .Y(n22328)
         );
  MAJx2_ASAP7_75t_SL U26436 ( .A(mult_x_1196_n1974), .B(n23934), .C(n18930), 
        .Y(n22330) );
  AND2x2_ASAP7_75t_SL U26437 ( .A(n23656), .B(mult_x_1196_n2633), .Y(n22331)
         );
  AND2x2_ASAP7_75t_SL U26438 ( .A(mult_x_1196_n2004), .B(n23624), .Y(n22333)
         );
  MAJx2_ASAP7_75t_SL U26439 ( .A(mult_x_1196_n2035), .B(mult_x_1196_n2031), 
        .C(n22490), .Y(n22334) );
  XNOR2x1_ASAP7_75t_SL U26440 ( .A(n22689), .B(n22638), .Y(n22336) );
  XNOR2x1_ASAP7_75t_SL U26441 ( .A(n22577), .B(n22575), .Y(mult_x_1196_n1173)
         );
  MAJx2_ASAP7_75t_SL U26442 ( .A(mult_x_1196_n1216), .B(mult_x_1196_n1222), 
        .C(mult_x_1196_n1218), .Y(n22337) );
  XNOR2x2_ASAP7_75t_SL U26443 ( .A(mult_x_1196_n1148), .B(n22561), .Y(
        mult_x_1196_n1142) );
  MAJx2_ASAP7_75t_SL U26444 ( .A(mult_x_1196_n1110), .B(n23917), .C(
        mult_x_1196_n1141), .Y(n22339) );
  XOR2x2_ASAP7_75t_SL U26445 ( .A(mult_x_1196_n945), .B(n22558), .Y(n22340) );
  MAJx2_ASAP7_75t_SL U26446 ( .A(mult_x_1196_n1789), .B(n22868), .C(
        mult_x_1196_n1787), .Y(n22342) );
  XOR2x2_ASAP7_75t_SL U26447 ( .A(n23184), .B(mult_x_1196_n1637), .Y(n22343)
         );
  MAJIxp5_ASAP7_75t_SL U26448 ( .A(n23613), .B(n23611), .C(n23610), .Y(n22345)
         );
  XOR2x2_ASAP7_75t_SL U26449 ( .A(n24297), .B(n22942), .Y(n22346) );
  XOR2x1_ASAP7_75t_SL U26450 ( .A(n23197), .B(n23196), .Y(n22347) );
  MAJx2_ASAP7_75t_SL U26451 ( .A(mult_x_1196_n1346), .B(mult_x_1196_n1352), 
        .C(mult_x_1196_n1348), .Y(n22348) );
  MAJx2_ASAP7_75t_SL U26452 ( .A(mult_x_1196_n1509), .B(n22935), .C(n22761), 
        .Y(n22349) );
  XOR2xp5_ASAP7_75t_SL U26453 ( .A(n23308), .B(n23307), .Y(n22350) );
  XNOR2x2_ASAP7_75t_SL U26454 ( .A(n18558), .B(n22683), .Y(mult_x_1196_n1340)
         );
  MAJx2_ASAP7_75t_SL U26455 ( .A(mult_x_1196_n1424), .B(mult_x_1196_n1416), 
        .C(mult_x_1196_n1418), .Y(n22351) );
  OR2x2_ASAP7_75t_SL U26456 ( .A(mult_x_1196_n2924), .B(n24020), .Y(n22352) );
  MAJx2_ASAP7_75t_SL U26457 ( .A(mult_x_1196_n1140), .B(mult_x_1196_n1136), 
        .C(n18616), .Y(n22353) );
  OR2x2_ASAP7_75t_SL U26458 ( .A(mult_x_1196_n1653), .B(n22212), .Y(n22355) );
  MAJx2_ASAP7_75t_SL U26459 ( .A(mult_x_1196_n1686), .B(mult_x_1196_n1681), 
        .C(mult_x_1196_n1718), .Y(n22356) );
  MAJx2_ASAP7_75t_SL U26460 ( .A(mult_x_1196_n1767), .B(n22535), .C(
        mult_x_1196_n1763), .Y(n22357) );
  MAJx2_ASAP7_75t_SL U26461 ( .A(mult_x_1196_n1446), .B(mult_x_1196_n1435), 
        .C(n22486), .Y(n22358) );
  AND2x2_ASAP7_75t_SL U26462 ( .A(n22725), .B(n22723), .Y(n22359) );
  XOR2xp5_ASAP7_75t_SL U26463 ( .A(n23067), .B(n23066), .Y(n22360) );
  INVx2_ASAP7_75t_SL U26464 ( .A(mult_x_1196_n312), .Y(n23385) );
  AND2x2_ASAP7_75t_SL U26465 ( .A(mult_x_1196_n324), .B(mult_x_1196_n331), .Y(
        n22361) );
  MAJx2_ASAP7_75t_SL U26466 ( .A(mult_x_1196_n951), .B(mult_x_1196_n954), .C(
        n22360), .Y(n22362) );
  MAJx2_ASAP7_75t_SL U26467 ( .A(mult_x_1196_n1050), .B(mult_x_1196_n1029), 
        .C(n22364), .Y(n22363) );
  XNOR2xp5_ASAP7_75t_SL U26468 ( .A(n23086), .B(n23083), .Y(n22364) );
  HB1xp67_ASAP7_75t_SL U26469 ( .A(n23669), .Y(n22676) );
  INVx2_ASAP7_75t_SL U26470 ( .A(n23669), .Y(n23387) );
  XOR2x1_ASAP7_75t_SL U26471 ( .A(n22675), .B(n22673), .Y(n22365) );
  AND2x2_ASAP7_75t_SL U26472 ( .A(mult_x_1196_n398), .B(mult_x_1196_n784), .Y(
        n22366) );
  AND2x2_ASAP7_75t_SL U26473 ( .A(mult_x_1196_n407), .B(mult_x_1196_n785), .Y(
        n22367) );
  NOR2x1p5_ASAP7_75t_SL U26474 ( .A(n23575), .B(n23572), .Y(mult_x_1196_n385)
         );
  INVxp33_ASAP7_75t_SRAM U26475 ( .A(mult_x_1196_n1650), .Y(n22744) );
  INVx1_ASAP7_75t_SL U26476 ( .A(mult_x_1196_n1447), .Y(n22369) );
  INVx2_ASAP7_75t_SL U26477 ( .A(n22369), .Y(n22370) );
  HB1xp67_ASAP7_75t_SL U26478 ( .A(mult_x_1196_n1288), .Y(n22439) );
  HB1xp67_ASAP7_75t_SL U26479 ( .A(mult_x_1196_n1371), .Y(n22739) );
  XNOR2x1_ASAP7_75t_SL U26480 ( .A(n24056), .B(n24231), .Y(mult_x_1196_n2953)
         );
  BUFx6f_ASAP7_75t_SL U26481 ( .A(u0_0_leon3x0_p0_muli[28]), .Y(n24056) );
  HB1xp67_ASAP7_75t_SL U26482 ( .A(n28848), .Y(n22952) );
  XOR2xp5_ASAP7_75t_SL U26483 ( .A(mult_x_1196_n2262), .B(mult_x_1196_n2604), 
        .Y(n22557) );
  XNOR2xp5_ASAP7_75t_SL U26484 ( .A(mult_x_1196_n2640), .B(mult_x_1196_n2512), 
        .Y(n23070) );
  NOR2x1_ASAP7_75t_SL U26485 ( .A(n24012), .B(mult_x_1196_n2998), .Y(n23880)
         );
  HB1xp67_ASAP7_75t_SL U26486 ( .A(mult_x_1196_n1483), .Y(n22648) );
  NAND2x1p5_ASAP7_75t_SL U26487 ( .A(n23296), .B(n23294), .Y(mult_x_1196_n1320) );
  HB1xp67_ASAP7_75t_SL U26488 ( .A(mult_x_1196_n1341), .Y(n23060) );
  INVx1_ASAP7_75t_SL U26489 ( .A(mult_x_1196_n1043), .Y(n22371) );
  INVx2_ASAP7_75t_SL U26490 ( .A(n22371), .Y(n22372) );
  OAI21xp5_ASAP7_75t_SL U26491 ( .A1(n30899), .A2(n22399), .B(n30896), .Y(
        timer0_v_TIMERS__1__VALUE__27_) );
  OAI21xp5_ASAP7_75t_SL U26492 ( .A1(n31852), .A2(n22399), .B(n31846), .Y(
        timer0_v_TIMERS__1__VALUE__21_) );
  OAI21xp5_ASAP7_75t_SL U26493 ( .A1(n26654), .A2(n22399), .B(n26653), .Y(
        timer0_v_TIMERS__1__VALUE__0_) );
  OAI21xp5_ASAP7_75t_SL U26494 ( .A1(n26646), .A2(n22399), .B(n26645), .Y(
        timer0_v_TIMERS__1__VALUE__2_) );
  AOI21xp5_ASAP7_75t_SL U26495 ( .A1(n31845), .A2(timer0_res_27_), .B(n30895), 
        .Y(n30896) );
  AOI21xp5_ASAP7_75t_SL U26496 ( .A1(n31845), .A2(timer0_res_21_), .B(n31844), 
        .Y(n31846) );
  INVx1_ASAP7_75t_SL U26497 ( .A(mult_x_1196_n456), .Y(mult_x_1196_n454) );
  AOI21xp5_ASAP7_75t_SL U26498 ( .A1(n31845), .A2(n22430), .B(n26652), .Y(
        n26653) );
  AOI21xp5_ASAP7_75t_SL U26499 ( .A1(n31845), .A2(timer0_res_2_), .B(n26644), 
        .Y(n26645) );
  OAI21xp5_ASAP7_75t_SL U26500 ( .A1(n24646), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N21), .B(n29095), .Y(n4273) );
  OAI22xp33_ASAP7_75t_SL U26501 ( .A1(n32380), .A2(n24637), .B1(n32379), .B2(
        n22383), .Y(n26330) );
  OAI22xp33_ASAP7_75t_SL U26502 ( .A1(n32308), .A2(n24637), .B1(n32307), .B2(
        n22383), .Y(n25870) );
  OAI22xp33_ASAP7_75t_SL U26503 ( .A1(n31378), .A2(n24637), .B1(n32395), .B2(
        n22383), .Y(n28407) );
  OAI22xp33_ASAP7_75t_SL U26504 ( .A1(n32354), .A2(n24637), .B1(n32360), .B2(
        n22383), .Y(n26663) );
  OAI22xp33_ASAP7_75t_SL U26505 ( .A1(n32371), .A2(n24637), .B1(n32375), .B2(
        n22383), .Y(n26538) );
  OAI22xp33_ASAP7_75t_SL U26506 ( .A1(n30904), .A2(n24637), .B1(n32402), .B2(
        n22383), .Y(n26343) );
  OAI22xp33_ASAP7_75t_SL U26507 ( .A1(n32391), .A2(n24637), .B1(n32392), .B2(
        n22383), .Y(n26510) );
  OAI22xp33_ASAP7_75t_SL U26508 ( .A1(n32377), .A2(n24637), .B1(n32376), .B2(
        n22383), .Y(n26963) );
  OAI22xp33_ASAP7_75t_SL U26509 ( .A1(n32301), .A2(n24637), .B1(n32300), .B2(
        n22383), .Y(n27490) );
  OAI22xp33_ASAP7_75t_SL U26510 ( .A1(n32297), .A2(n24637), .B1(n32293), .B2(
        n22383), .Y(n28101) );
  OAI22xp33_ASAP7_75t_SL U26511 ( .A1(n32399), .A2(n24637), .B1(n32401), .B2(
        n22383), .Y(n26232) );
  INVxp67_ASAP7_75t_SL U26512 ( .A(mult_x_1196_n486), .Y(mult_x_1196_n484) );
  OAI22xp33_ASAP7_75t_SL U26513 ( .A1(n29861), .A2(n24637), .B1(n29847), .B2(
        n22383), .Y(n25427) );
  INVxp67_ASAP7_75t_SL U26514 ( .A(n31587), .Y(n31593) );
  OAI21xp33_ASAP7_75t_SL U26515 ( .A1(n22421), .A2(u0_0_leon3x0_p0_ici[60]), 
        .B(n28909), .Y(n3202) );
  NAND2xp5_ASAP7_75t_SL U26516 ( .A(mult_x_1196_n793), .B(mult_x_1196_n795), 
        .Y(n22492) );
  NOR2xp67_ASAP7_75t_SL U26517 ( .A(n25587), .B(n31257), .Y(n25591) );
  AOI21xp33_ASAP7_75t_SL U26518 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__9_), .B(n32579), .Y(n2958)
         );
  AOI21xp33_ASAP7_75t_SL U26519 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__8_), .B(n32576), .Y(n2959)
         );
  AOI21xp33_ASAP7_75t_SL U26520 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__7_), .B(n32573), .Y(n2960)
         );
  AOI21xp33_ASAP7_75t_SL U26521 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[25]), .B(n32554), .Y(n2939) );
  AOI21xp33_ASAP7_75t_SL U26522 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__28_), .B(n32554), .Y(n2940)
         );
  AOI21xp33_ASAP7_75t_SL U26523 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__24_), .B(n32544), .Y(n2466)
         );
  INVx2_ASAP7_75t_SL U26524 ( .A(n23576), .Y(n22404) );
  INVx1_ASAP7_75t_SL U26525 ( .A(mult_x_1196_n781), .Y(n22406) );
  INVxp67_ASAP7_75t_SL U26526 ( .A(mult_x_1196_n398), .Y(mult_x_1196_n396) );
  INVxp33_ASAP7_75t_SL U26527 ( .A(n27280), .Y(n27286) );
  INVxp67_ASAP7_75t_SL U26528 ( .A(mult_x_1196_n354), .Y(mult_x_1196_n781) );
  AOI21xp5_ASAP7_75t_SL U26529 ( .A1(n30495), .A2(n31342), .B(n27221), .Y(
        n30490) );
  INVxp67_ASAP7_75t_SL U26530 ( .A(n30646), .Y(n30647) );
  AOI21xp33_ASAP7_75t_SL U26531 ( .A1(n29867), .A2(n31342), .B(n28281), .Y(
        n29615) );
  BUFx2_ASAP7_75t_SL U26532 ( .A(mult_x_1196_n1400), .Y(n22570) );
  AOI21xp5_ASAP7_75t_SL U26533 ( .A1(n28608), .A2(n31342), .B(n27190), .Y(
        n29618) );
  AOI21xp5_ASAP7_75t_SL U26534 ( .A1(n30972), .A2(n31342), .B(n29840), .Y(
        n31053) );
  AOI21xp5_ASAP7_75t_SL U26535 ( .A1(n30736), .A2(n31342), .B(n29931), .Y(
        n30732) );
  AOI21xp5_ASAP7_75t_SL U26536 ( .A1(n27174), .A2(n31342), .B(n27173), .Y(
        n30733) );
  OAI21xp5_ASAP7_75t_SL U26537 ( .A1(DP_OP_5187J1_124_3275_n290), .A2(
        DP_OP_5187J1_124_3275_n262), .B(DP_OP_5187J1_124_3275_n263), .Y(
        DP_OP_5187J1_124_3275_n261) );
  NOR2xp33_ASAP7_75t_SL U26538 ( .A(mult_x_1196_n859), .B(mult_x_1196_n852), 
        .Y(mult_x_1196_n316) );
  OAI21xp33_ASAP7_75t_SL U26539 ( .A1(n2925), .A2(n22408), .B(n25326), .Y(
        n17887) );
  INVx4_ASAP7_75t_SL U26540 ( .A(n24424), .Y(n22408) );
  INVxp67_ASAP7_75t_SL U26541 ( .A(DP_OP_5187J1_124_3275_n169), .Y(
        DP_OP_5187J1_124_3275_n320) );
  NOR2xp33_ASAP7_75t_SL U26542 ( .A(timer0_N72), .B(n18861), .Y(n24351) );
  OAI21xp5_ASAP7_75t_SL U26543 ( .A1(DP_OP_5187J1_124_3275_n159), .A2(
        DP_OP_5187J1_124_3275_n151), .B(DP_OP_5187J1_124_3275_n152), .Y(
        DP_OP_5187J1_124_3275_n146) );
  OAI22xp33_ASAP7_75t_SL U26544 ( .A1(n32988), .A2(n22386), .B1(n33053), .B2(
        n32987), .Y(n32989) );
  NOR3xp33_ASAP7_75t_SL U26545 ( .A(n24341), .B(timer0_N74), .C(timer0_N75), 
        .Y(n24347) );
  INVxp67_ASAP7_75t_SL U26546 ( .A(n28675), .Y(n27161) );
  NAND2xp33_ASAP7_75t_SL U26547 ( .A(n29987), .B(n29976), .Y(n29983) );
  NAND2xp33_ASAP7_75t_SL U26548 ( .A(n30632), .B(n29604), .Y(n26904) );
  INVxp67_ASAP7_75t_SL U26549 ( .A(n30021), .Y(n30022) );
  INVxp67_ASAP7_75t_SL U26550 ( .A(n28854), .Y(n28876) );
  INVxp67_ASAP7_75t_SL U26551 ( .A(add_x_746_n153), .Y(add_x_746_n152) );
  INVx3_ASAP7_75t_SL U26552 ( .A(n29937), .Y(n31631) );
  INVx1_ASAP7_75t_SL U26553 ( .A(n31364), .Y(n30575) );
  NAND2xp5_ASAP7_75t_SL U26554 ( .A(n30632), .B(n28498), .Y(n27079) );
  INVxp67_ASAP7_75t_SL U26555 ( .A(mult_x_1196_n928), .Y(n22527) );
  AOI21xp33_ASAP7_75t_SL U26556 ( .A1(n28974), .A2(n28977), .B(n26300), .Y(
        n28913) );
  OAI21xp33_ASAP7_75t_SL U26557 ( .A1(n28975), .A2(n25464), .B(n25203), .Y(
        n29602) );
  INVx1_ASAP7_75t_SL U26558 ( .A(n31054), .Y(n32110) );
  INVxp67_ASAP7_75t_SL U26559 ( .A(add_x_735_n3), .Y(add_x_735_n77) );
  INVxp67_ASAP7_75t_SL U26560 ( .A(mult_x_1196_n929), .Y(n22795) );
  OAI22xp33_ASAP7_75t_SL U26561 ( .A1(n2924), .A2(n33023), .B1(n32761), .B2(
        n33011), .Y(n32756) );
  AOI21xp33_ASAP7_75t_SL U26562 ( .A1(n28873), .A2(n28977), .B(n26280), .Y(
        n28858) );
  INVx1_ASAP7_75t_SL U26563 ( .A(n32776), .Y(n31737) );
  NAND2xp5_ASAP7_75t_SL U26564 ( .A(n24681), .B(n31967), .Y(n30706) );
  NAND2xp5_ASAP7_75t_SL U26565 ( .A(n24575), .B(n27090), .Y(n27095) );
  INVxp67_ASAP7_75t_SL U26566 ( .A(n27089), .Y(n27096) );
  OAI21xp33_ASAP7_75t_SL U26567 ( .A1(apbi[9]), .A2(n31840), .B(n26620), .Y(
        n1793) );
  OAI21xp33_ASAP7_75t_SL U26568 ( .A1(apbi[1]), .A2(n31840), .B(n26647), .Y(
        n2845) );
  OAI21xp33_ASAP7_75t_SL U26569 ( .A1(n31761), .A2(n22415), .B(n25247), .Y(
        n33039) );
  OAI21xp33_ASAP7_75t_SL U26570 ( .A1(apbi[19]), .A2(n31840), .B(n26543), .Y(
        n2347) );
  OAI21xp33_ASAP7_75t_SL U26571 ( .A1(apbi[28]), .A2(n31840), .B(n31495), .Y(
        n1776) );
  OAI21xp33_ASAP7_75t_SL U26572 ( .A1(apbi[3]), .A2(n31840), .B(n26640), .Y(
        n2841) );
  OAI21xp33_ASAP7_75t_SL U26573 ( .A1(apbi[0]), .A2(n31840), .B(n26651), .Y(
        n2847) );
  INVx1_ASAP7_75t_SL U26574 ( .A(n28849), .Y(n27090) );
  OAI21xp33_ASAP7_75t_SL U26575 ( .A1(apbi[29]), .A2(n31840), .B(n26491), .Y(
        n1751) );
  OAI21xp33_ASAP7_75t_SL U26576 ( .A1(n31768), .A2(n22415), .B(n25254), .Y(
        n33029) );
  NOR2x1_ASAP7_75t_SL U26577 ( .A(n23781), .B(n23780), .Y(n23779) );
  OAI21xp33_ASAP7_75t_SL U26578 ( .A1(apbi[16]), .A2(n31840), .B(n26451), .Y(
        n1772) );
  OAI21xp33_ASAP7_75t_SL U26579 ( .A1(apbi[6]), .A2(n31840), .B(n26630), .Y(
        n1729) );
  OAI21xp33_ASAP7_75t_SL U26580 ( .A1(apbi[14]), .A2(n31840), .B(n26594), .Y(
        n2323) );
  OAI21xp33_ASAP7_75t_SL U26581 ( .A1(apbi[2]), .A2(n31840), .B(n26643), .Y(
        n2843) );
  OAI21xp33_ASAP7_75t_SL U26582 ( .A1(apbi[5]), .A2(n31840), .B(n26633), .Y(
        n2839) );
  AOI22xp33_ASAP7_75t_SL U26583 ( .A1(n28979), .A2(n23665), .B1(n22999), .B2(
        n28980), .Y(n28984) );
  OAI21xp33_ASAP7_75t_SL U26584 ( .A1(apbi[30]), .A2(n31840), .B(n26478), .Y(
        n1640) );
  OAI21xp33_ASAP7_75t_SL U26585 ( .A1(apbi[12]), .A2(n31840), .B(n26607), .Y(
        n1635) );
  OAI21xp33_ASAP7_75t_SL U26586 ( .A1(apbi[4]), .A2(n31840), .B(n26636), .Y(
        n1631) );
  OAI21xp33_ASAP7_75t_SL U26587 ( .A1(apbi[27]), .A2(n31840), .B(n30893), .Y(
        n2232) );
  OAI21xp33_ASAP7_75t_SL U26588 ( .A1(apbi[7]), .A2(n31840), .B(n26627), .Y(
        n1627) );
  NAND2xp33_ASAP7_75t_SL U26589 ( .A(n25436), .B(n25435), .Y(n25437) );
  OAI21xp33_ASAP7_75t_SL U26590 ( .A1(apbi[26]), .A2(n31840), .B(n26497), .Y(
        n2828) );
  OAI21xp33_ASAP7_75t_SL U26591 ( .A1(apbi[11]), .A2(n31840), .B(n25969), .Y(
        n2234) );
  OAI21xp33_ASAP7_75t_SL U26592 ( .A1(apbi[23]), .A2(n31840), .B(n26529), .Y(
        n2830) );
  OAI21xp33_ASAP7_75t_SL U26593 ( .A1(apbi[22]), .A2(n31840), .B(n31640), .Y(
        n2831) );
  OAI21xp33_ASAP7_75t_SL U26594 ( .A1(apbi[18]), .A2(n31840), .B(n25847), .Y(
        n2834) );
  NAND2xp5_ASAP7_75t_SL U26595 ( .A(n28132), .B(n28404), .Y(n27089) );
  INVxp67_ASAP7_75t_SL U26596 ( .A(n30307), .Y(n30316) );
  OAI21xp33_ASAP7_75t_SL U26597 ( .A1(apbi[31]), .A2(n31840), .B(n26461), .Y(
        n2827) );
  NAND2xp33_ASAP7_75t_SL U26598 ( .A(n26919), .B(n26918), .Y(n26935) );
  NAND2xp33_ASAP7_75t_SL U26599 ( .A(n31646), .B(n31840), .Y(n31640) );
  NAND2xp33_ASAP7_75t_SL U26600 ( .A(n31373), .B(n31840), .Y(n31367) );
  NAND2xp33_ASAP7_75t_SL U26601 ( .A(n31532), .B(n31840), .Y(n31525) );
  NOR2x1_ASAP7_75t_SL U26602 ( .A(n23812), .B(n23811), .Y(n23810) );
  NAND2xp33_ASAP7_75t_SL U26603 ( .A(n31852), .B(n31840), .Y(n31839) );
  NAND2xp33_ASAP7_75t_SL U26604 ( .A(n29573), .B(n31840), .Y(n25847) );
  NAND2xp33_ASAP7_75t_SL U26605 ( .A(n31975), .B(n31840), .Y(n26529) );
  NAND2xp33_ASAP7_75t_SL U26606 ( .A(n26477), .B(n31840), .Y(n26461) );
  NAND2xp33_ASAP7_75t_SL U26607 ( .A(n28121), .B(n31840), .Y(n25969) );
  NAND2xp33_ASAP7_75t_SL U26608 ( .A(n26639), .B(n31840), .Y(n26636) );
  NAND2xp33_ASAP7_75t_SL U26609 ( .A(n26610), .B(n31840), .Y(n26607) );
  INVxp33_ASAP7_75t_SRAM U26610 ( .A(n28692), .Y(n26903) );
  AOI22xp33_ASAP7_75t_SL U26611 ( .A1(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DCS__1_), .A2(n30995), .B1(ic_q[3]), 
        .B2(n22387), .Y(n30879) );
  NAND2xp33_ASAP7_75t_SL U26612 ( .A(ic_q[8]), .B(n22387), .Y(n29759) );
  NAND2xp33_ASAP7_75t_SL U26613 ( .A(n30899), .B(n31840), .Y(n30893) );
  OAI21xp33_ASAP7_75t_SL U26614 ( .A1(n28829), .A2(n25198), .B(n25091), .Y(
        n26423) );
  O2A1O1Ixp5_ASAP7_75t_SL U26615 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[2]), .A2(
        n22396), .B(n31304), .C(n31464), .Y(n31305) );
  NAND2x1_ASAP7_75t_SL U26616 ( .A(n26473), .B(n31841), .Y(n31843) );
  NAND2xp33_ASAP7_75t_SL U26617 ( .A(n30803), .B(n31840), .Y(n26604) );
  AOI22xp33_ASAP7_75t_SL U26618 ( .A1(u0_0_leon3x0_p0_c0mmu_mcii[25]), .A2(
        n31877), .B1(u0_0_leon3x0_p0_c0mmu_mcdi[61]), .B2(n24583), .Y(n32751)
         );
  NAND2xp33_ASAP7_75t_SL U26619 ( .A(n26650), .B(n31840), .Y(n26647) );
  NAND2xp33_ASAP7_75t_SL U26620 ( .A(ic_q[10]), .B(n22387), .Y(n30999) );
  OAI21xp33_ASAP7_75t_SL U26621 ( .A1(n30391), .A2(n29595), .B(n27115), .Y(
        n27116) );
  NAND2xp33_ASAP7_75t_SL U26622 ( .A(n26659), .B(n31840), .Y(n26451) );
  NAND2xp33_ASAP7_75t_SL U26623 ( .A(n26654), .B(n31840), .Y(n26651) );
  NAND2xp33_ASAP7_75t_SL U26624 ( .A(n31504), .B(n31840), .Y(n31495) );
  AOI22xp33_ASAP7_75t_SL U26625 ( .A1(it_q[27]), .A2(n24636), .B1(n32659), 
        .B2(n30130), .Y(n25034) );
  INVxp67_ASAP7_75t_SL U26626 ( .A(n22389), .Y(n23195) );
  INVxp33_ASAP7_75t_SL U26627 ( .A(n28978), .Y(n28985) );
  BUFx3_ASAP7_75t_SL U26628 ( .A(DP_OP_1196_128_7433_n2), .Y(n23941) );
  INVxp67_ASAP7_75t_SL U26629 ( .A(n23980), .Y(n23291) );
  INVxp67_ASAP7_75t_SL U26630 ( .A(add_x_735_n225), .Y(add_x_735_n295) );
  OAI22xp33_ASAP7_75t_SL U26631 ( .A1(n30219), .A2(n29595), .B1(n30220), .B2(
        n29594), .Y(n29596) );
  AOI22xp33_ASAP7_75t_SL U26632 ( .A1(n25200), .A2(n22999), .B1(n23665), .B2(
        n22416), .Y(n25096) );
  INVxp67_ASAP7_75t_SL U26633 ( .A(add_x_735_n92), .Y(add_x_735_n279) );
  OAI211xp5_ASAP7_75t_SRAM U26634 ( .A1(n24572), .A2(n29146), .B(
        u0_0_leon3x0_p0_divi[26]), .C(n24580), .Y(n26893) );
  INVxp67_ASAP7_75t_SL U26635 ( .A(n28742), .Y(n30628) );
  OAI21xp33_ASAP7_75t_SL U26636 ( .A1(n28829), .A2(n24469), .B(n25759), .Y(
        n27100) );
  NAND2xp33_ASAP7_75t_SL U26637 ( .A(n22999), .B(n22416), .Y(n26145) );
  INVxp67_ASAP7_75t_SL U26638 ( .A(n31880), .Y(n32452) );
  OAI21xp33_ASAP7_75t_SL U26639 ( .A1(n30366), .A2(n26176), .B(n26175), .Y(
        n26177) );
  OAI22xp33_ASAP7_75t_SL U26640 ( .A1(n30291), .A2(n29595), .B1(n30292), .B2(
        n29594), .Y(n26997) );
  INVx2_ASAP7_75t_SL U26641 ( .A(n24426), .Y(n24636) );
  OAI21xp33_ASAP7_75t_SL U26642 ( .A1(add_x_735_n251), .A2(add_x_735_n247), 
        .B(add_x_735_n248), .Y(add_x_735_n246) );
  AOI22xp33_ASAP7_75t_SL U26643 ( .A1(n28835), .A2(n30383), .B1(
        u0_0_leon3x0_p0_divi[42]), .B2(n28782), .Y(n28688) );
  AOI22xp33_ASAP7_75t_SL U26644 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__12_), 
        .A2(n28935), .B1(n28737), .B2(n28620), .Y(n28641) );
  OAI21xp33_ASAP7_75t_SL U26645 ( .A1(n27521), .A2(n31940), .B(n27514), .Y(
        n27523) );
  INVxp67_ASAP7_75t_SL U26646 ( .A(n29564), .Y(n25820) );
  AOI22xp33_ASAP7_75t_SL U26647 ( .A1(n28835), .A2(n30423), .B1(
        u0_0_leon3x0_p0_divi[36]), .B2(n28782), .Y(n26311) );
  NAND2xp5_ASAP7_75t_SL U26648 ( .A(n29585), .B(n30619), .Y(n28426) );
  INVxp33_ASAP7_75t_SRAM U26649 ( .A(n30656), .Y(n30657) );
  INVx3_ASAP7_75t_SL U26650 ( .A(n31469), .Y(n22387) );
  INVxp67_ASAP7_75t_SL U26651 ( .A(add_x_735_n173), .Y(add_x_735_n288) );
  NAND2xp33_ASAP7_75t_SRAM U26652 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__4_), 
        .B(n26854), .Y(n26864) );
  AOI21xp33_ASAP7_75t_SL U26653 ( .A1(n30611), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__WIM__2_), .B(n28994), .Y(n28938) );
  INVx1_ASAP7_75t_SL U26654 ( .A(DP_OP_1196_128_7433_n206), .Y(
        DP_OP_1196_128_7433_n204) );
  AOI22xp33_ASAP7_75t_SL U26655 ( .A1(u0_0_leon3x0_p0_iu_r_E__ET_), .A2(n30621), .B1(n27294), .B2(n28779), .Y(n26312) );
  AOI21xp33_ASAP7_75t_SL U26656 ( .A1(n28167), .A2(uart1_uarto_SCALER__10_), 
        .B(n22419), .Y(n28143) );
  AOI21xp33_ASAP7_75t_SL U26657 ( .A1(n28167), .A2(uart1_uarto_SCALER__1_), 
        .B(n22419), .Y(n28168) );
  AOI21xp33_ASAP7_75t_SL U26658 ( .A1(n28167), .A2(uart1_uarto_SCALER__2_), 
        .B(n22419), .Y(n28163) );
  AOI21xp33_ASAP7_75t_SL U26659 ( .A1(n28167), .A2(uart1_uarto_SCALER__3_), 
        .B(n22419), .Y(n28159) );
  AOI22xp33_ASAP7_75t_SL U26660 ( .A1(n30697), .A2(n30621), .B1(
        u0_0_leon3x0_p0_iu_r_W__S__TT__6_), .B2(n28779), .Y(n27149) );
  AOI21xp33_ASAP7_75t_SL U26661 ( .A1(n28167), .A2(uart1_uarto_SCALER__4_), 
        .B(n22419), .Y(n28155) );
  NAND2x1p5_ASAP7_75t_SL U26662 ( .A(n25848), .B(n31956), .Y(n31840) );
  OAI21xp33_ASAP7_75t_SL U26663 ( .A1(n27144), .A2(n22392), .B(n25496), .Y(
        n27155) );
  NOR2xp33_ASAP7_75t_SRAM U26664 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[26]), 
        .Y(n26891) );
  AOI22xp33_ASAP7_75t_SL U26665 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__8_), 
        .A2(n24581), .B1(u0_0_leon3x0_p0_iu_r_W__S__TT__4_), .B2(n28779), .Y(
        n28726) );
  INVx1_ASAP7_75t_SL U26666 ( .A(DP_OP_1196_128_7433_n178), .Y(
        DP_OP_1196_128_7433_n176) );
  AOI22xp33_ASAP7_75t_SRAM U26667 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__18_), 
        .A2(n22375), .B1(n28540), .B2(n28403), .Y(n25712) );
  NAND2xp5_ASAP7_75t_SL U26668 ( .A(sr1_r_MCFG1__IOWS__2_), .B(n32003), .Y(
        n31644) );
  AOI22xp33_ASAP7_75t_SRAM U26669 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__16_), 
        .A2(n22375), .B1(n28554), .B2(n28403), .Y(n26445) );
  HB1xp67_ASAP7_75t_SL U26670 ( .A(n18610), .Y(n23154) );
  NAND2xp5_ASAP7_75t_SL U26671 ( .A(sr1_r_MCFG1__IOWS__3_), .B(n32003), .Y(
        n31972) );
  AOI21xp33_ASAP7_75t_SL U26672 ( .A1(n28167), .A2(uart1_uarto_SCALER__9_), 
        .B(n22419), .Y(n28147) );
  INVx1_ASAP7_75t_SL U26673 ( .A(DP_OP_1196_128_7433_n353), .Y(
        DP_OP_1196_128_7433_n352) );
  INVxp67_ASAP7_75t_SL U26674 ( .A(u0_0_leon3x0_p0_divi[5]), .Y(n22417) );
  INVxp67_ASAP7_75t_SL U26675 ( .A(u0_0_leon3x0_p0_divi[12]), .Y(n26168) );
  NAND2xp5_ASAP7_75t_SL U26676 ( .A(n31398), .B(n28601), .Y(n29617) );
  NAND2xp5_ASAP7_75t_SL U26677 ( .A(n26055), .B(n26053), .Y(n31171) );
  NOR2x1_ASAP7_75t_SL U26678 ( .A(n31402), .B(n24511), .Y(n31403) );
  XNOR2xp5_ASAP7_75t_SL U26679 ( .A(n24054), .B(n23089), .Y(n23394) );
  NAND2xp5_ASAP7_75t_SL U26680 ( .A(n26036), .B(n26066), .Y(n31139) );
  NAND2xp5_ASAP7_75t_SL U26681 ( .A(n26032), .B(n26066), .Y(n31143) );
  XNOR2xp5_ASAP7_75t_SL U26682 ( .A(n23969), .B(n24048), .Y(mult_x_1196_n2911)
         );
  NAND2xp5_ASAP7_75t_SL U26683 ( .A(n26068), .B(n26053), .Y(n31059) );
  OAI21xp33_ASAP7_75t_SRAM U26684 ( .A1(irqctrl0_r_IFORCE__0__7_), .A2(n29282), 
        .B(n24694), .Y(n29284) );
  INVx1_ASAP7_75t_SL U26685 ( .A(n30616), .Y(n28994) );
  NAND2xp5_ASAP7_75t_SL U26686 ( .A(n26049), .B(n26053), .Y(n31167) );
  OAI21xp33_ASAP7_75t_SL U26687 ( .A1(n27464), .A2(n30134), .B(n24694), .Y(
        n29514) );
  OAI21xp33_ASAP7_75t_SL U26688 ( .A1(n28931), .A2(n22999), .B(n24632), .Y(
        n26740) );
  NAND2xp5_ASAP7_75t_SL U26689 ( .A(n26045), .B(n26053), .Y(n31131) );
  NAND2xp5_ASAP7_75t_SL U26690 ( .A(n26036), .B(n26053), .Y(n31151) );
  NAND2xp5_ASAP7_75t_SL U26691 ( .A(n26062), .B(n26066), .Y(n31163) );
  NAND2xp5_ASAP7_75t_SL U26692 ( .A(n22906), .B(n28982), .Y(n26253) );
  NOR2xp33_ASAP7_75t_SRAM U26693 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__19_), 
        .B(n28637), .Y(n25766) );
  AOI21xp33_ASAP7_75t_SRAM U26694 ( .A1(n29697), .A2(n29224), .B(n29223), .Y(
        n29226) );
  NAND2xp33_ASAP7_75t_SL U26695 ( .A(n31336), .B(n28554), .Y(n27242) );
  BUFx2_ASAP7_75t_SL U26696 ( .A(n22423), .Y(n22556) );
  AOI21xp33_ASAP7_75t_SL U26697 ( .A1(n28888), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__16_), .B(n28887), .Y(n26676) );
  BUFx3_ASAP7_75t_SL U26698 ( .A(n29018), .Y(n24629) );
  AOI21xp33_ASAP7_75t_SL U26699 ( .A1(n28888), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__10_), .B(n27148), .Y(n27150) );
  AOI21xp33_ASAP7_75t_SL U26700 ( .A1(n24582), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__20_), .B(n28887), .Y(n26994) );
  INVx1_ASAP7_75t_SL U26701 ( .A(n26947), .Y(n28272) );
  OAI21xp33_ASAP7_75t_SL U26702 ( .A1(n31574), .A2(n25398), .B(n24684), .Y(
        n25400) );
  INVx3_ASAP7_75t_SL U26703 ( .A(n26338), .Y(n22392) );
  OAI21xp5_ASAP7_75t_SL U26704 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__26_), 
        .A2(n24652), .B(n28394), .Y(n3258) );
  NOR2xp33_ASAP7_75t_SL U26705 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__19_), 
        .B(n26762), .Y(n26796) );
  AOI22xp33_ASAP7_75t_SL U26706 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__14_), .B1(u0_0_leon3x0_p0_divo[14]), .B2(
        n28371), .Y(n28331) );
  OAI21xp5_ASAP7_75t_SL U26707 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__14_), 
        .A2(n24650), .B(n27184), .Y(n3206) );
  OAI21xp5_ASAP7_75t_SL U26708 ( .A1(u0_0_leon3x0_p0_ici[54]), .A2(n24652), 
        .B(n28390), .Y(n3262) );
  OAI21xp5_ASAP7_75t_SL U26709 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__26_), 
        .A2(n24652), .B(n28392), .Y(n3260) );
  AOI22xp33_ASAP7_75t_SL U26710 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__20_), .B1(u0_0_leon3x0_p0_divo[20]), .B2(
        n28371), .Y(n28317) );
  OAI21xp5_ASAP7_75t_SL U26711 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__21_), 
        .A2(n24651), .B(n27048), .Y(n3234) );
  OAI21xp5_ASAP7_75t_SL U26712 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__16_), 
        .A2(n24651), .B(n27236), .Y(n2619) );
  OAI21xp5_ASAP7_75t_SL U26713 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__26_), 
        .A2(n24652), .B(n28396), .Y(n3256) );
  AOI22xp33_ASAP7_75t_SL U26714 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__22_), .B1(u0_0_leon3x0_p0_divo[22]), .B2(
        n28371), .Y(n28314) );
  AOI22xp33_ASAP7_75t_SL U26715 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__16_), .B1(u0_0_leon3x0_p0_divo[16]), .B2(
        n28371), .Y(n28325) );
  INVxp33_ASAP7_75t_SL U26716 ( .A(DP_OP_1196_128_7433_n108), .Y(
        DP_OP_1196_128_7433_n365) );
  NAND2xp33_ASAP7_75t_SL U26717 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__9_), 
        .B(n28888), .Y(n27113) );
  AOI22xp33_ASAP7_75t_SL U26718 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__7_), .B1(u0_0_leon3x0_p0_divo[7]), .B2(
        n28371), .Y(n28348) );
  AOI22xp33_ASAP7_75t_SL U26719 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__9_), .B1(u0_0_leon3x0_p0_divo[9]), .B2(
        n28371), .Y(n28342) );
  NOR2xp33_ASAP7_75t_SL U26720 ( .A(n25989), .B(n25988), .Y(n27473) );
  INVx3_ASAP7_75t_SL U26721 ( .A(n32270), .Y(n22396) );
  AOI22xp33_ASAP7_75t_SL U26722 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__8_), .B1(u0_0_leon3x0_p0_divo[8]), .B2(
        n28371), .Y(n28345) );
  AOI22xp33_ASAP7_75t_SL U26723 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__11_), .B1(u0_0_leon3x0_p0_divo[11]), .B2(
        n28371), .Y(n28338) );
  INVx2_ASAP7_75t_SL U26724 ( .A(n31676), .Y(n31421) );
  AOI22xp33_ASAP7_75t_SL U26725 ( .A1(n22431), .A2(n28295), .B1(
        u0_0_leon3x0_p0_divo[33]), .B2(n28371), .Y(n28296) );
  INVx2_ASAP7_75t_SL U26726 ( .A(n24491), .Y(n22374) );
  AOI22xp33_ASAP7_75t_SL U26727 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__30_), .B1(u0_0_leon3x0_p0_divo[30]), .B2(
        n28371), .Y(n28299) );
  AOI22xp33_ASAP7_75t_SL U26728 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__10_), .B1(u0_0_leon3x0_p0_divo[10]), .B2(
        n28371), .Y(n28340) );
  NAND2xp33_ASAP7_75t_SL U26729 ( .A(n29734), .B(n32075), .Y(n29735) );
  AOI22xp33_ASAP7_75t_SL U26730 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__6_), .B1(u0_0_leon3x0_p0_divo[6]), .B2(
        n28371), .Y(n28350) );
  INVx4_ASAP7_75t_SL U26731 ( .A(n31677), .Y(n31662) );
  NAND2xp33_ASAP7_75t_SL U26732 ( .A(n26482), .B(n27065), .Y(n26394) );
  INVx1_ASAP7_75t_SL U26733 ( .A(n31398), .Y(n31340) );
  INVxp33_ASAP7_75t_SL U26734 ( .A(n22421), .Y(n23589) );
  AOI22xp33_ASAP7_75t_SL U26735 ( .A1(uart1_r_RHOLD__27__6_), .A2(n31230), 
        .B1(n31229), .B2(uart1_r_RHOLD__22__6_), .Y(n31231) );
  AOI22xp33_ASAP7_75t_SL U26736 ( .A1(u0_0_leon3x0_p0_divi[32]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[31]), .B2(n28367), .Y(n28369) );
  AOI22xp33_ASAP7_75t_SL U26737 ( .A1(uart1_r_RHOLD__31__1_), .A2(n31221), 
        .B1(n31220), .B2(uart1_r_RHOLD__13__1_), .Y(n27440) );
  NAND2xp33_ASAP7_75t_SL U26738 ( .A(n27526), .B(n27525), .Y(n27533) );
  AOI22xp33_ASAP7_75t_SL U26739 ( .A1(n31205), .A2(uart1_r_RHOLD__16__1_), 
        .B1(uart1_r_RHOLD__9__1_), .B2(n31204), .Y(n27435) );
  INVxp67_ASAP7_75t_SL U26740 ( .A(n32430), .Y(n32659) );
  AOI22xp33_ASAP7_75t_SL U26741 ( .A1(n31229), .A2(uart1_r_RHOLD__22__1_), 
        .B1(uart1_r_RHOLD__27__1_), .B2(n31230), .Y(n27452) );
  AOI22xp33_ASAP7_75t_SL U26742 ( .A1(uart1_r_RHOLD__6__1_), .A2(n31226), .B1(
        n31225), .B2(uart1_r_RHOLD__10__1_), .Y(n27454) );
  AOI22xp33_ASAP7_75t_SL U26743 ( .A1(uart1_r_RHOLD__4__1_), .A2(n31224), .B1(
        n31223), .B2(uart1_r_RHOLD__2__1_), .Y(n27455) );
  NAND2x1_ASAP7_75t_SL U26744 ( .A(n22397), .B(n32888), .Y(n31638) );
  INVx2_ASAP7_75t_SL U26745 ( .A(n24682), .Y(n24679) );
  AOI22xp33_ASAP7_75t_SL U26746 ( .A1(ahbso_0__HRDATA__23_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__23_), .Y(n32384) );
  INVx5_ASAP7_75t_SL U26747 ( .A(n24423), .Y(n22431) );
  NOR2x1_ASAP7_75t_SL U26748 ( .A(n25210), .B(n25209), .Y(n31392) );
  INVxp33_ASAP7_75t_SL U26749 ( .A(n28481), .Y(n28935) );
  OR2x4_ASAP7_75t_SL U26750 ( .A(n24899), .B(n31420), .Y(n28371) );
  INVx3_ASAP7_75t_SL U26751 ( .A(n24428), .Y(n24638) );
  INVxp67_ASAP7_75t_SL U26752 ( .A(n32888), .Y(n32909) );
  NOR2xp33_ASAP7_75t_SL U26753 ( .A(n5061), .B(n1634), .Y(timer0_N79) );
  INVxp67_ASAP7_75t_SL U26754 ( .A(n33054), .Y(n32077) );
  NAND2xp33_ASAP7_75t_SL U26755 ( .A(uart1_uarto_SCALER__0_), .B(n28172), .Y(
        n28173) );
  INVx3_ASAP7_75t_SL U26756 ( .A(n24427), .Y(n24634) );
  INVx2_ASAP7_75t_SL U26757 ( .A(n30637), .Y(n22398) );
  NAND2xp33_ASAP7_75t_SL U26758 ( .A(n31380), .B(n32091), .Y(n32101) );
  INVx3_ASAP7_75t_SL U26759 ( .A(n31639), .Y(n22397) );
  INVx2_ASAP7_75t_SL U26760 ( .A(n24632), .Y(n24631) );
  A2O1A1Ixp33_ASAP7_75t_SL U26761 ( .A1(n31904), .A2(n32677), .B(n31903), .C(
        u0_0_leon3x0_p0_ici[62]), .Y(n31905) );
  INVxp33_ASAP7_75t_SL U26762 ( .A(n32237), .Y(n25008) );
  INVx1_ASAP7_75t_SL U26763 ( .A(DP_OP_1196_128_7433_n336), .Y(
        DP_OP_1196_128_7433_n334) );
  INVxp33_ASAP7_75t_SL U26764 ( .A(n26352), .Y(n26353) );
  INVx1_ASAP7_75t_SL U26765 ( .A(DP_OP_1196_128_7433_n277), .Y(
        DP_OP_1196_128_7433_n378) );
  NAND2xp5_ASAP7_75t_SL U26766 ( .A(u0_0_leon3x0_p0_iu_r_X__NPC__0_), .B(
        n25736), .Y(n25738) );
  NAND2xp5_ASAP7_75t_SL U26767 ( .A(u0_0_leon3x0_p0_iu_r_X__NPC__1_), .B(
        n25733), .Y(n25734) );
  NOR2x1_ASAP7_75t_SL U26768 ( .A(n25031), .B(n32037), .Y(n29999) );
  INVxp67_ASAP7_75t_SL U26769 ( .A(uart1_r_TRADDR__0_), .Y(n27411) );
  INVxp67_ASAP7_75t_SL U26770 ( .A(n25151), .Y(n25153) );
  NOR2xp33_ASAP7_75t_SRAM U26771 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_), .B(n32250), .Y(n32241) );
  NOR2x1_ASAP7_75t_SL U26772 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__0_), .B(
        n26731), .Y(n30640) );
  OR2x2_ASAP7_75t_SL U26773 ( .A(n3725), .B(n28291), .Y(n24423) );
  INVxp33_ASAP7_75t_SRAM U26774 ( .A(n32084), .Y(n31859) );
  NAND2xp33_ASAP7_75t_SL U26775 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), 
        .B(n25695), .Y(n25693) );
  INVxp33_ASAP7_75t_SL U26776 ( .A(n25697), .Y(n25699) );
  NAND2xp5_ASAP7_75t_SL U26777 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__2_), .B(
        n26729), .Y(n26730) );
  NAND2xp33_ASAP7_75t_SL U26778 ( .A(it_q[7]), .B(u0_0_leon3x0_p0_ici[60]), 
        .Y(n31902) );
  INVxp67_ASAP7_75t_SL U26779 ( .A(u0_0_leon3x0_p0_divi[47]), .Y(n30334) );
  INVxp67_ASAP7_75t_SL U26780 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__2_), .Y(
        n25894) );
  INVx1_ASAP7_75t_SL U26781 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .Y(n26482) );
  INVx1_ASAP7_75t_SL U26782 ( .A(u0_0_leon3x0_p0_ici[62]), .Y(n29481) );
  INVxp67_ASAP7_75t_SL U26783 ( .A(ramsn[2]), .Y(n32805) );
  INVx1_ASAP7_75t_SL U26784 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TT__4_), .Y(n29734) );
  INVxp67_ASAP7_75t_SL U26785 ( .A(u0_0_leon3x0_p0_div0_r_CNT__1_), .Y(n24902)
         );
  NAND2xp5_ASAP7_75t_SL U26786 ( .A(u0_0_leon3x0_p0_iu_r_X__NPC__1_), .B(
        u0_0_leon3x0_p0_iu_r_X__NPC__0_), .Y(n25735) );
  INVxp33_ASAP7_75t_SL U26787 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PV_), .Y(
        n30685) );
  INVxp67_ASAP7_75t_SL U26788 ( .A(u0_0_leon3x0_p0_divi[54]), .Y(n30265) );
  INVxp33_ASAP7_75t_SL U26789 ( .A(n3897), .Y(n25569) );
  INVxp67_ASAP7_75t_SL U26790 ( .A(n4391), .Y(n25031) );
  INVxp67_ASAP7_75t_SL U26791 ( .A(uart1_r_BRATE__9_), .Y(n28148) );
  INVxp33_ASAP7_75t_SL U26792 ( .A(u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__1_), .Y(
        n24972) );
  INVxp67_ASAP7_75t_SL U26793 ( .A(u0_0_leon3x0_p0_divi[53]), .Y(n30273) );
  INVx1_ASAP7_75t_SL U26794 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__2_), .Y(n26733) );
  NAND2xp5_ASAP7_75t_SL U26795 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .Y(n28931) );
  INVxp67_ASAP7_75t_SL U26796 ( .A(ramsn[0]), .Y(n32794) );
  INVx1_ASAP7_75t_SL U26797 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__15_), .Y(
        n30339) );
  INVxp33_ASAP7_75t_SL U26798 ( .A(n4927), .Y(n26820) );
  INVx1_ASAP7_75t_SL U26799 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__0_), .Y(n26747)
         );
  INVxp33_ASAP7_75t_SRAM U26800 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__LD_), .Y(
        n31864) );
  INVx1_ASAP7_75t_SL U26801 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__20_), .Y(
        n30285) );
  INVxp67_ASAP7_75t_SL U26802 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__18_), .Y(
        n30309) );
  INVxp67_ASAP7_75t_SL U26803 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__6_), .Y(
        n26260) );
  INVxp67_ASAP7_75t_SL U26804 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__19_), .Y(
        n30300) );
  INVxp67_ASAP7_75t_SL U26805 ( .A(u0_0_leon3x0_p0_divi[55]), .Y(n30258) );
  INVxp67_ASAP7_75t_SL U26806 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_), 
        .Y(n32137) );
  INVxp67_ASAP7_75t_SL U26807 ( .A(uart1_r_RHOLD__24__0_), .Y(n28093) );
  INVxp67_ASAP7_75t_SL U26808 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__13_), .Y(
        n30363) );
  INVx1_ASAP7_75t_SL U26809 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__22_), .Y(
        n30267) );
  INVxp67_ASAP7_75t_SL U26810 ( .A(u0_0_leon3x0_p0_iu_r_E__SHCNT__2_), .Y(
        n25082) );
  INVxp67_ASAP7_75t_SL U26811 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__15_), .Y(
        n30342) );
  INVxp67_ASAP7_75t_SL U26812 ( .A(uart1_r_BRATE__1_), .Y(n28169) );
  INVxp67_ASAP7_75t_SL U26813 ( .A(uart1_r_BRATE__10_), .Y(n28144) );
  INVx1_ASAP7_75t_SL U26814 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[26]), .Y(n25250)
         );
  INVxp33_ASAP7_75t_SL U26815 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__27_), .Y(
        n26956) );
  INVxp33_ASAP7_75t_SL U26816 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__30_), .Y(n25621) );
  INVxp33_ASAP7_75t_SL U26817 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__15_), .Y(
        n27243) );
  INVxp67_ASAP7_75t_SL U26818 ( .A(uart1_r_RHOLD__0__0_), .Y(n28095) );
  INVxp67_ASAP7_75t_SL U26819 ( .A(n2356), .Y(n31719) );
  INVx1_ASAP7_75t_SL U26820 ( .A(sr1_r_MCFG1__BRDYEN_), .Y(n31696) );
  INVxp67_ASAP7_75t_SL U26821 ( .A(uart1_r_BRATE__2_), .Y(n28164) );
  INVxp67_ASAP7_75t_SL U26822 ( .A(u0_0_leon3x0_p0_divo[6]), .Y(n28352) );
  INVxp67_ASAP7_75t_SL U26823 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[53]), .Y(n31770)
         );
  INVx1_ASAP7_75t_SL U26824 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__0_), .Y(
        n32094) );
  NAND2xp5_ASAP7_75t_SL U26825 ( .A(u0_0_leon3x0_p0_iu_r_A__BP_), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__29_), .Y(n24847) );
  INVxp67_ASAP7_75t_SL U26826 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__5_), .Y(
        n30421) );
  INVxp67_ASAP7_75t_SL U26827 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__6_), .Y(
        n30409) );
  INVxp67_ASAP7_75t_SL U26828 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__7_), .Y(
        n30399) );
  INVxp67_ASAP7_75t_SL U26829 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[56]), .Y(n31763)
         );
  INVxp67_ASAP7_75t_SL U26830 ( .A(u0_0_leon3x0_p0_iu_r_A__CTRL__WREG_), .Y(
        n24816) );
  INVxp33_ASAP7_75t_SL U26831 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__6_), .Y(n29903) );
  NAND2xp5_ASAP7_75t_SL U26832 ( .A(n2389), .B(n4715), .Y(n27444) );
  INVxp33_ASAP7_75t_SL U26833 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__7_), .Y(n29928) );
  INVxp67_ASAP7_75t_SL U26834 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__21_), .Y(
        n30279) );
  INVxp67_ASAP7_75t_SL U26835 ( .A(sr1_r_MCFG1__ROMWIDTH__0_), .Y(n32876) );
  INVxp33_ASAP7_75t_SL U26836 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__25_), .Y(
        n29805) );
  INVxp33_ASAP7_75t_SL U26837 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_), 
        .Y(n32130) );
  INVxp33_ASAP7_75t_SL U26838 ( .A(n4929), .Y(n26827) );
  INVxp67_ASAP7_75t_SL U26839 ( .A(u0_0_leon3x0_p0_iu_r_A__CTRL__ANNUL_), .Y(
        n32066) );
  INVx1_ASAP7_75t_SL U26840 ( .A(dt_q[17]), .Y(n31278) );
  OAI21xp5_ASAP7_75t_SL U26841 ( .A1(n22428), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N42), .B(n25282), .Y(n4231) );
  OAI21xp5_ASAP7_75t_SL U26842 ( .A1(n26520), .A2(n22399), .B(n26519), .Y(
        timer0_v_TIMERS__1__VALUE__24_) );
  OAI21xp5_ASAP7_75t_SL U26843 ( .A1(n26626), .A2(n22399), .B(n26625), .Y(
        timer0_v_TIMERS__1__VALUE__8_) );
  OAI21xp5_ASAP7_75t_SL U26844 ( .A1(n29988), .A2(n22399), .B(n26494), .Y(
        timer0_v_TIMERS__1__VALUE__29_) );
  OAI21xp5_ASAP7_75t_SL U26845 ( .A1(n26550), .A2(n22399), .B(n26549), .Y(
        timer0_v_TIMERS__1__VALUE__17_) );
  OAI21xp5_ASAP7_75t_SL U26846 ( .A1(n26639), .A2(n22399), .B(n26638), .Y(
        timer0_v_TIMERS__1__VALUE__4_) );
  OAI21xp5_ASAP7_75t_SL U26847 ( .A1(n30151), .A2(n22399), .B(n26622), .Y(
        timer0_v_TIMERS__1__VALUE__9_) );
  OAI21xp5_ASAP7_75t_SL U26848 ( .A1(n31021), .A2(n22399), .B(n26593), .Y(
        timer0_v_TIMERS__1__VALUE__15_) );
  OAI21xp5_ASAP7_75t_SL U26849 ( .A1(n26610), .A2(n22399), .B(n26609), .Y(
        timer0_v_TIMERS__1__VALUE__12_) );
  OAI21xp5_ASAP7_75t_SL U26850 ( .A1(n31532), .A2(n22399), .B(n31528), .Y(
        timer0_v_TIMERS__1__VALUE__20_) );
  OAI21xp5_ASAP7_75t_SL U26851 ( .A1(n31328), .A2(n22399), .B(n26500), .Y(
        timer0_v_TIMERS__1__VALUE__26_) );
  OAI21xp5_ASAP7_75t_SL U26852 ( .A1(n31244), .A2(n22399), .B(n26632), .Y(
        timer0_v_TIMERS__1__VALUE__6_) );
  OAI21xp5_ASAP7_75t_SL U26853 ( .A1(n32005), .A2(n22399), .B(n26546), .Y(
        timer0_v_TIMERS__1__VALUE__19_) );
  OAI21xp5_ASAP7_75t_SL U26854 ( .A1(n29573), .A2(n22399), .B(n29572), .Y(
        timer0_v_TIMERS__1__VALUE__18_) );
  OAI21xp5_ASAP7_75t_SL U26855 ( .A1(n30549), .A2(n22399), .B(n26596), .Y(
        timer0_v_TIMERS__1__VALUE__14_) );
  OAI21xp5_ASAP7_75t_SL U26856 ( .A1(n31975), .A2(n22399), .B(n26532), .Y(
        timer0_v_TIMERS__1__VALUE__23_) );
  OAI21xp5_ASAP7_75t_SL U26857 ( .A1(n30106), .A2(n22399), .B(n26635), .Y(
        timer0_v_TIMERS__1__VALUE__5_) );
  OAI21xp5_ASAP7_75t_SL U26858 ( .A1(n31646), .A2(n22399), .B(n31643), .Y(
        timer0_v_TIMERS__1__VALUE__22_) );
  OAI21xp5_ASAP7_75t_SL U26859 ( .A1(n31941), .A2(n22399), .B(n26481), .Y(
        timer0_v_TIMERS__1__VALUE__30_) );
  OAI21xp5_ASAP7_75t_SL U26860 ( .A1(n22427), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N29), .B(n29087), .Y(n4257) );
  OAI21xp5_ASAP7_75t_SL U26861 ( .A1(n28121), .A2(n22399), .B(n28118), .Y(
        timer0_v_TIMERS__1__VALUE__11_) );
  OAI21xp5_ASAP7_75t_SL U26862 ( .A1(n30874), .A2(n22399), .B(n26629), .Y(
        timer0_v_TIMERS__1__VALUE__7_) );
  OAI21xp5_ASAP7_75t_SL U26863 ( .A1(n26619), .A2(n22399), .B(n26618), .Y(
        timer0_v_TIMERS__1__VALUE__10_) );
  OAI21xp5_ASAP7_75t_SL U26864 ( .A1(n26650), .A2(n22399), .B(n26649), .Y(
        timer0_v_TIMERS__1__VALUE__1_) );
  OAI21xp5_ASAP7_75t_SL U26865 ( .A1(n31504), .A2(n22399), .B(n31498), .Y(
        timer0_v_TIMERS__1__VALUE__28_) );
  OAI21xp5_ASAP7_75t_SL U26866 ( .A1(n31373), .A2(n22399), .B(n31370), .Y(
        timer0_v_TIMERS__1__VALUE__25_) );
  OAI21xp5_ASAP7_75t_SL U26867 ( .A1(n26659), .A2(n22399), .B(n26657), .Y(
        timer0_v_TIMERS__1__VALUE__16_) );
  OAI21xp5_ASAP7_75t_SL U26868 ( .A1(n26477), .A2(n22399), .B(n26476), .Y(
        timer0_v_TIMERS__1__VALUE__31_) );
  OAI21xp5_ASAP7_75t_SL U26869 ( .A1(n30803), .A2(n22399), .B(n26606), .Y(
        timer0_v_TIMERS__1__VALUE__13_) );
  AOI21xp5_ASAP7_75t_SL U26870 ( .A1(n31845), .A2(timer0_res_17_), .B(n26548), 
        .Y(n26549) );
  AOI21xp5_ASAP7_75t_SL U26871 ( .A1(n31845), .A2(timer0_res_8_), .B(n26624), 
        .Y(n26625) );
  AOI21xp5_ASAP7_75t_SL U26872 ( .A1(n31845), .A2(timer0_res_1_), .B(n26648), 
        .Y(n26649) );
  AOI21xp5_ASAP7_75t_SL U26873 ( .A1(n31845), .A2(timer0_res_3_), .B(n26641), 
        .Y(n26642) );
  OAI21xp5_ASAP7_75t_SL U26874 ( .A1(n22427), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N27), .B(n29089), .Y(n4261) );
  AOI21xp5_ASAP7_75t_SL U26875 ( .A1(n31845), .A2(timer0_res_28_), .B(n31497), 
        .Y(n31498) );
  AOI21xp5_ASAP7_75t_SL U26876 ( .A1(n31845), .A2(timer0_res_15_), .B(n26592), 
        .Y(n26593) );
  AOI21xp5_ASAP7_75t_SL U26877 ( .A1(n31845), .A2(timer0_res_25_), .B(n31369), 
        .Y(n31370) );
  INVx1_ASAP7_75t_SL U26878 ( .A(mult_x_1196_n418), .Y(n22517) );
  AOI21xp5_ASAP7_75t_SL U26879 ( .A1(n31845), .A2(timer0_res_10_), .B(n26617), 
        .Y(n26618) );
  AOI21xp5_ASAP7_75t_SL U26880 ( .A1(n31845), .A2(timer0_res_20_), .B(n31527), 
        .Y(n31528) );
  AOI21xp5_ASAP7_75t_SL U26881 ( .A1(n31845), .A2(timer0_res_22_), .B(n31642), 
        .Y(n31643) );
  AOI21xp5_ASAP7_75t_SL U26882 ( .A1(n31845), .A2(timer0_res_11_), .B(n28117), 
        .Y(n28118) );
  AOI21xp5_ASAP7_75t_SL U26883 ( .A1(n31845), .A2(timer0_res_16_), .B(n26656), 
        .Y(n26657) );
  AOI21xp5_ASAP7_75t_SL U26884 ( .A1(n31845), .A2(timer0_res_9_), .B(n26621), 
        .Y(n26622) );
  AOI21xp5_ASAP7_75t_SL U26885 ( .A1(n31845), .A2(timer0_res_18_), .B(n29571), 
        .Y(n29572) );
  AOI21xp33_ASAP7_75t_SL U26886 ( .A1(n31845), .A2(n18882), .B(n26475), .Y(
        n26476) );
  OAI21xp5_ASAP7_75t_SL U26887 ( .A1(n22427), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N20), .B(n27266), .Y(n4275) );
  AOI21xp33_ASAP7_75t_SL U26888 ( .A1(n22254), .A2(mult_x_1196_n813), .B(
        mult_x_1196_n644), .Y(mult_x_1196_n642) );
  AOI22xp33_ASAP7_75t_SL U26889 ( .A1(n30186), .A2(n30178), .B1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__5_), .B2(n30182), .Y(n3047) );
  OAI22xp33_ASAP7_75t_SL U26890 ( .A1(n30808), .A2(n24637), .B1(n29993), .B2(
        n23893), .Y(n29994) );
  OAI22xp33_ASAP7_75t_SL U26891 ( .A1(n32328), .A2(n24637), .B1(n32329), .B2(
        n23893), .Y(n30994) );
  OAI22xp33_ASAP7_75t_SL U26892 ( .A1(n32419), .A2(n24637), .B1(n32418), .B2(
        n23893), .Y(n30572) );
  AOI21xp33_ASAP7_75t_SL U26893 ( .A1(n30182), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__0_), .B(n30164), .Y(n3052) );
  OAI22xp33_ASAP7_75t_SL U26894 ( .A1(n32306), .A2(n24637), .B1(n32305), .B2(
        n23893), .Y(n29506) );
  INVxp67_ASAP7_75t_SL U26895 ( .A(n30182), .Y(n30162) );
  OAI22xp33_ASAP7_75t_SL U26896 ( .A1(n31032), .A2(n24637), .B1(n31031), .B2(
        n23893), .Y(n31033) );
  OAI22xp33_ASAP7_75t_SL U26897 ( .A1(n32430), .A2(n24637), .B1(n32432), .B2(
        n23893), .Y(n31041) );
  AOI22xp33_ASAP7_75t_SL U26898 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[30]), .A2(
        n24644), .B1(n31999), .B2(n23885), .Y(n32001) );
  OAI22xp33_ASAP7_75t_SL U26899 ( .A1(n30876), .A2(n24637), .B1(n32317), .B2(
        n23893), .Y(n29911) );
  OAI21xp33_ASAP7_75t_SL U26900 ( .A1(n24645), .A2(n30918), .B(n30917), .Y(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__3_) );
  OAI22xp33_ASAP7_75t_SL U26901 ( .A1(n30557), .A2(n24637), .B1(n30556), .B2(
        n23893), .Y(n30558) );
  OAI22xp33_ASAP7_75t_SL U26902 ( .A1(n32303), .A2(n24637), .B1(n32302), .B2(
        n23893), .Y(n29565) );
  NAND2xp5_ASAP7_75t_SL U26903 ( .A(n31305), .B(n31599), .Y(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_XADDRESS__2_) );
  OAI22xp33_ASAP7_75t_SL U26904 ( .A1(n32322), .A2(n24637), .B1(n32320), .B2(
        n23893), .Y(n29758) );
  OAI22xp33_ASAP7_75t_SL U26905 ( .A1(n32311), .A2(n24637), .B1(n32310), .B2(
        n23893), .Y(n30011) );
  OAI21xp5_ASAP7_75t_SL U26906 ( .A1(n22427), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N18), .B(n28564), .Y(n4279) );
  OAI22xp33_ASAP7_75t_SL U26907 ( .A1(n32384), .A2(n24637), .B1(n32387), .B2(
        n23893), .Y(n29908) );
  OAI22xp33_ASAP7_75t_SL U26908 ( .A1(n30829), .A2(n24645), .B1(n32636), .B2(
        n32729), .Y(n30830) );
  OAI22xp33_ASAP7_75t_SL U26909 ( .A1(n31770), .A2(n24645), .B1(n32638), .B2(
        n32729), .Y(n31771) );
  OAI22xp33_ASAP7_75t_SL U26910 ( .A1(n31774), .A2(n24645), .B1(n32642), .B2(
        n32729), .Y(n31775) );
  INVxp67_ASAP7_75t_SL U26911 ( .A(mult_x_1196_n487), .Y(mult_x_1196_n485) );
  OAI22xp33_ASAP7_75t_SL U26912 ( .A1(n31763), .A2(n24645), .B1(n32644), .B2(
        n32729), .Y(n31764) );
  OAI22xp33_ASAP7_75t_SL U26913 ( .A1(n31776), .A2(n24645), .B1(n32729), .B2(
        n32646), .Y(n31777) );
  OAI22xp33_ASAP7_75t_SL U26914 ( .A1(n31784), .A2(n24645), .B1(n32729), .B2(
        n32648), .Y(n31785) );
  OAI21xp33_ASAP7_75t_SL U26915 ( .A1(n3065), .A2(n31562), .B(n32545), .Y(
        n3063) );
  OAI22xp33_ASAP7_75t_SL U26916 ( .A1(n32714), .A2(n24645), .B1(n32713), .B2(
        n32735), .Y(n32715) );
  BUFx6f_ASAP7_75t_SL U26917 ( .A(n31637), .Y(n22382) );
  OAI22xp33_ASAP7_75t_SL U26918 ( .A1(n22422), .A2(n28377), .B1(n4949), .B2(
        n31672), .Y(n18171) );
  OAI21xp5_ASAP7_75t_SL U26919 ( .A1(n22427), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N16), .B(n27178), .Y(n4283) );
  OAI21xp33_ASAP7_75t_SL U26920 ( .A1(n22379), .A2(u0_0_leon3x0_p0_ici[64]), 
        .B(n26240), .Y(n3944) );
  OAI21xp33_ASAP7_75t_SL U26921 ( .A1(n23229), .A2(u0_0_leon3x0_p0_ici[69]), 
        .B(n28662), .Y(n4478) );
  INVxp67_ASAP7_75t_SL U26922 ( .A(n24088), .Y(n24087) );
  NOR2x1_ASAP7_75t_SL U26923 ( .A(n32198), .B(n25591), .Y(n31568) );
  OAI21xp5_ASAP7_75t_SL U26924 ( .A1(n22427), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N14), .B(n28658), .Y(n4287) );
  NOR2x1_ASAP7_75t_SL U26925 ( .A(n30509), .B(n32025), .Y(n25592) );
  INVx1_ASAP7_75t_SL U26926 ( .A(mult_x_1196_n636), .Y(n23450) );
  OAI21xp5_ASAP7_75t_SL U26927 ( .A1(n32301), .A2(n22402), .B(n26824), .Y(
        n18212) );
  OAI21xp5_ASAP7_75t_SL U26928 ( .A1(n32297), .A2(n22402), .B(n26821), .Y(
        n18213) );
  OAI21xp5_ASAP7_75t_SL U26929 ( .A1(n32303), .A2(n22402), .B(n26828), .Y(
        n18211) );
  OAI21xp5_ASAP7_75t_SL U26930 ( .A1(n32306), .A2(n22402), .B(n28256), .Y(
        n18210) );
  NOR2xp33_ASAP7_75t_SL U26931 ( .A(mult_x_1196_n361), .B(n22406), .Y(n23672)
         );
  OAI21xp33_ASAP7_75t_SL U26932 ( .A1(n22427), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N13), .B(n26189), .Y(n4289) );
  OR3x1_ASAP7_75t_SL U26933 ( .A(n31257), .B(n25587), .C(n32198), .Y(n24549)
         );
  AOI21xp5_ASAP7_75t_SL U26934 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_6_), .A2(n31833), .B(n26239), .Y(n32572) );
  OAI21xp5_ASAP7_75t_SL U26935 ( .A1(n32640), .A2(n18851), .B(n31546), .Y(
        n31548) );
  NAND2xp5_ASAP7_75t_SL U26936 ( .A(n24684), .B(n18851), .Y(n30190) );
  INVxp33_ASAP7_75t_SL U26937 ( .A(mult_x_1196_n481), .Y(mult_x_1196_n792) );
  OA21x2_ASAP7_75t_SL U26938 ( .A1(n22405), .A2(n31778), .B(n32550), .Y(n31779) );
  OA21x2_ASAP7_75t_SL U26939 ( .A1(n22405), .A2(n31761), .B(n32539), .Y(n31762) );
  OAI21xp33_ASAP7_75t_SL U26940 ( .A1(n22427), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N12), .B(n27126), .Y(n4291) );
  OA21x2_ASAP7_75t_SL U26941 ( .A1(n22405), .A2(n31782), .B(n32547), .Y(n31783) );
  AND2x2_ASAP7_75t_SL U26942 ( .A(n22421), .B(n22366), .Y(n23328) );
  OA21x2_ASAP7_75t_SL U26943 ( .A1(n22405), .A2(n31997), .B(n32556), .Y(n31998) );
  OA21x2_ASAP7_75t_SL U26944 ( .A1(n22405), .A2(n32535), .B(n32533), .Y(n32534) );
  OA21x2_ASAP7_75t_SL U26945 ( .A1(n22405), .A2(n31768), .B(n32533), .Y(n31769) );
  OA21x2_ASAP7_75t_SL U26946 ( .A1(n22405), .A2(n32541), .B(n32539), .Y(n32540) );
  NAND2xp5_ASAP7_75t_SL U26947 ( .A(u0_0_leon3x0_p0_ici[78]), .B(n22405), .Y(
        n32533) );
  NAND2xp5_ASAP7_75t_SL U26948 ( .A(u0_0_leon3x0_p0_ici[88]), .B(n22405), .Y(
        n32556) );
  NAND2xp5_ASAP7_75t_SL U26949 ( .A(u0_0_leon3x0_p0_ici[83]), .B(n22405), .Y(
        n32547) );
  NAND2xp5_ASAP7_75t_SL U26950 ( .A(u0_0_leon3x0_p0_ici[62]), .B(n22405), .Y(
        n32683) );
  NAND2xp5_ASAP7_75t_SL U26951 ( .A(u0_0_leon3x0_p0_ici[61]), .B(n22405), .Y(
        n32675) );
  NAND2xp5_ASAP7_75t_SL U26952 ( .A(u0_0_leon3x0_p0_ici[84]), .B(n22405), .Y(
        n32550) );
  NAND2xp5_ASAP7_75t_SL U26953 ( .A(u0_0_leon3x0_p0_ici[81]), .B(n22405), .Y(
        n32539) );
  NAND2xp33_ASAP7_75t_SL U26954 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[1]), .B(
        n31429), .Y(n26784) );
  INVxp67_ASAP7_75t_SL U26955 ( .A(mult_x_1196_n683), .Y(mult_x_1196_n819) );
  OAI21xp33_ASAP7_75t_SL U26956 ( .A1(n22379), .A2(
        u0_0_leon3x0_p0_iu_r_D__ANNUL_), .B(n31816), .Y(n4173) );
  OAI21xp33_ASAP7_75t_SL U26957 ( .A1(n22379), .A2(
        u0_0_leon3x0_p0_iu_r_A__CTRL__ANNUL_), .B(n32104), .Y(n3739) );
  INVx1_ASAP7_75t_SL U26958 ( .A(n23600), .Y(n23231) );
  OAI21xp33_ASAP7_75t_SL U26959 ( .A1(n29844), .A2(n29843), .B(n29842), .Y(
        n4461) );
  OAI21xp33_ASAP7_75t_SL U26960 ( .A1(n32110), .A2(n29905), .B(n26326), .Y(
        n4380) );
  OA21x2_ASAP7_75t_SL U26961 ( .A1(n22379), .A2(n32661), .B(n26452), .Y(n26453) );
  AOI21xp5_ASAP7_75t_SL U26962 ( .A1(n26955), .A2(n31342), .B(n26954), .Y(
        n29802) );
  INVx1_ASAP7_75t_SL U26963 ( .A(n24252), .Y(n22407) );
  OAI21xp33_ASAP7_75t_SL U26964 ( .A1(n22427), .A2(n29800), .B(n25510), .Y(
        n4121) );
  OAI21xp33_ASAP7_75t_SL U26965 ( .A1(n22427), .A2(n30597), .B(n30596), .Y(
        n4113) );
  AOI21xp33_ASAP7_75t_SL U26966 ( .A1(n28578), .A2(n22432), .B(n28577), .Y(
        n28581) );
  OAI21xp33_ASAP7_75t_SL U26967 ( .A1(n22427), .A2(n28578), .B(n26584), .Y(
        n3984) );
  AOI21xp33_ASAP7_75t_SL U26968 ( .A1(n29767), .A2(n22432), .B(n28466), .Y(
        n28469) );
  AOI21xp5_ASAP7_75t_SL U26969 ( .A1(n29078), .A2(n22432), .B(n28512), .Y(
        n28516) );
  AOI21xp33_ASAP7_75t_SL U26970 ( .A1(n31875), .A2(n22432), .B(n28557), .Y(
        n28560) );
  AOI21xp33_ASAP7_75t_SL U26971 ( .A1(n28608), .A2(n22432), .B(n28607), .Y(
        n28611) );
  AOI21xp33_ASAP7_75t_SL U26972 ( .A1(n30820), .A2(n22432), .B(n28531), .Y(
        n28534) );
  INVxp67_ASAP7_75t_SL U26973 ( .A(DP_OP_5187J1_124_3275_n4), .Y(
        DP_OP_5187J1_124_3275_n123) );
  INVx1_ASAP7_75t_SL U26974 ( .A(DP_OP_5187J1_124_3275_n3), .Y(
        DP_OP_5187J1_124_3275_n124) );
  AOI21xp33_ASAP7_75t_SL U26975 ( .A1(n30799), .A2(n22432), .B(n28798), .Y(
        n28803) );
  AOI21xp5_ASAP7_75t_SL U26976 ( .A1(n27032), .A2(n22432), .B(n27012), .Y(
        n27016) );
  AOI21xp33_ASAP7_75t_SL U26977 ( .A1(n30736), .A2(n22432), .B(n28753), .Y(
        n28757) );
  AOI21xp33_ASAP7_75t_SL U26978 ( .A1(n27174), .A2(n22432), .B(n27132), .Y(
        n27135) );
  INVxp67_ASAP7_75t_SL U26979 ( .A(mult_x_1196_n870), .Y(mult_x_1196_n866) );
  INVxp67_ASAP7_75t_SL U26980 ( .A(mult_x_1196_n891), .Y(mult_x_1196_n887) );
  OAI21xp33_ASAP7_75t_SL U26981 ( .A1(apbi[38]), .A2(n22408), .B(n30525), .Y(
        n2662) );
  OAI21xp33_ASAP7_75t_SL U26982 ( .A1(n2931), .A2(n22408), .B(n25329), .Y(
        n17885) );
  OAI21xp33_ASAP7_75t_SL U26983 ( .A1(n2929), .A2(n22408), .B(n25337), .Y(
        n17886) );
  INVxp33_ASAP7_75t_SL U26984 ( .A(u0_0_leon3x0_p0_dci[31]), .Y(n28386) );
  OAI21xp33_ASAP7_75t_SL U26985 ( .A1(apbi[42]), .A2(n22408), .B(n30539), .Y(
        n2614) );
  OAI21xp33_ASAP7_75t_SL U26986 ( .A1(n4371), .A2(n22408), .B(n25264), .Y(
        n17889) );
  OAI21xp33_ASAP7_75t_SL U26987 ( .A1(n30659), .A2(u0_0_leon3x0_p0_dci[36]), 
        .B(n30656), .Y(n27021) );
  OAI21xp33_ASAP7_75t_SL U26988 ( .A1(apbi[39]), .A2(n22408), .B(n30532), .Y(
        n2638) );
  OAI21xp33_ASAP7_75t_SL U26989 ( .A1(apbi[41]), .A2(n22408), .B(n30523), .Y(
        n2947) );
  OAI21xp33_ASAP7_75t_SL U26990 ( .A1(apbi[40]), .A2(n22408), .B(n30516), .Y(
        n2950) );
  AOI21xp33_ASAP7_75t_SL U26991 ( .A1(n31947), .A2(n22432), .B(n28814), .Y(
        n28818) );
  OAI21xp33_ASAP7_75t_SL U26992 ( .A1(apbi[43]), .A2(n22408), .B(n30546), .Y(
        n2590) );
  OAI21xp33_ASAP7_75t_SL U26993 ( .A1(n22408), .A2(n2992), .B(n25262), .Y(
        n17890) );
  INVxp33_ASAP7_75t_SL U26994 ( .A(u0_0_leon3x0_p0_dci[25]), .Y(n26972) );
  OAI21xp33_ASAP7_75t_SL U26995 ( .A1(apbi[33]), .A2(n22408), .B(n25266), .Y(
        n2994) );
  OAI21xp33_ASAP7_75t_SL U26996 ( .A1(apbi[34]), .A2(n22408), .B(n25268), .Y(
        n4433) );
  OAI21xp33_ASAP7_75t_SL U26997 ( .A1(apbi[37]), .A2(n22408), .B(n25271), .Y(
        n2989) );
  NAND2xp33_ASAP7_75t_SL U26998 ( .A(n32996), .B(n22408), .Y(n25268) );
  NAND2xp33_ASAP7_75t_SL U26999 ( .A(n33002), .B(n22408), .Y(n25271) );
  XNOR2xp5_ASAP7_75t_SL U27000 ( .A(add_x_735_n15), .B(add_x_735_n143), .Y(
        u0_0_leon3x0_p0_dci[25]) );
  XNOR2xp5_ASAP7_75t_SL U27001 ( .A(add_x_735_n9), .B(add_x_735_n87), .Y(
        u0_0_leon3x0_p0_dci[31]) );
  NAND2xp33_ASAP7_75t_SL U27002 ( .A(n32992), .B(n22408), .Y(n25266) );
  INVxp67_ASAP7_75t_SL U27003 ( .A(mult_x_1196_n1025), .Y(n24144) );
  XNOR2xp5_ASAP7_75t_SL U27004 ( .A(add_x_735_n6), .B(add_x_735_n58), .Y(
        u0_0_leon3x0_p0_dci[34]) );
  NAND2xp33_ASAP7_75t_SL U27005 ( .A(n30545), .B(n22408), .Y(n30546) );
  NAND2xp33_ASAP7_75t_SL U27006 ( .A(n32995), .B(n22408), .Y(n25262) );
  NAND2xp5_ASAP7_75t_SL U27007 ( .A(n31695), .B(n22408), .Y(n31837) );
  NAND2xp33_ASAP7_75t_SL U27008 ( .A(n30522), .B(n22408), .Y(n30523) );
  INVxp67_ASAP7_75t_SL U27009 ( .A(DP_OP_5187J1_124_3275_n71), .Y(
        DP_OP_5187J1_124_3275_n69) );
  NAND2xp33_ASAP7_75t_SL U27010 ( .A(n30531), .B(n22408), .Y(n30532) );
  NAND2xp33_ASAP7_75t_SL U27011 ( .A(n32994), .B(n22408), .Y(n25264) );
  NAND2xp33_ASAP7_75t_SL U27012 ( .A(n30538), .B(n22408), .Y(n30539) );
  NAND2xp33_ASAP7_75t_SL U27013 ( .A(n31321), .B(n22408), .Y(n25326) );
  NAND2xp33_ASAP7_75t_SL U27014 ( .A(n32985), .B(n22408), .Y(n25337) );
  NAND2xp33_ASAP7_75t_SL U27015 ( .A(n32984), .B(n22408), .Y(n25329) );
  NAND2xp33_ASAP7_75t_SL U27016 ( .A(n33004), .B(n22408), .Y(n30525) );
  INVxp67_ASAP7_75t_SL U27017 ( .A(u0_0_leon3x0_p0_dci[16]), .Y(n25344) );
  NAND2xp33_ASAP7_75t_SL U27018 ( .A(n30515), .B(n22408), .Y(n30516) );
  INVxp67_ASAP7_75t_SL U27019 ( .A(mult_x_1196_n302), .Y(n23390) );
  INVxp67_ASAP7_75t_SL U27020 ( .A(DP_OP_5187J1_124_3275_n80), .Y(
        DP_OP_5187J1_124_3275_n311) );
  INVxp67_ASAP7_75t_SL U27021 ( .A(DP_OP_5187J1_124_3275_n131), .Y(
        DP_OP_5187J1_124_3275_n316) );
  INVxp67_ASAP7_75t_SL U27022 ( .A(DP_OP_5187J1_124_3275_n138), .Y(
        DP_OP_5187J1_124_3275_n317) );
  INVxp67_ASAP7_75t_SL U27023 ( .A(DP_OP_5187J1_124_3275_n177), .Y(
        DP_OP_5187J1_124_3275_n175) );
  INVxp67_ASAP7_75t_SL U27024 ( .A(DP_OP_5187J1_124_3275_n176), .Y(
        DP_OP_5187J1_124_3275_n321) );
  INVxp67_ASAP7_75t_SL U27025 ( .A(DP_OP_5187J1_124_3275_n113), .Y(
        DP_OP_5187J1_124_3275_n314) );
  INVxp67_ASAP7_75t_SL U27026 ( .A(DP_OP_5187J1_124_3275_n158), .Y(
        DP_OP_5187J1_124_3275_n319) );
  INVxp67_ASAP7_75t_SL U27027 ( .A(DP_OP_5187J1_124_3275_n151), .Y(
        DP_OP_5187J1_124_3275_n318) );
  INVx1_ASAP7_75t_SL U27028 ( .A(DP_OP_5187J1_124_3275_n62), .Y(
        DP_OP_5187J1_124_3275_n60) );
  INVxp67_ASAP7_75t_SL U27029 ( .A(n30014), .Y(n30013) );
  AOI22xp33_ASAP7_75t_SL U27030 ( .A1(n29603), .A2(n26914), .B1(n28742), .B2(
        n25475), .Y(n25506) );
  INVxp67_ASAP7_75t_SL U27031 ( .A(DP_OP_5187J1_124_3275_n100), .Y(
        DP_OP_5187J1_124_3275_n313) );
  INVxp67_ASAP7_75t_SL U27032 ( .A(n28799), .Y(n28809) );
  INVxp67_ASAP7_75t_SL U27033 ( .A(mult_x_1196_n872), .Y(n22530) );
  NAND2xp5_ASAP7_75t_SL U27034 ( .A(n24347), .B(n24399), .Y(n24349) );
  NAND2xp5_ASAP7_75t_SL U27035 ( .A(n25438), .B(n25053), .Y(n25072) );
  INVxp67_ASAP7_75t_SL U27036 ( .A(n28443), .Y(n25475) );
  O2A1O1Ixp33_ASAP7_75t_SL U27037 ( .A1(n28176), .A2(n28179), .B(n28175), .C(
        n22419), .Y(n28177) );
  XNOR2xp5_ASAP7_75t_SL U27038 ( .A(mult_x_1196_n1248), .B(n23738), .Y(
        mult_x_1196_n1202) );
  OAI22xp33_ASAP7_75t_SL U27039 ( .A1(n31730), .A2(n31731), .B1(read), .B2(
        n32875), .Y(n31707) );
  NAND2xp33_ASAP7_75t_SL U27040 ( .A(n24681), .B(n24890), .Y(n24891) );
  INVxp67_ASAP7_75t_SL U27041 ( .A(n28615), .Y(n26151) );
  NOR2xp33_ASAP7_75t_SL U27042 ( .A(n27017), .B(n26751), .Y(n30648) );
  INVxp33_ASAP7_75t_SL U27043 ( .A(add_x_746_n103), .Y(add_x_746_n104) );
  OAI21xp33_ASAP7_75t_SL U27044 ( .A1(n28977), .A2(n25912), .B(n25911), .Y(
        n29604) );
  AOI22xp33_ASAP7_75t_SL U27045 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__12_), 
        .A2(n31364), .B1(n31477), .B2(n31043), .Y(n25446) );
  AOI22xp33_ASAP7_75t_SL U27046 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__8_), 
        .A2(n31364), .B1(n30479), .B2(n31043), .Y(n29763) );
  OAI22xp33_ASAP7_75t_SL U27047 ( .A1(n29641), .A2(n30706), .B1(n23229), .B2(
        n29640), .Y(n29644) );
  XNOR2xp5_ASAP7_75t_SL U27048 ( .A(n22852), .B(mult_x_1196_n2519), .Y(n23533)
         );
  INVxp33_ASAP7_75t_SL U27049 ( .A(n29918), .Y(n25441) );
  OAI21xp33_ASAP7_75t_SL U27050 ( .A1(n31001), .A2(n25621), .B(n25620), .Y(
        n30573) );
  AOI22xp33_ASAP7_75t_SL U27051 ( .A1(n26893), .A2(n26892), .B1(n24572), .B2(
        n26902), .Y(n30241) );
  INVxp67_ASAP7_75t_SL U27052 ( .A(mult_x_1196_n2466), .Y(n23722) );
  NOR2x1_ASAP7_75t_SL U27053 ( .A(n23635), .B(n24202), .Y(n24203) );
  NAND2xp33_ASAP7_75t_SL U27054 ( .A(n28894), .B(n30261), .Y(n26404) );
  INVxp67_ASAP7_75t_SL U27055 ( .A(n33020), .Y(n30545) );
  OAI21xp33_ASAP7_75t_SL U27056 ( .A1(n22379), .A2(
        u0_0_leon3x0_p0_iu_r_E__MULSTEP_), .B(n31343), .Y(n3574) );
  INVx1_ASAP7_75t_SL U27057 ( .A(u0_0_leon3x0_p0_iu_fe_pc_21_), .Y(
        add_x_746_n63) );
  INVxp67_ASAP7_75t_SL U27058 ( .A(n33014), .Y(n30522) );
  INVx1_ASAP7_75t_SL U27059 ( .A(u0_0_leon3x0_p0_iu_fe_pc_29_), .Y(
        add_x_746_n15) );
  INVx1_ASAP7_75t_SL U27060 ( .A(n30276), .Y(n29167) );
  INVxp67_ASAP7_75t_SL U27061 ( .A(n33008), .Y(n30531) );
  NAND2xp33_ASAP7_75t_SL U27062 ( .A(n31001), .B(n25619), .Y(n25620) );
  NOR2x1_ASAP7_75t_SL U27063 ( .A(n28167), .B(n28141), .Y(n28174) );
  INVx1_ASAP7_75t_SL U27064 ( .A(n31343), .Y(n31542) );
  AOI21xp5_ASAP7_75t_SL U27065 ( .A1(n30266), .A2(n30671), .B(n29813), .Y(
        n29814) );
  INVxp67_ASAP7_75t_SL U27066 ( .A(mult_x_1196_n2506), .Y(n23653) );
  NOR3xp33_ASAP7_75t_SL U27067 ( .A(n29143), .B(n30326), .C(n30380), .Y(n29153) );
  INVxp67_ASAP7_75t_SL U27068 ( .A(u0_0_leon3x0_p0_iu_fe_pc_10_), .Y(
        add_x_746_n123) );
  INVx1_ASAP7_75t_SL U27069 ( .A(u0_0_leon3x0_p0_iu_fe_pc_6_), .Y(
        add_x_746_n143) );
  INVxp67_ASAP7_75t_SL U27070 ( .A(u0_0_leon3x0_p0_iu_fe_pc_7_), .Y(
        add_x_746_n139) );
  INVxp33_ASAP7_75t_SL U27071 ( .A(n25439), .Y(n25445) );
  AOI21xp5_ASAP7_75t_SL U27072 ( .A1(add_x_735_n118), .A2(add_x_735_n90), .B(
        add_x_735_n91), .Y(add_x_735_n89) );
  INVx1_ASAP7_75t_SL U27073 ( .A(u0_0_leon3x0_p0_iu_fe_pc_12_), .Y(
        add_x_746_n113) );
  INVx1_ASAP7_75t_SL U27074 ( .A(n33052), .Y(n31798) );
  AOI21xp33_ASAP7_75t_SL U27075 ( .A1(n31157), .A2(uart1_r_RHOLD__7__1_), .B(
        n26119), .Y(n2449) );
  AOI21xp33_ASAP7_75t_SL U27076 ( .A1(n31061), .A2(uart1_r_RHOLD__0__0_), .B(
        n25982), .Y(n2448) );
  AOI21xp33_ASAP7_75t_SL U27077 ( .A1(n31187), .A2(uart1_r_RHOLD__16__7_), .B(
        n30867), .Y(n2059) );
  AOI21xp33_ASAP7_75t_SL U27078 ( .A1(n31077), .A2(uart1_r_RHOLD__31__0_), .B(
        n26008), .Y(n2447) );
  AOI21xp33_ASAP7_75t_SL U27079 ( .A1(n31157), .A2(uart1_r_RHOLD__7__0_), .B(
        n26040), .Y(n2450) );
  OAI21xp33_ASAP7_75t_SL U27080 ( .A1(n32761), .A2(n33040), .B(
        sr1_r_MCFG2__RAMBANKSZ__1_), .Y(n32759) );
  AOI22xp33_ASAP7_75t_SL U27081 ( .A1(n24576), .A2(n27097), .B1(n28847), .B2(
        n27100), .Y(n25762) );
  AOI21xp33_ASAP7_75t_SL U27082 ( .A1(n31077), .A2(uart1_r_RHOLD__31__3_), .B(
        n28197), .Y(n2198) );
  AOI21xp33_ASAP7_75t_SL U27083 ( .A1(n31169), .A2(uart1_r_RHOLD__5__2_), .B(
        n29551), .Y(n2203) );
  AOI21xp33_ASAP7_75t_SL U27084 ( .A1(n31153), .A2(uart1_r_RHOLD__4__2_), .B(
        n29547), .Y(n2202) );
  AOI21xp33_ASAP7_75t_SL U27085 ( .A1(n31141), .A2(uart1_r_RHOLD__20__7_), .B(
        n30854), .Y(n2063) );
  AOI21xp33_ASAP7_75t_SL U27086 ( .A1(n31173), .A2(uart1_r_RHOLD__2__2_), .B(
        n29552), .Y(n2200) );
  OAI21xp33_ASAP7_75t_SRAM U27087 ( .A1(n31001), .A2(n29760), .B(n29759), .Y(
        n29762) );
  OAI21xp5_ASAP7_75t_SL U27088 ( .A1(n30426), .A2(n28964), .B(n26749), .Y(
        n28365) );
  AOI21xp33_ASAP7_75t_SL U27089 ( .A1(n31161), .A2(uart1_r_RHOLD__30__3_), .B(
        n28218), .Y(n2197) );
  AOI21xp33_ASAP7_75t_SL U27090 ( .A1(n31069), .A2(uart1_r_RHOLD__27__3_), .B(
        n28195), .Y(n2194) );
  AOI21xp33_ASAP7_75t_SL U27091 ( .A1(n31137), .A2(uart1_r_RHOLD__25__3_), .B(
        n28212), .Y(n2192) );
  AOI21xp33_ASAP7_75t_SL U27092 ( .A1(n31141), .A2(uart1_r_RHOLD__20__3_), .B(
        n28213), .Y(n2187) );
  AOI21xp33_ASAP7_75t_SL U27093 ( .A1(n31145), .A2(uart1_r_RHOLD__19__3_), .B(
        n28214), .Y(n2186) );
  AOI21xp33_ASAP7_75t_SL U27094 ( .A1(n31165), .A2(uart1_r_RHOLD__17__3_), .B(
        n28219), .Y(n2184) );
  AOI21xp33_ASAP7_75t_SL U27095 ( .A1(n31187), .A2(uart1_r_RHOLD__16__3_), .B(
        n28226), .Y(n2183) );
  AOI21xp33_ASAP7_75t_SL U27096 ( .A1(n31149), .A2(uart1_r_RHOLD__10__3_), .B(
        n28215), .Y(n2177) );
  AOI21xp33_ASAP7_75t_SL U27097 ( .A1(n31181), .A2(uart1_r_RHOLD__9__3_), .B(
        n28223), .Y(n2176) );
  AOI21xp33_ASAP7_75t_SL U27098 ( .A1(n31177), .A2(uart1_r_RHOLD__8__3_), .B(
        n28222), .Y(n2175) );
  AOI21xp33_ASAP7_75t_SL U27099 ( .A1(n31157), .A2(uart1_r_RHOLD__7__3_), .B(
        n28217), .Y(n2174) );
  AOI21xp33_ASAP7_75t_SL U27100 ( .A1(n31165), .A2(uart1_r_RHOLD__17__7_), .B(
        n30860), .Y(n2060) );
  AOI21xp33_ASAP7_75t_SL U27101 ( .A1(n31077), .A2(uart1_r_RHOLD__31__2_), .B(
        n29528), .Y(n2229) );
  AOI21xp33_ASAP7_75t_SL U27102 ( .A1(n31161), .A2(uart1_r_RHOLD__30__2_), .B(
        n29549), .Y(n2228) );
  INVxp67_ASAP7_75t_SL U27103 ( .A(add_x_735_n74), .Y(add_x_735_n72) );
  AOI21xp33_ASAP7_75t_SL U27104 ( .A1(n31069), .A2(uart1_r_RHOLD__27__2_), .B(
        n29526), .Y(n2225) );
  AOI21xp33_ASAP7_75t_SL U27105 ( .A1(n31137), .A2(uart1_r_RHOLD__25__2_), .B(
        n29543), .Y(n2223) );
  AOI21xp33_ASAP7_75t_SL U27106 ( .A1(n31141), .A2(uart1_r_RHOLD__20__2_), .B(
        n29544), .Y(n2218) );
  AOI21xp33_ASAP7_75t_SL U27107 ( .A1(n31145), .A2(uart1_r_RHOLD__19__2_), .B(
        n29545), .Y(n2217) );
  AOI21xp33_ASAP7_75t_SL U27108 ( .A1(n31165), .A2(uart1_r_RHOLD__17__2_), .B(
        n29550), .Y(n2215) );
  AOI21xp33_ASAP7_75t_SL U27109 ( .A1(n31187), .A2(uart1_r_RHOLD__16__2_), .B(
        n29557), .Y(n2214) );
  AOI21xp33_ASAP7_75t_SL U27110 ( .A1(n31149), .A2(uart1_r_RHOLD__10__2_), .B(
        n29546), .Y(n2208) );
  OAI21xp33_ASAP7_75t_SL U27111 ( .A1(add_x_735_n75), .A2(add_x_735_n67), .B(
        add_x_735_n68), .Y(add_x_735_n62) );
  AOI21xp33_ASAP7_75t_SL U27112 ( .A1(n31181), .A2(uart1_r_RHOLD__9__2_), .B(
        n29554), .Y(n2207) );
  AOI21xp33_ASAP7_75t_SL U27113 ( .A1(n31177), .A2(uart1_r_RHOLD__8__2_), .B(
        n29553), .Y(n2206) );
  AOI21xp33_ASAP7_75t_SL U27114 ( .A1(n31145), .A2(uart1_r_RHOLD__19__7_), .B(
        n30855), .Y(n2062) );
  AOI21xp33_ASAP7_75t_SL U27115 ( .A1(n31157), .A2(uart1_r_RHOLD__7__2_), .B(
        n29548), .Y(n2205) );
  AOI21xp33_ASAP7_75t_SL U27116 ( .A1(n31061), .A2(uart1_r_RHOLD__0__6_), .B(
        n31060), .Y(n1736) );
  AOI21xp33_ASAP7_75t_SL U27117 ( .A1(n31061), .A2(uart1_r_RHOLD__0__5_), .B(
        n30031), .Y(n1737) );
  AOI21xp33_ASAP7_75t_SL U27118 ( .A1(n31061), .A2(uart1_r_RHOLD__0__4_), .B(
        n30740), .Y(n1738) );
  AOI21xp33_ASAP7_75t_SL U27119 ( .A1(n31173), .A2(uart1_r_RHOLD__2__0_), .B(
        n26056), .Y(n2393) );
  AOI21xp33_ASAP7_75t_SL U27120 ( .A1(n31173), .A2(uart1_r_RHOLD__2__1_), .B(
        n26123), .Y(n2392) );
  AOI21xp33_ASAP7_75t_SL U27121 ( .A1(n31141), .A2(uart1_r_RHOLD__20__0_), .B(
        n26030), .Y(n2425) );
  AOI21xp33_ASAP7_75t_SL U27122 ( .A1(n31187), .A2(uart1_r_RHOLD__16__0_), .B(
        n26070), .Y(n2417) );
  AOI21xp33_ASAP7_75t_SL U27123 ( .A1(n31187), .A2(uart1_r_RHOLD__16__1_), .B(
        n26128), .Y(n2416) );
  AOI21xp33_ASAP7_75t_SL U27124 ( .A1(n31165), .A2(uart1_r_RHOLD__17__1_), .B(
        n26121), .Y(n2418) );
  AOI21xp33_ASAP7_75t_SL U27125 ( .A1(n31165), .A2(uart1_r_RHOLD__17__0_), .B(
        n26047), .Y(n2419) );
  AOI21xp33_ASAP7_75t_SL U27126 ( .A1(n29598), .A2(n29778), .B(n28729), .Y(
        n26402) );
  AOI21xp33_ASAP7_75t_SL U27127 ( .A1(n31149), .A2(uart1_r_RHOLD__10__0_), .B(
        n26034), .Y(n2407) );
  AOI21xp33_ASAP7_75t_SL U27128 ( .A1(n31149), .A2(uart1_r_RHOLD__10__1_), .B(
        n26117), .Y(n2406) );
  AOI21xp33_ASAP7_75t_SL U27129 ( .A1(n31181), .A2(uart1_r_RHOLD__9__0_), .B(
        n26063), .Y(n2405) );
  AOI21xp33_ASAP7_75t_SL U27130 ( .A1(n31181), .A2(uart1_r_RHOLD__9__1_), .B(
        n26125), .Y(n2404) );
  AOI21xp33_ASAP7_75t_SL U27131 ( .A1(n31177), .A2(uart1_r_RHOLD__8__0_), .B(
        n26057), .Y(n2403) );
  AOI21xp33_ASAP7_75t_SL U27132 ( .A1(n31177), .A2(uart1_r_RHOLD__8__1_), .B(
        n26124), .Y(n2402) );
  AOI21xp33_ASAP7_75t_SL U27133 ( .A1(n31169), .A2(uart1_r_RHOLD__5__0_), .B(
        n26050), .Y(n2399) );
  AOI21xp33_ASAP7_75t_SL U27134 ( .A1(n31169), .A2(uart1_r_RHOLD__5__1_), .B(
        n26122), .Y(n2398) );
  AOI21xp33_ASAP7_75t_SL U27135 ( .A1(n31061), .A2(uart1_r_RHOLD__0__7_), .B(
        n30834), .Y(n1735) );
  AOI21xp33_ASAP7_75t_SL U27136 ( .A1(n31145), .A2(uart1_r_RHOLD__19__1_), .B(
        n26116), .Y(n2422) );
  AOI21xp33_ASAP7_75t_SL U27137 ( .A1(n31153), .A2(uart1_r_RHOLD__4__0_), .B(
        n26037), .Y(n2397) );
  AOI21xp33_ASAP7_75t_SL U27138 ( .A1(n31145), .A2(uart1_r_RHOLD__19__0_), .B(
        n26033), .Y(n2423) );
  AOI21xp33_ASAP7_75t_SL U27139 ( .A1(n31141), .A2(uart1_r_RHOLD__20__1_), .B(
        n26115), .Y(n2424) );
  AOI21xp33_ASAP7_75t_SL U27140 ( .A1(n31153), .A2(uart1_r_RHOLD__4__1_), .B(
        n26118), .Y(n2396) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U27141 ( .A1(n25901), .A2(n27155), .B(n25499), 
        .C(n24634), .Y(n25500) );
  AOI21xp33_ASAP7_75t_SL U27142 ( .A1(n31157), .A2(uart1_r_RHOLD__7__7_), .B(
        n30858), .Y(n2050) );
  AOI21xp33_ASAP7_75t_SL U27143 ( .A1(n25133), .A2(n28830), .B(n25132), .Y(
        n25134) );
  AOI21xp33_ASAP7_75t_SL U27144 ( .A1(n31177), .A2(uart1_r_RHOLD__8__7_), .B(
        n30863), .Y(n2051) );
  AOI21xp33_ASAP7_75t_SL U27145 ( .A1(n31181), .A2(uart1_r_RHOLD__9__7_), .B(
        n30864), .Y(n2052) );
  INVx2_ASAP7_75t_SL U27146 ( .A(n23810), .Y(n22411) );
  AOI21xp33_ASAP7_75t_SL U27147 ( .A1(n31149), .A2(uart1_r_RHOLD__10__7_), .B(
        n30856), .Y(n2053) );
  AOI21xp33_ASAP7_75t_SL U27148 ( .A1(u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__0_), 
        .A2(n30017), .B(n25049), .Y(n29915) );
  INVxp67_ASAP7_75t_SL U27149 ( .A(n26423), .Y(n25468) );
  AOI21xp33_ASAP7_75t_SL U27150 ( .A1(n31161), .A2(uart1_r_RHOLD__30__1_), .B(
        n26120), .Y(n2444) );
  NAND2xp33_ASAP7_75t_SL U27151 ( .A(n24576), .B(n26424), .Y(n25471) );
  AOI21xp33_ASAP7_75t_SL U27152 ( .A1(n31161), .A2(uart1_r_RHOLD__30__0_), .B(
        n26046), .Y(n2445) );
  AOI21xp33_ASAP7_75t_SL U27153 ( .A1(n31077), .A2(uart1_r_RHOLD__31__1_), .B(
        n26101), .Y(n2446) );
  AOI21xp33_ASAP7_75t_SL U27154 ( .A1(n31137), .A2(uart1_r_RHOLD__25__1_), .B(
        n26114), .Y(n2434) );
  AOI21xp33_ASAP7_75t_SL U27155 ( .A1(n31137), .A2(uart1_r_RHOLD__25__0_), .B(
        n26029), .Y(n2435) );
  OAI21xp33_ASAP7_75t_SL U27156 ( .A1(n31778), .A2(n22415), .B(n25255), .Y(
        n33049) );
  HB1xp67_ASAP7_75t_SL U27157 ( .A(mult_x_1196_n2485), .Y(n23922) );
  AOI21xp33_ASAP7_75t_SL U27158 ( .A1(n31069), .A2(uart1_r_RHOLD__27__1_), .B(
        n26099), .Y(n2438) );
  AOI21xp33_ASAP7_75t_SL U27159 ( .A1(n31173), .A2(uart1_r_RHOLD__2__7_), .B(
        n30862), .Y(n2045) );
  AOI21xp33_ASAP7_75t_SL U27160 ( .A1(n31069), .A2(uart1_r_RHOLD__27__0_), .B(
        n26002), .Y(n2439) );
  AOI21xp33_ASAP7_75t_SL U27161 ( .A1(n31153), .A2(uart1_r_RHOLD__4__7_), .B(
        n30857), .Y(n2047) );
  AOI21xp33_ASAP7_75t_SL U27162 ( .A1(n31169), .A2(uart1_r_RHOLD__5__7_), .B(
        n30861), .Y(n2048) );
  INVxp67_ASAP7_75t_SL U27163 ( .A(n28544), .Y(n28545) );
  OAI21xp33_ASAP7_75t_SL U27164 ( .A1(n22379), .A2(
        u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .B(n24951), .Y(n3560) );
  AOI21xp33_ASAP7_75t_SL U27165 ( .A1(n31149), .A2(uart1_r_RHOLD__10__6_), .B(
        n31148), .Y(n2084) );
  NAND2xp5_ASAP7_75t_SL U27166 ( .A(n29990), .B(n29989), .Y(n29992) );
  AOI21xp33_ASAP7_75t_SL U27167 ( .A1(n31181), .A2(uart1_r_RHOLD__9__6_), .B(
        n31180), .Y(n2083) );
  AOI21xp33_ASAP7_75t_SL U27168 ( .A1(n31145), .A2(uart1_r_RHOLD__19__6_), .B(
        n31144), .Y(n2093) );
  AOI21xp33_ASAP7_75t_SL U27169 ( .A1(n31187), .A2(uart1_r_RHOLD__16__4_), .B(
        n30773), .Y(n2152) );
  AOI21xp33_ASAP7_75t_SL U27170 ( .A1(n31165), .A2(uart1_r_RHOLD__17__4_), .B(
        n30766), .Y(n2153) );
  AOI21xp33_ASAP7_75t_SL U27171 ( .A1(n31177), .A2(uart1_r_RHOLD__8__6_), .B(
        n31176), .Y(n2082) );
  AOI21xp33_ASAP7_75t_SL U27172 ( .A1(n31141), .A2(uart1_r_RHOLD__20__6_), .B(
        n31140), .Y(n2094) );
  AOI21xp33_ASAP7_75t_SL U27173 ( .A1(n31165), .A2(uart1_r_RHOLD__17__5_), .B(
        n30057), .Y(n2122) );
  AOI21xp33_ASAP7_75t_SL U27174 ( .A1(n31145), .A2(uart1_r_RHOLD__19__4_), .B(
        n30761), .Y(n2155) );
  AOI21xp33_ASAP7_75t_SL U27175 ( .A1(n31141), .A2(uart1_r_RHOLD__20__4_), .B(
        n30760), .Y(n2156) );
  NAND2xp33_ASAP7_75t_SRAM U27176 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__5_), 
        .B(n32184), .Y(n30933) );
  AOI21xp33_ASAP7_75t_SL U27177 ( .A1(n31077), .A2(uart1_r_RHOLD__31__5_), .B(
        n30035), .Y(n2136) );
  AOI21xp33_ASAP7_75t_SL U27178 ( .A1(n31157), .A2(uart1_r_RHOLD__7__6_), .B(
        n31156), .Y(n2081) );
  OAI21xp33_ASAP7_75t_SL U27179 ( .A1(n22379), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__CWP__0_), .B(n31431), .Y(n2806) );
  INVxp33_ASAP7_75t_SL U27180 ( .A(n24869), .Y(n24738) );
  AOI21xp33_ASAP7_75t_SL U27181 ( .A1(n31069), .A2(uart1_r_RHOLD__27__6_), .B(
        n31068), .Y(n2101) );
  AOI21xp33_ASAP7_75t_SL U27182 ( .A1(n31169), .A2(uart1_r_RHOLD__5__6_), .B(
        n31168), .Y(n2079) );
  AOI21xp33_ASAP7_75t_SL U27183 ( .A1(n31149), .A2(uart1_r_RHOLD__10__5_), .B(
        n30053), .Y(n2115) );
  AOI21xp33_ASAP7_75t_SL U27184 ( .A1(n31153), .A2(uart1_r_RHOLD__4__6_), .B(
        n31152), .Y(n2078) );
  AOI21xp33_ASAP7_75t_SL U27185 ( .A1(n31153), .A2(uart1_r_RHOLD__4__4_), .B(
        n30763), .Y(n2140) );
  AOI21xp33_ASAP7_75t_SL U27186 ( .A1(n31165), .A2(uart1_r_RHOLD__17__6_), .B(
        n31164), .Y(n2091) );
  AOI21xp33_ASAP7_75t_SL U27187 ( .A1(n31173), .A2(uart1_r_RHOLD__2__4_), .B(
        n30768), .Y(n2138) );
  AOI21xp33_ASAP7_75t_SL U27188 ( .A1(n31169), .A2(uart1_r_RHOLD__5__4_), .B(
        n30767), .Y(n2141) );
  OAI21xp33_ASAP7_75t_SL U27189 ( .A1(n22379), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__29_), .B(n30226), .Y(n1784) );
  AOI21xp33_ASAP7_75t_SL U27190 ( .A1(n31157), .A2(uart1_r_RHOLD__7__4_), .B(
        n30764), .Y(n2143) );
  NAND2xp5_ASAP7_75t_SL U27191 ( .A(n24423), .B(n29017), .Y(n28961) );
  AOI21xp33_ASAP7_75t_SL U27192 ( .A1(n31177), .A2(uart1_r_RHOLD__8__4_), .B(
        n30769), .Y(n2144) );
  AOI21xp33_ASAP7_75t_SL U27193 ( .A1(n31187), .A2(uart1_r_RHOLD__16__5_), .B(
        n30064), .Y(n2121) );
  AOI21xp33_ASAP7_75t_SL U27194 ( .A1(n31161), .A2(uart1_r_RHOLD__30__6_), .B(
        n31160), .Y(n2104) );
  AOI21xp33_ASAP7_75t_SL U27195 ( .A1(n31181), .A2(uart1_r_RHOLD__9__4_), .B(
        n30770), .Y(n2145) );
  NAND2xp33_ASAP7_75t_SL U27196 ( .A(n31298), .B(n24644), .Y(n32735) );
  AOI21xp33_ASAP7_75t_SL U27197 ( .A1(n31149), .A2(uart1_r_RHOLD__10__4_), .B(
        n30762), .Y(n2146) );
  AOI21xp33_ASAP7_75t_SL U27198 ( .A1(n31077), .A2(uart1_r_RHOLD__31__6_), .B(
        n31076), .Y(n2105) );
  AOI21xp33_ASAP7_75t_SL U27199 ( .A1(n31069), .A2(uart1_r_RHOLD__27__5_), .B(
        n30033), .Y(n2132) );
  OAI21xp33_ASAP7_75t_SL U27200 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_X__ICC__2_), .B(n29171), .Y(n1789) );
  AOI21xp33_ASAP7_75t_SL U27201 ( .A1(n31161), .A2(uart1_r_RHOLD__30__4_), .B(
        n30765), .Y(n2166) );
  AOI21xp33_ASAP7_75t_SL U27202 ( .A1(n31177), .A2(uart1_r_RHOLD__8__5_), .B(
        n30060), .Y(n2113) );
  AOI21xp33_ASAP7_75t_SL U27203 ( .A1(n31077), .A2(uart1_r_RHOLD__31__4_), .B(
        n30744), .Y(n2167) );
  AOI21xp33_ASAP7_75t_SL U27204 ( .A1(n31069), .A2(uart1_r_RHOLD__27__7_), .B(
        n30836), .Y(n2070) );
  INVxp33_ASAP7_75t_SL U27205 ( .A(n26162), .Y(n26167) );
  AOI21xp33_ASAP7_75t_SL U27206 ( .A1(n31173), .A2(uart1_r_RHOLD__2__3_), .B(
        n28221), .Y(n2169) );
  AOI21xp33_ASAP7_75t_SL U27207 ( .A1(n31153), .A2(uart1_r_RHOLD__4__5_), .B(
        n30054), .Y(n2109) );
  NAND2xp5_ASAP7_75t_SL U27208 ( .A(n24681), .B(n27241), .Y(n31343) );
  AOI21xp33_ASAP7_75t_SL U27209 ( .A1(n31137), .A2(uart1_r_RHOLD__25__7_), .B(
        n30853), .Y(n2068) );
  AOI21xp33_ASAP7_75t_SL U27210 ( .A1(n31169), .A2(uart1_r_RHOLD__5__5_), .B(
        n30058), .Y(n2110) );
  AOI21xp33_ASAP7_75t_SL U27211 ( .A1(n31157), .A2(uart1_r_RHOLD__7__5_), .B(
        n30055), .Y(n2112) );
  AOI21xp33_ASAP7_75t_SL U27212 ( .A1(n31137), .A2(uart1_r_RHOLD__25__5_), .B(
        n30050), .Y(n2130) );
  AOI21xp33_ASAP7_75t_SL U27213 ( .A1(n31153), .A2(uart1_r_RHOLD__4__3_), .B(
        n28216), .Y(n2171) );
  AOI21xp33_ASAP7_75t_SL U27214 ( .A1(n31137), .A2(uart1_r_RHOLD__25__6_), .B(
        n31136), .Y(n2099) );
  AOI21xp33_ASAP7_75t_SL U27215 ( .A1(n31169), .A2(uart1_r_RHOLD__5__3_), .B(
        n28220), .Y(n2172) );
  OAI21xp33_ASAP7_75t_SRAM U27216 ( .A1(n31001), .A2(n31000), .B(n30999), .Y(
        n31003) );
  AOI21xp33_ASAP7_75t_SL U27217 ( .A1(n31181), .A2(uart1_r_RHOLD__9__5_), .B(
        n30061), .Y(n2114) );
  AOI21xp33_ASAP7_75t_SL U27218 ( .A1(n31145), .A2(uart1_r_RHOLD__19__5_), .B(
        n30052), .Y(n2124) );
  AOI21xp33_ASAP7_75t_SL U27219 ( .A1(n31187), .A2(uart1_r_RHOLD__16__6_), .B(
        n31186), .Y(n2090) );
  AOI21xp33_ASAP7_75t_SL U27220 ( .A1(n31069), .A2(uart1_r_RHOLD__27__4_), .B(
        n30742), .Y(n2163) );
  AOI21xp33_ASAP7_75t_SL U27221 ( .A1(n31173), .A2(uart1_r_RHOLD__2__6_), .B(
        n31172), .Y(n2076) );
  AOI21xp33_ASAP7_75t_SL U27222 ( .A1(n31077), .A2(uart1_r_RHOLD__31__7_), .B(
        n30838), .Y(n2074) );
  AOI21xp33_ASAP7_75t_SL U27223 ( .A1(n31141), .A2(uart1_r_RHOLD__20__5_), .B(
        n30051), .Y(n2125) );
  AOI21xp33_ASAP7_75t_SL U27224 ( .A1(n31161), .A2(uart1_r_RHOLD__30__5_), .B(
        n30056), .Y(n2135) );
  AOI21xp33_ASAP7_75t_SL U27225 ( .A1(n31161), .A2(uart1_r_RHOLD__30__7_), .B(
        n30859), .Y(n2073) );
  AOI21xp33_ASAP7_75t_SL U27226 ( .A1(n31137), .A2(uart1_r_RHOLD__25__4_), .B(
        n30759), .Y(n2161) );
  AOI21xp33_ASAP7_75t_SL U27227 ( .A1(n31173), .A2(uart1_r_RHOLD__2__5_), .B(
        n30059), .Y(n2107) );
  INVxp33_ASAP7_75t_SL U27228 ( .A(n29664), .Y(n29879) );
  AOI22xp33_ASAP7_75t_SL U27229 ( .A1(dc_q[20]), .A2(n31004), .B1(dt_q[16]), 
        .B2(n29991), .Y(n26966) );
  AOI21xp33_ASAP7_75t_SL U27230 ( .A1(n30423), .A2(n30453), .B(n30422), .Y(
        n30424) );
  OAI21xp33_ASAP7_75t_SL U27231 ( .A1(n29108), .A2(n29114), .B(n24532), .Y(
        n2369) );
  AOI22xp33_ASAP7_75t_SL U27232 ( .A1(dc_q[22]), .A2(n31004), .B1(dt_q[18]), 
        .B2(n29991), .Y(n26223) );
  INVxp67_ASAP7_75t_SL U27233 ( .A(n32164), .Y(n24761) );
  AOI21xp33_ASAP7_75t_SL U27234 ( .A1(n30302), .A2(n30453), .B(n30301), .Y(
        n30303) );
  AOI21xp33_ASAP7_75t_SL U27235 ( .A1(n25966), .A2(n25965), .B(n24695), .Y(
        n25967) );
  NOR2xp33_ASAP7_75t_SL U27236 ( .A(n23163), .B(n25486), .Y(n25503) );
  OAI21xp33_ASAP7_75t_SL U27237 ( .A1(n22902), .A2(n25198), .B(n25114), .Y(
        n26389) );
  NAND2xp33_ASAP7_75t_SL U27238 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[60]), .B(
        n24583), .Y(n25256) );
  AOI22xp33_ASAP7_75t_SL U27239 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__31_), .B1(u0_0_leon3x0_p0_ici[59]), 
        .B2(n29059), .Y(n25885) );
  OAI21xp33_ASAP7_75t_SL U27240 ( .A1(n18806), .A2(n32661), .B(n29810), .Y(
        n31681) );
  INVxp67_ASAP7_75t_SL U27241 ( .A(n30340), .Y(n30345) );
  INVxp67_ASAP7_75t_SL U27242 ( .A(add_x_735_n136), .Y(add_x_735_n134) );
  OAI21xp33_ASAP7_75t_SL U27243 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_E__SHLEFT_), .B(n25007), .Y(n3568) );
  NAND2xp33_ASAP7_75t_SL U27244 ( .A(n26482), .B(n28825), .Y(n26915) );
  NAND2xp33_ASAP7_75t_SL U27245 ( .A(n30614), .B(n30452), .Y(n28937) );
  INVxp67_ASAP7_75t_SL U27246 ( .A(n26430), .Y(n26432) );
  NAND2xp33_ASAP7_75t_SL U27247 ( .A(n24681), .B(n25897), .Y(n30226) );
  NOR2xp33_ASAP7_75t_SL U27248 ( .A(n23365), .B(u0_0_leon3x0_p0_divi[29]), .Y(
        add_x_735_n47) );
  AOI22xp33_ASAP7_75t_SL U27249 ( .A1(dc_q[18]), .A2(n31004), .B1(dt_q[14]), 
        .B2(n29991), .Y(n25717) );
  NAND2xp5_ASAP7_75t_SL U27250 ( .A(n31999), .B(n24583), .Y(n25253) );
  INVxp67_ASAP7_75t_SL U27251 ( .A(add_x_735_n67), .Y(add_x_735_n276) );
  AOI22xp33_ASAP7_75t_SL U27252 ( .A1(u0_0_leon3x0_p0_c0mmu_mcii[18]), .A2(
        n31877), .B1(u0_0_leon3x0_p0_c0mmu_mcdi[54]), .B2(n24583), .Y(n32780)
         );
  AOI21xp33_ASAP7_75t_SL U27253 ( .A1(n29245), .A2(n29244), .B(n24695), .Y(
        n29246) );
  OAI21xp33_ASAP7_75t_SL U27254 ( .A1(n22419), .A2(uart1_r_BRATE__9_), .B(
        n28149), .Y(n1800) );
  AND2x2_ASAP7_75t_SL U27255 ( .A(n23960), .B(n22416), .Y(n25791) );
  NAND2xp5_ASAP7_75t_SL U27256 ( .A(dt_q[27]), .B(n24573), .Y(n25037) );
  NAND2xp33_ASAP7_75t_SL U27257 ( .A(add_x_735_A_9_), .B(n22416), .Y(n25757)
         );
  INVxp67_ASAP7_75t_SL U27258 ( .A(mult_x_1196_n3238), .Y(n22706) );
  NAND2xp33_ASAP7_75t_SL U27259 ( .A(n22721), .B(n22416), .Y(n25465) );
  AND2x2_ASAP7_75t_SL U27260 ( .A(n22939), .B(n22416), .Y(n26142) );
  AOI211xp5_ASAP7_75t_SRAM U27261 ( .A1(n29322), .A2(n29321), .B(n24695), .C(
        n29320), .Y(n29323) );
  OAI21xp33_ASAP7_75t_SL U27262 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__WIM__4_), .B(n29625), .Y(n2725) );
  NAND2xp33_ASAP7_75t_SL U27263 ( .A(n18610), .B(n22416), .Y(n25457) );
  AOI211xp5_ASAP7_75t_SRAM U27264 ( .A1(n29300), .A2(n29299), .B(n24695), .C(
        n29298), .Y(n29301) );
  INVxp67_ASAP7_75t_SL U27265 ( .A(add_x_735_n241), .Y(add_x_735_n297) );
  AOI21xp33_ASAP7_75t_SL U27266 ( .A1(n22416), .A2(n22837), .B(n26155), .Y(
        n25796) );
  AOI21xp33_ASAP7_75t_SL U27267 ( .A1(n26278), .A2(n23969), .B(n26155), .Y(
        n25797) );
  OR2x2_ASAP7_75t_SL U27268 ( .A(n23651), .B(n25198), .Y(n23649) );
  AOI21xp33_ASAP7_75t_SL U27269 ( .A1(n22416), .A2(n23161), .B(n18813), .Y(
        n25091) );
  OAI21xp33_ASAP7_75t_SL U27270 ( .A1(n22419), .A2(uart1_r_BRATE__10_), .B(
        n28145), .Y(n2885) );
  NAND2xp33_ASAP7_75t_SL U27271 ( .A(n27275), .B(n29598), .Y(n26706) );
  OAI21xp33_ASAP7_75t_SL U27272 ( .A1(n22419), .A2(uart1_r_BRATE__8_), .B(
        n28151), .Y(n2886) );
  OAI21xp33_ASAP7_75t_SL U27273 ( .A1(n22419), .A2(uart1_r_BRATE__7_), .B(
        n28152), .Y(n2887) );
  OAI21xp33_ASAP7_75t_SL U27274 ( .A1(n22419), .A2(uart1_r_BRATE__6_), .B(
        n28153), .Y(n2888) );
  AOI21xp33_ASAP7_75t_SL U27275 ( .A1(n22417), .A2(n29150), .B(n22902), .Y(
        n26262) );
  NOR2xp33_ASAP7_75t_SL U27276 ( .A(n22417), .B(n23447), .Y(n24486) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27277 ( .A1(u0_0_leon3x0_p0_divi[6]), .A2(n28931), 
        .B(n28772), .C(n18394), .Y(n28773) );
  INVxp67_ASAP7_75t_SL U27278 ( .A(add_x_735_n112), .Y(add_x_735_n281) );
  INVxp67_ASAP7_75t_SL U27279 ( .A(add_x_735_n105), .Y(add_x_735_n280) );
  AOI21xp33_ASAP7_75t_SL U27280 ( .A1(n29738), .A2(u0_0_dbgo_SU_), .B(n29209), 
        .Y(n29210) );
  OAI21xp5_ASAP7_75t_SL U27281 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__7_), .A2(
        n29216), .B(n29215), .Y(n29218) );
  INVxp67_ASAP7_75t_SL U27282 ( .A(u0_0_leon3x0_p0_divi[30]), .Y(n31418) );
  AOI211xp5_ASAP7_75t_SRAM U27283 ( .A1(n28243), .A2(n28242), .B(n24695), .C(
        n28241), .Y(n28244) );
  OAI21xp33_ASAP7_75t_SL U27284 ( .A1(n22419), .A2(uart1_r_BRATE__5_), .B(
        n28154), .Y(n2889) );
  NAND2xp33_ASAP7_75t_SL U27285 ( .A(n23965), .B(n22416), .Y(n25189) );
  OAI21xp33_ASAP7_75t_SL U27286 ( .A1(n22419), .A2(uart1_r_BRATE__4_), .B(
        n28157), .Y(n2890) );
  NAND2xp5_ASAP7_75t_SL U27287 ( .A(n31398), .B(n29866), .Y(n29614) );
  OAI21xp33_ASAP7_75t_SL U27288 ( .A1(n22419), .A2(uart1_r_BRATE__3_), .B(
        n28161), .Y(n2891) );
  OAI21xp33_ASAP7_75t_SL U27289 ( .A1(n22419), .A2(uart1_r_BRATE__2_), .B(
        n28165), .Y(n2892) );
  OAI21xp33_ASAP7_75t_SL U27290 ( .A1(n22419), .A2(uart1_r_BRATE__1_), .B(
        n28170), .Y(n2893) );
  AOI211xp5_ASAP7_75t_SRAM U27291 ( .A1(n29267), .A2(n29266), .B(n24695), .C(
        n29265), .Y(n29268) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27292 ( .A1(apbi[1]), .A2(n24695), .B(n29522), 
        .C(n26132), .Y(n2900) );
  AOI22xp33_ASAP7_75t_SL U27293 ( .A1(dc_q[17]), .A2(n31473), .B1(dt_q[13]), 
        .B2(n24573), .Y(n27253) );
  INVxp67_ASAP7_75t_SL U27294 ( .A(add_x_735_n198), .Y(add_x_735_n291) );
  AOI21xp33_ASAP7_75t_SL U27295 ( .A1(n26383), .A2(n29150), .B(n22418), .Y(
        n26385) );
  NAND2xp5_ASAP7_75t_SL U27296 ( .A(n26534), .B(n28878), .Y(n26535) );
  AOI21xp5_ASAP7_75t_SL U27297 ( .A1(n26429), .A2(n29150), .B(n22493), .Y(
        n26430) );
  AOI211xp5_ASAP7_75t_SRAM U27298 ( .A1(n18299), .A2(n29148), .B(n24631), .C(
        u0_0_leon3x0_p0_divi[14]), .Y(n26570) );
  OAI21xp33_ASAP7_75t_SL U27299 ( .A1(n22379), .A2(u0_0_leon3x0_p0_dci[5]), 
        .B(n24981), .Y(n3590) );
  INVxp67_ASAP7_75t_SL U27300 ( .A(add_x_735_n181), .Y(add_x_735_n179) );
  AOI211xp5_ASAP7_75t_SRAM U27301 ( .A1(n29313), .A2(n29312), .B(n24695), .C(
        n29311), .Y(n29314) );
  INVxp67_ASAP7_75t_SL U27302 ( .A(add_x_735_n130), .Y(add_x_735_n283) );
  AND2x2_ASAP7_75t_SL U27303 ( .A(n23964), .B(n22416), .Y(n25477) );
  AOI21xp33_ASAP7_75t_SL U27304 ( .A1(n29379), .A2(n29378), .B(n24695), .Y(
        n29380) );
  INVxp67_ASAP7_75t_SL U27305 ( .A(n27316), .Y(n28046) );
  INVxp67_ASAP7_75t_SL U27306 ( .A(n29603), .Y(n28790) );
  AOI21xp33_ASAP7_75t_SL U27307 ( .A1(n29211), .A2(
        u0_0_leon3x0_p0_iu_r_X__RESULT__0_), .B(n24679), .Y(n26774) );
  NAND2xp33_ASAP7_75t_SL U27308 ( .A(n31302), .B(n31605), .Y(n32193) );
  NAND2xp5_ASAP7_75t_SL U27309 ( .A(n29074), .B(n28403), .Y(n28489) );
  AOI21xp33_ASAP7_75t_SL U27310 ( .A1(n28403), .A2(n27027), .B(n30006), .Y(
        n26961) );
  INVxp33_ASAP7_75t_SRAM U27311 ( .A(u0_0_leon3x0_p0_divi[24]), .Y(n28431) );
  INVxp67_ASAP7_75t_SL U27312 ( .A(n30593), .Y(n30651) );
  OAI21xp33_ASAP7_75t_SL U27313 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_X__ICC__0_), .B(n27019), .Y(n2279) );
  AOI22xp33_ASAP7_75t_SL U27314 ( .A1(dataout[30]), .A2(n22433), .B1(n32972), 
        .B2(n32963), .Y(n32965) );
  AOI22xp33_ASAP7_75t_SL U27315 ( .A1(dataout[29]), .A2(n22433), .B1(n32972), 
        .B2(n32955), .Y(n32957) );
  AOI22xp33_ASAP7_75t_SL U27316 ( .A1(dataout[28]), .A2(n22433), .B1(n32972), 
        .B2(n32947), .Y(n32949) );
  INVxp33_ASAP7_75t_SL U27317 ( .A(u0_0_leon3x0_p0_divi[15]), .Y(n26682) );
  OA21x2_ASAP7_75t_SL U27318 ( .A1(n23964), .A2(n28827), .B(
        u0_0_leon3x0_p0_divi[14]), .Y(n26566) );
  NOR2xp33_ASAP7_75t_SL U27319 ( .A(n23161), .B(u0_0_leon3x0_p0_divi[19]), .Y(
        add_x_735_n141) );
  AOI21xp5_ASAP7_75t_SL U27320 ( .A1(n25725), .A2(
        u0_0_leon3x0_p0_iu_r_X__NPC__1_), .B(n25724), .Y(n3703) );
  AOI22xp33_ASAP7_75t_SL U27321 ( .A1(dataout[27]), .A2(n22433), .B1(n32972), 
        .B2(n32939), .Y(n32941) );
  AOI22xp33_ASAP7_75t_SL U27322 ( .A1(dataout[25]), .A2(n22433), .B1(n32972), 
        .B2(n32923), .Y(n32925) );
  NOR2x1_ASAP7_75t_SL U27323 ( .A(n22436), .B(u0_0_leon3x0_p0_divi[21]), .Y(
        add_x_735_n123) );
  AOI22xp33_ASAP7_75t_SL U27324 ( .A1(dataout[24]), .A2(n22433), .B1(n32972), 
        .B2(n32911), .Y(n32915) );
  AOI22xp33_ASAP7_75t_SL U27325 ( .A1(dataout[31]), .A2(n22433), .B1(n32972), 
        .B2(n32971), .Y(n32975) );
  NOR2xp33_ASAP7_75t_SL U27326 ( .A(n22556), .B(u0_0_leon3x0_p0_divi[25]), .Y(
        add_x_735_n85) );
  OAI21xp33_ASAP7_75t_SL U27327 ( .A1(n23229), .A2(n28956), .B(n30593), .Y(
        n28958) );
  OAI21xp33_ASAP7_75t_SL U27328 ( .A1(n22421), .A2(n28904), .B(n30593), .Y(
        n28906) );
  NAND2xp33_ASAP7_75t_SL U27329 ( .A(u0_0_leon3x0_p0_divi[39]), .B(n22373), 
        .Y(n30393) );
  INVxp33_ASAP7_75t_SL U27330 ( .A(n29211), .Y(n29216) );
  NAND2xp33_ASAP7_75t_SL U27331 ( .A(n23964), .B(n24577), .Y(n26146) );
  OAI21xp33_ASAP7_75t_SL U27332 ( .A1(n22379), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__TT__0_), .B(n29227), .Y(n29228) );
  OAI21xp33_ASAP7_75t_SL U27333 ( .A1(n22427), .A2(DP_OP_1196_128_7433_n455), 
        .B(n30816), .Y(n3542) );
  OAI21xp5_ASAP7_75t_SL U27334 ( .A1(n3916), .A2(n29738), .B(n29730), .Y(
        n18053) );
  NAND2xp5_ASAP7_75t_SL U27335 ( .A(sr1_r_MCFG1__BEXCEN_), .B(n32003), .Y(
        n31371) );
  OAI21xp33_ASAP7_75t_SL U27336 ( .A1(n23229), .A2(n23837), .B(n30593), .Y(
        n28866) );
  OAI21xp33_ASAP7_75t_SL U27337 ( .A1(n22428), .A2(DP_OP_1196_128_7433_n452), 
        .B(n28963), .Y(n3470) );
  NAND2xp33_ASAP7_75t_SL U27338 ( .A(n29744), .B(n22419), .Y(n28151) );
  AOI21xp33_ASAP7_75t_SL U27339 ( .A1(n32003), .A2(sr1_r_MCFG1__ROMWIDTH__0_), 
        .B(n31849), .Y(n29747) );
  NAND2xp33_ASAP7_75t_SL U27340 ( .A(n30978), .B(n22419), .Y(n28145) );
  INVxp33_ASAP7_75t_SL U27341 ( .A(u0_0_leon3x0_p0_divi[21]), .Y(n28491) );
  NAND2xp33_ASAP7_75t_SL U27342 ( .A(apbi[11]), .B(n22419), .Y(n28138) );
  NAND2xp33_ASAP7_75t_SL U27343 ( .A(n31197), .B(n22419), .Y(n28153) );
  INVxp33_ASAP7_75t_SRAM U27344 ( .A(u0_0_leon3x0_p0_divi[17]), .Y(n25822) );
  NAND2xp33_ASAP7_75t_SL U27345 ( .A(n30833), .B(n22419), .Y(n28152) );
  NAND2xp33_ASAP7_75t_SL U27346 ( .A(n30073), .B(n22419), .Y(n28154) );
  INVx1_ASAP7_75t_SL U27347 ( .A(u0_0_leon3x0_p0_divi[4]), .Y(n26307) );
  INVxp67_ASAP7_75t_SL U27348 ( .A(u0_0_leon3x0_p0_divi[6]), .Y(n28770) );
  NAND2xp33_ASAP7_75t_SL U27349 ( .A(n27493), .B(n22419), .Y(n28170) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U27350 ( .A1(n29199), .A2(n22379), .B(n30472), 
        .C(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .Y(n29200) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27351 ( .A1(apbi[9]), .A2(n31501), .B(n30138), 
        .C(n24695), .Y(n1802) );
  NAND2xp33_ASAP7_75t_SL U27352 ( .A(n30139), .B(n22419), .Y(n28149) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27353 ( .A1(apbi[6]), .A2(n31501), .B(n31196), 
        .C(n24695), .Y(n2903) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27354 ( .A1(apbi[7]), .A2(n31501), .B(n30869), 
        .C(n24695), .Y(n2902) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27355 ( .A1(apbi[3]), .A2(n31501), .B(n28237), 
        .C(n24695), .Y(n2898) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27356 ( .A1(apbi[0]), .A2(n31501), .B(n28058), 
        .C(n24695), .Y(n2901) );
  NAND2xp33_ASAP7_75t_SL U27357 ( .A(n30780), .B(n22419), .Y(n28157) );
  NAND2xp33_ASAP7_75t_SL U27358 ( .A(n29568), .B(n22419), .Y(n28165) );
  INVxp33_ASAP7_75t_SL U27359 ( .A(n31248), .Y(n30983) );
  NAND2xp33_ASAP7_75t_SL U27360 ( .A(n29510), .B(n22419), .Y(n28161) );
  NOR2xp33_ASAP7_75t_SL U27361 ( .A(n23375), .B(u0_0_leon3x0_p0_divi[5]), .Y(
        add_x_735_n247) );
  NAND2xp5_ASAP7_75t_SL U27362 ( .A(n24694), .B(n27291), .Y(n29649) );
  AOI21xp33_ASAP7_75t_SL U27363 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__18_), .B(n30310), .Y(n30311) );
  NAND2xp5_ASAP7_75t_SL U27364 ( .A(n26062), .B(n26053), .Y(n31111) );
  NAND2xp33_ASAP7_75t_SL U27365 ( .A(n22556), .B(n24578), .Y(n25479) );
  OAI21xp33_ASAP7_75t_SL U27366 ( .A1(n31396), .A2(n26413), .B(n26412), .Y(
        n26414) );
  NAND2xp5_ASAP7_75t_SL U27367 ( .A(n26032), .B(n26053), .Y(n31103) );
  INVxp33_ASAP7_75t_SL U27368 ( .A(n31250), .Y(n30982) );
  AOI21xp33_ASAP7_75t_SL U27369 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__15_), .B(n30343), .Y(n30344) );
  INVxp67_ASAP7_75t_SL U27370 ( .A(add_x_735_n259), .Y(add_x_735_n301) );
  AOI21xp33_ASAP7_75t_SL U27371 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__21_), .B(n30280), .Y(n30281) );
  AOI21xp33_ASAP7_75t_SL U27372 ( .A1(n22429), .A2(
        u0_0_leon3x0_p0_iu_r_X__Y__13_), .B(n30364), .Y(n30365) );
  INVxp67_ASAP7_75t_SL U27373 ( .A(DP_OP_1196_128_7433_n137), .Y(
        DP_OP_1196_128_7433_n139) );
  NAND2xp5_ASAP7_75t_SL U27374 ( .A(n30872), .B(n29949), .Y(n27316) );
  AOI22xp33_ASAP7_75t_SL U27375 ( .A1(u0_0_leon3x0_p0_ici[23]), .A2(n30722), 
        .B1(n29796), .B2(n32162), .Y(n28399) );
  OAI21xp33_ASAP7_75t_SL U27376 ( .A1(n31396), .A2(n26287), .B(n26286), .Y(
        n26288) );
  AOI22xp33_ASAP7_75t_SL U27377 ( .A1(u0_0_leon3x0_p0_ici[25]), .A2(n30722), 
        .B1(n28272), .B2(n32162), .Y(n28270) );
  AOI22xp33_ASAP7_75t_SL U27378 ( .A1(u0_0_leon3x0_p0_ici[26]), .A2(n30722), 
        .B1(n29579), .B2(n32162), .Y(n29582) );
  AOI22xp33_ASAP7_75t_SL U27379 ( .A1(u0_0_leon3x0_p0_ici[27]), .A2(n30722), 
        .B1(n30591), .B2(n32162), .Y(n30589) );
  AOI22xp33_ASAP7_75t_SL U27380 ( .A1(u0_0_leon3x0_p0_ici[28]), .A2(n30722), 
        .B1(n26725), .B2(n32162), .Y(n26728) );
  INVx2_ASAP7_75t_SL U27381 ( .A(n23991), .Y(n22388) );
  INVxp33_ASAP7_75t_SL U27382 ( .A(n31238), .Y(n30870) );
  AOI22xp33_ASAP7_75t_SL U27383 ( .A1(u0_0_leon3x0_p0_ici[7]), .A2(n30722), 
        .B1(n28714), .B2(n32162), .Y(n28712) );
  AOI22xp33_ASAP7_75t_SL U27384 ( .A1(u0_0_leon3x0_p0_ici[5]), .A2(n30722), 
        .B1(n30721), .B2(n32162), .Y(n30729) );
  AOI22xp33_ASAP7_75t_SL U27385 ( .A1(u0_0_leon3x0_p0_ici[9]), .A2(n30722), 
        .B1(n29832), .B2(n32162), .Y(n29835) );
  AOI22xp33_ASAP7_75t_SL U27386 ( .A1(u0_0_leon3x0_p0_ici[4]), .A2(n30722), 
        .B1(n29899), .B2(n32162), .Y(n29897) );
  AOI22xp33_ASAP7_75t_SL U27387 ( .A1(u0_0_leon3x0_p0_ici[10]), .A2(n30722), 
        .B1(n28602), .B2(n32162), .Y(n28600) );
  AOI22xp33_ASAP7_75t_SL U27388 ( .A1(u0_0_leon3x0_p0_ici[11]), .A2(n30722), 
        .B1(n28586), .B2(n32162), .Y(n27187) );
  NAND2xp33_ASAP7_75t_SRAM U27389 ( .A(uart1_r_TRADDR__0_), .B(n27702), .Y(
        n27710) );
  BUFx6f_ASAP7_75t_SL U27390 ( .A(mult_x_1196_n6), .Y(n22389) );
  AOI22xp33_ASAP7_75t_SL U27391 ( .A1(u0_0_leon3x0_p0_ici[2]), .A2(n30722), 
        .B1(n29680), .B2(n32162), .Y(n29683) );
  AOI22xp33_ASAP7_75t_SL U27392 ( .A1(u0_0_leon3x0_p0_ici[13]), .A2(n30722), 
        .B1(n28554), .B2(n32162), .Y(n27239) );
  AOI22xp33_ASAP7_75t_SL U27393 ( .A1(u0_0_leon3x0_p0_ici[14]), .A2(n30722), 
        .B1(n27275), .B2(n32162), .Y(n27278) );
  AOI22xp33_ASAP7_75t_SL U27394 ( .A1(u0_0_leon3x0_p0_ici[1]), .A2(n30722), 
        .B1(n29482), .B2(n32162), .Y(n29485) );
  AOI22xp33_ASAP7_75t_SL U27395 ( .A1(u0_0_leon3x0_p0_ici[0]), .A2(n30722), 
        .B1(n29490), .B2(n32162), .Y(n29493) );
  AOI22xp33_ASAP7_75t_SL U27396 ( .A1(u0_0_leon3x0_p0_ici[15]), .A2(n30722), 
        .B1(n28540), .B2(n32162), .Y(n25741) );
  AOI22xp33_ASAP7_75t_SL U27397 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__PC__2_), 
        .A2(n30722), .B1(n30465), .B2(n32162), .Y(n28912) );
  AOI22xp33_ASAP7_75t_SL U27398 ( .A1(u0_0_leon3x0_p0_ici[16]), .A2(n30722), 
        .B1(n28529), .B2(n32162), .Y(n25756) );
  AOI22xp33_ASAP7_75t_SL U27399 ( .A1(u0_0_leon3x0_p0_ici[17]), .A2(n30722), 
        .B1(n27027), .B2(n32162), .Y(n26985) );
  AOI22xp33_ASAP7_75t_SL U27400 ( .A1(u0_0_leon3x0_p0_ici[18]), .A2(n30722), 
        .B1(n28521), .B2(n32162), .Y(n27055) );
  AOI22xp33_ASAP7_75t_SL U27401 ( .A1(u0_0_leon3x0_p0_ici[20]), .A2(n30722), 
        .B1(n29067), .B2(n32162), .Y(n29070) );
  AOI22xp33_ASAP7_75t_SL U27402 ( .A1(u0_0_leon3x0_p0_ici[21]), .A2(n30722), 
        .B1(n29778), .B2(n32162), .Y(n29781) );
  AOI22xp33_ASAP7_75t_SL U27403 ( .A1(u0_0_leon3x0_p0_ici[22]), .A2(n30722), 
        .B1(n29783), .B2(n32162), .Y(n28459) );
  NAND2xp5_ASAP7_75t_SL U27404 ( .A(n27895), .B(n27400), .Y(n27425) );
  INVx1_ASAP7_75t_SL U27405 ( .A(DP_OP_1196_128_7433_n339), .Y(
        DP_OP_1196_128_7433_n4) );
  INVx1_ASAP7_75t_SL U27406 ( .A(n25033), .Y(n25025) );
  A2O1A1Ixp33_ASAP7_75t_SL U27407 ( .A1(uart1_r_BRATE__11_), .A2(n28172), .B(
        uart1_uarto_SCALER__11_), .C(n24531), .Y(n28139) );
  INVx2_ASAP7_75t_SL U27408 ( .A(n18798), .Y(n29060) );
  AOI21xp33_ASAP7_75t_SRAM U27409 ( .A1(n24932), .A2(n30955), .B(n24964), .Y(
        n24933) );
  NAND2xp5_ASAP7_75t_SL U27410 ( .A(n26049), .B(n26066), .Y(n31127) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27411 ( .A1(n27995), .A2(n27994), .B(
        uart1_r_TRADDR__0_), .C(n27993), .Y(n28026) );
  NAND2xp33_ASAP7_75t_SL U27412 ( .A(uart1_r_RCNT__0_), .B(n31238), .Y(n27495)
         );
  OAI21xp33_ASAP7_75t_SL U27413 ( .A1(n31396), .A2(n29785), .B(n29784), .Y(
        n29786) );
  OAI21xp33_ASAP7_75t_SL U27414 ( .A1(n31396), .A2(n29495), .B(n29494), .Y(
        n29496) );
  OAI21xp33_ASAP7_75t_SL U27415 ( .A1(n31396), .A2(n27189), .B(n27188), .Y(
        n27190) );
  INVxp33_ASAP7_75t_SL U27416 ( .A(n28631), .Y(n28632) );
  NAND2xp5_ASAP7_75t_SL U27417 ( .A(n24681), .B(n28536), .Y(n30593) );
  AOI21xp33_ASAP7_75t_SL U27418 ( .A1(n22375), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__6_), .B(n30006), .Y(n25857) );
  AOI21xp33_ASAP7_75t_SL U27419 ( .A1(n22375), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__4_), .B(n30006), .Y(n25871) );
  INVxp67_ASAP7_75t_SL U27420 ( .A(n22968), .Y(n24690) );
  AOI21xp33_ASAP7_75t_SL U27421 ( .A1(n22429), .A2(u0_0_leon3x0_p0_muli[7]), 
        .B(n30400), .Y(n30401) );
  OAI21xp33_ASAP7_75t_SL U27422 ( .A1(n31396), .A2(n29798), .B(n29797), .Y(
        n29799) );
  NAND2xp33_ASAP7_75t_SRAM U27423 ( .A(n22721), .B(n26338), .Y(n25424) );
  AOI21xp33_ASAP7_75t_SL U27424 ( .A1(n22429), .A2(u0_0_leon3x0_p0_muli[6]), 
        .B(n30410), .Y(n30411) );
  AOI21xp33_ASAP7_75t_SL U27425 ( .A1(n22375), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__2_), .B(n30006), .Y(n29560) );
  NOR2x1p5_ASAP7_75t_SL U27426 ( .A(n25125), .B(n25126), .Y(
        u0_0_leon3x0_p0_divi[30]) );
  OAI21xp33_ASAP7_75t_SL U27427 ( .A1(n22379), .A2(u0_0_leon3x0_p0_muli[10]), 
        .B(n30680), .Y(n3728) );
  NOR2x1_ASAP7_75t_SL U27428 ( .A(n24463), .B(n26988), .Y(
        u0_0_leon3x0_p0_divi[19]) );
  INVx1_ASAP7_75t_SL U27429 ( .A(n29563), .Y(n30010) );
  OAI21xp33_ASAP7_75t_SL U27430 ( .A1(n31396), .A2(n30467), .B(n30466), .Y(
        n30468) );
  NAND2xp33_ASAP7_75t_SL U27431 ( .A(n26521), .B(n22375), .Y(n26438) );
  OA21x2_ASAP7_75t_SL U27432 ( .A1(u0_0_leon3x0_p0_divo[31]), .A2(n26188), .B(
        n22422), .Y(n26187) );
  OAI21xp5_ASAP7_75t_SL U27433 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__16_), 
        .A2(n24651), .B(n27234), .Y(n2621) );
  NOR2x1_ASAP7_75t_SL U27434 ( .A(n25084), .B(n28926), .Y(n28977) );
  NAND2xp33_ASAP7_75t_SL U27435 ( .A(n26956), .B(n22375), .Y(n26906) );
  AOI21xp33_ASAP7_75t_SL U27436 ( .A1(n24581), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__5_), .B(n28887), .Y(n26313) );
  INVxp67_ASAP7_75t_SL U27437 ( .A(n30721), .Y(n29930) );
  AOI22xp33_ASAP7_75t_SL U27438 ( .A1(irqctrl0_r_IMASK__0__15_), .A2(n31249), 
        .B1(irqctrl0_r_IFORCE__0__15_), .B2(n31251), .Y(n31022) );
  OAI21xp5_ASAP7_75t_SL U27439 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__17_), 
        .A2(n24651), .B(n27272), .Y(n2597) );
  OAI21xp5_ASAP7_75t_SL U27440 ( .A1(u0_0_leon3x0_p0_ici[45]), .A2(n24651), 
        .B(n27259), .Y(n2601) );
  OAI21xp5_ASAP7_75t_SL U27441 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__17_), 
        .A2(n24651), .B(n27261), .Y(n2599) );
  NAND2xp33_ASAP7_75t_SL U27442 ( .A(n27175), .B(n22375), .Y(n27122) );
  OAI21xp33_ASAP7_75t_SL U27443 ( .A1(n31396), .A2(n29864), .B(n28280), .Y(
        n28281) );
  NAND2xp33_ASAP7_75t_SL U27444 ( .A(n29841), .B(n22375), .Y(n28693) );
  NAND2xp33_ASAP7_75t_SL U27445 ( .A(n26318), .B(n22375), .Y(n26319) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U27446 ( .A1(n25688), .A2(n25687), .B(n31980), 
        .C(n25686), .Y(n25706) );
  NAND2xp33_ASAP7_75t_SL U27447 ( .A(n26692), .B(n22375), .Y(n26693) );
  NAND2xp33_ASAP7_75t_SL U27448 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__28_), .B(
        n22375), .Y(n26945) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27449 ( .A1(u0_0_leon3x0_p0_iu_r_E__JMPL_), .A2(
        n27067), .B(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__21_), .C(n27148), .Y(
        n27068) );
  OAI21xp33_ASAP7_75t_SL U27450 ( .A1(n31396), .A2(n26947), .B(n26946), .Y(
        n26948) );
  NAND2xp5_ASAP7_75t_SL U27451 ( .A(n25957), .B(n25963), .Y(n27293) );
  INVxp67_ASAP7_75t_SL U27452 ( .A(n29783), .Y(n29785) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27453 ( .A1(n29946), .A2(n28036), .B(n4518), .C(
        n28035), .Y(n28040) );
  INVxp67_ASAP7_75t_SL U27454 ( .A(n30666), .Y(n30674) );
  NAND2xp33_ASAP7_75t_SL U27455 ( .A(n27243), .B(n22375), .Y(n26580) );
  NAND2xp33_ASAP7_75t_SL U27456 ( .A(n26181), .B(n22375), .Y(n26182) );
  INVxp67_ASAP7_75t_SL U27457 ( .A(n29778), .Y(n26413) );
  NAND2xp33_ASAP7_75t_SL U27458 ( .A(n29619), .B(n22375), .Y(n28643) );
  OAI21xp5_ASAP7_75t_SL U27459 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__17_), 
        .A2(n24651), .B(n27274), .Y(n2595) );
  OAI21xp5_ASAP7_75t_SL U27460 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__16_), 
        .A2(n24651), .B(n27232), .Y(n2623) );
  NOR2xp33_ASAP7_75t_SL U27461 ( .A(n28769), .B(n28941), .Y(n28631) );
  NAND2xp33_ASAP7_75t_SL U27462 ( .A(n29805), .B(n22375), .Y(n28444) );
  HB1xp67_ASAP7_75t_SL U27463 ( .A(n18604), .Y(n22493) );
  OAI21xp5_ASAP7_75t_SL U27464 ( .A1(u0_0_leon3x0_p0_ici[44]), .A2(n24650), 
        .B(n27230), .Y(n2625) );
  NAND2xp33_ASAP7_75t_SL U27465 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__29_), .B(
        n22375), .Y(n26484) );
  AOI22xp33_ASAP7_75t_SL U27466 ( .A1(u0_0_leon3x0_p0_ici[35]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__7_), .B2(n30723), .Y(n29896) );
  AOI22xp33_ASAP7_75t_SL U27467 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__7_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__7_), 
        .Y(n29895) );
  NAND2xp5_ASAP7_75t_SL U27468 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__8_), .B(
        n22375), .Y(n28748) );
  OAI22xp33_ASAP7_75t_SL U27469 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__11_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__21_), .Y(
        n28519) );
  AOI22xp33_ASAP7_75t_SL U27470 ( .A1(u0_0_leon3x0_p0_ici[36]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__8_), .B2(n30723), .Y(n30728) );
  AOI22xp33_ASAP7_75t_SL U27471 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__8_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__8_), 
        .Y(n30727) );
  AOI22xp33_ASAP7_75t_SL U27472 ( .A1(u0_0_leon3x0_p0_ici[38]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__10_), .B2(n30723), .Y(n28711) );
  AOI22xp33_ASAP7_75t_SL U27473 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__10_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__10_), 
        .Y(n28710) );
  AOI22xp33_ASAP7_75t_SL U27474 ( .A1(u0_0_leon3x0_p0_ici[8]), .A2(n30722), 
        .B1(n29837), .B2(n32162), .Y(n28665) );
  INVx1_ASAP7_75t_SL U27475 ( .A(n29490), .Y(n29495) );
  AOI22xp33_ASAP7_75t_SL U27476 ( .A1(u0_0_leon3x0_p0_ici[39]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__11_), .B2(n30723), .Y(n28664) );
  AOI22xp33_ASAP7_75t_SL U27477 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__11_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__11_), 
        .Y(n28663) );
  AOI22xp33_ASAP7_75t_SL U27478 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__31_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__31_), 
        .Y(n26726) );
  AOI22xp33_ASAP7_75t_SL U27479 ( .A1(u0_0_leon3x0_p0_ici[40]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__12_), .B2(n30723), .Y(n29834) );
  AOI22xp33_ASAP7_75t_SL U27480 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__12_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__12_), 
        .Y(n29833) );
  NAND2xp33_ASAP7_75t_SL U27481 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__22_), .B(
        n22375), .Y(n28506) );
  AOI22xp33_ASAP7_75t_SL U27482 ( .A1(u0_0_leon3x0_p0_ici[41]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__13_), .B2(n30723), .Y(n28599) );
  AOI22xp33_ASAP7_75t_SL U27483 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__13_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__13_), 
        .Y(n28598) );
  OAI21xp33_ASAP7_75t_SL U27484 ( .A1(n31396), .A2(n29499), .B(n29498), .Y(
        n29500) );
  NAND2xp33_ASAP7_75t_SL U27485 ( .A(n27284), .B(n22375), .Y(n26712) );
  OAI21xp5_ASAP7_75t_SL U27486 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__14_), 
        .A2(n24650), .B(n27182), .Y(n3208) );
  NAND2xp5_ASAP7_75t_SL U27487 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__1_), .B(
        n22375), .Y(n30639) );
  NAND2xp5_ASAP7_75t_SL U27488 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__26_), .B(
        n28769), .Y(n25487) );
  NAND2xp5_ASAP7_75t_SL U27489 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__25_), .B(
        n28769), .Y(n28430) );
  AOI22xp33_ASAP7_75t_SL U27490 ( .A1(u0_0_leon3x0_p0_ici[30]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__2_), .B2(n30725), .Y(n28911) );
  AOI22xp33_ASAP7_75t_SL U27491 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__2_), 
        .A2(n30726), .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__2_), .B2(n30723), 
        .Y(n28910) );
  AOI22xp33_ASAP7_75t_SL U27492 ( .A1(u0_0_leon3x0_p0_ici[31]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__3_), .B2(n30723), .Y(n29492) );
  AOI22xp33_ASAP7_75t_SL U27493 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__3_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__3_), 
        .Y(n29491) );
  AOI22xp33_ASAP7_75t_SL U27494 ( .A1(u0_0_leon3x0_p0_ici[32]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__4_), .B2(n30723), .Y(n29484) );
  AOI22xp33_ASAP7_75t_SL U27495 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__4_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__4_), 
        .Y(n29483) );
  AOI22xp33_ASAP7_75t_SL U27496 ( .A1(u0_0_leon3x0_p0_ici[33]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__5_), .B2(n30723), .Y(n29682) );
  INVxp67_ASAP7_75t_SL U27497 ( .A(n28253), .Y(n26661) );
  AOI22xp33_ASAP7_75t_SL U27498 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__5_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__5_), 
        .Y(n29681) );
  AOI22xp33_ASAP7_75t_SL U27499 ( .A1(u0_0_leon3x0_p0_ici[57]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__29_), .B2(n30723), .Y(n29581) );
  AOI21xp33_ASAP7_75t_SL U27500 ( .A1(n24582), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__7_), .B(n28887), .Y(n28780) );
  INVxp33_ASAP7_75t_SL U27501 ( .A(n29864), .Y(n29579) );
  OAI21xp5_ASAP7_75t_SL U27502 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__28_), 
        .A2(n24652), .B(n28267), .Y(n3270) );
  AOI22xp33_ASAP7_75t_SL U27503 ( .A1(u0_0_leon3x0_p0_ici[47]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__19_), .B2(n30723), .Y(n25755) );
  INVx1_ASAP7_75t_SL U27504 ( .A(n22952), .Y(n23161) );
  NAND2xp33_ASAP7_75t_SL U27505 ( .A(n29928), .B(n22375), .Y(n28791) );
  AOI22xp33_ASAP7_75t_SL U27506 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__19_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__19_), 
        .Y(n25754) );
  AOI22xp33_ASAP7_75t_SL U27507 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__28_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__28_), 
        .Y(n28268) );
  AOI22xp33_ASAP7_75t_SL U27508 ( .A1(u0_0_leon3x0_p0_ici[48]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__20_), .B2(n30723), .Y(n26984) );
  INVx2_ASAP7_75t_SL U27509 ( .A(n31402), .Y(n22390) );
  AOI22xp33_ASAP7_75t_SL U27510 ( .A1(u0_0_leon3x0_p0_ici[56]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__28_), .B2(n30723), .Y(n28269) );
  AOI22xp33_ASAP7_75t_SL U27511 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__20_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__20_), 
        .Y(n26983) );
  AOI22xp33_ASAP7_75t_SL U27512 ( .A1(u0_0_leon3x0_p0_ici[49]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__21_), .B2(n30723), .Y(n27054) );
  AOI22xp33_ASAP7_75t_SL U27513 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__21_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__21_), 
        .Y(n27053) );
  OAI21xp5_ASAP7_75t_SL U27514 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__28_), 
        .A2(n24652), .B(n28265), .Y(n3272) );
  AOI22xp33_ASAP7_75t_SL U27515 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__26_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__26_), 
        .Y(n28397) );
  INVxp67_ASAP7_75t_SL U27516 ( .A(n26523), .Y(n29067) );
  AOI22xp33_ASAP7_75t_SL U27517 ( .A1(u0_0_leon3x0_p0_ici[51]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__23_), .B2(n30723), .Y(n29069) );
  AOI22xp33_ASAP7_75t_SL U27518 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__23_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__23_), 
        .Y(n29068) );
  AOI22xp33_ASAP7_75t_SL U27519 ( .A1(u0_0_leon3x0_p0_ici[54]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__26_), .B2(n30723), .Y(n28398) );
  AOI22xp33_ASAP7_75t_SL U27520 ( .A1(u0_0_leon3x0_p0_ici[52]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__24_), .B2(n30723), .Y(n29780) );
  AOI22xp33_ASAP7_75t_SL U27521 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__24_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__24_), 
        .Y(n29779) );
  AOI22xp33_ASAP7_75t_SL U27522 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__25_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__25_), 
        .Y(n28457) );
  AOI22xp33_ASAP7_75t_SL U27523 ( .A1(u0_0_leon3x0_p0_ici[53]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__25_), .B2(n30723), .Y(n28458) );
  AOI22xp33_ASAP7_75t_SL U27524 ( .A1(u0_0_leon3x0_p0_ici[59]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__31_), .B2(n30723), .Y(n26727) );
  AOI22xp33_ASAP7_75t_SL U27525 ( .A1(u0_0_leon3x0_p0_ici[42]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__14_), .B2(n30723), .Y(n27186) );
  AOI22xp33_ASAP7_75t_SL U27526 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__14_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__14_), 
        .Y(n27185) );
  NAND2xp33_ASAP7_75t_SL U27527 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__21_), .B(
        n22375), .Y(n27085) );
  AOI22xp33_ASAP7_75t_SL U27528 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__30_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__30_), 
        .Y(n30587) );
  INVxp33_ASAP7_75t_SL U27529 ( .A(n32068), .Y(n30680) );
  AOI22xp33_ASAP7_75t_SL U27530 ( .A1(u0_0_leon3x0_p0_ici[58]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__30_), .B2(n30723), .Y(n30588) );
  AOI22xp33_ASAP7_75t_SL U27531 ( .A1(u0_0_leon3x0_p0_ici[44]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__16_), .B2(n30723), .Y(n27238) );
  AOI22xp33_ASAP7_75t_SL U27532 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__16_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__16_), 
        .Y(n27237) );
  NAND2xp33_ASAP7_75t_SL U27533 ( .A(n27088), .B(n22375), .Y(n27002) );
  AOI22xp33_ASAP7_75t_SL U27534 ( .A1(u0_0_leon3x0_p0_ici[45]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__17_), .B2(n30723), .Y(n27277) );
  OAI21xp33_ASAP7_75t_SL U27535 ( .A1(n22379), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__8_), .B(n24523), .Y(n3666) );
  AOI22xp33_ASAP7_75t_SL U27536 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__17_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__17_), 
        .Y(n27276) );
  INVxp67_ASAP7_75t_SL U27537 ( .A(n31585), .Y(n31575) );
  OAI21xp5_ASAP7_75t_SL U27538 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__28_), 
        .A2(n24652), .B(n28263), .Y(n3274) );
  AOI22xp33_ASAP7_75t_SL U27539 ( .A1(u0_0_leon3x0_p0_ici[46]), .A2(n30724), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__18_), .B2(n30723), .Y(n25740) );
  AOI22xp33_ASAP7_75t_SL U27540 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__29_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__29_), 
        .Y(n29580) );
  AOI22xp33_ASAP7_75t_SL U27541 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__18_), 
        .A2(n30726), .B1(n30725), .B2(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__18_), 
        .Y(n25739) );
  NAND2xp5_ASAP7_75t_SL U27542 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__18_), .B(
        n28769), .Y(n25821) );
  NAND2xp5_ASAP7_75t_SL U27543 ( .A(n2931), .B(n26130), .Y(n31501) );
  NAND2xp5_ASAP7_75t_SL U27544 ( .A(n31661), .B(n33056), .Y(n31659) );
  AND2x2_ASAP7_75t_SL U27545 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__21_), 
        .B(n18806), .Y(n24491) );
  NAND2xp5_ASAP7_75t_SL U27546 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__10_), .B(
        n22375), .Y(n27164) );
  OAI31xp33_ASAP7_75t_SL U27547 ( .A1(n24989), .A2(n30956), .A3(n24922), .B(
        n24927), .Y(n24924) );
  NAND2xp5_ASAP7_75t_SL U27548 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__27_), .B(
        n28769), .Y(n26890) );
  INVx5_ASAP7_75t_SL U27549 ( .A(n24036), .Y(n22391) );
  AOI22xp33_ASAP7_75t_SL U27550 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__18_), .A2(
        n30641), .B1(rf_do_b[18]), .B2(n30640), .Y(n28537) );
  AOI22xp33_ASAP7_75t_SL U27551 ( .A1(n31391), .A2(rf_do_a[17]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__17_), .B2(n31392), .Y(n26717) );
  AOI22xp33_ASAP7_75t_SL U27552 ( .A1(u0_0_leon3x0_p0_divi[33]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[32]), .B2(n28367), .Y(n28363) );
  INVxp33_ASAP7_75t_SL U27553 ( .A(n25232), .Y(n26191) );
  AOI22xp33_ASAP7_75t_SL U27554 ( .A1(u0_0_leon3x0_p0_divi[34]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[33]), .B2(n28367), .Y(n28361) );
  OAI21xp33_ASAP7_75t_SL U27555 ( .A1(n25687), .A2(n25695), .B(n24947), .Y(
        n24948) );
  NAND2xp33_ASAP7_75t_SL U27556 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__0_), .B(
        n31392), .Y(n31393) );
  NAND2xp33_ASAP7_75t_SL U27557 ( .A(n27271), .B(n22427), .Y(n27272) );
  NAND2xp5_ASAP7_75t_SL U27558 ( .A(n28180), .B(n26015), .Y(n26014) );
  INVxp67_ASAP7_75t_SL U27559 ( .A(n31553), .Y(n31555) );
  NAND2xp33_ASAP7_75t_SL U27560 ( .A(n27260), .B(n22427), .Y(n27261) );
  AOI22xp33_ASAP7_75t_SL U27561 ( .A1(n31391), .A2(rf_do_a[27]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__27_), .B2(n31392), .Y(n26952) );
  NAND2xp33_ASAP7_75t_SL U27562 ( .A(n27258), .B(n22427), .Y(n27259) );
  INVxp67_ASAP7_75t_SL U27563 ( .A(n31556), .Y(n31557) );
  AOI22xp33_ASAP7_75t_SL U27564 ( .A1(u0_0_leon3x0_p0_divi[62]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[61]), .B2(n28367), .Y(n28300) );
  AOI22xp33_ASAP7_75t_SL U27565 ( .A1(n31391), .A2(rf_do_a[7]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__7_), .B2(n31392), .Y(n29901) );
  AOI22xp33_ASAP7_75t_SL U27566 ( .A1(u0_0_leon3x0_p0_divi[46]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[45]), .B2(n28367), .Y(n28332) );
  AOI22xp33_ASAP7_75t_SL U27567 ( .A1(n31391), .A2(rf_do_a[4]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__4_), .B2(n31392), .Y(n29498) );
  AOI22xp33_ASAP7_75t_SL U27568 ( .A1(n31391), .A2(rf_do_a[3]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__3_), .B2(n31392), .Y(n29494) );
  AOI22xp33_ASAP7_75t_SL U27569 ( .A1(u0_0_leon3x0_p0_divi[48]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[47]), .B2(n28367), .Y(n28326) );
  AOI22xp33_ASAP7_75t_SL U27570 ( .A1(u0_0_leon3x0_p0_divi[62]), .A2(n28367), 
        .B1(n28378), .B2(n28294), .Y(n28297) );
  INVxp33_ASAP7_75t_SL U27571 ( .A(n32380), .Y(n32639) );
  AOI22xp33_ASAP7_75t_SL U27572 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__16_), .A2(
        n30641), .B1(rf_do_b[16]), .B2(n30640), .Y(n28551) );
  AOI22xp33_ASAP7_75t_SL U27573 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__8_), .A2(
        n30641), .B1(rf_do_b[8]), .B2(n30640), .Y(n28750) );
  AOI21xp5_ASAP7_75t_SL U27574 ( .A1(n22429), .A2(u0_0_leon3x0_p0_muli[0]), 
        .B(n26748), .Y(n26749) );
  AOI22xp33_ASAP7_75t_SL U27575 ( .A1(n31391), .A2(rf_do_a[5]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__5_), .B2(n31392), .Y(n26323) );
  AOI22xp33_ASAP7_75t_SL U27576 ( .A1(n31201), .A2(uart1_r_RHOLD__30__1_), 
        .B1(uart1_r_RHOLD__5__1_), .B2(n31200), .Y(n27434) );
  AOI22xp33_ASAP7_75t_SL U27577 ( .A1(u0_0_leon3x0_p0_iu_r_W__RESULT__11_), 
        .A2(n31392), .B1(rf_do_a[11]), .B2(n31391), .Y(n29839) );
  AOI22xp33_ASAP7_75t_SL U27578 ( .A1(n31391), .A2(rf_do_a[24]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__24_), .B2(n31392), .Y(n26412) );
  INVxp67_ASAP7_75t_SL U27579 ( .A(n24985), .Y(n24967) );
  NAND2xp33_ASAP7_75t_SL U27580 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__16_), .B(
        n22429), .Y(n30330) );
  AOI22xp33_ASAP7_75t_SL U27581 ( .A1(n31391), .A2(rf_do_a[8]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__8_), .B2(n31392), .Y(n29929) );
  AOI21xp33_ASAP7_75t_SL U27582 ( .A1(n31824), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__6_), .B(n24680), .Y(n31825) );
  NAND2xp5_ASAP7_75t_SL U27583 ( .A(n29090), .B(n22378), .Y(n29091) );
  AOI22xp33_ASAP7_75t_SL U27584 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__15_), .A2(
        n30641), .B1(rf_do_b[15]), .B2(n30640), .Y(n28571) );
  NAND2xp33_ASAP7_75t_SL U27585 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__14_), .B(
        n22429), .Y(n30353) );
  NAND2xp33_ASAP7_75t_SL U27586 ( .A(n27273), .B(n22427), .Y(n27274) );
  AOI22xp33_ASAP7_75t_SL U27587 ( .A1(n31391), .A2(rf_do_a[6]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__6_), .B2(n31392), .Y(n26286) );
  NAND2xp33_ASAP7_75t_SL U27588 ( .A(n27233), .B(n22427), .Y(n27234) );
  NAND2xp33_ASAP7_75t_SL U27589 ( .A(u0_0_leon3x0_p0_muli[4]), .B(n22429), .Y(
        n30432) );
  AOI22xp33_ASAP7_75t_SL U27590 ( .A1(u0_0_leon3x0_p0_divi[41]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[40]), .B2(n28367), .Y(n28343) );
  NAND2xp33_ASAP7_75t_SL U27591 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__24_), .B(
        n22429), .Y(n30254) );
  NOR2x1_ASAP7_75t_SL U27592 ( .A(n24679), .B(n28291), .Y(n31676) );
  NAND2xp33_ASAP7_75t_SL U27593 ( .A(n25311), .B(n24672), .Y(n25310) );
  AOI22xp33_ASAP7_75t_SL U27594 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__24_), .A2(
        n30641), .B1(rf_do_b[24]), .B2(n30640), .Y(n28463) );
  AOI22xp33_ASAP7_75t_SL U27595 ( .A1(n31391), .A2(rf_do_a[9]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__9_), .B2(n31392), .Y(n27171) );
  AOI22xp33_ASAP7_75t_SL U27596 ( .A1(u0_0_leon3x0_p0_divi[40]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[39]), .B2(n28367), .Y(n28346) );
  AOI22xp33_ASAP7_75t_SL U27597 ( .A1(n31391), .A2(rf_do_a[22]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__22_), .B2(n31392), .Y(n29076) );
  NAND2xp5_ASAP7_75t_SL U27598 ( .A(n25321), .B(n24671), .Y(n25320) );
  AOI22xp33_ASAP7_75t_SL U27599 ( .A1(u0_0_leon3x0_p0_divi[39]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[38]), .B2(n28367), .Y(n28349) );
  NOR2xp33_ASAP7_75t_SL U27600 ( .A(n24427), .B(n28827), .Y(n29588) );
  AOI22xp33_ASAP7_75t_SL U27601 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__4_), .A2(
        n30641), .B1(rf_do_b[4]), .B2(n30640), .Y(n28862) );
  AOI22xp33_ASAP7_75t_SL U27602 ( .A1(rf_do_a[19]), .A2(n31391), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__19_), .B2(n31392), .Y(n25807) );
  OAI21xp33_ASAP7_75t_SRAM U27603 ( .A1(n26781), .A2(n18844), .B(n26780), .Y(
        n26782) );
  AOI22xp33_ASAP7_75t_SL U27604 ( .A1(u0_0_leon3x0_p0_divi[43]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[42]), .B2(n28367), .Y(n28339) );
  AOI22xp33_ASAP7_75t_SL U27605 ( .A1(u0_0_leon3x0_p0_divi[41]), .A2(n28367), 
        .B1(u0_0_leon3x0_p0_divi[42]), .B2(n28378), .Y(n28341) );
  AOI22xp33_ASAP7_75t_SL U27606 ( .A1(u0_0_leon3x0_p0_divi[36]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[35]), .B2(n28367), .Y(n28355) );
  AOI22xp33_ASAP7_75t_SL U27607 ( .A1(n31391), .A2(rf_do_a[12]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__12_), .B2(n31392), .Y(n29616) );
  AOI22xp33_ASAP7_75t_SL U27608 ( .A1(u0_0_leon3x0_p0_divi[35]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[34]), .B2(n28367), .Y(n28359) );
  AOI22xp33_ASAP7_75t_SL U27609 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__20_), .A2(
        n30641), .B1(rf_do_b[20]), .B2(n30640), .Y(n27008) );
  AOI22xp33_ASAP7_75t_SL U27610 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__19_), .A2(
        n30641), .B1(rf_do_b[19]), .B2(n30640), .Y(n28526) );
  AOI22xp33_ASAP7_75t_SL U27611 ( .A1(n31391), .A2(rf_do_a[13]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__13_), .B2(n31392), .Y(n27188) );
  NAND2xp33_ASAP7_75t_SL U27612 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__19_), .B(
        n22429), .Y(n30299) );
  NAND2xp33_ASAP7_75t_SL U27613 ( .A(n32632), .B(n22427), .Y(n27262) );
  AOI22xp33_ASAP7_75t_SL U27614 ( .A1(n31391), .A2(rf_do_a[10]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__10_), .B2(n31392), .Y(n27165) );
  NAND2xp33_ASAP7_75t_SL U27615 ( .A(n32654), .B(n22427), .Y(n28274) );
  AOI22xp33_ASAP7_75t_SL U27616 ( .A1(u0_0_leon3x0_p0_divi[38]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[37]), .B2(n28367), .Y(n28351) );
  AOI22xp33_ASAP7_75t_SL U27617 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__22_), .A2(
        n30641), .B1(rf_do_b[22]), .B2(n30640), .Y(n28508) );
  AOI22xp33_ASAP7_75t_SL U27618 ( .A1(n31391), .A2(rf_do_a[28]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__28_), .B2(n31392), .Y(n26946) );
  NAND2xp5_ASAP7_75t_SL U27619 ( .A(n26371), .B(n24669), .Y(n26372) );
  AOI22xp33_ASAP7_75t_SL U27620 ( .A1(n31391), .A2(rf_do_a[29]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__29_), .B2(n31392), .Y(n28280) );
  NAND2xp5_ASAP7_75t_SL U27621 ( .A(n25317), .B(n24671), .Y(n25316) );
  AOI21xp33_ASAP7_75t_SL U27622 ( .A1(n31824), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__3_), .B(n24680), .Y(n28565) );
  NAND2xp33_ASAP7_75t_SL U27623 ( .A(n28262), .B(n22427), .Y(n28263) );
  AOI22xp33_ASAP7_75t_SL U27624 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__5_), .A2(
        n30641), .B1(rf_do_b[5]), .B2(n30640), .Y(n28811) );
  NOR2xp33_ASAP7_75t_SL U27625 ( .A(n32131), .B(n26269), .Y(n28480) );
  AOI22xp33_ASAP7_75t_SL U27626 ( .A1(n31391), .A2(rf_do_a[20]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__20_), .B2(n31392), .Y(n27029) );
  NOR3xp33_ASAP7_75t_SL U27627 ( .A(n29347), .B(n31188), .C(n29346), .Y(n29348) );
  AOI22xp33_ASAP7_75t_SL U27628 ( .A1(n31391), .A2(rf_do_a[25]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__25_), .B2(n31392), .Y(n29784) );
  NAND2xp33_ASAP7_75t_SL U27629 ( .A(u0_0_leon3x0_p0_muli[5]), .B(n22429), .Y(
        n30420) );
  AND2x2_ASAP7_75t_SL U27630 ( .A(n27224), .B(n22427), .Y(n27225) );
  AOI22xp33_ASAP7_75t_SL U27631 ( .A1(n31391), .A2(rf_do_a[14]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__14_), .B2(n31392), .Y(n27220) );
  INVx8_ASAP7_75t_SL U27632 ( .A(n23961), .Y(n22394) );
  NAND2xp33_ASAP7_75t_SL U27633 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__29_), .B(
        n22429), .Y(n30227) );
  AOI21xp33_ASAP7_75t_SL U27634 ( .A1(n31824), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__0_), .B(n24680), .Y(n29819) );
  AND2x2_ASAP7_75t_SL U27635 ( .A(n28277), .B(n22427), .Y(n28278) );
  INVxp67_ASAP7_75t_SL U27636 ( .A(n26394), .Y(n29585) );
  NOR2xp33_ASAP7_75t_SL U27637 ( .A(apbi[9]), .B(n24695), .Y(n29258) );
  NAND2xp33_ASAP7_75t_SL U27638 ( .A(n27181), .B(n22427), .Y(n27182) );
  NOR2x1p5_ASAP7_75t_SL U27639 ( .A(n23153), .B(n22273), .Y(n23155) );
  AOI22xp33_ASAP7_75t_SL U27640 ( .A1(rf_do_a[2]), .A2(n31391), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__2_), .B2(n31392), .Y(n30466) );
  NAND2xp33_ASAP7_75t_SL U27641 ( .A(n24681), .B(n30958), .Y(n30959) );
  AOI22xp33_ASAP7_75t_SL U27642 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__12_), .A2(
        n30641), .B1(rf_do_b[12]), .B2(n30640), .Y(n28650) );
  AOI22xp33_ASAP7_75t_SL U27643 ( .A1(n31391), .A2(rf_do_a[26]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__26_), .B2(n31392), .Y(n29797) );
  AOI22xp33_ASAP7_75t_SL U27644 ( .A1(n31391), .A2(rf_do_a[31]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__31_), .B2(n31392), .Y(n25211) );
  INVx1_ASAP7_75t_SL U27645 ( .A(n30207), .Y(n31001) );
  AOI22xp33_ASAP7_75t_SL U27646 ( .A1(timer0_N91), .A2(n24416), .B1(timer0_N90), .B2(n22430), .Y(timer0_res_1_) );
  AOI22xp33_ASAP7_75t_SL U27647 ( .A1(n31391), .A2(rf_do_a[1]), .B1(
        u0_0_leon3x0_p0_iu_r_W__RESULT__1_), .B2(n31392), .Y(n31338) );
  NOR2xp33_ASAP7_75t_SL U27648 ( .A(n25082), .B(n18997), .Y(n25084) );
  NAND2xp33_ASAP7_75t_SL U27649 ( .A(n28266), .B(n22427), .Y(n28267) );
  INVxp67_ASAP7_75t_SL U27650 ( .A(DP_OP_1196_128_7433_n70), .Y(
        DP_OP_1196_128_7433_n361) );
  AOI22xp33_ASAP7_75t_SL U27651 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__7_), .A2(
        n30641), .B1(rf_do_b[7]), .B2(n30640), .Y(n28795) );
  NAND2xp33_ASAP7_75t_SL U27652 ( .A(n27229), .B(n22427), .Y(n27230) );
  AOI22xp33_ASAP7_75t_SL U27653 ( .A1(u0_0_leon3x0_p0_divi[51]), .A2(n28367), 
        .B1(u0_0_leon3x0_p0_divi[52]), .B2(n28378), .Y(n28318) );
  AOI22xp33_ASAP7_75t_SL U27654 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__9_), .A2(
        n30641), .B1(rf_do_b[9]), .B2(n30640), .Y(n27128) );
  AOI22xp33_ASAP7_75t_SL U27655 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__13_), .A2(
        n30641), .B1(rf_do_b[13]), .B2(n30640), .Y(n28605) );
  AOI22xp33_ASAP7_75t_SL U27656 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__2_), .A2(
        n30641), .B1(rf_do_b[2]), .B2(n30640), .Y(n28951) );
  NAND2xp33_ASAP7_75t_SL U27657 ( .A(n27231), .B(n22427), .Y(n27232) );
  NAND2xp33_ASAP7_75t_SL U27658 ( .A(n28264), .B(n22427), .Y(n28265) );
  AOI21xp33_ASAP7_75t_SL U27659 ( .A1(n32860), .A2(ahbso_0__HRDATA__10_), .B(
        n22433), .Y(n32862) );
  AOI22xp33_ASAP7_75t_SL U27660 ( .A1(u0_0_leon3x0_p0_divi[54]), .A2(n28378), 
        .B1(u0_0_leon3x0_p0_divi[53]), .B2(n28367), .Y(n28315) );
  INVx1_ASAP7_75t_SL U27661 ( .A(n31868), .Y(n30645) );
  NAND2xp33_ASAP7_75t_SL U27662 ( .A(n24634), .B(n28482), .Y(n27066) );
  NAND2xp5_ASAP7_75t_SL U27663 ( .A(n24634), .B(n29144), .Y(n28941) );
  NAND2xp33_ASAP7_75t_SRAM U27664 ( .A(n32074), .B(n25565), .Y(n25566) );
  INVx1_ASAP7_75t_SL U27665 ( .A(n24681), .Y(n24670) );
  NAND3xp33_ASAP7_75t_SRAM U27666 ( .A(n22431), .B(n29111), .C(n29110), .Y(
        n29113) );
  A2O1A1Ixp33_ASAP7_75t_SL U27667 ( .A1(n30118), .A2(n30117), .B(n30116), .C(
        n31981), .Y(n30123) );
  AOI21xp5_ASAP7_75t_SL U27668 ( .A1(n25231), .A2(n25230), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__LD_), .Y(n24864) );
  AOI22xp33_ASAP7_75t_SL U27669 ( .A1(uart1_r_RHOLD__14__1_), .A2(n31203), 
        .B1(n31202), .B2(uart1_r_RHOLD__12__1_), .Y(n27436) );
  OAI22xp5_ASAP7_75t_SL U27670 ( .A1(n26747), .A2(n24638), .B1(n26746), .B2(
        n31404), .Y(n26748) );
  NAND2xp33_ASAP7_75t_SRAM U27671 ( .A(n3730), .B(n26791), .Y(n25606) );
  NAND2xp33_ASAP7_75t_SL U27672 ( .A(ahbso_1__HRDATA__24_), .B(n30002), .Y(
        n26506) );
  AOI22xp33_ASAP7_75t_SL U27673 ( .A1(ahbso_0__HRDATA__25_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__25_), .Y(n31378) );
  AOI22xp33_ASAP7_75t_SL U27674 ( .A1(ahbso_0__HRDATA__3_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__3_), .Y(n32306) );
  AOI22xp33_ASAP7_75t_SL U27675 ( .A1(ahbso_0__HRDATA__2_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__2_), .Y(n32303) );
  AOI22xp33_ASAP7_75t_SL U27676 ( .A1(ahbso_0__HRDATA__27_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__27_), .Y(n30904) );
  NAND2xp33_ASAP7_75t_SL U27677 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__18_), 
        .B(n22376), .Y(n25711) );
  AOI22xp33_ASAP7_75t_SL U27678 ( .A1(ahbso_0__HRDATA__28_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__28_), .Y(n31509) );
  AOI22xp33_ASAP7_75t_SL U27679 ( .A1(ahbso_0__HRDATA__0_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__0_), .Y(n32297) );
  NAND2xp33_ASAP7_75t_SL U27680 ( .A(ahbso_1__HRDATA__12_), .B(n30002), .Y(
        n25419) );
  OAI21xp33_ASAP7_75t_SL U27681 ( .A1(n29963), .A2(n31188), .B(n29962), .Y(
        n29970) );
  OAI22xp33_ASAP7_75t_SL U27682 ( .A1(n28183), .A2(n31188), .B1(n24695), .B2(
        n30774), .Y(uart1_v_RXCLK__2_) );
  INVx1_ASAP7_75t_SL U27683 ( .A(n28821), .Y(n28827) );
  NAND2xp33_ASAP7_75t_SL U27684 ( .A(n25634), .B(n25941), .Y(n25954) );
  AOI22xp33_ASAP7_75t_SL U27685 ( .A1(ahbso_0__HRDATA__18_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__18_), .Y(n32367) );
  AOI22xp33_ASAP7_75t_SL U27686 ( .A1(ahbso_0__HRDATA__19_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__19_), .Y(n32371) );
  NAND2xp33_ASAP7_75t_SL U27687 ( .A(ahbso_1__HRDATA__6_), .B(n30002), .Y(
        n25852) );
  AOI22xp33_ASAP7_75t_SL U27688 ( .A1(ahbso_0__HRDATA__20_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__20_), .Y(n32377) );
  NOR2xp33_ASAP7_75t_SL U27689 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .B(
        n23933), .Y(n30614) );
  AOI22xp33_ASAP7_75t_SL U27690 ( .A1(ahbso_0__HRDATA__21_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__21_), .Y(n32380) );
  INVx1_ASAP7_75t_SL U27691 ( .A(n27460), .Y(n30555) );
  NAND2xp33_ASAP7_75t_SL U27692 ( .A(ahbso_1__HRDATA__5_), .B(n30002), .Y(
        n30003) );
  AOI22xp33_ASAP7_75t_SL U27693 ( .A1(ahbso_0__HRDATA__22_), .A2(n29999), .B1(
        n30002), .B2(ahbso_1__HRDATA__22_), .Y(n32382) );
  NOR2x1_ASAP7_75t_SL U27694 ( .A(n25734), .B(n25737), .Y(n30723) );
  NAND2xp33_ASAP7_75t_SL U27695 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__8_), .B(
        n22376), .Y(n25519) );
  NAND2xp33_ASAP7_75t_SRAM U27696 ( .A(n26804), .B(n31862), .Y(n26780) );
  NOR2x1_ASAP7_75t_SL U27697 ( .A(n25735), .B(n25737), .Y(n30726) );
  NOR2x1_ASAP7_75t_SL U27698 ( .A(n25738), .B(n25737), .Y(n30725) );
  OAI21x1_ASAP7_75t_SL U27699 ( .A1(n25732), .A2(n25737), .B(n32153), .Y(
        n30722) );
  OAI21xp5_ASAP7_75t_SL U27700 ( .A1(n4774), .A2(n30694), .B(n25373), .Y(
        n25374) );
  OAI22xp5_ASAP7_75t_SL U27701 ( .A1(n24698), .A2(n24697), .B1(n24474), .B2(
        n24697), .Y(n24699) );
  NAND2xp5_ASAP7_75t_SL U27702 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__3_), 
        .B(n31554), .Y(n31553) );
  AOI31xp33_ASAP7_75t_SL U27703 ( .A1(irqctrl0_r_ILEVEL__2_), .A2(
        irqctrl0_r_IMASK__0__2_), .A3(n29417), .B(n29447), .Y(n29444) );
  INVx1_ASAP7_75t_SL U27704 ( .A(n24856), .Y(n24874) );
  NAND2xp5_ASAP7_75t_SL U27705 ( .A(irqctrl0_r_ILEVEL__4_), .B(n29421), .Y(
        n29448) );
  INVxp33_ASAP7_75t_SL U27706 ( .A(n29456), .Y(n29459) );
  INVxp67_ASAP7_75t_SL U27707 ( .A(n29945), .Y(n28038) );
  NAND2xp33_ASAP7_75t_SL U27708 ( .A(n29147), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__WY_), .Y(n23933) );
  INVxp67_ASAP7_75t_SL U27709 ( .A(n25998), .Y(n25999) );
  NAND2xp33_ASAP7_75t_SL U27710 ( .A(n30115), .B(n26353), .Y(n26355) );
  INVx1_ASAP7_75t_SL U27711 ( .A(n27380), .Y(n27388) );
  INVxp33_ASAP7_75t_SL U27712 ( .A(n25379), .Y(n25380) );
  INVx1_ASAP7_75t_SL U27713 ( .A(n25366), .Y(n30687) );
  INVx2_ASAP7_75t_SL U27714 ( .A(n32564), .Y(n32660) );
  NOR2x1_ASAP7_75t_SL U27715 ( .A(n32012), .B(n28292), .Y(n28367) );
  NOR2x1p5_ASAP7_75t_SL U27716 ( .A(n22919), .B(n28292), .Y(n28378) );
  NAND2xp5_ASAP7_75t_SL U27717 ( .A(n27411), .B(n27997), .Y(n27986) );
  NOR2x1_ASAP7_75t_SL U27718 ( .A(n26482), .B(n28830), .Y(n29144) );
  INVx1_ASAP7_75t_SL U27719 ( .A(n28894), .Y(n30625) );
  INVxp33_ASAP7_75t_SL U27720 ( .A(n31420), .Y(n31654) );
  OR2x2_ASAP7_75t_SL U27721 ( .A(n18864), .B(n4614), .Y(timer0_N65) );
  OAI21xp5_ASAP7_75t_SL U27722 ( .A1(address[0]), .A2(address[1]), .B(n32886), 
        .Y(n32913) );
  INVxp67_ASAP7_75t_SL U27723 ( .A(n30195), .Y(n25582) );
  INVx1_ASAP7_75t_SL U27724 ( .A(n30446), .Y(n30453) );
  NOR2x1_ASAP7_75t_SL U27725 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__0_), .B(
        n26730), .Y(n30641) );
  INVxp67_ASAP7_75t_SL U27726 ( .A(n25488), .Y(n25624) );
  INVx1_ASAP7_75t_SL U27727 ( .A(n28830), .Y(n29146) );
  NAND4xp25_ASAP7_75t_SRAM U27728 ( .A(n25691), .B(n25690), .C(n25689), .D(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__26_), .Y(n25696) );
  NAND2xp33_ASAP7_75t_SL U27729 ( .A(n25970), .B(n27536), .Y(n27535) );
  NAND2xp5_ASAP7_75t_SL U27730 ( .A(n4371), .B(n25952), .Y(n1637) );
  NOR2xp33_ASAP7_75t_SL U27731 ( .A(n31848), .B(n31529), .Y(n25940) );
  NAND3xp33_ASAP7_75t_SRAM U27732 ( .A(n32730), .B(n3055), .C(
        u0_0_leon3x0_p0_dci[5]), .Y(n32195) );
  OR2x2_ASAP7_75t_SL U27733 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__ANNUL_), .B(
        n25152), .Y(n24425) );
  NAND2xp33_ASAP7_75t_SL U27734 ( .A(sr1_r_SRHSEL_), .B(n32832), .Y(n31749) );
  INVxp33_ASAP7_75t_SRAM U27735 ( .A(n32710), .Y(n31713) );
  NOR2xp33_ASAP7_75t_SRAM U27736 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__21_), 
        .B(n29708), .Y(n25357) );
  NOR2xp33_ASAP7_75t_SL U27737 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_), 
        .B(n31943), .Y(n24921) );
  INVxp33_ASAP7_75t_SL U27738 ( .A(n32832), .Y(n31739) );
  INVxp33_ASAP7_75t_SL U27739 ( .A(n28167), .Y(n28172) );
  INVxp67_ASAP7_75t_SL U27740 ( .A(DP_OP_1196_128_7433_n147), .Y(
        DP_OP_1196_128_7433_n368) );
  NAND2xp33_ASAP7_75t_SL U27741 ( .A(n29632), .B(n29631), .Y(n29661) );
  NOR2xp67_ASAP7_75t_SL U27742 ( .A(n3704), .B(n25607), .Y(n33054) );
  INVxp67_ASAP7_75t_SL U27743 ( .A(n29432), .Y(n29413) );
  INVxp67_ASAP7_75t_SL U27744 ( .A(n24979), .Y(n31565) );
  INVxp67_ASAP7_75t_SL U27745 ( .A(n28045), .Y(n28047) );
  INVx1_ASAP7_75t_SL U27746 ( .A(DP_OP_1196_128_7433_n167), .Y(
        DP_OP_1196_128_7433_n370) );
  INVx1_ASAP7_75t_SL U27747 ( .A(DP_OP_1196_128_7433_n221), .Y(
        DP_OP_1196_128_7433_n374) );
  INVx1_ASAP7_75t_SL U27748 ( .A(DP_OP_1196_128_7433_n251), .Y(
        DP_OP_1196_128_7433_n376) );
  NAND2xp5_ASAP7_75t_SL U27749 ( .A(n22919), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_), .Y(n32131) );
  INVx1_ASAP7_75t_SL U27750 ( .A(DP_OP_1196_128_7433_n128), .Y(
        DP_OP_1196_128_7433_n367) );
  INVxp33_ASAP7_75t_SL U27751 ( .A(n29000), .Y(n29001) );
  NAND2x1_ASAP7_75t_SL U27752 ( .A(n31658), .B(n28291), .Y(n31660) );
  OA21x2_ASAP7_75t_SL U27753 ( .A1(n24879), .A2(n24878), .B(n18820), .Y(n24880) );
  NOR2x1_ASAP7_75t_SL U27754 ( .A(n4391), .B(n32037), .Y(n30002) );
  INVx1_ASAP7_75t_SL U27755 ( .A(DP_OP_1196_128_7433_n307), .Y(
        DP_OP_1196_128_7433_n380) );
  NOR2xp33_ASAP7_75t_SRAM U27756 ( .A(n4316), .B(n32236), .Y(n24956) );
  NAND2xp33_ASAP7_75t_SL U27757 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .B(
        n29147), .Y(n28481) );
  O2A1O1Ixp5_ASAP7_75t_SL U27758 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), 
        .A2(n29166), .B(n29165), .C(n30667), .Y(n29170) );
  INVx1_ASAP7_75t_SL U27759 ( .A(DP_OP_1196_128_7433_n195), .Y(
        DP_OP_1196_128_7433_n372) );
  INVxp67_ASAP7_75t_SL U27760 ( .A(u0_0_leon3x0_p0_divi[60]), .Y(n30230) );
  INVx1_ASAP7_75t_SL U27761 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__26_), .Y(
        n30242) );
  INVx1_ASAP7_75t_SL U27762 ( .A(n2389), .Y(n25990) );
  INVxp33_ASAP7_75t_SL U27763 ( .A(n1741), .Y(n29752) );
  INVx1_ASAP7_75t_SL U27764 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__27_), .Y(
        n30239) );
  INVxp67_ASAP7_75t_SL U27765 ( .A(u0_0_leon3x0_p0_iu_r_E__CTRL__ANNUL_), .Y(
        n32069) );
  INVxp67_ASAP7_75t_SL U27766 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__7_), .Y(
        n32160) );
  INVx1_ASAP7_75t_SL U27767 ( .A(apbi[2]), .Y(n29568) );
  INVx2_ASAP7_75t_SL U27768 ( .A(uart1_r_RSHIFT__2_), .Y(n29555) );
  INVx1_ASAP7_75t_SL U27769 ( .A(u0_0_leon3x0_p0_iu_r_A__CTRL__WICC_), .Y(
        n24719) );
  NAND2xp33_ASAP7_75t_SL U27770 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_OVERRUN_), 
        .B(u0_0_leon3x0_p0_ici[29]), .Y(n32126) );
  INVxp67_ASAP7_75t_SL U27771 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_ASI__0_), 
        .Y(n32598) );
  INVx1_ASAP7_75t_SL U27772 ( .A(n2235), .Y(n29412) );
  INVx1_ASAP7_75t_SL U27773 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__21_), .Y(
        n30277) );
  OAI21xp5_ASAP7_75t_SL U27774 ( .A1(irqctrl0_r_IPEND__10_), .A2(
        irqctrl0_r_IFORCE__0__10_), .B(irqctrl0_r_IMASK__0__10_), .Y(n29432)
         );
  INVxp67_ASAP7_75t_SL U27775 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__0_), .Y(
        n25074) );
  INVxp33_ASAP7_75t_SL U27776 ( .A(n2233), .Y(n28125) );
  INVx1_ASAP7_75t_SL U27777 ( .A(apbi[1]), .Y(n27493) );
  INVx1_ASAP7_75t_SL U27778 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__4_), .Y(
        n30705) );
  INVx1_ASAP7_75t_SL U27779 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__17_), .Y(
        n30317) );
  INVx1_ASAP7_75t_SL U27780 ( .A(apbi[27]), .Y(n30894) );
  INVx1_ASAP7_75t_SL U27781 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__16_), .Y(
        n30328) );
  INVx1_ASAP7_75t_SL U27782 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__18_), .Y(
        n30306) );
  NAND2xp5_ASAP7_75t_SL U27783 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__20_), 
        .B(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), .Y(n30156) );
  INVxp67_ASAP7_75t_SL U27784 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__26_), 
        .Y(n25553) );
  INVx1_ASAP7_75t_SL U27785 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__19_), .Y(
        n30297) );
  NAND3xp33_ASAP7_75t_SL U27786 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__30_), 
        .B(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__31_), .C(
        u0_0_leon3x0_p0_iu_v_X__CTRL__PV_), .Y(n25392) );
  INVxp67_ASAP7_75t_SL U27787 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_), 
        .Y(n25549) );
  NAND2xp5_ASAP7_75t_SL U27788 ( .A(n3071), .B(n3132), .Y(n24979) );
  INVxp67_ASAP7_75t_SL U27789 ( .A(u0_0_leon3x0_p0_iu_r_X__NPC__1_), .Y(n25736) );
  INVx2_ASAP7_75t_SL U27790 ( .A(uart1_r_RSHIFT__6_), .Y(n31182) );
  INVxp67_ASAP7_75t_SL U27791 ( .A(u0_0_leon3x0_p0_iu_r_D__ANNUL_), .Y(n24855)
         );
  INVx1_ASAP7_75t_SL U27792 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .Y(
        n24879) );
  INVx2_ASAP7_75t_SL U27793 ( .A(uart1_r_RSHIFT__7_), .Y(n30865) );
  INVxp67_ASAP7_75t_SL U27794 ( .A(uart1_r_TRADDR__4_), .Y(n27391) );
  INVx2_ASAP7_75t_SL U27795 ( .A(uart1_r_RSHIFT__1_), .Y(n26126) );
  INVxp67_ASAP7_75t_SL U27796 ( .A(u0_0_leon3x0_p0_iu_r_X__NPC__0_), .Y(n25733) );
  INVx2_ASAP7_75t_SL U27797 ( .A(uart1_r_RSHIFT__4_), .Y(n30771) );
  INVxp33_ASAP7_75t_SL U27798 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_), 
        .Y(n25359) );
  INVx1_ASAP7_75t_SL U27799 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__24_), .Y(
        n30252) );
  OAI21xp33_ASAP7_75t_SL U27800 ( .A1(irqctrl0_r_IPEND__3_), .A2(
        irqctrl0_r_IFORCE__0__3_), .B(irqctrl0_r_IMASK__0__3_), .Y(n29415) );
  BUFx3_ASAP7_75t_SL U27801 ( .A(u0_0_leon3x0_p0_muli[9]), .Y(n22919) );
  INVx2_ASAP7_75t_SL U27802 ( .A(uart1_r_RSHIFT__5_), .Y(n30062) );
  INVx2_ASAP7_75t_SL U27803 ( .A(uart1_r_RSHIFT__3_), .Y(n28224) );
  INVxp67_ASAP7_75t_SL U27804 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[14]), .Y(n26614)
         );
  NAND2xp5_ASAP7_75t_SL U27805 ( .A(apbi[46]), .B(apb0_r_PSEL_), .Y(n25986) );
  INVxp33_ASAP7_75t_SL U27806 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__30_), .Y(
        n30598) );
  INVxp67_ASAP7_75t_SL U27807 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__25_), .Y(
        n28425) );
  INVx1_ASAP7_75t_SL U27808 ( .A(n2811), .Y(n28379) );
  INVxp67_ASAP7_75t_SL U27809 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__30_), .Y(
        n30213) );
  INVxp67_ASAP7_75t_SL U27810 ( .A(n3068), .Y(n31448) );
  INVxp67_ASAP7_75t_SL U27811 ( .A(u0_0_leon3x0_p0_iu_r_E__CTRL__WREG_), .Y(
        n24755) );
  INVx1_ASAP7_75t_SL U27812 ( .A(u0_0_leon3x0_p0_divo[3]), .Y(n28903) );
  INVx1_ASAP7_75t_SL U27813 ( .A(sr1_sdi_HWRITE_), .Y(n31708) );
  INVxp33_ASAP7_75t_SL U27814 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__11_), .Y(
        n29841) );
  INVxp67_ASAP7_75t_SL U27815 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__1_), .Y(
        n25948) );
  INVxp33_ASAP7_75t_SL U27816 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__30_), 
        .Y(n31943) );
  INVxp67_ASAP7_75t_SL U27817 ( .A(sr1_r_MCFG2__RAMBANKSZ__3_), .Y(n32762) );
  NOR2xp33_ASAP7_75t_SL U27818 ( .A(uart1_r_RXSTATE__0_), .B(
        uart1_r_RXSTATE__1_), .Y(n27536) );
  INVxp67_ASAP7_75t_SL U27819 ( .A(u0_0_leon3x0_p0_divi[57]), .Y(n30245) );
  INVx1_ASAP7_75t_SL U27820 ( .A(u0_0_leon3x0_p0_muli[9]), .Y(n32012) );
  INVx1_ASAP7_75t_SL U27821 ( .A(u0_0_leon3x0_p0_div0_r_CNT__2_), .Y(n24884)
         );
  INVx1_ASAP7_75t_SL U27822 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__22_), .Y(n22599)
         );
  INVxp67_ASAP7_75t_SL U27823 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[60]), .Y(n31787)
         );
  INVxp67_ASAP7_75t_SL U27824 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__2_), .Y(
        n24819) );
  INVxp67_ASAP7_75t_SL U27825 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__3_), .Y(
        n24818) );
  INVxp67_ASAP7_75t_SL U27826 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[61]), .Y(n31772)
         );
  INVxp33_ASAP7_75t_SL U27827 ( .A(n4316), .Y(n32253) );
  INVx1_ASAP7_75t_SL U27828 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__28_), .Y(n23833)
         );
  INVxp67_ASAP7_75t_SL U27829 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__1_), 
        .Y(n32142) );
  INVxp67_ASAP7_75t_SL U27830 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[59]), .Y(n31780)
         );
  INVx1_ASAP7_75t_SL U27831 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__6_), .Y(
        n24829) );
  OAI21xp5_ASAP7_75t_SL U27832 ( .A1(n24646), .A2(n23735), .B(n25320), .Y(
        n4187) );
  OAI21xp5_ASAP7_75t_SL U27833 ( .A1(n24646), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N28), .B(n28450), .Y(n4259) );
  OAI21xp5_ASAP7_75t_SL U27834 ( .A1(n24646), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N26), .B(n29091), .Y(n4263) );
  OAI211xp5_ASAP7_75t_SRAM U27835 ( .A1(n2962), .A2(n32443), .B(n32442), .C(
        n32441), .Y(dc_address[1]) );
  OAI211xp5_ASAP7_75t_SRAM U27836 ( .A1(n2963), .A2(n32443), .B(n32440), .C(
        n32439), .Y(dc_address[0]) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U27837 ( .A1(n32284), .A2(n32283), .B(n32282), .C(
        n33067), .Y(dc_wren) );
  INVxp67_ASAP7_75t_SL U27838 ( .A(n28113), .Y(n28114) );
  AOI21xp33_ASAP7_75t_SL U27839 ( .A1(n31845), .A2(timer0_res_12_), .B(n26608), 
        .Y(n26609) );
  NAND2xp33_ASAP7_75t_SL U27840 ( .A(n24694), .B(n30739), .Y(n2346) );
  AOI21xp33_ASAP7_75t_SL U27841 ( .A1(n31845), .A2(timer0_res_6_), .B(n26631), 
        .Y(n26632) );
  OAI21xp33_ASAP7_75t_SL U27842 ( .A1(n18877), .A2(n32841), .B(n28106), .Y(
        n28107) );
  OAI21xp33_ASAP7_75t_SL U27843 ( .A1(n18877), .A2(n32857), .B(n29940), .Y(
        n29941) );
  AOI21xp33_ASAP7_75t_SL U27844 ( .A1(n31845), .A2(timer0_res_14_), .B(n26595), 
        .Y(n26596) );
  OAI21xp33_ASAP7_75t_SL U27845 ( .A1(n18877), .A2(n32853), .B(n25861), .Y(
        n25862) );
  OAI21xp33_ASAP7_75t_SL U27846 ( .A1(n18877), .A2(n32849), .B(n25875), .Y(
        n25876) );
  AOI21xp33_ASAP7_75t_SL U27847 ( .A1(n31845), .A2(timer0_res_5_), .B(n26634), 
        .Y(n26635) );
  AOI21xp33_ASAP7_75t_SL U27848 ( .A1(n31845), .A2(timer0_res_7_), .B(n26628), 
        .Y(n26629) );
  XNOR2xp5_ASAP7_75t_SL U27849 ( .A(mult_x_1196_n266), .B(n23902), .Y(n23895)
         );
  AOI21xp33_ASAP7_75t_SL U27850 ( .A1(n31845), .A2(timer0_res_13_), .B(n26605), 
        .Y(n26606) );
  AOI21xp33_ASAP7_75t_SL U27851 ( .A1(n31845), .A2(timer0_res_4_), .B(n26637), 
        .Y(n26638) );
  INVxp67_ASAP7_75t_SL U27852 ( .A(n25594), .Y(n25595) );
  OAI21xp33_ASAP7_75t_SL U27853 ( .A1(n30189), .A2(n30188), .B(n30187), .Y(
        u0_0_leon3x0_p0_c0mmu_dcache0_v_FLUSH_) );
  INVx1_ASAP7_75t_SL U27854 ( .A(mult_x_1196_n455), .Y(mult_x_1196_n453) );
  NAND2xp5_ASAP7_75t_SL U27855 ( .A(n31580), .B(n31596), .Y(n31588) );
  OAI211xp5_ASAP7_75t_SRAM U27856 ( .A1(n32392), .A2(n32232), .B(n32221), .C(
        n32220), .Y(dt_data[20]) );
  OAI211xp5_ASAP7_75t_SRAM U27857 ( .A1(n32395), .A2(n32232), .B(n32223), .C(
        n32222), .Y(dt_data[21]) );
  OAI211xp5_ASAP7_75t_SRAM U27858 ( .A1(n32401), .A2(n32232), .B(n32225), .C(
        n32224), .Y(dt_data[22]) );
  OAI211xp5_ASAP7_75t_SRAM U27859 ( .A1(n32402), .A2(n32232), .B(n32227), .C(
        n32226), .Y(dt_data[23]) );
  OAI21xp33_ASAP7_75t_SL U27860 ( .A1(n3063), .A2(n22380), .B(n24684), .Y(
        n24555) );
  OAI22xp33_ASAP7_75t_SL U27861 ( .A1(n31766), .A2(n24645), .B1(n32640), .B2(
        n32729), .Y(n31767) );
  OAI22xp33_ASAP7_75t_SL U27862 ( .A1(n32636), .A2(n31632), .B1(n32375), .B2(
        n31631), .Y(n26541) );
  OAI22xp33_ASAP7_75t_SL U27863 ( .A1(n32648), .A2(n31632), .B1(n32395), .B2(
        n31631), .Y(n31366) );
  OAI22xp33_ASAP7_75t_SL U27864 ( .A1(n32644), .A2(n31632), .B1(n32387), .B2(
        n31631), .Y(n26528) );
  OAI22xp33_ASAP7_75t_SL U27865 ( .A1(n32604), .A2(n31632), .B1(n32305), .B2(
        n31631), .Y(n29508) );
  OAI22xp33_ASAP7_75t_SL U27866 ( .A1(n32614), .A2(n31632), .B1(n32320), .B2(
        n31631), .Y(n25524) );
  OAI22xp33_ASAP7_75t_SL U27867 ( .A1(n32650), .A2(n31632), .B1(n32401), .B2(
        n31631), .Y(n26496) );
  INVxp67_ASAP7_75t_SL U27868 ( .A(n22553), .Y(mult_x_1196_n568) );
  OAI22xp33_ASAP7_75t_SL U27869 ( .A1(n32602), .A2(n31632), .B1(n32302), .B2(
        n31631), .Y(n29567) );
  OAI22xp33_ASAP7_75t_SL U27870 ( .A1(n32640), .A2(n31632), .B1(n32379), .B2(
        n31631), .Y(n29293) );
  OAI22xp33_ASAP7_75t_SL U27871 ( .A1(n32626), .A2(n31632), .B1(n30556), .B2(
        n31631), .Y(n25633) );
  OAI22xp33_ASAP7_75t_SL U27872 ( .A1(n32734), .A2(n31632), .B1(n32300), .B2(
        n31631), .Y(n27492) );
  OAI22xp33_ASAP7_75t_SL U27873 ( .A1(n31780), .A2(n24645), .B1(n32729), .B2(
        n32650), .Y(n31781) );
  OAI22xp33_ASAP7_75t_SL U27874 ( .A1(n32620), .A2(n31632), .B1(n32332), .B2(
        n31631), .Y(n28137) );
  OAI22xp33_ASAP7_75t_SL U27875 ( .A1(n32616), .A2(n31632), .B1(n32325), .B2(
        n31631), .Y(n30133) );
  OAI22xp33_ASAP7_75t_SL U27876 ( .A1(n31787), .A2(n24645), .B1(n32729), .B2(
        n32652), .Y(n31788) );
  OAI22xp33_ASAP7_75t_SL U27877 ( .A1(n32646), .A2(n31632), .B1(n32392), .B2(
        n31631), .Y(n26516) );
  OAI22xp33_ASAP7_75t_SL U27878 ( .A1(n32658), .A2(n31632), .B1(n32418), .B2(
        n31631), .Y(n25647) );
  OAI22xp33_ASAP7_75t_SL U27879 ( .A1(n31688), .A2(n24645), .B1(n32729), .B2(
        n32661), .Y(n31689) );
  OAI22xp33_ASAP7_75t_SL U27880 ( .A1(n31772), .A2(n24645), .B1(n32729), .B2(
        n32654), .Y(n31773) );
  AOI21xp33_ASAP7_75t_SL U27881 ( .A1(n22553), .A2(mult_x_1196_n801), .B(
        mult_x_1196_n563), .Y(mult_x_1196_n561) );
  OAI22xp33_ASAP7_75t_SL U27882 ( .A1(n31691), .A2(n24645), .B1(n32656), .B2(
        n32729), .Y(n31692) );
  OAI22xp33_ASAP7_75t_SL U27883 ( .A1(n32642), .A2(n31632), .B1(n32383), .B2(
        n31631), .Y(n31636) );
  OAI22xp33_ASAP7_75t_SL U27884 ( .A1(n32608), .A2(n31632), .B1(n32310), .B2(
        n31631), .Y(n30028) );
  OAI22xp33_ASAP7_75t_SL U27885 ( .A1(n32622), .A2(n31632), .B1(n29847), .B2(
        n31631), .Y(n29850) );
  OAI22xp33_ASAP7_75t_SL U27886 ( .A1(n32652), .A2(n31632), .B1(n32402), .B2(
        n31631), .Y(n30892) );
  OAI22xp33_ASAP7_75t_SL U27887 ( .A1(n32737), .A2(n24645), .B1(n32735), .B2(
        n32734), .Y(n32738) );
  NAND2xp5_ASAP7_75t_SL U27888 ( .A(n31550), .B(n32545), .Y(n3058) );
  OAI22xp33_ASAP7_75t_SL U27889 ( .A1(n32661), .A2(n31632), .B1(n32432), .B2(
        n31631), .Y(n26460) );
  AOI22xp33_ASAP7_75t_SL U27890 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[3]), .A2(
        n31314), .B1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__3_), .B2(n31313), .Y(
        n30917) );
  NAND2xp5_ASAP7_75t_SL U27891 ( .A(n31552), .B(n32545), .Y(n3059) );
  OAI22xp33_ASAP7_75t_SL U27892 ( .A1(n30511), .A2(n24645), .B1(n32626), .B2(
        n32729), .Y(n30512) );
  OAI21xp33_ASAP7_75t_SL U27893 ( .A1(n31445), .A2(n32272), .B(n24684), .Y(
        n3042) );
  OAI22xp33_ASAP7_75t_SL U27894 ( .A1(n32630), .A2(n31632), .B1(n32360), .B2(
        n31631), .Y(n26450) );
  OAI22xp33_ASAP7_75t_SL U27895 ( .A1(n32624), .A2(n31632), .B1(n29993), .B2(
        n31631), .Y(n26603) );
  OAI22xp33_ASAP7_75t_SL U27896 ( .A1(n32634), .A2(n31632), .B1(n32366), .B2(
        n31631), .Y(n25845) );
  OAI22xp33_ASAP7_75t_SL U27897 ( .A1(n32628), .A2(n31632), .B1(n31031), .B2(
        n31631), .Y(n26591) );
  OAI22xp33_ASAP7_75t_SL U27898 ( .A1(n32632), .A2(n31632), .B1(n32365), .B2(
        n31631), .Y(n27289) );
  OAI22xp33_ASAP7_75t_SL U27899 ( .A1(n31835), .A2(n24645), .B1(n32634), .B2(
        n32729), .Y(n31836) );
  AOI211xp5_ASAP7_75t_SRAM U27900 ( .A1(u0_0_leon3x0_p0_dco_HIT_), .A2(n32273), 
        .B(n32251), .C(n32274), .Y(n32252) );
  OAI22xp33_ASAP7_75t_SL U27901 ( .A1(n32656), .A2(n31632), .B1(n32417), .B2(
        n31631), .Y(n26490) );
  OAI22xp33_ASAP7_75t_SL U27902 ( .A1(n30527), .A2(n24645), .B1(n32624), .B2(
        n32729), .Y(n30528) );
  OAI22xp33_ASAP7_75t_SL U27903 ( .A1(n30534), .A2(n24645), .B1(n32630), .B2(
        n32729), .Y(n30535) );
  OAI22xp33_ASAP7_75t_SL U27904 ( .A1(n32654), .A2(n31632), .B1(n32405), .B2(
        n31631), .Y(n31493) );
  OAI22xp33_ASAP7_75t_SL U27905 ( .A1(n32618), .A2(n31632), .B1(n32329), .B2(
        n31631), .Y(n26616) );
  OAI22xp33_ASAP7_75t_SL U27906 ( .A1(n32638), .A2(n31632), .B1(n32376), .B2(
        n31631), .Y(n31524) );
  OAI22xp33_ASAP7_75t_SL U27907 ( .A1(n30518), .A2(n24645), .B1(n32628), .B2(
        n32729), .Y(n30519) );
  AOI22xp33_ASAP7_75t_SL U27908 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[4]), .A2(
        n31314), .B1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__4_), .B2(n31313), .Y(
        n31315) );
  OAI22xp33_ASAP7_75t_SL U27909 ( .A1(n30541), .A2(n24645), .B1(n32632), .B2(
        n32729), .Y(n30542) );
  AOI21xp5_ASAP7_75t_SL U27910 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_26_), .A2(
        n31996), .B(n28388), .Y(n3266) );
  AOI21xp5_ASAP7_75t_SL U27911 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_30_), .A2(
        n31996), .B(n31995), .Y(n4319) );
  AOI21xp5_ASAP7_75t_SL U27912 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_14_), .A2(
        n31996), .B(n30501), .Y(n3216) );
  AOI22xp33_ASAP7_75t_SL U27913 ( .A1(n32121), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_NOFLUSH_), .B1(
        u0_0_leon3x0_p0_c0mmu_mmudci[30]), .B2(n32120), .Y(n3056) );
  AOI21xp5_ASAP7_75t_SL U27914 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_24_), .A2(
        n31996), .B(n29772), .Y(n2479) );
  AOI21xp5_ASAP7_75t_SL U27915 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_28_), .A2(
        n31996), .B(n28261), .Y(n3280) );
  AOI22xp33_ASAP7_75t_SL U27916 ( .A1(n32121), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__BURST_), .B1(
        u0_0_leon3x0_p0_c0mmu_mmudci[16]), .B2(n32120), .Y(n2964) );
  INVxp67_ASAP7_75t_SL U27917 ( .A(n31609), .Y(n31309) );
  AOI21xp5_ASAP7_75t_SL U27918 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_13_), .A2(
        n31996), .B(n28592), .Y(n2653) );
  AOI22xp33_ASAP7_75t_SL U27919 ( .A1(n32121), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__0_), .B1(
        u0_0_leon3x0_p0_c0mmu_mmudci[0]), .B2(n32120), .Y(n3907) );
  AOI21xp5_ASAP7_75t_SL U27920 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_20_), .A2(
        n31996), .B(n26974), .Y(n2533) );
  NAND2xp5_ASAP7_75t_SL U27921 ( .A(n30916), .B(n31609), .Y(n32028) );
  AOI21xp5_ASAP7_75t_SL U27922 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_23_), .A2(
        n31996), .B(n29065), .Y(n3252) );
  AOI21xp5_ASAP7_75t_SL U27923 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_17_), .A2(
        n31996), .B(n27270), .Y(n2605) );
  NOR2xp33_ASAP7_75t_SRAM U27924 ( .A(n32234), .B(n33067), .Y(n32202) );
  AOI21xp5_ASAP7_75t_SL U27925 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_16_), .A2(
        n31996), .B(n27228), .Y(n2629) );
  INVxp33_ASAP7_75t_SL U27926 ( .A(n25592), .Y(n25593) );
  INVxp67_ASAP7_75t_SL U27927 ( .A(n22541), .Y(mult_x_1196_n802) );
  AOI21xp5_ASAP7_75t_SL U27928 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_25_), .A2(
        n31996), .B(n28416), .Y(n4599) );
  AOI21xp5_ASAP7_75t_SL U27929 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_22_), .A2(
        n31996), .B(n28477), .Y(n2506) );
  INVxp67_ASAP7_75t_SL U27930 ( .A(n23165), .Y(mult_x_1196_n606) );
  INVxp67_ASAP7_75t_SL U27931 ( .A(n31563), .Y(n32524) );
  AOI22xp33_ASAP7_75t_SL U27932 ( .A1(n32060), .A2(ic_q[14]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__14_), .B2(n22384), .Y(n28461) );
  OAI22xp33_ASAP7_75t_SL U27933 ( .A1(n32602), .A2(n30191), .B1(n3046), .B2(
        n30190), .Y(u0_0_leon3x0_p0_c0mmu_dcache0_v_CCTRL__DCS__0_) );
  AOI22xp33_ASAP7_75t_SL U27934 ( .A1(n32060), .A2(ic_q[30]), .B1(n18839), 
        .B2(n22384), .Y(n31942) );
  AOI22xp33_ASAP7_75t_SL U27935 ( .A1(n32060), .A2(ic_q[21]), .B1(n18842), 
        .B2(n22384), .Y(n31856) );
  AOI22xp33_ASAP7_75t_SL U27936 ( .A1(n32060), .A2(ic_q[20]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), .B2(n22384), .Y(n31536) );
  AOI22xp33_ASAP7_75t_SL U27937 ( .A1(n32060), .A2(ic_q[25]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_), .B2(n22384), .Y(n31377) );
  AOI22xp33_ASAP7_75t_SL U27938 ( .A1(n32060), .A2(ic_q[26]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_), .B2(n22384), .Y(n31332) );
  INVx1_ASAP7_75t_SL U27939 ( .A(n22592), .Y(n22401) );
  AOI22xp33_ASAP7_75t_SL U27940 ( .A1(n32060), .A2(ic_q[22]), .B1(n18819), 
        .B2(n22384), .Y(n31650) );
  NAND2xp33_ASAP7_75t_SL U27941 ( .A(n22379), .B(n32572), .Y(n26240) );
  INVxp33_ASAP7_75t_SL U27942 ( .A(mult_x_1196_n564), .Y(mult_x_1196_n801) );
  AOI22xp33_ASAP7_75t_SL U27943 ( .A1(n32060), .A2(ic_q[15]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__15_), .B2(n22384), .Y(n28412) );
  OAI21xp33_ASAP7_75t_SL U27944 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[5]), .A2(
        n18851), .B(n29998), .Y(n2965) );
  OAI21xp33_ASAP7_75t_SL U27945 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[4]), .A2(
        n18851), .B(n31351), .Y(n2967) );
  AOI22xp33_ASAP7_75t_SL U27946 ( .A1(ic_q[1]), .A2(n32060), .B1(n26823), .B2(
        n22384), .Y(n26824) );
  AOI22xp33_ASAP7_75t_SL U27947 ( .A1(n32060), .A2(ic_q[29]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_), .B2(n22384), .Y(n32061) );
  NAND2xp33_ASAP7_75t_SL U27948 ( .A(n24681), .B(n32596), .Y(n28662) );
  AOI22xp33_ASAP7_75t_SL U27949 ( .A1(n32060), .A2(ic_q[8]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__8_), .B2(n22384), .Y(n25573) );
  AOI22xp33_ASAP7_75t_SL U27950 ( .A1(ic_q[0]), .A2(n32060), .B1(n26820), .B2(
        n22384), .Y(n26821) );
  INVxp67_ASAP7_75t_SL U27951 ( .A(n22441), .Y(mult_x_1196_n644) );
  AOI21xp33_ASAP7_75t_SL U27952 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[24]), .B(n32553), .Y(n4393) );
  AOI21xp33_ASAP7_75t_SL U27953 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__15_), .B(n32528), .Y(n2949)
         );
  AOI21xp33_ASAP7_75t_SL U27954 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[16]), .B(n32532), .Y(n2542) );
  OAI21xp33_ASAP7_75t_SL U27955 ( .A1(mult_x_1196_n714), .A2(mult_x_1196_n716), 
        .B(mult_x_1196_n715), .Y(mult_x_1196_n713) );
  AOI21xp33_ASAP7_75t_SL U27956 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[12]), .B(n32528), .Y(n2948) );
  AOI21xp33_ASAP7_75t_SL U27957 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__11_), .B(n32589), .Y(n2957)
         );
  AOI21xp33_ASAP7_75t_SL U27958 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__21_), .B(n32536), .Y(n2946)
         );
  AOI21xp5_ASAP7_75t_SL U27959 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_11_), .A2(
        n31833), .B(n28661), .Y(n32596) );
  AOI21xp33_ASAP7_75t_SL U27960 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[7]), .B(n32582), .Y(n2953) );
  AOI21xp33_ASAP7_75t_SL U27961 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__14_), .B(n32527), .Y(n2952)
         );
  AOI21xp33_ASAP7_75t_SL U27962 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[11]), .B(n32527), .Y(n2951) );
  AOI21xp33_ASAP7_75t_SL U27963 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__19_), .B(n32532), .Y(n2543)
         );
  AOI21xp33_ASAP7_75t_SL U27964 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__10_), .B(n32582), .Y(n2954)
         );
  OAI21xp33_ASAP7_75t_SL U27965 ( .A1(n31992), .A2(n26972), .B(n26971), .Y(
        n26973) );
  AOI21xp33_ASAP7_75t_SL U27966 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__27_), .B(n32553), .Y(n2955)
         );
  AOI21xp33_ASAP7_75t_SL U27967 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__5_), .B(n32560), .Y(n2961)
         );
  XNOR2xp5_ASAP7_75t_SL U27968 ( .A(mult_x_1196_n275), .B(mult_x_1196_n716), 
        .Y(n23881) );
  NAND2xp33_ASAP7_75t_SL U27969 ( .A(n30012), .B(n18851), .Y(n29998) );
  AOI21xp33_ASAP7_75t_SL U27970 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__13_), .B(n32526), .Y(n2640)
         );
  NAND2xp33_ASAP7_75t_SL U27971 ( .A(n31467), .B(n18851), .Y(n31351) );
  AOI21xp33_ASAP7_75t_SL U27972 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[8]), .B(n32589), .Y(n4477) );
  NAND2xp5_ASAP7_75t_SL U27973 ( .A(n31684), .B(n31683), .Y(n31686) );
  AOI21xp33_ASAP7_75t_SL U27974 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[10]), .B(n32526), .Y(n2639) );
  AOI21xp33_ASAP7_75t_SL U27975 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[6]), .B(n32579), .Y(n4561) );
  OAI21xp33_ASAP7_75t_SL U27976 ( .A1(n31992), .A2(n28259), .B(n28258), .Y(
        n28260) );
  NAND2xp5_ASAP7_75t_SL U27977 ( .A(n30825), .B(n30824), .Y(n30827) );
  NAND2xp5_ASAP7_75t_SL U27978 ( .A(n29028), .B(n29027), .Y(n29030) );
  AOI21xp33_ASAP7_75t_SL U27979 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[15]), .B(n32531), .Y(n2570) );
  AOI21xp33_ASAP7_75t_SL U27980 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__18_), .B(n32531), .Y(n2571)
         );
  AOI21xp33_ASAP7_75t_SL U27981 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[5]), .B(n32576), .Y(n4645) );
  OAI21xp5_ASAP7_75t_SL U27982 ( .A1(n30499), .A2(n30533), .B(n27226), .Y(
        n27227) );
  NAND2xp5_ASAP7_75t_SL U27983 ( .A(n28568), .B(n28567), .Y(n28570) );
  OAI21xp5_ASAP7_75t_SL U27984 ( .A1(n30499), .A2(n30506), .B(n30498), .Y(
        n30500) );
  AOI21xp33_ASAP7_75t_SL U27985 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[14]), .B(n32530), .Y(n2591) );
  AOI21xp33_ASAP7_75t_SL U27986 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__17_), .B(n32530), .Y(n2592)
         );
  NOR2x1_ASAP7_75t_SL U27987 ( .A(n18928), .B(mult_x_1196_n1745), .Y(
        mult_x_1196_n640) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U27988 ( .A1(n32686), .A2(n32679), .B(n32678), 
        .C(n14803), .Y(n32680) );
  NAND2xp33_ASAP7_75t_SL U27989 ( .A(n31618), .B(n31622), .Y(n31445) );
  OAI21xp5_ASAP7_75t_SL U27990 ( .A1(n30499), .A2(n30540), .B(n27268), .Y(
        n27269) );
  AOI21xp33_ASAP7_75t_SL U27991 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__16_), .B(n32529), .Y(n2616)
         );
  AOI21xp33_ASAP7_75t_SL U27992 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[13]), .B(n32529), .Y(n2615) );
  AOI21xp33_ASAP7_75t_SL U27993 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[4]), .B(n32573), .Y(n4759) );
  OAI22xp33_ASAP7_75t_SL U27994 ( .A1(n26786), .A2(n26785), .B1(n22421), .B2(
        u0_0_leon3x0_p0_iu_v_A__CWP__1_), .Y(n2802) );
  NAND2xp5_ASAP7_75t_SL U27995 ( .A(n26876), .B(n26875), .Y(n26878) );
  AOI21xp33_ASAP7_75t_SL U27996 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__31_), .B(n32558), .Y(n2365)
         );
  AOI21xp33_ASAP7_75t_SL U27997 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[28]), .B(n32558), .Y(n2364) );
  NAND2xp5_ASAP7_75t_SL U27998 ( .A(n27042), .B(n27041), .Y(n27044) );
  OAI21xp33_ASAP7_75t_SL U27999 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(n31436), .Y(n2788) );
  OAI21xp33_ASAP7_75t_SL U28000 ( .A1(n31992), .A2(n29063), .B(n29062), .Y(
        n29064) );
  OAI21xp33_ASAP7_75t_SL U28001 ( .A1(n31992), .A2(n28414), .B(n28413), .Y(
        n28415) );
  AOI21xp33_ASAP7_75t_SL U28002 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__6_), .B(n32569), .Y(n2687)
         );
  AOI21xp33_ASAP7_75t_SL U28003 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[3]), .B(n32569), .Y(n2686) );
  NAND2xp5_ASAP7_75t_SL U28004 ( .A(n29822), .B(n29821), .Y(n29824) );
  OAI21xp33_ASAP7_75t_SL U28005 ( .A1(n31992), .A2(n29770), .B(n29769), .Y(
        n29771) );
  AOI21xp33_ASAP7_75t_SL U28006 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__12_), .B(n32523), .Y(n2664)
         );
  AOI21xp33_ASAP7_75t_SL U28007 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[9]), .B(n32523), .Y(n2663) );
  INVxp67_ASAP7_75t_SL U28008 ( .A(n32664), .Y(n30912) );
  OAI21xp5_ASAP7_75t_SL U28009 ( .A1(n30499), .A2(n30526), .B(n28590), .Y(
        n28591) );
  OAI21xp33_ASAP7_75t_SL U28010 ( .A1(n31992), .A2(n28386), .B(n28385), .Y(
        n28387) );
  AOI21xp33_ASAP7_75t_SL U28011 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[18]), .B(n32536), .Y(n2945) );
  AOI21xp33_ASAP7_75t_SL U28012 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[26]), .B(n32555), .Y(n2937) );
  AOI21xp33_ASAP7_75t_SL U28013 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[2]), .B(n32560), .Y(n4748) );
  AOI21xp33_ASAP7_75t_SL U28014 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__29_), .B(n32555), .Y(n2938)
         );
  OAI21xp33_ASAP7_75t_SL U28015 ( .A1(n31992), .A2(n28475), .B(n28474), .Y(
        n28476) );
  OAI21xp33_ASAP7_75t_SL U28016 ( .A1(n31992), .A2(n31991), .B(n31990), .Y(
        n31993) );
  AOI21xp33_ASAP7_75t_SL U28017 ( .A1(u0_0_leon3x0_p0_iu_N5472), .A2(n31830), 
        .B(n30711), .Y(n30713) );
  AOI22xp33_ASAP7_75t_SL U28018 ( .A1(n32060), .A2(ic_q[27]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__27_), .B2(n18901), .Y(n30903) );
  AOI22xp33_ASAP7_75t_SL U28019 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__13_), 
        .A2(n31989), .B1(u0_0_leon3x0_p0_ici[83]), .B2(n31988), .Y(n28413) );
  OAI21xp33_ASAP7_75t_SL U28020 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_E__ALUCIN_), .B(n30964), .Y(n2276) );
  AOI22xp33_ASAP7_75t_SL U28021 ( .A1(ic_q[3]), .A2(n32060), .B1(n28255), .B2(
        n18901), .Y(n28256) );
  AOI22xp33_ASAP7_75t_SL U28022 ( .A1(ic_q[4]), .A2(n32060), .B1(n30791), .B2(
        n18900), .Y(n30792) );
  AOI22xp33_ASAP7_75t_SL U28023 ( .A1(ic_q[2]), .A2(n32060), .B1(n26827), .B2(
        n18901), .Y(n26828) );
  INVxp33_ASAP7_75t_SL U28024 ( .A(u0_0_leon3x0_p0_div0_addout_32_), .Y(n25920) );
  AOI22xp33_ASAP7_75t_SL U28025 ( .A1(n32060), .A2(ic_q[19]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .B2(n18901), .Y(n32009) );
  AOI22xp33_ASAP7_75t_SL U28026 ( .A1(n32060), .A2(ic_q[28]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__28_), .B2(n18900), .Y(n31508) );
  AOI21xp33_ASAP7_75t_SL U28027 ( .A1(u0_0_leon3x0_p0_iu_N5473), .A2(n31830), 
        .B(n26201), .Y(n26207) );
  AOI21xp33_ASAP7_75t_SL U28028 ( .A1(u0_0_leon3x0_p0_iu_N5471), .A2(n31830), 
        .B(n29892), .Y(n29894) );
  O2A1O1Ixp33_ASAP7_75t_SL U28029 ( .A1(n26813), .A2(n26807), .B(n26784), .C(
        n31428), .Y(n26785) );
  OAI22xp33_ASAP7_75t_SL U28030 ( .A1(n26777), .A2(n31435), .B1(n31427), .B2(
        n26776), .Y(n26786) );
  OAI21xp33_ASAP7_75t_SL U28031 ( .A1(n18829), .A2(u0_0_leon3x0_p0_ici[58]), 
        .B(n25886), .Y(n2382) );
  AOI22xp33_ASAP7_75t_SL U28032 ( .A1(n32060), .A2(ic_q[31]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__31_), .B2(n18900), .Y(n31957) );
  AOI22xp33_ASAP7_75t_SL U28033 ( .A1(n32060), .A2(ic_q[17]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_), .B2(n18901), .Y(n30919) );
  AOI22xp33_ASAP7_75t_SL U28034 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__11_), 
        .A2(n31989), .B1(u0_0_leon3x0_p0_ici[81]), .B2(n31988), .Y(n29062) );
  AOI22xp33_ASAP7_75t_SL U28035 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__14_), 
        .A2(n31989), .B1(u0_0_leon3x0_p0_ici[84]), .B2(n31988), .Y(n28385) );
  AOI22xp33_ASAP7_75t_SL U28036 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__16_), 
        .A2(n31989), .B1(u0_0_leon3x0_p0_ici[86]), .B2(n31988), .Y(n28258) );
  NAND2xp33_ASAP7_75t_SL U28037 ( .A(n22242), .B(mult_x_1196_n815), .Y(
        mult_x_1196_n265) );
  OAI21xp33_ASAP7_75t_SL U28038 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_M__DIVZ_), .B(n29871), .Y(n4093) );
  AOI22xp33_ASAP7_75t_SL U28039 ( .A1(n32060), .A2(ic_q[16]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__16_), .B2(n18900), .Y(n28383) );
  AOI22xp33_ASAP7_75t_SL U28040 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__10_), 
        .A2(n31989), .B1(u0_0_leon3x0_p0_ici[80]), .B2(n31988), .Y(n28474) );
  AOI22xp33_ASAP7_75t_SL U28041 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__8_), 
        .A2(n31989), .B1(u0_0_leon3x0_p0_ici[78]), .B2(n31988), .Y(n26971) );
  AOI22xp33_ASAP7_75t_SL U28042 ( .A1(n32060), .A2(ic_q[12]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__12_), .B2(n18900), .Y(n29860) );
  AOI22xp33_ASAP7_75t_SL U28043 ( .A1(n32060), .A2(ic_q[13]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_), .B2(n18900), .Y(n30807) );
  AOI21xp33_ASAP7_75t_SL U28044 ( .A1(u0_0_leon3x0_p0_div0_addout_20_), .A2(
        n31679), .B(n27024), .Y(n2539) );
  AOI21xp33_ASAP7_75t_SL U28045 ( .A1(u0_0_leon3x0_p0_div0_addout_22_), .A2(
        n24639), .B(n28313), .Y(n2512) );
  AOI22xp33_ASAP7_75t_SL U28046 ( .A1(n32060), .A2(ic_q[7]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__7_), .B2(n18901), .Y(n30875) );
  AOI22xp33_ASAP7_75t_SL U28047 ( .A1(n32060), .A2(ic_q[18]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_), .B2(n18900), .Y(n29574) );
  AOI22xp33_ASAP7_75t_SL U28048 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__18_), 
        .A2(n31989), .B1(u0_0_leon3x0_p0_ici[88]), .B2(n31988), .Y(n31990) );
  AOI22xp33_ASAP7_75t_SL U28049 ( .A1(n32060), .A2(ic_q[24]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), .B2(n18901), .Y(n32047) );
  AOI21xp33_ASAP7_75t_SL U28050 ( .A1(u0_0_leon3x0_p0_iu_N5474), .A2(n31830), 
        .B(n28703), .Y(n28705) );
  AOI22xp33_ASAP7_75t_SL U28051 ( .A1(n32060), .A2(ic_q[11]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__11_), .B2(n18900), .Y(n28518) );
  AOI22xp33_ASAP7_75t_SL U28052 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__12_), 
        .A2(n31989), .B1(u0_0_leon3x0_p0_ici[82]), .B2(n31988), .Y(n29769) );
  AOI21xp33_ASAP7_75t_SL U28053 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[19]), .B(n32537), .Y(n2492) );
  NAND2xp33_ASAP7_75t_SL U28054 ( .A(n31804), .B(n18901), .Y(n31805) );
  AOI22xp33_ASAP7_75t_SL U28055 ( .A1(n32060), .A2(ic_q[23]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), .B2(n18901), .Y(n31979) );
  AOI22xp33_ASAP7_75t_SL U28056 ( .A1(n32060), .A2(ic_q[9]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__9_), .B2(n18900), .Y(n30154) );
  AOI22xp33_ASAP7_75t_SL U28057 ( .A1(n32060), .A2(ic_q[10]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__10_), .B2(n18901), .Y(n26969) );
  AOI21xp33_ASAP7_75t_SL U28058 ( .A1(n22385), .A2(
        u0_0_leon3x0_p0_c0mmu_mcii[21]), .B(n32544), .Y(n2465) );
  AOI22xp33_ASAP7_75t_SL U28059 ( .A1(n32060), .A2(ic_q[6]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__6_), .B2(n18900), .Y(n31253) );
  AOI21xp33_ASAP7_75t_SL U28060 ( .A1(u0_0_leon3x0_p0_div0_addout_24_), .A2(
        n24639), .B(n28308), .Y(n2485) );
  AOI22xp33_ASAP7_75t_SL U28061 ( .A1(n32060), .A2(ic_q[5]), .B1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__5_), .B2(n18901), .Y(n30113) );
  OAI21xp33_ASAP7_75t_SL U28062 ( .A1(n32110), .A2(n26958), .B(n26957), .Y(
        n4404) );
  OAI21xp33_ASAP7_75t_SL U28063 ( .A1(n30828), .A2(n24585), .B(n30822), .Y(
        n30823) );
  OAI21xp33_ASAP7_75t_SL U28064 ( .A1(n24585), .A2(n32577), .B(n30710), .Y(
        n30711) );
  OAI21xp33_ASAP7_75t_SL U28065 ( .A1(n31786), .A2(n24585), .B(n26873), .Y(
        n26874) );
  OAI21xp33_ASAP7_75t_SL U28066 ( .A1(n31765), .A2(n24585), .B(n27039), .Y(
        n27040) );
  NAND2xp33_ASAP7_75t_SL U28067 ( .A(n25890), .B(n18829), .Y(n25886) );
  NAND2x1p5_ASAP7_75t_SL U28068 ( .A(mult_x_1196_n815), .B(mult_x_1196_n816), 
        .Y(mult_x_1196_n654) );
  OAI21xp33_ASAP7_75t_SL U28069 ( .A1(n31834), .A2(n24585), .B(n31825), .Y(
        n31827) );
  AOI21xp33_ASAP7_75t_SL U28070 ( .A1(u0_0_leon3x0_p0_iu_r_A__CTRL__WREG_), 
        .A2(n22378), .B(n32106), .Y(n2714) );
  OAI21xp33_ASAP7_75t_SL U28071 ( .A1(n24585), .A2(n32567), .B(n29677), .Y(
        n29678) );
  OAI21xp33_ASAP7_75t_SL U28072 ( .A1(n24585), .A2(n32677), .B(n30910), .Y(
        n30911) );
  OAI21xp33_ASAP7_75t_SL U28073 ( .A1(n31690), .A2(n24585), .B(n29025), .Y(
        n29026) );
  NAND2xp5_ASAP7_75t_SL U28074 ( .A(n23785), .B(n23787), .Y(n23786) );
  OAI21xp33_ASAP7_75t_SL U28075 ( .A1(n24585), .A2(n30974), .B(n28659), .Y(
        n28660) );
  AOI22xp33_ASAP7_75t_SL U28076 ( .A1(u0_0_leon3x0_p0_iu_r_A__BP_), .A2(n24648), .B1(n26191), .B2(n25233), .Y(n3298) );
  OAI21xp33_ASAP7_75t_SL U28077 ( .A1(n24585), .A2(n32580), .B(n26200), .Y(
        n26201) );
  AOI21xp33_ASAP7_75t_SL U28078 ( .A1(u0_0_leon3x0_p0_iu_r_A__NOBP_), .A2(
        n22378), .B(n32058), .Y(n3300) );
  INVxp67_ASAP7_75t_SL U28079 ( .A(mult_x_1196_n423), .Y(mult_x_1196_n425) );
  OAI21xp33_ASAP7_75t_SL U28080 ( .A1(n30524), .A2(n24585), .B(n29819), .Y(
        n29820) );
  INVxp67_ASAP7_75t_SL U28081 ( .A(mult_x_1196_n692), .Y(mult_x_1196_n821) );
  AOI22xp33_ASAP7_75t_SL U28082 ( .A1(n31432), .A2(n31431), .B1(n31430), .B2(
        n31429), .Y(n31433) );
  OAI21xp33_ASAP7_75t_SL U28083 ( .A1(n24585), .A2(n32574), .B(n29891), .Y(
        n29892) );
  AOI22xp33_ASAP7_75t_SL U28084 ( .A1(u0_0_leon3x0_p0_iu_r_A__CTRL__WICC_), 
        .A2(n24649), .B1(n25229), .B2(n31387), .Y(n4410) );
  OAI21xp33_ASAP7_75t_SL U28085 ( .A1(n24585), .A2(n32586), .B(n28702), .Y(
        n28703) );
  OAI21xp33_ASAP7_75t_SL U28086 ( .A1(n24585), .A2(n31018), .B(n26237), .Y(
        n26238) );
  OAI21xp33_ASAP7_75t_SL U28087 ( .A1(n30517), .A2(n24585), .B(n28565), .Y(
        n28566) );
  INVxp67_ASAP7_75t_SL U28088 ( .A(n23215), .Y(n23213) );
  INVxp67_ASAP7_75t_SL U28089 ( .A(n22726), .Y(n22725) );
  INVx1_ASAP7_75t_SL U28090 ( .A(mult_x_1196_n416), .Y(n23225) );
  NAND2xp33_ASAP7_75t_SL U28091 ( .A(n31830), .B(u0_0_leon3x0_p0_iu_N5491), 
        .Y(n26875) );
  NAND2xp5_ASAP7_75t_SL U28092 ( .A(n25603), .B(n25602), .Y(n31815) );
  INVxp67_ASAP7_75t_SL U28093 ( .A(mult_x_1196_n1327), .Y(n23787) );
  NAND2xp33_ASAP7_75t_SL U28094 ( .A(n31830), .B(u0_0_leon3x0_p0_iu_N5476), 
        .Y(n29821) );
  OAI21xp33_ASAP7_75t_SL U28095 ( .A1(n32482), .A2(n31894), .B(n31882), .Y(
        n31937) );
  NAND2xp33_ASAP7_75t_SL U28096 ( .A(n31833), .B(u0_0_leon3x0_p0_iu_fe_npc_9_), 
        .Y(n26206) );
  NAND2xp33_ASAP7_75t_SL U28097 ( .A(n31830), .B(u0_0_leon3x0_p0_iu_N5479), 
        .Y(n28567) );
  AOI21xp33_ASAP7_75t_SL U28098 ( .A1(n31426), .A2(n31425), .B(
        u0_0_leon3x0_p0_iu_v_A__CWP__0_), .Y(n31434) );
  OAI21xp33_ASAP7_75t_SL U28099 ( .A1(n32110), .A2(n27035), .B(n25842), .Y(
        n4358) );
  OAI21xp33_ASAP7_75t_SL U28100 ( .A1(n32114), .A2(n32113), .B(n32112), .Y(
        n2762) );
  AOI22xp33_ASAP7_75t_SL U28101 ( .A1(u0_0_leon3x0_p0_iu_r_E__SARI_), .A2(
        n24648), .B1(n25078), .B2(n30949), .Y(n3572) );
  AOI21xp5_ASAP7_75t_SL U28102 ( .A1(n30963), .A2(n30960), .B(n30959), .Y(
        n30961) );
  OAI21xp33_ASAP7_75t_SL U28103 ( .A1(n30794), .A2(n28866), .B(n28865), .Y(
        n2753) );
  NAND2xp33_ASAP7_75t_SL U28104 ( .A(n31833), .B(u0_0_leon3x0_p0_iu_fe_npc_7_), 
        .Y(n29893) );
  AND2x2_ASAP7_75t_SL U28105 ( .A(n23229), .B(mult_x_1196_n227), .Y(n23236) );
  NAND2xp33_ASAP7_75t_SL U28106 ( .A(n31830), .B(u0_0_leon3x0_p0_iu_N5493), 
        .Y(n29027) );
  OAI21xp33_ASAP7_75t_SL U28107 ( .A1(n31343), .A2(n27286), .B(n27285), .Y(
        n4036) );
  AOI22xp33_ASAP7_75t_SL U28108 ( .A1(u0_0_leon3x0_p0_ici[29]), .A2(n24649), 
        .B1(n33056), .B2(n31896), .Y(n3296) );
  INVxp67_ASAP7_75t_SL U28109 ( .A(n32104), .Y(n25233) );
  NAND2xp33_ASAP7_75t_SL U28110 ( .A(n31830), .B(u0_0_leon3x0_p0_iu_N5495), 
        .Y(n31683) );
  NAND2xp33_ASAP7_75t_SL U28111 ( .A(n30648), .B(n29014), .Y(n29016) );
  NAND2xp33_ASAP7_75t_SL U28112 ( .A(n31830), .B(u0_0_leon3x0_p0_iu_N5485), 
        .Y(n27041) );
  AOI22xp33_ASAP7_75t_SL U28113 ( .A1(n24647), .A2(n26956), .B1(n31542), .B2(
        n29802), .Y(n26957) );
  OR2x2_ASAP7_75t_SL U28114 ( .A(mult_x_1196_n932), .B(n22221), .Y(n24305) );
  INVxp33_ASAP7_75t_SL U28115 ( .A(u0_0_leon3x0_p0_div0_addout_15_), .Y(n25927) );
  INVxp67_ASAP7_75t_SL U28116 ( .A(mult_x_1196_n368), .Y(mult_x_1196_n366) );
  NAND2xp33_ASAP7_75t_SL U28117 ( .A(n31833), .B(u0_0_leon3x0_p0_iu_fe_npc_8_), 
        .Y(n30712) );
  NAND2xp33_ASAP7_75t_SL U28118 ( .A(n31833), .B(u0_0_leon3x0_p0_iu_fe_npc_10_), .Y(n28704) );
  NAND2xp5_ASAP7_75t_SL U28119 ( .A(n24307), .B(n24276), .Y(mult_x_1196_n718)
         );
  OAI21xp33_ASAP7_75t_SL U28120 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[18]), .B(n31822), .Y(n4000) );
  NAND2xp33_ASAP7_75t_SL U28121 ( .A(n31830), .B(u0_0_leon3x0_p0_iu_N5483), 
        .Y(n30824) );
  NAND2xp33_ASAP7_75t_SL U28122 ( .A(n31830), .B(u0_0_leon3x0_p0_iu_N5468), 
        .Y(n29478) );
  NOR2xp33_ASAP7_75t_SL U28123 ( .A(n24646), .B(mult_x_1196_n229), .Y(n23215)
         );
  AOI21xp33_ASAP7_75t_SL U28124 ( .A1(u0_0_leon3x0_p0_iu_de_icc_1_), .A2(
        n30946), .B(n30945), .Y(n30947) );
  OAI22xp33_ASAP7_75t_SL U28125 ( .A1(n32110), .A2(n31540), .B1(n23229), .B2(
        n31539), .Y(n31541) );
  NAND2xp5_ASAP7_75t_SL U28126 ( .A(n29934), .B(n29933), .Y(n3965) );
  OAI21xp33_ASAP7_75t_SL U28127 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__4_), 
        .A2(n31491), .B(n31490), .Y(n2966) );
  INVxp67_ASAP7_75t_SL U28128 ( .A(n28279), .Y(n26958) );
  NAND2xp33_ASAP7_75t_SL U28129 ( .A(n31054), .B(n27280), .Y(n26719) );
  INVxp67_ASAP7_75t_SL U28130 ( .A(n31821), .Y(n31822) );
  NAND2xp5_ASAP7_75t_SL U28131 ( .A(n30954), .B(n30953), .Y(n30963) );
  OAI21xp33_ASAP7_75t_SL U28132 ( .A1(n32819), .A2(n32821), .B(n32818), .Y(
        n1643) );
  OAI21xp33_ASAP7_75t_SL U28133 ( .A1(n31400), .A2(n29789), .B(n29788), .Y(
        n29806) );
  AOI22xp33_ASAP7_75t_SL U28134 ( .A1(n24647), .A2(n27284), .B1(n27283), .B2(
        n27282), .Y(n27285) );
  INVxp67_ASAP7_75t_SL U28135 ( .A(n29013), .Y(n29014) );
  OAI21xp33_ASAP7_75t_SL U28136 ( .A1(n24646), .A2(n26955), .B(n26911), .Y(
        n4119) );
  AOI22xp33_ASAP7_75t_SL U28137 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__1_), 
        .A2(n31364), .B1(n31491), .B2(n31363), .Y(n3912) );
  AOI22xp33_ASAP7_75t_SL U28138 ( .A1(n24647), .A2(n25841), .B1(n25840), .B2(
        n27282), .Y(n25842) );
  O2A1O1Ixp33_ASAP7_75t_SL U28139 ( .A1(n30595), .A2(n28818), .B(n28817), .C(
        n28816), .Y(n2688) );
  NAND2xp33_ASAP7_75t_SL U28140 ( .A(n30648), .B(n30647), .Y(n30650) );
  NAND2xp33_ASAP7_75t_SL U28141 ( .A(n32689), .B(n32127), .Y(n32046) );
  OAI21xp33_ASAP7_75t_SL U28142 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__6_), 
        .A2(n31491), .B(n30571), .Y(n3034) );
  OAI21xp33_ASAP7_75t_SL U28143 ( .A1(n24541), .A2(n29845), .B(n28652), .Y(
        n28656) );
  OAI21xp33_ASAP7_75t_SL U28144 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__3_), 
        .A2(n31491), .B(n30890), .Y(n3036) );
  AOI21xp33_ASAP7_75t_SL U28145 ( .A1(n31542), .A2(n27035), .B(n27034), .Y(
        n4040) );
  OAI21xp33_ASAP7_75t_SL U28146 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__2_), 
        .A2(n31491), .B(n31011), .Y(n3040) );
  OAI21xp33_ASAP7_75t_SL U28147 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__0_), 
        .A2(n31491), .B(n30486), .Y(n3041) );
  NAND2xp33_ASAP7_75t_SL U28148 ( .A(n30593), .B(n28516), .Y(n28515) );
  OAI21xp33_ASAP7_75t_SL U28149 ( .A1(n31400), .A2(n29845), .B(n24539), .Y(
        n29843) );
  OAI21xp33_ASAP7_75t_SL U28150 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_E__SHCNT__4_), .B(n30795), .Y(n2755) );
  OAI22xp33_ASAP7_75t_SL U28151 ( .A1(n32808), .A2(n32807), .B1(n32821), .B2(
        n32806), .Y(n1647) );
  INVxp67_ASAP7_75t_SL U28152 ( .A(n32111), .Y(n32112) );
  NAND2xp33_ASAP7_75t_SL U28153 ( .A(n31542), .B(n30490), .Y(n30494) );
  OAI21xp33_ASAP7_75t_SL U28154 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_r_E__YMSB_), .B(n32113), .Y(n2764) );
  OAI22xp33_ASAP7_75t_SL U28155 ( .A1(n32816), .A2(n32807), .B1(n32821), .B2(
        n32795), .Y(n1655) );
  OAI21xp33_ASAP7_75t_SL U28156 ( .A1(n32800), .A2(n32821), .B(n32799), .Y(
        n1651) );
  NAND2xp33_ASAP7_75t_SL U28157 ( .A(n30648), .B(n30794), .Y(n28865) );
  OAI21xp33_ASAP7_75t_SL U28158 ( .A1(n31343), .A2(n29905), .B(n29904), .Y(
        n3930) );
  OAI21xp33_ASAP7_75t_SL U28159 ( .A1(n24646), .A2(n27263), .B(n27262), .Y(
        n4038) );
  OAI22xp33_ASAP7_75t_SL U28160 ( .A1(n31343), .A2(n32109), .B1(n22421), .B2(
        u0_0_leon3x0_p0_iu_r_E__OP1__1_), .Y(n31344) );
  NAND2xp33_ASAP7_75t_SL U28161 ( .A(n30593), .B(n28818), .Y(n28817) );
  OAI21xp33_ASAP7_75t_SL U28162 ( .A1(n31343), .A2(n30469), .B(n29502), .Y(
        n3961) );
  OAI21xp33_ASAP7_75t_SL U28163 ( .A1(n30818), .A2(n28906), .B(n28905), .Y(
        n3957) );
  NAND2xp5_ASAP7_75t_SL U28164 ( .A(n32811), .B(n32817), .Y(n32807) );
  OAI21xp33_ASAP7_75t_SL U28165 ( .A1(n31013), .A2(n28958), .B(n28957), .Y(
        n3951) );
  AOI21xp33_ASAP7_75t_SL U28166 ( .A1(n30946), .A2(
        u0_0_leon3x0_p0_iu_de_icc_3_), .B(n30944), .Y(n30948) );
  OAI21xp33_ASAP7_75t_SL U28167 ( .A1(n32119), .A2(n31400), .B(n31399), .Y(
        n32113) );
  OAI22xp33_ASAP7_75t_SL U28168 ( .A1(n32110), .A2(n32109), .B1(n23229), .B2(
        u0_0_leon3x0_p0_iu_r_E__OP1__0_), .Y(n32111) );
  AOI22xp33_ASAP7_75t_SL U28169 ( .A1(n24647), .A2(n29903), .B1(n31054), .B2(
        n29927), .Y(n29904) );
  OAI22xp33_ASAP7_75t_SL U28170 ( .A1(n31873), .A2(n30794), .B1(n31872), .B2(
        n30793), .Y(n30795) );
  AOI21xp33_ASAP7_75t_SL U28171 ( .A1(n27263), .A2(n31342), .B(n26718), .Y(
        n27280) );
  AOI21xp33_ASAP7_75t_SL U28172 ( .A1(n29800), .A2(n31342), .B(n29799), .Y(
        n29804) );
  AOI22xp33_ASAP7_75t_SL U28173 ( .A1(n24647), .A2(n29928), .B1(n31542), .B2(
        n29927), .Y(n29934) );
  OAI21xp33_ASAP7_75t_SL U28174 ( .A1(n31400), .A2(n28807), .B(n26289), .Y(
        n29905) );
  OAI21xp33_ASAP7_75t_SL U28175 ( .A1(n24646), .A2(n29867), .B(n25918), .Y(
        n4115) );
  OAI21xp33_ASAP7_75t_SL U28176 ( .A1(n24646), .A2(n28275), .B(n28274), .Y(
        n4117) );
  INVxp67_ASAP7_75t_SL U28177 ( .A(n22332), .Y(n23607) );
  NOR2x1_ASAP7_75t_SL U28178 ( .A(mult_x_1196_n323), .B(mult_x_1196_n316), .Y(
        n23474) );
  OAI21xp33_ASAP7_75t_SL U28179 ( .A1(u0_0_leon3x0_p0_c0mmu_icache0_r_OVERRUN_), .A2(n32123), .B(n31893), .Y(n32127) );
  OAI22xp33_ASAP7_75t_SL U28180 ( .A1(n31051), .A2(n31050), .B1(n23229), .B2(
        u0_0_leon3x0_p0_iu_r_E__OP1__10_), .Y(n31052) );
  NAND2xp33_ASAP7_75t_SL U28181 ( .A(n30593), .B(n27016), .Y(n27015) );
  AOI22xp5_ASAP7_75t_SL U28182 ( .A1(n30671), .A2(n30295), .B1(n30666), .B2(
        n27022), .Y(n30953) );
  AOI21xp33_ASAP7_75t_SL U28183 ( .A1(n29078), .A2(n31342), .B(n29077), .Y(
        n31540) );
  OAI22xp33_ASAP7_75t_SL U28184 ( .A1(n32110), .A2(n27087), .B1(n22421), .B2(
        n27033), .Y(n27034) );
  AOI22xp33_ASAP7_75t_SL U28185 ( .A1(n24647), .A2(n29841), .B1(n31542), .B2(
        n31053), .Y(n29842) );
  NAND2xp33_ASAP7_75t_SL U28186 ( .A(n31054), .B(n30733), .Y(n30734) );
  AOI21xp5_ASAP7_75t_SL U28187 ( .A1(n31486), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__6_), .B(n30567), .Y(n30568)
         );
  OAI22xp33_ASAP7_75t_SL U28188 ( .A1(n32811), .A2(n32810), .B1(ramsn[3]), 
        .B2(n32809), .Y(n1645) );
  NAND2xp5_ASAP7_75t_SL U28189 ( .A(n28506), .B(n28505), .Y(n29078) );
  AOI21xp5_ASAP7_75t_SL U28190 ( .A1(n27032), .A2(n31342), .B(n27031), .Y(
        n27087) );
  NAND2xp5_ASAP7_75t_SL U28191 ( .A(n26185), .B(n26184), .Y(n28608) );
  OAI21xp33_ASAP7_75t_SL U28192 ( .A1(n24646), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N8), .B(n29103), .Y(n4299) );
  NAND2xp5_ASAP7_75t_SL U28193 ( .A(n29612), .B(n29611), .Y(n30597) );
  AOI21xp33_ASAP7_75t_SL U28194 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__1_), .A2(n31486), .B(n31360), .Y(n31361) );
  AOI21xp33_ASAP7_75t_SL U28195 ( .A1(n30799), .A2(n31342), .B(n29902), .Y(
        n29927) );
  OAI21xp33_ASAP7_75t_SL U28196 ( .A1(DP_OP_5187J1_124_3275_n296), .A2(
        DP_OP_5187J1_124_3275_n298), .B(DP_OP_5187J1_124_3275_n297), .Y(
        DP_OP_5187J1_124_3275_n295) );
  AOI21xp5_ASAP7_75t_SL U28197 ( .A1(n31486), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__4_), .B(n31485), .Y(n31487)
         );
  NAND2xp33_ASAP7_75t_SL U28198 ( .A(n30648), .B(n31013), .Y(n28957) );
  AOI21xp5_ASAP7_75t_SL U28199 ( .A1(n31486), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__0_), .B(n30483), .Y(n30484)
         );
  OAI22xp33_ASAP7_75t_SL U28200 ( .A1(n32811), .A2(n32796), .B1(ramsn[1]), 
        .B2(n32809), .Y(n1653) );
  MAJx2_ASAP7_75t_SL U28201 ( .A(n22523), .B(mult_x_1196_n924), .C(n22362), 
        .Y(mult_x_1196_n918) );
  AOI21xp5_ASAP7_75t_SL U28202 ( .A1(n31486), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__2_), .B(n31008), .Y(n31009)
         );
  OAI22xp33_ASAP7_75t_SL U28203 ( .A1(n32110), .A2(n30469), .B1(n22421), .B2(
        u0_0_leon3x0_p0_iu_r_E__OP1__2_), .Y(n30470) );
  OAI21xp33_ASAP7_75t_SL U28204 ( .A1(n1723), .A2(n33053), .B(n32740), .Y(
        sr1_v_ADDRESS__1_) );
  OAI22xp33_ASAP7_75t_SL U28205 ( .A1(n32815), .A2(n32810), .B1(ramsn[2]), 
        .B2(n32809), .Y(n1649) );
  NAND2xp33_ASAP7_75t_SL U28206 ( .A(n30648), .B(n30818), .Y(n28905) );
  AOI21xp5_ASAP7_75t_SL U28207 ( .A1(n31486), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__3_), .B(n30888), .Y(n30889)
         );
  OAI21xp33_ASAP7_75t_SL U28208 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[3]), .B(n30967), .Y(n3959) );
  INVx1_ASAP7_75t_SL U28209 ( .A(mult_x_1196_n947), .Y(n24208) );
  OAI22xp33_ASAP7_75t_SL U28210 ( .A1(n30659), .A2(n30658), .B1(
        u0_0_leon3x0_p0_dci[36]), .B2(n30657), .Y(n30676) );
  OAI21xp33_ASAP7_75t_SL U28211 ( .A1(n1724), .A2(n33053), .B(n32720), .Y(
        sr1_v_ADDRESS__0_) );
  NAND2xp5_ASAP7_75t_SL U28212 ( .A(n26696), .B(n26695), .Y(n31875) );
  INVxp67_ASAP7_75t_SL U28213 ( .A(n28645), .Y(n28646) );
  OAI22xp33_ASAP7_75t_SL U28214 ( .A1(n32815), .A2(n32796), .B1(ramsn[0]), 
        .B2(n32809), .Y(n1657) );
  NAND2xp5_ASAP7_75t_SL U28215 ( .A(n28748), .B(n28747), .Y(n30736) );
  INVxp67_ASAP7_75t_SL U28216 ( .A(mult_x_1196_n1147), .Y(n23508) );
  AOI21xp33_ASAP7_75t_SL U28217 ( .A1(n32991), .A2(n32990), .B(n32989), .Y(
        n1684) );
  AOI22xp33_ASAP7_75t_SL U28218 ( .A1(n22386), .A2(address[6]), .B1(n32994), 
        .B2(n33053), .Y(n1683) );
  OAI21xp33_ASAP7_75t_SL U28219 ( .A1(n22386), .A2(n33049), .B(n33048), .Y(
        n1664) );
  AOI22xp33_ASAP7_75t_SL U28220 ( .A1(n22386), .A2(address[11]), .B1(n33003), 
        .B2(n33053), .Y(n1679) );
  AOI21xp33_ASAP7_75t_SL U28221 ( .A1(n24424), .A2(ahbso_1__HREADY_), .B(
        n32041), .Y(n4392) );
  AOI22xp33_ASAP7_75t_SL U28222 ( .A1(n22386), .A2(address[10]), .B1(n33001), 
        .B2(n33053), .Y(n1680) );
  AOI22xp33_ASAP7_75t_SL U28223 ( .A1(n22386), .A2(address[8]), .B1(n32997), 
        .B2(n33053), .Y(n1682) );
  AOI22xp33_ASAP7_75t_SL U28224 ( .A1(n22386), .A2(address[3]), .B1(n32985), 
        .B2(n33053), .Y(n1685) );
  AOI22xp33_ASAP7_75t_SL U28225 ( .A1(n22386), .A2(address[7]), .B1(n32995), 
        .B2(n33053), .Y(n1632) );
  AOI22xp33_ASAP7_75t_SL U28226 ( .A1(n31989), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__5_), .B1(n30497), .B2(
        u0_0_leon3x0_p0_dci[22]), .Y(n27268) );
  NAND2xp5_ASAP7_75t_SL U28227 ( .A(n27164), .B(n27163), .Y(n31055) );
  AOI22xp33_ASAP7_75t_SL U28228 ( .A1(n22386), .A2(address[9]), .B1(n32999), 
        .B2(n33053), .Y(n1681) );
  OAI21xp33_ASAP7_75t_SL U28229 ( .A1(n22386), .A2(n33046), .B(n33045), .Y(
        n1665) );
  AOI22xp33_ASAP7_75t_SL U28230 ( .A1(n22386), .A2(address[2]), .B1(n32984), 
        .B2(n33053), .Y(n1686) );
  INVx1_ASAP7_75t_SL U28231 ( .A(n25447), .Y(n31047) );
  OAI21xp33_ASAP7_75t_SL U28232 ( .A1(n22386), .A2(n33017), .B(n33016), .Y(
        n1674) );
  OAI21xp33_ASAP7_75t_SL U28233 ( .A1(n22386), .A2(n33020), .B(n33019), .Y(
        n1673) );
  OAI21xp33_ASAP7_75t_SL U28234 ( .A1(n31359), .A2(n31483), .B(n31358), .Y(
        n31360) );
  OAI21xp33_ASAP7_75t_SL U28235 ( .A1(n22386), .A2(n33023), .B(n33022), .Y(
        n1672) );
  NAND2xp33_ASAP7_75t_SL U28236 ( .A(n22398), .B(u0_0_leon3x0_p0_dci[29]), .Y(
        n26411) );
  OAI21xp33_ASAP7_75t_SL U28237 ( .A1(n22386), .A2(n33026), .B(n33025), .Y(
        n1671) );
  INVxp33_ASAP7_75t_SL U28238 ( .A(u0_0_leon3x0_p0_dci[29]), .Y(n29770) );
  OAI21xp33_ASAP7_75t_SL U28239 ( .A1(n22386), .A2(n33039), .B(n33038), .Y(
        n1667) );
  OAI21xp33_ASAP7_75t_SL U28240 ( .A1(n22386), .A2(n33029), .B(n33028), .Y(
        n1670) );
  INVxp33_ASAP7_75t_SL U28241 ( .A(u0_0_leon3x0_p0_dci[28]), .Y(n29063) );
  OAI21xp33_ASAP7_75t_SL U28242 ( .A1(n22386), .A2(n33032), .B(n33031), .Y(
        n1669) );
  INVxp33_ASAP7_75t_SL U28243 ( .A(u0_0_leon3x0_p0_dci[36]), .Y(n30658) );
  INVxp33_ASAP7_75t_SL U28244 ( .A(u0_0_leon3x0_p0_dci[33]), .Y(n28259) );
  INVxp33_ASAP7_75t_SL U28245 ( .A(u0_0_leon3x0_p0_dci[30]), .Y(n28414) );
  NAND2xp33_ASAP7_75t_SL U28246 ( .A(n24681), .B(n30966), .Y(n30967) );
  AOI21xp33_ASAP7_75t_SL U28247 ( .A1(n29626), .A2(n31342), .B(n29500), .Y(
        n29688) );
  NAND2xp33_ASAP7_75t_SL U28248 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[37]), .B(
        n32991), .Y(n32740) );
  INVxp67_ASAP7_75t_SL U28249 ( .A(DP_OP_5187J1_124_3275_n162), .Y(
        DP_OP_5187J1_124_3275_n164) );
  AOI21xp33_ASAP7_75t_SL U28250 ( .A1(n31947), .A2(n31342), .B(n26324), .Y(
        n29686) );
  INVxp67_ASAP7_75t_SL U28251 ( .A(DP_OP_5187J1_124_3275_n161), .Y(
        DP_OP_5187J1_124_3275_n163) );
  OAI21xp33_ASAP7_75t_SL U28252 ( .A1(n22386), .A2(n33036), .B(n33035), .Y(
        n1668) );
  NAND2xp33_ASAP7_75t_SL U28253 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[36]), .B(
        n32991), .Y(n32720) );
  OAI21xp33_ASAP7_75t_SL U28254 ( .A1(n31400), .A2(n30966), .B(n29497), .Y(
        n30469) );
  AOI22xp33_ASAP7_75t_SL U28255 ( .A1(n31989), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__1_), .B1(u0_0_leon3x0_p0_dci[18]), 
        .B2(n30497), .Y(n28590) );
  INVxp33_ASAP7_75t_SL U28256 ( .A(u0_0_leon3x0_p0_dci[27]), .Y(n28475) );
  INVxp67_ASAP7_75t_SL U28257 ( .A(n22525), .Y(n22523) );
  NAND2xp5_ASAP7_75t_SL U28258 ( .A(n27125), .B(n27124), .Y(n27174) );
  OAI21xp33_ASAP7_75t_SL U28259 ( .A1(n22386), .A2(n33007), .B(n33006), .Y(
        n1678) );
  INVxp67_ASAP7_75t_SL U28260 ( .A(mult_x_1196_n734), .Y(mult_x_1196_n732) );
  OAI21xp33_ASAP7_75t_SL U28261 ( .A1(n30482), .A2(n31045), .B(n29763), .Y(
        n29764) );
  OAI21xp33_ASAP7_75t_SL U28262 ( .A1(n30970), .A2(n31045), .B(n30969), .Y(
        n30971) );
  NAND2xp5_ASAP7_75t_SL U28263 ( .A(n24142), .B(n24144), .Y(n24145) );
  OAI21xp33_ASAP7_75t_SL U28264 ( .A1(n22386), .A2(n33043), .B(n33042), .Y(
        n1666) );
  OAI21xp33_ASAP7_75t_SL U28265 ( .A1(n31484), .A2(n31045), .B(n25446), .Y(
        n25448) );
  AOI22xp33_ASAP7_75t_SL U28266 ( .A1(n31989), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__4_), .B1(n30497), .B2(
        u0_0_leon3x0_p0_dci[21]), .Y(n27226) );
  AOI22xp33_ASAP7_75t_SL U28267 ( .A1(n31989), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__2_), .B1(n30497), .B2(
        u0_0_leon3x0_p0_dci[19]), .Y(n30498) );
  AOI22xp33_ASAP7_75t_SL U28268 ( .A1(n22386), .A2(address[5]), .B1(n32993), 
        .B2(n33053), .Y(n1636) );
  OAI21xp33_ASAP7_75t_SL U28269 ( .A1(n22386), .A2(n33014), .B(n33013), .Y(
        n1675) );
  AOI21xp33_ASAP7_75t_SL U28270 ( .A1(u0_0_leon3x0_p0_dci[23]), .A2(n22398), 
        .B(n25837), .Y(n25839) );
  OAI21xp33_ASAP7_75t_SL U28271 ( .A1(n22386), .A2(n33011), .B(n33010), .Y(
        n1676) );
  INVxp67_ASAP7_75t_SL U28272 ( .A(DP_OP_5187J1_124_3275_n6), .Y(
        DP_OP_5187J1_124_3275_n87) );
  OAI21xp33_ASAP7_75t_SL U28273 ( .A1(n31037), .A2(n31045), .B(n31036), .Y(
        n31038) );
  OAI21xp33_ASAP7_75t_SL U28274 ( .A1(n22386), .A2(n33052), .B(n33051), .Y(
        n1663) );
  INVxp67_ASAP7_75t_SL U28275 ( .A(DP_OP_5187J1_124_3275_n5), .Y(
        DP_OP_5187J1_124_3275_n88) );
  OAI21xp33_ASAP7_75t_SL U28276 ( .A1(datadir[3]), .A2(n32831), .B(n32830), 
        .Y(n2293) );
  NAND2xp33_ASAP7_75t_SL U28277 ( .A(n33050), .B(n22386), .Y(n33051) );
  INVxp33_ASAP7_75t_SL U28278 ( .A(DP_OP_5187J1_124_3275_n108), .Y(
        DP_OP_5187J1_124_3275_n110) );
  INVxp67_ASAP7_75t_SL U28279 ( .A(n32880), .Y(n32881) );
  OAI21xp33_ASAP7_75t_SL U28280 ( .A1(datadir[1]), .A2(n32831), .B(n32830), 
        .Y(n2297) );
  INVxp33_ASAP7_75t_SL U28281 ( .A(DP_OP_5187J1_124_3275_n107), .Y(
        DP_OP_5187J1_124_3275_n109) );
  OAI21xp33_ASAP7_75t_SL U28282 ( .A1(datadir[2]), .A2(n32831), .B(n32830), 
        .Y(n2295) );
  XNOR2xp5_ASAP7_75t_SL U28283 ( .A(n22350), .B(mult_x_1196_n1368), .Y(n24154)
         );
  OAI21xp33_ASAP7_75t_SL U28284 ( .A1(n2356), .A2(n32875), .B(n31693), .Y(
        n17904) );
  NAND2xp33_ASAP7_75t_SL U28285 ( .A(n33005), .B(n22386), .Y(n33006) );
  NAND2xp33_ASAP7_75t_SL U28286 ( .A(n33009), .B(n22386), .Y(n33010) );
  NAND2xp33_ASAP7_75t_SL U28287 ( .A(n33012), .B(n22386), .Y(n33013) );
  NAND2xp33_ASAP7_75t_SL U28288 ( .A(n33015), .B(n22386), .Y(n33016) );
  NAND2xp33_ASAP7_75t_SL U28289 ( .A(n33018), .B(n22386), .Y(n33019) );
  NAND2xp33_ASAP7_75t_SL U28290 ( .A(n33021), .B(n22386), .Y(n33022) );
  NAND2xp33_ASAP7_75t_SL U28291 ( .A(n33024), .B(n22386), .Y(n33025) );
  INVx1_ASAP7_75t_SL U28292 ( .A(mult_x_1196_n1661), .Y(n22759) );
  NAND2xp33_ASAP7_75t_SL U28293 ( .A(n33027), .B(n22386), .Y(n33028) );
  OAI21xp33_ASAP7_75t_SL U28294 ( .A1(n29816), .A2(n29868), .B(n29172), .Y(
        n29175) );
  NAND2xp33_ASAP7_75t_SL U28295 ( .A(n33030), .B(n22386), .Y(n33031) );
  NAND2xp33_ASAP7_75t_SL U28296 ( .A(n33034), .B(n22386), .Y(n33035) );
  XNOR2xp5_ASAP7_75t_SL U28297 ( .A(add_x_735_n11), .B(add_x_735_n107), .Y(
        u0_0_leon3x0_p0_dci[29]) );
  AOI21xp33_ASAP7_75t_SL U28298 ( .A1(n31478), .A2(n31477), .B(n31476), .Y(
        n31482) );
  NAND2xp33_ASAP7_75t_SL U28299 ( .A(n22398), .B(u0_0_leon3x0_p0_dci[24]), .Y(
        n25805) );
  XNOR2xp5_ASAP7_75t_SL U28300 ( .A(add_x_735_n5), .B(add_x_735_n49), .Y(
        u0_0_leon3x0_p0_dci[35]) );
  NAND2xp33_ASAP7_75t_SL U28301 ( .A(n33037), .B(n22386), .Y(n33038) );
  XNOR2xp5_ASAP7_75t_SL U28302 ( .A(add_x_735_n14), .B(add_x_735_n132), .Y(
        u0_0_leon3x0_p0_dci[26]) );
  XNOR2xp5_ASAP7_75t_SL U28303 ( .A(add_x_735_n23), .B(add_x_735_n211), .Y(
        u0_0_leon3x0_p0_dci[17]) );
  NAND2xp33_ASAP7_75t_SL U28304 ( .A(n33041), .B(n22386), .Y(n33042) );
  NAND2xp33_ASAP7_75t_SL U28305 ( .A(n33044), .B(n22386), .Y(n33045) );
  NAND2xp5_ASAP7_75t_SL U28306 ( .A(n30575), .B(n29913), .Y(n31045) );
  NAND2xp33_ASAP7_75t_SL U28307 ( .A(n33047), .B(n22386), .Y(n33048) );
  AOI22xp33_ASAP7_75t_SL U28308 ( .A1(n31478), .A2(n31357), .B1(n31356), .B2(
        n31479), .Y(n31358) );
  XNOR2xp5_ASAP7_75t_SL U28309 ( .A(add_x_735_n21), .B(add_x_735_n193), .Y(
        u0_0_leon3x0_p0_dci[19]) );
  INVxp67_ASAP7_75t_SL U28310 ( .A(n32725), .Y(n32726) );
  OAI21xp33_ASAP7_75t_SL U28311 ( .A1(n22421), .A2(u0_0_leon3x0_p0_dci[3]), 
        .B(n31970), .Y(n3304) );
  INVxp33_ASAP7_75t_SL U28312 ( .A(DP_OP_5187J1_124_3275_n145), .Y(
        DP_OP_5187J1_124_3275_n147) );
  INVxp33_ASAP7_75t_SL U28313 ( .A(DP_OP_5187J1_124_3275_n146), .Y(
        DP_OP_5187J1_124_3275_n148) );
  AOI21xp5_ASAP7_75t_SL U28314 ( .A1(n31742), .A2(n32703), .B(n31741), .Y(
        n32789) );
  NOR2x1_ASAP7_75t_SL U28315 ( .A(n24867), .B(n24868), .Y(n25214) );
  INVxp33_ASAP7_75t_SL U28316 ( .A(DP_OP_5187J1_124_3275_n181), .Y(
        DP_OP_5187J1_124_3275_n179) );
  INVxp67_ASAP7_75t_SL U28317 ( .A(DP_OP_5187J1_124_3275_n182), .Y(
        DP_OP_5187J1_124_3275_n180) );
  INVxp67_ASAP7_75t_SL U28318 ( .A(mult_x_1196_n758), .Y(mult_x_1196_n756) );
  AOI21xp33_ASAP7_75t_SL U28319 ( .A1(n30473), .A2(n31342), .B(n30468), .Y(
        n31345) );
  INVxp33_ASAP7_75t_SL U28320 ( .A(DP_OP_5187J1_124_3275_n277), .Y(
        DP_OP_5187J1_124_3275_n279) );
  INVxp33_ASAP7_75t_SL U28321 ( .A(DP_OP_5187J1_124_3275_n276), .Y(
        DP_OP_5187J1_124_3275_n278) );
  INVxp67_ASAP7_75t_SL U28322 ( .A(DP_OP_5187J1_124_3275_n72), .Y(
        DP_OP_5187J1_124_3275_n70) );
  INVxp67_ASAP7_75t_SL U28323 ( .A(DP_OP_5187J1_124_3275_n93), .Y(
        DP_OP_5187J1_124_3275_n312) );
  INVxp33_ASAP7_75t_SL U28324 ( .A(DP_OP_5187J1_124_3275_n282), .Y(
        DP_OP_5187J1_124_3275_n334) );
  INVxp67_ASAP7_75t_SL U28325 ( .A(add_x_746_n2), .Y(add_x_746_n34) );
  INVxp67_ASAP7_75t_SL U28326 ( .A(DP_OP_5187J1_124_3275_n121), .Y(
        DP_OP_5187J1_124_3275_n119) );
  INVxp67_ASAP7_75t_SL U28327 ( .A(DP_OP_5187J1_124_3275_n120), .Y(
        DP_OP_5187J1_124_3275_n315) );
  BUFx2_ASAP7_75t_SL U28328 ( .A(n22609), .Y(n22513) );
  INVx1_ASAP7_75t_SL U28329 ( .A(n32829), .Y(n32830) );
  NAND2xp33_ASAP7_75t_SL U28330 ( .A(n30885), .B(n31479), .Y(n30887) );
  INVxp67_ASAP7_75t_SL U28331 ( .A(DP_OP_5187J1_124_3275_n159), .Y(
        DP_OP_5187J1_124_3275_n157) );
  OAI22xp33_ASAP7_75t_SL U28332 ( .A1(n30577), .A2(n30576), .B1(n30575), .B2(
        n30574), .Y(n30579) );
  BUFx2_ASAP7_75t_SL U28333 ( .A(mult_x_1196_n1407), .Y(n22581) );
  AOI22xp33_ASAP7_75t_SL U28334 ( .A1(u0_0_leon3x0_p0_iu_v_E__RFE2_), .A2(
        n24648), .B1(n32175), .B2(n32174), .Y(n2463) );
  NAND2xp33_ASAP7_75t_SL U28335 ( .A(n22379), .B(n31969), .Y(n31970) );
  INVxp67_ASAP7_75t_SL U28336 ( .A(DP_OP_5187J1_124_3275_n63), .Y(
        DP_OP_5187J1_124_3275_n61) );
  INVxp67_ASAP7_75t_SL U28337 ( .A(DP_OP_5187J1_124_3275_n288), .Y(
        DP_OP_5187J1_124_3275_n286) );
  NAND2xp33_ASAP7_75t_SL U28338 ( .A(n31005), .B(n31479), .Y(n31007) );
  INVxp33_ASAP7_75t_SL U28339 ( .A(DP_OP_5187J1_124_3275_n293), .Y(
        DP_OP_5187J1_124_3275_n336) );
  OAI21xp5_ASAP7_75t_SL U28340 ( .A1(n25065), .A2(n29921), .B(n25064), .Y(
        n25071) );
  INVxp67_ASAP7_75t_SL U28341 ( .A(mult_x_1196_n294), .Y(mult_x_1196_n775) );
  NAND2xp33_ASAP7_75t_SL U28342 ( .A(n31740), .B(n32707), .Y(n31741) );
  INVxp67_ASAP7_75t_SL U28343 ( .A(DP_OP_5187J1_124_3275_n51), .Y(
        DP_OP_5187J1_124_3275_n308) );
  AOI22xp33_ASAP7_75t_SL U28344 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__15_), 
        .A2(n31364), .B1(n31035), .B2(n31043), .Y(n31036) );
  OAI21xp33_ASAP7_75t_SL U28345 ( .A1(n28055), .A2(n28054), .B(n28053), .Y(
        n5591) );
  OAI21xp33_ASAP7_75t_SL U28346 ( .A1(DP_OP_5187J1_124_3275_n227), .A2(
        DP_OP_5187J1_124_3275_n219), .B(DP_OP_5187J1_124_3275_n220), .Y(
        DP_OP_5187J1_124_3275_n214) );
  OAI21xp33_ASAP7_75t_SL U28347 ( .A1(DP_OP_5187J1_124_3275_n245), .A2(
        DP_OP_5187J1_124_3275_n237), .B(DP_OP_5187J1_124_3275_n238), .Y(
        DP_OP_5187J1_124_3275_n236) );
  AOI21xp5_ASAP7_75t_SL U28348 ( .A1(n30018), .A2(n31034), .B(n25048), .Y(
        n25073) );
  AOI22xp33_ASAP7_75t_SL U28349 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__11_), 
        .A2(n31364), .B1(n30968), .B2(n31043), .Y(n30969) );
  INVxp67_ASAP7_75t_SL U28350 ( .A(n29642), .Y(n29643) );
  NAND2xp5_ASAP7_75t_SL U28351 ( .A(n28950), .B(n28949), .Y(n30473) );
  AOI22xp33_ASAP7_75t_SL U28352 ( .A1(n31824), .A2(n29648), .B1(n31828), .B2(
        u0_0_leon3x0_p0_dci[11]), .Y(n26237) );
  AOI21xp33_ASAP7_75t_SL U28353 ( .A1(u0_0_leon3x0_p0_dci[12]), .A2(n31828), 
        .B(n29890), .Y(n29891) );
  NAND2xp33_ASAP7_75t_SL U28354 ( .A(n29919), .B(n31479), .Y(n29920) );
  NAND2xp33_ASAP7_75t_SL U28355 ( .A(n29979), .B(n29977), .Y(n29978) );
  AOI21xp33_ASAP7_75t_SL U28356 ( .A1(n28924), .A2(n26938), .B(n26888), .Y(
        n26909) );
  INVxp33_ASAP7_75t_SL U28357 ( .A(DP_OP_5187J1_124_3275_n266), .Y(
        DP_OP_5187J1_124_3275_n332) );
  OAI21xp33_ASAP7_75t_SL U28358 ( .A1(DP_OP_5187J1_124_3275_n121), .A2(
        DP_OP_5187J1_124_3275_n113), .B(DP_OP_5187J1_124_3275_n114), .Y(
        DP_OP_5187J1_124_3275_n108) );
  INVx1_ASAP7_75t_SL U28359 ( .A(n32108), .Y(n4406) );
  NAND2xp33_ASAP7_75t_SL U28360 ( .A(n30563), .B(n31479), .Y(n30564) );
  INVxp33_ASAP7_75t_SL U28361 ( .A(DP_OP_5187J1_124_3275_n287), .Y(
        DP_OP_5187J1_124_3275_n335) );
  XNOR2xp5_ASAP7_75t_SL U28362 ( .A(n22931), .B(n22930), .Y(mult_x_1196_n1153)
         );
  INVxp33_ASAP7_75t_SL U28363 ( .A(DP_OP_5187J1_124_3275_n226), .Y(
        DP_OP_5187J1_124_3275_n327) );
  INVxp67_ASAP7_75t_SL U28364 ( .A(DP_OP_5187J1_124_3275_n227), .Y(
        DP_OP_5187J1_124_3275_n225) );
  INVxp33_ASAP7_75t_SL U28365 ( .A(DP_OP_5187J1_124_3275_n187), .Y(
        DP_OP_5187J1_124_3275_n322) );
  NAND2xp33_ASAP7_75t_SL U28366 ( .A(n31480), .B(n31479), .Y(n31481) );
  AOI22xp33_ASAP7_75t_SL U28367 ( .A1(u0_0_leon3x0_p0_iu_r_A__RSEL2__1_), .A2(
        n24648), .B1(n32172), .B2(n32174), .Y(n4051) );
  NAND2xp5_ASAP7_75t_SL U28368 ( .A(n32824), .B(n32770), .Y(n32802) );
  NAND2xp33_ASAP7_75t_SL U28369 ( .A(n22398), .B(u0_0_leon3x0_p0_dci[11]), .Y(
        n26284) );
  OAI21xp33_ASAP7_75t_SL U28370 ( .A1(n28790), .A2(n28789), .B(n28788), .Y(
        n28792) );
  INVxp33_ASAP7_75t_SL U28371 ( .A(DP_OP_5187J1_124_3275_n190), .Y(
        DP_OP_5187J1_124_3275_n323) );
  AOI21xp5_ASAP7_75t_SL U28372 ( .A1(n26292), .A2(n28924), .B(n26291), .Y(
        n26322) );
  OAI21xp33_ASAP7_75t_SL U28373 ( .A1(n32698), .A2(n22393), .B(n32770), .Y(
        n32701) );
  INVxp33_ASAP7_75t_SL U28374 ( .A(DP_OP_5187J1_124_3275_n255), .Y(
        DP_OP_5187J1_124_3275_n330) );
  INVxp33_ASAP7_75t_SL U28375 ( .A(DP_OP_5187J1_124_3275_n244), .Y(
        DP_OP_5187J1_124_3275_n329) );
  INVx1_ASAP7_75t_SL U28376 ( .A(add_x_746_n125), .Y(add_x_746_n124) );
  AOI21xp33_ASAP7_75t_SL U28377 ( .A1(sr1_r_AREA__0_), .A2(n32722), .B(n32698), 
        .Y(n2355) );
  INVx1_ASAP7_75t_SL U28378 ( .A(n32883), .Y(n31693) );
  NAND2xp33_ASAP7_75t_SL U28379 ( .A(n30478), .B(n31479), .Y(n30481) );
  INVxp33_ASAP7_75t_SL U28380 ( .A(DP_OP_5187J1_124_3275_n219), .Y(
        DP_OP_5187J1_124_3275_n326) );
  OAI21xp33_ASAP7_75t_SL U28381 ( .A1(n27208), .A2(n28789), .B(n26275), .Y(
        n26276) );
  INVxp67_ASAP7_75t_SL U28382 ( .A(DP_OP_5187J1_124_3275_n73), .Y(
        DP_OP_5187J1_124_3275_n310) );
  INVxp67_ASAP7_75t_SL U28383 ( .A(mult_x_1196_n1048), .Y(n23740) );
  INVx1_ASAP7_75t_SL U28384 ( .A(mult_x_1196_n301), .Y(n22409) );
  INVx1_ASAP7_75t_SL U28385 ( .A(n32228), .Y(n32417) );
  AOI22xp33_ASAP7_75t_SL U28386 ( .A1(n28762), .A2(n26986), .B1(n28764), .B2(
        n26697), .Y(n26715) );
  INVxp67_ASAP7_75t_SL U28387 ( .A(n25068), .Y(n25048) );
  XOR2xp5_ASAP7_75t_SL U28388 ( .A(n22987), .B(n23515), .Y(mult_x_1196_n1067)
         );
  NAND2xp5_ASAP7_75t_SL U28389 ( .A(n32786), .B(n32697), .Y(n32770) );
  INVxp67_ASAP7_75t_SL U28390 ( .A(n29914), .Y(n25065) );
  NAND2xp5_ASAP7_75t_SL U28391 ( .A(n28764), .B(n26292), .Y(n26281) );
  INVxp67_ASAP7_75t_SL U28392 ( .A(n28411), .Y(n30577) );
  OAI21xp33_ASAP7_75t_SL U28393 ( .A1(n28672), .A2(n28671), .B(n28670), .Y(
        n28673) );
  INVxp67_ASAP7_75t_SL U28394 ( .A(n30573), .Y(n30576) );
  AOI21xp33_ASAP7_75t_SL U28395 ( .A1(n28742), .A2(n28741), .B(n28740), .Y(
        n28743) );
  OAI22xp33_ASAP7_75t_SL U28396 ( .A1(n28921), .A2(n28854), .B1(n28914), .B2(
        n26290), .Y(n26291) );
  INVx1_ASAP7_75t_SL U28397 ( .A(n32336), .Y(n29847) );
  NOR2x1_ASAP7_75t_SL U28398 ( .A(n24678), .B(n30648), .Y(n30595) );
  OAI22xp33_ASAP7_75t_SL U28399 ( .A1(n28790), .A2(n26405), .B1(n27208), .B2(
        n28443), .Y(n26406) );
  NAND2xp33_ASAP7_75t_SL U28400 ( .A(n24343), .B(n24400), .Y(n24344) );
  AOI22xp33_ASAP7_75t_SL U28401 ( .A1(n29605), .A2(n28763), .B1(n30632), .B2(
        n28718), .Y(n28744) );
  INVxp67_ASAP7_75t_SL U28402 ( .A(add_x_746_n58), .Y(add_x_746_n59) );
  OAI22xp33_ASAP7_75t_SL U28403 ( .A1(n28921), .A2(n28420), .B1(n26887), .B2(
        n24427), .Y(n26888) );
  INVxp67_ASAP7_75t_SL U28404 ( .A(u0_0_leon3x0_p0_div0_b[0]), .Y(
        DP_OP_5187J1_124_3275_n306) );
  AOI22xp33_ASAP7_75t_SL U28405 ( .A1(n30632), .A2(n29602), .B1(n28742), .B2(
        n29604), .Y(n25913) );
  INVxp67_ASAP7_75t_SL U28406 ( .A(add_x_746_n145), .Y(add_x_746_n144) );
  OAI21xp33_ASAP7_75t_SL U28407 ( .A1(n29675), .A2(n29475), .B(n18845), .Y(
        n29642) );
  NAND2xp33_ASAP7_75t_SL U28408 ( .A(n29605), .B(n28741), .Y(n27120) );
  INVxp67_ASAP7_75t_SL U28409 ( .A(n28741), .Y(n28789) );
  AOI22xp33_ASAP7_75t_SL U28410 ( .A1(n31824), .A2(n29676), .B1(n31828), .B2(
        u0_0_leon3x0_p0_dci[10]), .Y(n29677) );
  NAND2xp5_ASAP7_75t_SL U28411 ( .A(n28054), .B(n28055), .Y(n28053) );
  AOI22xp33_ASAP7_75t_SL U28412 ( .A1(n28764), .A2(n28675), .B1(n28762), .B2(
        n28615), .Y(n28616) );
  INVx1_ASAP7_75t_SL U28413 ( .A(mult_x_1196_n1901), .Y(n24214) );
  AOI22xp33_ASAP7_75t_SL U28414 ( .A1(n28855), .A2(n26986), .B1(n28924), .B2(
        n27077), .Y(n27006) );
  NOR2xp33_ASAP7_75t_SRAM U28415 ( .A(n32189), .B(n32188), .Y(n32191) );
  OAI22xp33_ASAP7_75t_SL U28416 ( .A1(n28618), .A2(n26151), .B1(n26150), .B2(
        n28671), .Y(n26159) );
  INVxp67_ASAP7_75t_SL U28417 ( .A(n32711), .Y(n31756) );
  INVx1_ASAP7_75t_SL U28418 ( .A(n32339), .Y(n29993) );
  AOI22xp33_ASAP7_75t_SL U28419 ( .A1(n29605), .A2(n28761), .B1(n28742), .B2(
        n28718), .Y(n27159) );
  OAI22xp33_ASAP7_75t_SL U28420 ( .A1(n28914), .A2(n28420), .B1(n28419), .B2(
        n24427), .Y(n28448) );
  AOI21xp33_ASAP7_75t_SL U28421 ( .A1(n28764), .A2(n26986), .B(n25801), .Y(
        n25802) );
  NAND2xp33_ASAP7_75t_SL U28422 ( .A(n29605), .B(n29604), .Y(n29606) );
  INVxp67_ASAP7_75t_SL U28423 ( .A(n25069), .Y(n25053) );
  AOI22xp33_ASAP7_75t_SL U28424 ( .A1(n29603), .A2(n26986), .B1(n29605), .B2(
        n26697), .Y(n25835) );
  OAI21xp33_ASAP7_75t_SL U28425 ( .A1(n32875), .A2(n2292), .B(n31709), .Y(
        n17903) );
  O2A1O1Ixp33_ASAP7_75t_SL U28426 ( .A1(n28990), .A2(n28989), .B(n28988), .C(
        n28992), .Y(n28991) );
  OA21x2_ASAP7_75t_SL U28427 ( .A1(n28920), .A2(n28858), .B(n28765), .Y(n28766) );
  INVx1_ASAP7_75t_SL U28428 ( .A(mult_x_1196_n884), .Y(mult_x_1196_n878) );
  AOI21xp33_ASAP7_75t_SL U28429 ( .A1(n29605), .A2(n28440), .B(n25504), .Y(
        n25505) );
  OAI22xp33_ASAP7_75t_SL U28430 ( .A1(n28914), .A2(n28667), .B1(n28920), .B2(
        n28666), .Y(n28674) );
  OAI21xp33_ASAP7_75t_SL U28431 ( .A1(n32696), .A2(n32695), .B(n32704), .Y(
        n32697) );
  OR2x2_ASAP7_75t_SL U28432 ( .A(n32718), .B(n32875), .Y(n33053) );
  INVxp67_ASAP7_75t_SL U28433 ( .A(n28503), .Y(n27077) );
  AOI22xp33_ASAP7_75t_SL U28434 ( .A1(n28762), .A2(n28499), .B1(n28764), .B2(
        n27078), .Y(n27005) );
  XNOR2xp5_ASAP7_75t_SL U28435 ( .A(n23284), .B(n23283), .Y(mult_x_1196_n1027)
         );
  O2A1O1Ixp33_ASAP7_75t_SL U28436 ( .A1(n26903), .A2(n26902), .B(n24634), .C(
        n26901), .Y(n26905) );
  NAND2xp5_ASAP7_75t_SL U28437 ( .A(n32700), .B(n32703), .Y(n32702) );
  NAND2xp33_ASAP7_75t_SL U28438 ( .A(n32751), .B(n32703), .Y(n32699) );
  NAND2xp33_ASAP7_75t_SL U28439 ( .A(n32879), .B(n32824), .Y(n32788) );
  NAND2xp5_ASAP7_75t_SL U28440 ( .A(n24233), .B(n24235), .Y(n24236) );
  NAND2xp33_ASAP7_75t_SL U28441 ( .A(n29605), .B(n28499), .Y(n26435) );
  INVxp67_ASAP7_75t_SL U28442 ( .A(n30214), .Y(n30223) );
  INVxp33_ASAP7_75t_SL U28443 ( .A(add_x_746_n116), .Y(add_x_746_n115) );
  AOI22xp33_ASAP7_75t_SL U28444 ( .A1(n28855), .A2(n30631), .B1(n28924), .B2(
        n28876), .Y(n28856) );
  OAI21xp33_ASAP7_75t_SL U28445 ( .A1(n30625), .A2(n30214), .B(n29599), .Y(
        n29600) );
  INVx1_ASAP7_75t_SL U28446 ( .A(n26914), .Y(n28420) );
  NAND2xp33_ASAP7_75t_SL U28447 ( .A(n28742), .B(n28440), .Y(n28441) );
  OAI22xp33_ASAP7_75t_SL U28448 ( .A1(n28921), .A2(n28971), .B1(n28920), .B2(
        n30627), .Y(n28922) );
  AOI22xp33_ASAP7_75t_SL U28449 ( .A1(n28742), .A2(n28498), .B1(n30632), .B2(
        n28440), .Y(n26437) );
  AOI22xp33_ASAP7_75t_SL U28450 ( .A1(n28742), .A2(n28499), .B1(n29603), .B2(
        n28498), .Y(n28500) );
  NOR2x1_ASAP7_75t_SL U28451 ( .A(n22657), .B(n22656), .Y(mult_x_1196_n1044)
         );
  AOI22xp33_ASAP7_75t_SL U28452 ( .A1(n28764), .A2(n28763), .B1(n28762), .B2(
        n28761), .Y(n28765) );
  MAJx2_ASAP7_75t_SL U28453 ( .A(mult_x_1196_n945), .B(mult_x_1196_n958), .C(
        mult_x_1196_n943), .Y(mult_x_1196_n937) );
  NAND2xp33_ASAP7_75t_SL U28454 ( .A(n28987), .B(n28971), .Y(n28972) );
  NAND2xp33_ASAP7_75t_SL U28455 ( .A(n28764), .B(n28669), .Y(n28670) );
  NAND2xp33_ASAP7_75t_SL U28456 ( .A(n28987), .B(n30627), .Y(n28988) );
  OAI21xp33_ASAP7_75t_SL U28457 ( .A1(n23065), .A2(n23068), .B(n23066), .Y(
        n23064) );
  OAI22xp33_ASAP7_75t_SL U28458 ( .A1(n30691), .A2(n30690), .B1(n23229), .B2(
        u0_0_leon3x0_p0_iu_v_M__IRQEN2_), .Y(n3385) );
  NAND2xp33_ASAP7_75t_SL U28459 ( .A(n25440), .B(n25439), .Y(n29918) );
  OAI21xp33_ASAP7_75t_SL U28460 ( .A1(n28502), .A2(n28913), .B(n26317), .Y(
        n26320) );
  INVx1_ASAP7_75t_SL U28461 ( .A(n32233), .Y(n32432) );
  INVxp33_ASAP7_75t_SL U28462 ( .A(n31034), .Y(n31037) );
  OAI21xp33_ASAP7_75t_SL U28463 ( .A1(n27524), .A2(n27508), .B(n27499), .Y(
        n27509) );
  AND4x1_ASAP7_75t_SL U28464 ( .A(n31798), .B(n33033), .C(n33040), .D(n32751), 
        .Y(n25258) );
  OAI21xp33_ASAP7_75t_SL U28465 ( .A1(n27209), .A2(n27208), .B(n27207), .Y(
        n27212) );
  OAI22xp33_ASAP7_75t_SL U28466 ( .A1(n28914), .A2(n26670), .B1(n28921), .B2(
        n27210), .Y(n26560) );
  INVx1_ASAP7_75t_SL U28467 ( .A(n32342), .Y(n30556) );
  AOI21xp33_ASAP7_75t_SL U28468 ( .A1(n28669), .A2(n29603), .B(n27158), .Y(
        n27160) );
  AOI22xp33_ASAP7_75t_SL U28469 ( .A1(n27096), .A2(n24634), .B1(n28762), .B2(
        n28669), .Y(n27125) );
  INVxp33_ASAP7_75t_SL U28470 ( .A(n29979), .Y(n29986) );
  OAI22xp33_ASAP7_75t_SL U28471 ( .A1(n28503), .A2(n28914), .B1(n28618), .B2(
        n25800), .Y(n25801) );
  INVxp67_ASAP7_75t_SL U28472 ( .A(n26709), .Y(n25836) );
  INVxp67_ASAP7_75t_SL U28473 ( .A(n32190), .Y(n30943) );
  INVxp67_ASAP7_75t_SL U28474 ( .A(n26670), .Y(n26697) );
  AOI21xp33_ASAP7_75t_SL U28475 ( .A1(n28761), .A2(n28742), .B(n27119), .Y(
        n27121) );
  NAND2xp5_ASAP7_75t_SL U28476 ( .A(n23429), .B(n23427), .Y(n23426) );
  NAND2xp5_ASAP7_75t_SL U28477 ( .A(n24694), .B(n32824), .Y(n32711) );
  INVxp67_ASAP7_75t_SL U28478 ( .A(mult_x_1196_n912), .Y(n22911) );
  NAND2xp5_ASAP7_75t_SL U28479 ( .A(n25440), .B(n31035), .Y(n25068) );
  INVxp33_ASAP7_75t_SL U28480 ( .A(n28440), .Y(n26405) );
  INVxp67_ASAP7_75t_SL U28481 ( .A(n28761), .Y(n28745) );
  INVx1_ASAP7_75t_SL U28482 ( .A(n32343), .Y(n31031) );
  INVxp33_ASAP7_75t_SL U28483 ( .A(add_x_746_n71), .Y(add_x_746_n70) );
  NAND2xp33_ASAP7_75t_SL U28484 ( .A(n32879), .B(n32875), .Y(n31709) );
  NAND2xp5_ASAP7_75t_SL U28485 ( .A(n26144), .B(n26143), .Y(n28675) );
  OAI22xp33_ASAP7_75t_SL U28486 ( .A1(n28921), .A2(n28667), .B1(n28914), .B2(
        n27210), .Y(n26158) );
  INVxp33_ASAP7_75t_SL U28487 ( .A(n32875), .Y(n32722) );
  XNOR2xp5_ASAP7_75t_SL U28488 ( .A(n23192), .B(n23719), .Y(n23596) );
  NAND2xp33_ASAP7_75t_SL U28489 ( .A(n24684), .B(n30690), .Y(n31968) );
  NAND2xp33_ASAP7_75t_SL U28490 ( .A(n28855), .B(n28669), .Y(n28617) );
  INVxp67_ASAP7_75t_SL U28491 ( .A(n28666), .Y(n28718) );
  NAND2xp33_ASAP7_75t_SL U28492 ( .A(n29603), .B(n26709), .Y(n26710) );
  OAI22xp33_ASAP7_75t_SL U28493 ( .A1(n28618), .A2(n26670), .B1(n28920), .B2(
        n27210), .Y(n26671) );
  NAND2xp33_ASAP7_75t_SL U28494 ( .A(n31474), .B(n30021), .Y(n29917) );
  AOI21xp33_ASAP7_75t_SL U28495 ( .A1(sr1_sdi_HWRITE_), .A2(n32786), .B(n31705), .Y(n2363) );
  INVx1_ASAP7_75t_SL U28496 ( .A(n23719), .Y(n23108) );
  INVxp33_ASAP7_75t_SL U28497 ( .A(n30477), .Y(n30478) );
  INVxp67_ASAP7_75t_SL U28498 ( .A(n28763), .Y(n26290) );
  INVx1_ASAP7_75t_SL U28499 ( .A(n28858), .Y(n26292) );
  OAI22xp33_ASAP7_75t_SL U28500 ( .A1(n28502), .A2(n28667), .B1(n28790), .B2(
        n27210), .Y(n27211) );
  INVx1_ASAP7_75t_SL U28501 ( .A(mult_x_1196_n843), .Y(mult_x_1196_n840) );
  AOI21xp33_ASAP7_75t_SL U28502 ( .A1(n28894), .A2(n30672), .B(n27076), .Y(
        n27082) );
  NAND2xp33_ASAP7_75t_SL U28503 ( .A(n29605), .B(n27078), .Y(n27080) );
  INVx1_ASAP7_75t_SL U28504 ( .A(n29916), .Y(n25067) );
  OAI22xp33_ASAP7_75t_SL U28505 ( .A1(n2842), .A2(n31843), .B1(n29568), .B2(
        n24640), .Y(n26644) );
  INVxp67_ASAP7_75t_SL U28506 ( .A(mult_x_1196_n2213), .Y(n23068) );
  AOI21xp33_ASAP7_75t_SL U28507 ( .A1(n32776), .A2(n32775), .B(n32774), .Y(
        n32777) );
  AOI22xp33_ASAP7_75t_SL U28508 ( .A1(n32773), .A2(n33014), .B1(n32775), .B2(
        n33052), .Y(n32764) );
  INVx1_ASAP7_75t_SL U28509 ( .A(u0_0_leon3x0_p0_iu_fe_pc_14_), .Y(
        add_x_746_n99) );
  AOI21xp33_ASAP7_75t_SL U28510 ( .A1(n33029), .A2(n32753), .B(
        sr1_r_MCFG2__RAMBANKSZ__3_), .Y(n32754) );
  INVx1_ASAP7_75t_SL U28511 ( .A(n32210), .Y(n32365) );
  OAI22xp33_ASAP7_75t_SL U28512 ( .A1(n4497), .A2(n31843), .B1(n31526), .B2(
        n31841), .Y(n31527) );
  INVx1_ASAP7_75t_SL U28513 ( .A(n32211), .Y(n32366) );
  INVxp33_ASAP7_75t_SL U28514 ( .A(n24889), .Y(n24890) );
  AOI21xp33_ASAP7_75t_SL U28515 ( .A1(n33017), .A2(n2924), .B(n32774), .Y(
        n32755) );
  OAI22xp33_ASAP7_75t_SL U28516 ( .A1(n4385), .A2(n31843), .B1(n31842), .B2(
        n24640), .Y(n31844) );
  OAI22xp33_ASAP7_75t_SL U28517 ( .A1(n2844), .A2(n31843), .B1(n27493), .B2(
        n24640), .Y(n26648) );
  OAI22xp33_ASAP7_75t_SL U28518 ( .A1(n2846), .A2(n31843), .B1(n28108), .B2(
        n24640), .Y(n26652) );
  NAND2xp33_ASAP7_75t_SL U28519 ( .A(n28742), .B(n26938), .Y(n26939) );
  O2A1O1Ixp33_ASAP7_75t_SL U28520 ( .A1(n26936), .A2(n26935), .B(n24634), .C(
        n26934), .Y(n26941) );
  INVx1_ASAP7_75t_SL U28521 ( .A(u0_0_leon3x0_p0_iu_fe_pc_20_), .Y(
        add_x_746_n68) );
  INVx1_ASAP7_75t_SL U28522 ( .A(n29915), .Y(n25438) );
  INVx1_ASAP7_75t_SL U28523 ( .A(u0_0_leon3x0_p0_iu_fe_pc_27_), .Y(
        add_x_746_n27) );
  OAI22xp5_ASAP7_75t_SL U28524 ( .A1(n25396), .A2(n31967), .B1(n25395), .B2(
        n25394), .Y(n25397) );
  AOI22xp33_ASAP7_75t_SL U28525 ( .A1(n32772), .A2(n33039), .B1(n32771), .B2(
        n33026), .Y(n32763) );
  INVxp67_ASAP7_75t_SL U28526 ( .A(u0_0_leon3x0_p0_iu_fe_pc_9_), .Y(
        add_x_746_n129) );
  INVxp67_ASAP7_75t_SL U28527 ( .A(u0_0_leon3x0_p0_iu_fe_pc_15_), .Y(
        add_x_746_n96) );
  NAND2xp5_ASAP7_75t_SL U28528 ( .A(n31889), .B(n26203), .Y(n26205) );
  OAI22xp33_ASAP7_75t_SL U28529 ( .A1(n4363), .A2(n31843), .B1(n26544), .B2(
        n24640), .Y(n26545) );
  INVx1_ASAP7_75t_SL U28530 ( .A(n32212), .Y(n32375) );
  INVx1_ASAP7_75t_SL U28531 ( .A(u0_0_leon3x0_p0_iu_fe_pc_22_), .Y(
        add_x_746_n56) );
  INVxp33_ASAP7_75t_SL U28532 ( .A(n27078), .Y(n25800) );
  OAI22xp33_ASAP7_75t_SL U28533 ( .A1(n1792), .A2(n31843), .B1(n30139), .B2(
        n24640), .Y(n26621) );
  OAI22xp33_ASAP7_75t_SL U28534 ( .A1(n2840), .A2(n31843), .B1(n29510), .B2(
        n24640), .Y(n26641) );
  OAI22xp33_ASAP7_75t_SL U28535 ( .A1(n4669), .A2(n31843), .B1(n26492), .B2(
        n24640), .Y(n26493) );
  NAND2xp33_ASAP7_75t_SL U28536 ( .A(n29836), .B(n31542), .Y(n29622) );
  INVxp67_ASAP7_75t_SL U28537 ( .A(u0_0_leon3x0_p0_iu_fe_pc_11_), .Y(
        add_x_746_n120) );
  OAI22xp33_ASAP7_75t_SL U28538 ( .A1(n4354), .A2(n31843), .B1(n29570), .B2(
        n31841), .Y(n29571) );
  INVx1_ASAP7_75t_SL U28539 ( .A(u0_0_leon3x0_p0_iu_fe_pc_23_), .Y(
        add_x_746_n51) );
  OAI22xp33_ASAP7_75t_SL U28540 ( .A1(n4531), .A2(n31843), .B1(n30894), .B2(
        n31841), .Y(n30895) );
  OAI22xp33_ASAP7_75t_SL U28541 ( .A1(n4635), .A2(n31843), .B1(n29389), .B2(
        n24640), .Y(n26592) );
  INVxp67_ASAP7_75t_SL U28542 ( .A(n22480), .Y(n22479) );
  OAI22xp33_ASAP7_75t_SL U28543 ( .A1(n2838), .A2(n31843), .B1(n30073), .B2(
        n24640), .Y(n26634) );
  NAND2xp5_ASAP7_75t_SL U28544 ( .A(n30632), .B(n18794), .Y(n26940) );
  AOI22xp33_ASAP7_75t_SL U28545 ( .A1(n32775), .A2(n33046), .B1(n32771), .B2(
        n33020), .Y(n32766) );
  AOI21xp33_ASAP7_75t_SL U28546 ( .A1(n26316), .A2(n28894), .B(n26315), .Y(
        n26317) );
  AOI21xp33_ASAP7_75t_SL U28547 ( .A1(add_x_735_n186), .A2(add_x_735_n167), 
        .B(add_x_735_n168), .Y(add_x_735_n166) );
  AOI22xp33_ASAP7_75t_SL U28548 ( .A1(n32773), .A2(n33020), .B1(n32772), .B2(
        n33046), .Y(n32778) );
  NAND2xp5_ASAP7_75t_SL U28549 ( .A(n30937), .B(n30936), .Y(n32190) );
  INVxp67_ASAP7_75t_SL U28550 ( .A(mult_x_1196_n958), .Y(n22559) );
  NAND2xp5_ASAP7_75t_SL U28551 ( .A(n29152), .B(n29151), .Y(n30214) );
  NAND2xp5_ASAP7_75t_SL U28552 ( .A(n28762), .B(n27078), .Y(n25838) );
  INVx1_ASAP7_75t_SL U28553 ( .A(n32209), .Y(n32360) );
  AOI21xp33_ASAP7_75t_SL U28554 ( .A1(n33008), .A2(n32773), .B(
        sr1_r_MCFG2__RAMBANKSZ__1_), .Y(n32765) );
  NAND2xp33_ASAP7_75t_SL U28555 ( .A(n29916), .B(n29915), .Y(n30021) );
  INVx1_ASAP7_75t_SL U28556 ( .A(u0_0_leon3x0_p0_iu_fe_pc_25_), .Y(
        add_x_746_n39) );
  INVxp67_ASAP7_75t_SL U28557 ( .A(u0_0_leon3x0_p0_iu_fe_pc_8_), .Y(
        add_x_746_n133) );
  NAND2xp33_ASAP7_75t_SL U28558 ( .A(n27517), .B(n27516), .Y(n27518) );
  OAI22xp33_ASAP7_75t_SL U28559 ( .A1(n2233), .A2(n31843), .B1(n28116), .B2(
        n24640), .Y(n28117) );
  INVxp67_ASAP7_75t_SL U28560 ( .A(u0_0_leon3x0_p0_iu_fe_pc_19_), .Y(
        add_x_746_n75) );
  AND4x1_ASAP7_75t_SL U28561 ( .A(n33014), .B(n33026), .C(n33039), .D(n32776), 
        .Y(n31799) );
  NAND2xp33_ASAP7_75t_SL U28562 ( .A(n28132), .B(n26597), .Y(n26598) );
  INVxp67_ASAP7_75t_SL U28563 ( .A(n26938), .Y(n25915) );
  OAI22xp33_ASAP7_75t_SL U28564 ( .A1(n4741), .A2(n31843), .B1(n26479), .B2(
        n24640), .Y(n26480) );
  OAI22xp33_ASAP7_75t_SL U28565 ( .A1(n4573), .A2(n31843), .B1(n31641), .B2(
        n31841), .Y(n31642) );
  OAI22xp33_ASAP7_75t_SL U28566 ( .A1(n1626), .A2(n31843), .B1(n30833), .B2(
        n24640), .Y(n26628) );
  OAI22xp33_ASAP7_75t_SL U28567 ( .A1(n1771), .A2(n31843), .B1(n26655), .B2(
        n24640), .Y(n26656) );
  OAI22xp33_ASAP7_75t_SL U28568 ( .A1(n1728), .A2(n31843), .B1(n31197), .B2(
        n24640), .Y(n26631) );
  OAI22xp33_ASAP7_75t_SL U28569 ( .A1(n4624), .A2(n31843), .B1(n31368), .B2(
        n31841), .Y(n31369) );
  OAI21xp33_ASAP7_75t_SL U28570 ( .A1(n23229), .A2(u0_0_leon3x0_p0_divi[36]), 
        .B(n30427), .Y(n3920) );
  NOR2x1_ASAP7_75t_SL U28571 ( .A(n22380), .B(n32729), .Y(n29937) );
  INVx1_ASAP7_75t_SL U28572 ( .A(u0_0_leon3x0_p0_iu_fe_pc_30_), .Y(
        add_x_746_n8) );
  OAI22xp33_ASAP7_75t_SL U28573 ( .A1(n1775), .A2(n31843), .B1(n31496), .B2(
        n31841), .Y(n31497) );
  INVxp67_ASAP7_75t_SL U28574 ( .A(u0_0_leon3x0_p0_iu_fe_pc_5_), .Y(
        add_x_746_n148) );
  NAND2xp5_ASAP7_75t_SL U28575 ( .A(n28924), .B(n28497), .Y(n26441) );
  INVx1_ASAP7_75t_SL U28576 ( .A(mult_x_1196_n842), .Y(mult_x_1196_n837) );
  AOI21xp33_ASAP7_75t_SL U28577 ( .A1(n28405), .A2(n26597), .B(n26485), .Y(
        n26487) );
  OAI22xp33_ASAP7_75t_SL U28578 ( .A1(n1752), .A2(n31843), .B1(n29236), .B2(
        n24640), .Y(n26605) );
  INVxp33_ASAP7_75t_SL U28579 ( .A(n28619), .Y(n28642) );
  INVxp67_ASAP7_75t_SL U28580 ( .A(u0_0_leon3x0_p0_iu_fe_pc_13_), .Y(
        add_x_746_n108) );
  NOR2x1_ASAP7_75t_SL U28581 ( .A(n23110), .B(n23109), .Y(n23719) );
  INVxp33_ASAP7_75t_SL U28582 ( .A(u0_0_leon3x0_p0_iu_fe_pc_3_), .Y(
        add_x_746_n155) );
  NAND2xp33_ASAP7_75t_SL U28583 ( .A(n29836), .B(n31054), .Y(n29844) );
  NAND2xp33_ASAP7_75t_SL U28584 ( .A(n31049), .B(n31542), .Y(n31051) );
  INVx1_ASAP7_75t_SL U28585 ( .A(u0_0_leon3x0_p0_iu_fe_pc_16_), .Y(
        add_x_746_n89) );
  OAI21xp33_ASAP7_75t_SL U28586 ( .A1(n28692), .A2(n24427), .B(n28691), .Y(
        n28694) );
  OAI22xp33_ASAP7_75t_SL U28587 ( .A1(n4456), .A2(n31843), .B1(n30978), .B2(
        n24640), .Y(n26617) );
  INVxp67_ASAP7_75t_SL U28588 ( .A(n33017), .Y(n30538) );
  OAI22xp33_ASAP7_75t_SL U28589 ( .A1(n1741), .A2(n31843), .B1(n29744), .B2(
        n24640), .Y(n26624) );
  OAI22xp33_ASAP7_75t_SL U28590 ( .A1(n1630), .A2(n31843), .B1(n30780), .B2(
        n24640), .Y(n26637) );
  INVxp33_ASAP7_75t_SL U28591 ( .A(u0_0_leon3x0_p0_iu_fe_pc_4_), .Y(
        add_x_746_n151) );
  INVx1_ASAP7_75t_SL U28592 ( .A(u0_0_leon3x0_p0_iu_fe_pc_17_), .Y(
        add_x_746_n84) );
  OAI22xp33_ASAP7_75t_SL U28593 ( .A1(n1634), .A2(n31843), .B1(n29851), .B2(
        n24640), .Y(n26608) );
  NAND2xp33_ASAP7_75t_SL U28594 ( .A(n24335), .B(n24403), .Y(n24336) );
  OAI22xp33_ASAP7_75t_SL U28595 ( .A1(n4032), .A2(n31843), .B1(n26547), .B2(
        n24640), .Y(n26548) );
  OAI21xp33_ASAP7_75t_SL U28596 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__16_), .A2(n31001), .B(
        n26669), .Y(n30477) );
  OAI22xp33_ASAP7_75t_SL U28597 ( .A1(n28986), .A2(n25468), .B1(n28869), .B2(
        n25467), .Y(n25474) );
  OAI22xp33_ASAP7_75t_SL U28598 ( .A1(n4770), .A2(n31843), .B1(n24640), .B2(
        n26474), .Y(n26475) );
  INVxp67_ASAP7_75t_SL U28599 ( .A(n32735), .Y(n31314) );
  NAND2xp33_ASAP7_75t_SL U28600 ( .A(n31828), .B(
        u0_0_leon3x0_p0_iu_ex_jump_address_2_), .Y(n32666) );
  INVxp67_ASAP7_75t_SL U28601 ( .A(u0_0_leon3x0_p0_iu_fe_pc_18_), .Y(
        add_x_746_n78) );
  INVxp67_ASAP7_75t_SL U28602 ( .A(n33011), .Y(n30515) );
  AOI22xp33_ASAP7_75t_SL U28603 ( .A1(n31824), .A2(n29476), .B1(n31828), .B2(
        u0_0_leon3x0_p0_dci[9]), .Y(n29477) );
  OAI21xp33_ASAP7_75t_SL U28604 ( .A1(n30625), .A2(n29167), .B(n28494), .Y(
        n28495) );
  OAI22xp33_ASAP7_75t_SL U28605 ( .A1(n4614), .A2(n31843), .B1(n26498), .B2(
        n24640), .Y(n26499) );
  AOI21xp33_ASAP7_75t_SL U28606 ( .A1(n28967), .A2(n25910), .B(n25909), .Y(
        n25911) );
  NAND2xp5_ASAP7_75t_SL U28607 ( .A(n26149), .B(n26148), .Y(n28615) );
  NAND2xp33_ASAP7_75t_SL U28608 ( .A(n28742), .B(n29602), .Y(n25204) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U28609 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__28_), 
        .A2(n30007), .B(n25431), .C(n25430), .Y(n25433) );
  OAI22xp33_ASAP7_75t_SL U28610 ( .A1(n2271), .A2(n31843), .B1(n29277), .B2(
        n24640), .Y(n26518) );
  NAND2xp33_ASAP7_75t_SL U28611 ( .A(n25405), .B(n27089), .Y(n25408) );
  INVx1_ASAP7_75t_SL U28612 ( .A(n32215), .Y(n32379) );
  INVx1_ASAP7_75t_SL U28613 ( .A(u0_0_leon3x0_p0_iu_fe_pc_28_), .Y(
        add_x_746_n20) );
  OAI21xp33_ASAP7_75t_SL U28614 ( .A1(n32705), .A2(n2926), .B(n31322), .Y(
        ahb0_v_HADDR__4_) );
  NAND2xp33_ASAP7_75t_SL U28615 ( .A(n28894), .B(n30369), .Y(n26180) );
  OAI22xp33_ASAP7_75t_SL U28616 ( .A1(n4414), .A2(n31843), .B1(n26530), .B2(
        n24640), .Y(n26531) );
  INVxp33_ASAP7_75t_SL U28617 ( .A(n29975), .Y(n29976) );
  NAND2xp33_ASAP7_75t_SL U28618 ( .A(n30007), .B(n28619), .Y(n25432) );
  NAND2xp5_ASAP7_75t_SL U28619 ( .A(n29351), .B(n28043), .Y(n28049) );
  NAND2xp5_ASAP7_75t_SL U28620 ( .A(n32705), .B(n31743), .Y(n32824) );
  INVx1_ASAP7_75t_SL U28621 ( .A(u0_0_leon3x0_p0_iu_fe_pc_26_), .Y(
        add_x_746_n32) );
  INVxp67_ASAP7_75t_SL U28622 ( .A(n28896), .Y(n28897) );
  INVx1_ASAP7_75t_SL U28623 ( .A(u0_0_leon3x0_p0_iu_fe_pc_24_), .Y(
        add_x_746_n44) );
  INVx1_ASAP7_75t_SL U28624 ( .A(n32786), .Y(n32703) );
  AOI22xp33_ASAP7_75t_SL U28625 ( .A1(n28847), .A2(n26293), .B1(n24575), .B2(
        n26258), .Y(n26144) );
  NAND2xp33_ASAP7_75t_SL U28626 ( .A(n30212), .B(n30211), .Y(n30690) );
  INVxp33_ASAP7_75t_SL U28627 ( .A(n26597), .Y(n26150) );
  NOR2x1_ASAP7_75t_SL U28628 ( .A(n32036), .B(n31794), .Y(n32875) );
  INVxp67_ASAP7_75t_SL U28629 ( .A(mult_x_1196_n2090), .Y(mult_x_1196_n2088)
         );
  NAND2xp33_ASAP7_75t_SL U28630 ( .A(n28967), .B(n27090), .Y(n26256) );
  OAI21xp33_ASAP7_75t_SL U28631 ( .A1(n28148), .A2(n28179), .B(n28147), .Y(
        n28150) );
  INVxp67_ASAP7_75t_SL U28632 ( .A(add_x_735_n183), .Y(add_x_735_n185) );
  OAI21xp33_ASAP7_75t_SL U28633 ( .A1(n29675), .A2(n29674), .B(n30159), .Y(
        n30211) );
  OAI21xp33_ASAP7_75t_SL U28634 ( .A1(n18876), .A2(n30974), .B(n29052), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_11_) );
  NAND2xp33_ASAP7_75t_SL U28635 ( .A(n27513), .B(n27512), .Y(n29975) );
  OAI21xp33_ASAP7_75t_SL U28636 ( .A1(n18876), .A2(n32586), .B(n29053), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_10_) );
  O2A1O1Ixp33_ASAP7_75t_SL U28637 ( .A1(n25833), .A2(n25832), .B(n24634), .C(
        n25831), .Y(n25834) );
  AOI22xp33_ASAP7_75t_SL U28638 ( .A1(n28967), .A2(n27092), .B1(n27098), .B2(
        n27091), .Y(n27093) );
  OAI21xp33_ASAP7_75t_SL U28639 ( .A1(n18876), .A2(n32574), .B(n29055), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_7_) );
  OAI21xp33_ASAP7_75t_SL U28640 ( .A1(n18876), .A2(n25890), .B(n25889), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_30_) );
  OAI21xp33_ASAP7_75t_SL U28641 ( .A1(n18876), .A2(n31018), .B(n29056), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_6_) );
  OAI21xp33_ASAP7_75t_SL U28642 ( .A1(n23229), .A2(u0_0_leon3x0_p0_divi[50]), 
        .B(n30305), .Y(n4045) );
  OAI21xp33_ASAP7_75t_SL U28643 ( .A1(n32303), .A2(n31470), .B(n30996), .Y(
        n30997) );
  NAND2xp5_ASAP7_75t_SL U28644 ( .A(n28405), .B(n28404), .Y(n28419) );
  OAI21xp33_ASAP7_75t_SL U28645 ( .A1(n18876), .A2(n29032), .B(n29031), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_28_) );
  AOI22xp33_ASAP7_75t_SL U28646 ( .A1(n27098), .A2(n26425), .B1(n28847), .B2(
        n27101), .Y(n26148) );
  AOI21xp33_ASAP7_75t_SL U28647 ( .A1(n31473), .A2(dc_q[6]), .B(n30560), .Y(
        n30570) );
  INVxp33_ASAP7_75t_SL U28648 ( .A(n33004), .Y(n33007) );
  INVxp67_ASAP7_75t_SL U28649 ( .A(add_x_735_n184), .Y(add_x_735_n186) );
  NAND2xp5_ASAP7_75t_SL U28650 ( .A(n26554), .B(n26553), .Y(n26559) );
  INVxp67_ASAP7_75t_SL U28651 ( .A(mult_x_1196_n2370), .Y(n23413) );
  OAI21xp33_ASAP7_75t_SL U28652 ( .A1(n26557), .A2(n28869), .B(n26556), .Y(
        n26558) );
  OAI21xp5_ASAP7_75t_SL U28653 ( .A1(mult_x_1196_n2782), .A2(n18341), .B(
        n22284), .Y(n23414) );
  AOI21xp33_ASAP7_75t_SL U28654 ( .A1(n30360), .A2(n28894), .B(n27206), .Y(
        n27207) );
  OAI21xp33_ASAP7_75t_SL U28655 ( .A1(n18876), .A2(n29034), .B(n29033), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_26_) );
  OAI21xp33_ASAP7_75t_SL U28656 ( .A1(n28849), .A2(n28869), .B(n26156), .Y(
        n26157) );
  INVx1_ASAP7_75t_SL U28657 ( .A(n32780), .Y(n33032) );
  OAI22xp33_ASAP7_75t_SL U28658 ( .A1(n28850), .A2(n26152), .B1(n27107), .B2(
        n28986), .Y(n26153) );
  OAI22xp33_ASAP7_75t_SL U28659 ( .A1(n2322), .A2(n31843), .B1(n30547), .B2(
        n24640), .Y(n26595) );
  OAI21xp33_ASAP7_75t_SL U28660 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_A__RSEL1__2_), .B(n31333), .Y(n4171) );
  XNOR2xp5_ASAP7_75t_SL U28661 ( .A(mult_x_1196_n2168), .B(mult_x_1196_n2509), 
        .Y(n23138) );
  OAI21xp33_ASAP7_75t_SL U28662 ( .A1(n18876), .A2(n32677), .B(n29061), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_3_) );
  INVxp67_ASAP7_75t_SL U28663 ( .A(n32021), .Y(n32034) );
  INVx1_ASAP7_75t_SL U28664 ( .A(n31474), .Y(n25018) );
  OAI21xp33_ASAP7_75t_SL U28665 ( .A1(n18876), .A2(n32567), .B(n29057), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_5_) );
  OAI21xp33_ASAP7_75t_SL U28666 ( .A1(n18876), .A2(n29481), .B(n29058), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_4_) );
  OAI211xp5_ASAP7_75t_SRAM U28667 ( .A1(n32026), .A2(n32025), .B(n32024), .C(
        n32023), .Y(n32032) );
  OAI22xp33_ASAP7_75t_SL U28668 ( .A1(n28850), .A2(n26279), .B1(n28871), .B2(
        n27108), .Y(n26280) );
  NAND2xp5_ASAP7_75t_SL U28669 ( .A(n25612), .B(n25611), .Y(n25615) );
  NAND2xp5_ASAP7_75t_SL U28670 ( .A(n27103), .B(n27102), .Y(n27104) );
  INVxp33_ASAP7_75t_SL U28671 ( .A(n30425), .Y(n26316) );
  AOI21xp33_ASAP7_75t_SL U28672 ( .A1(u0_0_leon3x0_p0_iu_r_X__LADDR__0_), .A2(
        n30017), .B(n25054), .Y(n29916) );
  INVx1_ASAP7_75t_SL U28673 ( .A(n31734), .Y(n31794) );
  INVxp67_ASAP7_75t_SL U28674 ( .A(n26557), .Y(n26258) );
  NAND2xp33_ASAP7_75t_SL U28675 ( .A(n29504), .B(n26915), .Y(n28619) );
  OAI21xp33_ASAP7_75t_SL U28676 ( .A1(n32297), .A2(n31470), .B(n30474), .Y(
        n30475) );
  INVxp67_ASAP7_75t_SL U28677 ( .A(n30208), .Y(n31491) );
  OAI22xp33_ASAP7_75t_SL U28678 ( .A1(n26924), .A2(n26329), .B1(n26947), .B2(
        n26522), .Y(n25430) );
  OAI21xp33_ASAP7_75t_SL U28679 ( .A1(n28871), .A2(n28869), .B(n27099), .Y(
        n27105) );
  OAI21xp33_ASAP7_75t_SL U28680 ( .A1(n18876), .A2(n32577), .B(n29054), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_8_) );
  OAI21xp33_ASAP7_75t_SL U28681 ( .A1(n18876), .A2(n30524), .B(n29051), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_12_) );
  AOI21xp33_ASAP7_75t_SL U28682 ( .A1(n29598), .A2(n29796), .B(n27153), .Y(
        n25501) );
  INVxp67_ASAP7_75t_SL U28683 ( .A(add_x_735_n2), .Y(add_x_735_n78) );
  OAI21xp33_ASAP7_75t_SL U28684 ( .A1(n18876), .A2(n29066), .B(n29039), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_23_) );
  NAND2xp33_ASAP7_75t_SL U28685 ( .A(n27523), .B(n27515), .Y(n27519) );
  NAND2xp33_ASAP7_75t_SL U28686 ( .A(n28894), .B(n30266), .Y(n26434) );
  OAI22xp33_ASAP7_75t_SL U28687 ( .A1(n27108), .A2(n26299), .B1(n26557), .B2(
        n28850), .Y(n26300) );
  NAND2xp5_ASAP7_75t_SL U28688 ( .A(n26961), .B(n26960), .Y(n26962) );
  OAI21xp33_ASAP7_75t_SL U28689 ( .A1(n18876), .A2(n29036), .B(n29035), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_25_) );
  AOI22xp33_ASAP7_75t_SL U28690 ( .A1(n24576), .A2(n26376), .B1(n28847), .B2(
        n27091), .Y(n26379) );
  OAI21xp33_ASAP7_75t_SL U28691 ( .A1(n32752), .A2(n32751), .B(
        sr1_r_MCFG2__RAMBANKSZ__3_), .Y(n32758) );
  NAND2xp33_ASAP7_75t_SL U28692 ( .A(n32705), .B(n31321), .Y(n31322) );
  AOI21xp5_ASAP7_75t_SL U28693 ( .A1(n29143), .A2(n29135), .B(n28965), .Y(
        n29007) );
  AOI21xp33_ASAP7_75t_SL U28694 ( .A1(n30672), .A2(n30671), .B(n30670), .Y(
        n30673) );
  INVxp33_ASAP7_75t_SL U28695 ( .A(n26425), .Y(n25467) );
  NAND2xp5_ASAP7_75t_SL U28696 ( .A(n25472), .B(n25471), .Y(n25473) );
  INVxp67_ASAP7_75t_SL U28697 ( .A(mult_x_1196_n2219), .Y(n22612) );
  NAND2xp5_ASAP7_75t_SL U28698 ( .A(n26392), .B(n26391), .Y(n28497) );
  NAND2xp5_ASAP7_75t_SL U28699 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[1]), .B(n32021), 
        .Y(n31612) );
  AOI21xp33_ASAP7_75t_SL U28700 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__3_), 
        .A2(n24647), .B(n30702), .Y(n3346) );
  AOI22xp33_ASAP7_75t_SL U28701 ( .A1(ahb0_r_HADDR__2_), .A2(n22393), .B1(
        n32705), .B2(n32984), .Y(n2932) );
  XNOR2xp5_ASAP7_75t_SL U28702 ( .A(mult_x_1196_n2190), .B(mult_x_1196_n1080), 
        .Y(n24093) );
  OAI21xp33_ASAP7_75t_SL U28703 ( .A1(n18876), .A2(n30506), .B(n29048), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_14_) );
  AOI21xp33_ASAP7_75t_SL U28704 ( .A1(n30438), .A2(n28894), .B(n28838), .Y(
        n28839) );
  INVxp33_ASAP7_75t_SL U28705 ( .A(n33040), .Y(n33043) );
  OAI21xp33_ASAP7_75t_SL U28706 ( .A1(n18876), .A2(n30540), .B(n29046), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_17_) );
  OAI21xp33_ASAP7_75t_SL U28707 ( .A1(n18876), .A2(n30533), .B(n29047), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_16_) );
  INVxp33_ASAP7_75t_SL U28708 ( .A(n29982), .Y(n27516) );
  OAI21xp33_ASAP7_75t_SL U28709 ( .A1(n18876), .A2(n31834), .B(n29045), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_18_) );
  OAI21xp33_ASAP7_75t_SL U28710 ( .A1(n28916), .A2(n28986), .B(n28915), .Y(
        n28919) );
  OAI21xp33_ASAP7_75t_SL U28711 ( .A1(n30426), .A2(n30425), .B(n30424), .Y(
        n30427) );
  OAI21xp33_ASAP7_75t_SL U28712 ( .A1(n18876), .A2(n30828), .B(n29044), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_19_) );
  OAI21xp33_ASAP7_75t_SL U28713 ( .A1(n28975), .A2(n25460), .B(n25118), .Y(
        n25119) );
  OAI21xp33_ASAP7_75t_SL U28714 ( .A1(n28977), .A2(n25460), .B(n25459), .Y(
        n26938) );
  OAI21xp33_ASAP7_75t_SL U28715 ( .A1(n18876), .A2(n31765), .B(n29041), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_21_) );
  OAI21xp33_ASAP7_75t_SL U28716 ( .A1(n18876), .A2(n29043), .B(n29042), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_20_) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U28717 ( .A1(u0_0_leon3x0_p0_c0mmu_mcdi[1]), .A2(
        n32021), .B(n32197), .C(n31621), .Y(n31623) );
  OAI22xp33_ASAP7_75t_SL U28718 ( .A1(n27017), .A2(n31343), .B1(n23229), .B2(
        u0_0_leon3x0_p0_iu_r_E__ALUADD_), .Y(n3306) );
  NAND2xp33_ASAP7_75t_SL U28719 ( .A(n28894), .B(n30246), .Y(n25502) );
  OAI21xp33_ASAP7_75t_SL U28720 ( .A1(n28871), .A2(n28986), .B(n28870), .Y(
        n28872) );
  NAND2xp33_ASAP7_75t_SL U28721 ( .A(n24575), .B(n26425), .Y(n26426) );
  OAI22xp33_ASAP7_75t_SL U28722 ( .A1(n28366), .A2(n28365), .B1(n22421), .B2(
        u0_0_leon3x0_p0_divi[31]), .Y(n4089) );
  OAI22xp33_ASAP7_75t_SL U28723 ( .A1(n25908), .A2(n28986), .B1(n28869), .B2(
        n27107), .Y(n25792) );
  NAND2xp33_ASAP7_75t_SL U28724 ( .A(n28894), .B(n30337), .Y(n26690) );
  INVxp33_ASAP7_75t_SL U28725 ( .A(n33033), .Y(n33036) );
  AOI22xp33_ASAP7_75t_SL U28726 ( .A1(n28847), .A2(n27092), .B1(n24575), .B2(
        n27091), .Y(n25789) );
  NAND2xp5_ASAP7_75t_SL U28727 ( .A(n25799), .B(n25798), .Y(n27078) );
  NAND2xp5_ASAP7_75t_SL U28728 ( .A(n26482), .B(n26524), .Y(n26588) );
  OAI22xp33_ASAP7_75t_SL U28729 ( .A1(n25908), .A2(n28850), .B1(n27108), .B2(
        n27107), .Y(n25811) );
  OAI21xp33_ASAP7_75t_SL U28730 ( .A1(n28144), .A2(n28179), .B(n28143), .Y(
        n28146) );
  OAI22xp33_ASAP7_75t_SL U28731 ( .A1(n28986), .A2(n26152), .B1(n27106), .B2(
        n28869), .Y(n25810) );
  OAI21xp33_ASAP7_75t_SL U28732 ( .A1(n28169), .A2(n28179), .B(n28168), .Y(
        n28171) );
  NAND2xp33_ASAP7_75t_SL U28733 ( .A(n28894), .B(n30349), .Y(n26579) );
  OAI21xp33_ASAP7_75t_SL U28734 ( .A1(n28164), .A2(n28179), .B(n28163), .Y(
        n28166) );
  INVxp33_ASAP7_75t_SL U28735 ( .A(n32751), .Y(n32700) );
  OAI21xp33_ASAP7_75t_SL U28736 ( .A1(n28156), .A2(n28179), .B(n28155), .Y(
        n28158) );
  OAI21xp33_ASAP7_75t_SL U28737 ( .A1(n28160), .A2(n28179), .B(n28159), .Y(
        n28162) );
  NAND2xp5_ASAP7_75t_SL U28738 ( .A(n25391), .B(n25395), .Y(n31967) );
  INVxp33_ASAP7_75t_SL U28739 ( .A(add_x_735_n62), .Y(add_x_735_n64) );
  AOI21xp33_ASAP7_75t_SL U28740 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__4_), 
        .A2(n22378), .B(n30702), .Y(n3350) );
  OAI22xp33_ASAP7_75t_SL U28741 ( .A1(n32308), .A2(n31470), .B1(n32491), .B2(
        n24426), .Y(n31471) );
  OAI22xp33_ASAP7_75t_SL U28742 ( .A1(n28869), .A2(n25908), .B1(n27108), .B2(
        n25907), .Y(n25909) );
  NAND2xp33_ASAP7_75t_SL U28743 ( .A(n27098), .B(n25910), .Y(n25480) );
  OAI21xp5_ASAP7_75t_SL U28744 ( .A1(n23061), .A2(n26329), .B(n26328), .Y(
        n32215) );
  AOI21xp33_ASAP7_75t_SL U28745 ( .A1(n28894), .A2(n28690), .B(n28689), .Y(
        n28691) );
  INVxp33_ASAP7_75t_SL U28746 ( .A(mult_x_1196_n1080), .Y(n24094) );
  NAND2xp33_ASAP7_75t_SL U28747 ( .A(n28967), .B(n26425), .Y(n25761) );
  INVx1_ASAP7_75t_SL U28748 ( .A(mult_x_1196_n1183), .Y(n22931) );
  INVxp33_ASAP7_75t_SL U28749 ( .A(n29154), .Y(n29157) );
  AOI21xp33_ASAP7_75t_SL U28750 ( .A1(n31093), .A2(uart1_r_RHOLD__11__4_), .B(
        n30748), .Y(n2147) );
  AOI21xp33_ASAP7_75t_SL U28751 ( .A1(n31121), .A2(uart1_r_RHOLD__12__7_), .B(
        n30849), .Y(n2055) );
  AOI22xp33_ASAP7_75t_SL U28752 ( .A1(ic_q[30]), .A2(n22387), .B1(dc_q[30]), 
        .B2(n31473), .Y(n25616) );
  AOI21xp33_ASAP7_75t_SL U28753 ( .A1(n31105), .A2(uart1_r_RHOLD__3__4_), .B(
        n30751), .Y(n2139) );
  NAND2xp33_ASAP7_75t_SL U28754 ( .A(n22968), .B(n28402), .Y(n26486) );
  AOI31xp33_ASAP7_75t_SRAM U28755 ( .A1(n26013), .A2(n26039), .A3(n28191), .B(
        n25978), .Y(n2457) );
  NAND2xp33_ASAP7_75t_SL U28756 ( .A(n28847), .B(n25790), .Y(n25481) );
  AOI21xp33_ASAP7_75t_SL U28757 ( .A1(n31129), .A2(uart1_r_RHOLD__21__3_), .B(
        n28210), .Y(n2188) );
  AOI21xp33_ASAP7_75t_SL U28758 ( .A1(n31081), .A2(uart1_r_RHOLD__22__3_), .B(
        n28198), .Y(n2189) );
  AOI21xp33_ASAP7_75t_SL U28759 ( .A1(n31085), .A2(uart1_r_RHOLD__23__3_), .B(
        n28199), .Y(n2190) );
  AOI22xp33_ASAP7_75t_SL U28760 ( .A1(n30130), .A2(n32657), .B1(dt_q[26]), 
        .B2(n24573), .Y(n25618) );
  AOI21xp33_ASAP7_75t_SL U28761 ( .A1(n31105), .A2(uart1_r_RHOLD__3__2_), .B(
        n29535), .Y(n2201) );
  INVxp67_ASAP7_75t_SL U28762 ( .A(n32992), .Y(n32993) );
  NAND2xp33_ASAP7_75t_SL U28763 ( .A(n28967), .B(n25794), .Y(n25482) );
  AOI21xp33_ASAP7_75t_SL U28764 ( .A1(n31089), .A2(uart1_r_RHOLD__13__7_), .B(
        n30841), .Y(n2056) );
  AOI21xp33_ASAP7_75t_SL U28765 ( .A1(n31109), .A2(uart1_r_RHOLD__28__3_), .B(
        n28205), .Y(n2195) );
  OAI21xp33_ASAP7_75t_SL U28766 ( .A1(apbi[8]), .A2(n31840), .B(n26623), .Y(
        n1742) );
  AOI21xp33_ASAP7_75t_SL U28767 ( .A1(n31065), .A2(uart1_r_RHOLD__24__3_), .B(
        n28194), .Y(n2191) );
  OAI21xp33_ASAP7_75t_SL U28768 ( .A1(n31412), .A2(n30345), .B(n30344), .Y(
        n30348) );
  INVx1_ASAP7_75t_SL U28769 ( .A(n32729), .Y(n24644) );
  AOI21xp33_ASAP7_75t_SL U28770 ( .A1(n31097), .A2(uart1_r_RHOLD__14__7_), .B(
        n30843), .Y(n2057) );
  AOI21xp33_ASAP7_75t_SL U28771 ( .A1(n31113), .A2(uart1_r_RHOLD__1__2_), .B(
        n29537), .Y(n2199) );
  OAI21xp33_ASAP7_75t_SL U28772 ( .A1(n30250), .A2(n30625), .B(n28437), .Y(
        n28438) );
  NAND2xp5_ASAP7_75t_SL U28773 ( .A(n31604), .B(n32451), .Y(n32021) );
  AOI21xp33_ASAP7_75t_SL U28774 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__PS_), .A2(
        n24647), .B(n29222), .Y(n3369) );
  AOI22xp33_ASAP7_75t_SL U28775 ( .A1(n27098), .A2(n25470), .B1(n28975), .B2(
        n25469), .Y(n25472) );
  AOI21xp33_ASAP7_75t_SL U28776 ( .A1(n31117), .A2(uart1_r_RHOLD__15__7_), .B(
        n30848), .Y(n2058) );
  NAND2xp33_ASAP7_75t_SL U28777 ( .A(n23650), .B(n29935), .Y(n29938) );
  AOI22xp33_ASAP7_75t_SL U28778 ( .A1(n28967), .A2(n26390), .B1(n28981), .B2(
        n26555), .Y(n26391) );
  INVxp67_ASAP7_75t_SL U28779 ( .A(n24135), .Y(n24136) );
  AOI21xp33_ASAP7_75t_SL U28780 ( .A1(n31133), .A2(uart1_r_RHOLD__6__4_), .B(
        n30758), .Y(n2142) );
  AOI22xp33_ASAP7_75t_SL U28781 ( .A1(n27098), .A2(n26551), .B1(n28967), .B2(
        n26552), .Y(n26143) );
  AOI21xp33_ASAP7_75t_SL U28782 ( .A1(n31065), .A2(uart1_r_RHOLD__24__5_), .B(
        n30032), .Y(n2129) );
  AOI21xp33_ASAP7_75t_SL U28783 ( .A1(n31125), .A2(uart1_r_RHOLD__26__3_), .B(
        n28209), .Y(n2193) );
  AOI21xp33_ASAP7_75t_SL U28784 ( .A1(n31101), .A2(uart1_r_RHOLD__29__3_), .B(
        n28203), .Y(n2196) );
  AOI22xp33_ASAP7_75t_SL U28785 ( .A1(n27098), .A2(n26389), .B1(n28847), .B2(
        n26551), .Y(n26392) );
  AOI21xp33_ASAP7_75t_SL U28786 ( .A1(n31109), .A2(uart1_r_RHOLD__28__6_), .B(
        n31108), .Y(n2102) );
  AOI21xp33_ASAP7_75t_SL U28787 ( .A1(n31065), .A2(uart1_r_RHOLD__24__4_), .B(
        n30741), .Y(n2160) );
  AOI21xp33_ASAP7_75t_SL U28788 ( .A1(n31125), .A2(uart1_r_RHOLD__26__4_), .B(
        n30756), .Y(n2162) );
  OAI21xp33_ASAP7_75t_SL U28789 ( .A1(n26675), .A2(n26674), .B(n26673), .Y(
        n26679) );
  OAI21xp5_ASAP7_75t_SL U28790 ( .A1(n26454), .A2(n29910), .B(n27489), .Y(
        n26524) );
  AOI21xp33_ASAP7_75t_SL U28791 ( .A1(n31085), .A2(uart1_r_RHOLD__23__4_), .B(
        n30746), .Y(n2159) );
  AOI21xp33_ASAP7_75t_SL U28792 ( .A1(n31101), .A2(uart1_r_RHOLD__29__5_), .B(
        n30041), .Y(n2134) );
  INVx1_ASAP7_75t_SL U28793 ( .A(n30130), .Y(n31470) );
  AOI21xp33_ASAP7_75t_SL U28794 ( .A1(n31081), .A2(uart1_r_RHOLD__22__4_), .B(
        n30745), .Y(n2158) );
  INVxp67_ASAP7_75t_SL U28795 ( .A(n31048), .Y(n31049) );
  AOI21xp33_ASAP7_75t_SL U28796 ( .A1(n31109), .A2(uart1_r_RHOLD__28__4_), .B(
        n30752), .Y(n2164) );
  AOI21xp33_ASAP7_75t_SL U28797 ( .A1(n31101), .A2(uart1_r_RHOLD__29__4_), .B(
        n30750), .Y(n2165) );
  AOI21xp33_ASAP7_75t_SL U28798 ( .A1(n31129), .A2(uart1_r_RHOLD__21__4_), .B(
        n30757), .Y(n2157) );
  NOR2x1_ASAP7_75t_SL U28799 ( .A(n23581), .B(n23582), .Y(n23580) );
  AOI21xp33_ASAP7_75t_SL U28800 ( .A1(n31113), .A2(uart1_r_RHOLD__1__7_), .B(
        n30847), .Y(n2044) );
  INVxp67_ASAP7_75t_SL U28801 ( .A(n28402), .Y(n26329) );
  NAND2xp33_ASAP7_75t_SL U28802 ( .A(n27098), .B(n26424), .Y(n25760) );
  AOI22xp33_ASAP7_75t_SL U28803 ( .A1(u0_0_leon3x0_p0_c0mmu_a0_r_HLOCKEN_), 
        .A2(n32042), .B1(n25600), .B2(n32035), .Y(n3896) );
  AOI22xp33_ASAP7_75t_SL U28804 ( .A1(it_q[12]), .A2(n24636), .B1(n32629), 
        .B2(n30130), .Y(n26666) );
  AOI21xp33_ASAP7_75t_SL U28805 ( .A1(n31113), .A2(uart1_r_RHOLD__1__3_), .B(
        n28206), .Y(n2168) );
  AOI21xp33_ASAP7_75t_SL U28806 ( .A1(n31133), .A2(uart1_r_RHOLD__6__7_), .B(
        n30852), .Y(n2049) );
  INVxp33_ASAP7_75t_SL U28807 ( .A(n27241), .Y(n32114) );
  AOI21xp33_ASAP7_75t_SL U28808 ( .A1(n31109), .A2(uart1_r_RHOLD__28__5_), .B(
        n30043), .Y(n2133) );
  NAND2xp33_ASAP7_75t_SL U28809 ( .A(timer0_vtimers_1__RELOAD__12_), .B(n30993), .Y(n29854) );
  AOI21xp33_ASAP7_75t_SL U28810 ( .A1(n31105), .A2(uart1_r_RHOLD__3__3_), .B(
        n28204), .Y(n2170) );
  INVxp33_ASAP7_75t_SL U28811 ( .A(n29351), .Y(n29375) );
  AOI21xp33_ASAP7_75t_SL U28812 ( .A1(n31105), .A2(uart1_r_RHOLD__3__7_), .B(
        n30845), .Y(n2046) );
  AOI21xp33_ASAP7_75t_SL U28813 ( .A1(n31073), .A2(uart1_r_RHOLD__18__4_), .B(
        n30743), .Y(n2154) );
  AOI21xp33_ASAP7_75t_SL U28814 ( .A1(n31133), .A2(uart1_r_RHOLD__6__3_), .B(
        n28211), .Y(n2173) );
  OAI21xp33_ASAP7_75t_SL U28815 ( .A1(apbi[13]), .A2(n29383), .B(n29233), .Y(
        n1755) );
  OAI21xp33_ASAP7_75t_SL U28816 ( .A1(apbi[13]), .A2(n31840), .B(n26604), .Y(
        n1753) );
  OAI21xp33_ASAP7_75t_SL U28817 ( .A1(n1765), .A2(n24633), .B(n29333), .Y(
        n17812) );
  NAND2xp33_ASAP7_75t_SL U28818 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[50]), .B(
        n24583), .Y(n30543) );
  NAND2xp33_ASAP7_75t_SL U28819 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[46]), .B(
        n24583), .Y(n30529) );
  AOI21xp33_ASAP7_75t_SL U28820 ( .A1(n22387), .A2(ic_q[17]), .B(n27249), .Y(
        n27252) );
  INVx1_ASAP7_75t_SL U28821 ( .A(n31621), .Y(n30916) );
  AOI22xp33_ASAP7_75t_SL U28822 ( .A1(it_q[13]), .A2(n24636), .B1(n32631), 
        .B2(n30130), .Y(n27251) );
  NAND2xp33_ASAP7_75t_SL U28823 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[51]), .B(
        n24583), .Y(n31791) );
  NAND2xp33_ASAP7_75t_SL U28824 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[47]), .B(
        n24583), .Y(n30513) );
  AOI21xp33_ASAP7_75t_SL U28825 ( .A1(n31117), .A2(uart1_r_RHOLD__15__4_), .B(
        n30754), .Y(n2151) );
  NAND2xp33_ASAP7_75t_SL U28826 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[49]), .B(
        n24583), .Y(n30536) );
  AOI21xp33_ASAP7_75t_SL U28827 ( .A1(n31113), .A2(uart1_r_RHOLD__1__4_), .B(
        n30753), .Y(n2137) );
  AOI21xp33_ASAP7_75t_SL U28828 ( .A1(n31093), .A2(uart1_r_RHOLD__11__3_), .B(
        n28201), .Y(n2178) );
  AOI21xp33_ASAP7_75t_SL U28829 ( .A1(n31097), .A2(uart1_r_RHOLD__14__4_), .B(
        n30749), .Y(n2150) );
  AOI21xp33_ASAP7_75t_SL U28830 ( .A1(n31121), .A2(uart1_r_RHOLD__12__3_), .B(
        n28208), .Y(n2179) );
  AOI21xp33_ASAP7_75t_SL U28831 ( .A1(n31089), .A2(uart1_r_RHOLD__13__3_), .B(
        n28200), .Y(n2180) );
  OAI21xp33_ASAP7_75t_SL U28832 ( .A1(apbi[8]), .A2(n29383), .B(n29271), .Y(
        n1744) );
  AOI21xp33_ASAP7_75t_SL U28833 ( .A1(n31089), .A2(uart1_r_RHOLD__13__4_), .B(
        n30747), .Y(n2149) );
  NAND2xp33_ASAP7_75t_SL U28834 ( .A(n30507), .B(n32729), .Y(n30508) );
  AOI21xp33_ASAP7_75t_SL U28835 ( .A1(n31097), .A2(uart1_r_RHOLD__14__3_), .B(
        n28202), .Y(n2181) );
  AOI21xp33_ASAP7_75t_SL U28836 ( .A1(n31117), .A2(uart1_r_RHOLD__15__3_), .B(
        n28207), .Y(n2182) );
  NAND2xp33_ASAP7_75t_SL U28837 ( .A(n27098), .B(n27092), .Y(n26255) );
  AOI21xp33_ASAP7_75t_SL U28838 ( .A1(n31121), .A2(uart1_r_RHOLD__12__4_), .B(
        n30755), .Y(n2148) );
  INVxp33_ASAP7_75t_SL U28839 ( .A(n30384), .Y(n28690) );
  AOI21xp33_ASAP7_75t_SL U28840 ( .A1(n31125), .A2(uart1_r_RHOLD__26__5_), .B(
        n30047), .Y(n2131) );
  OAI21xp33_ASAP7_75t_SL U28841 ( .A1(n27315), .A2(n27314), .B(n27304), .Y(
        n2239) );
  AOI21xp33_ASAP7_75t_SL U28842 ( .A1(n26483), .A2(n26482), .B(n30006), .Y(
        n26600) );
  NAND2xp33_ASAP7_75t_SL U28843 ( .A(n29018), .B(n29017), .Y(
        u0_0_leon3x0_p0_div0_vaddsub) );
  AOI21xp33_ASAP7_75t_SL U28844 ( .A1(n31093), .A2(uart1_r_RHOLD__11__7_), .B(
        n30842), .Y(n2054) );
  AOI21xp33_ASAP7_75t_SL U28845 ( .A1(n31073), .A2(uart1_r_RHOLD__18__3_), .B(
        n28196), .Y(n2185) );
  NAND2xp5_ASAP7_75t_SL U28846 ( .A(n25514), .B(n31570), .Y(n32025) );
  NAND2xp33_ASAP7_75t_SL U28847 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[48]), .B(
        n24583), .Y(n30520) );
  OAI21xp33_ASAP7_75t_SL U28848 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_X__ICC__3_), .B(n29818), .Y(n2367) );
  AOI21xp33_ASAP7_75t_SL U28849 ( .A1(n31113), .A2(uart1_r_RHOLD__1__5_), .B(
        n30044), .Y(n2106) );
  OAI21xp33_ASAP7_75t_SL U28850 ( .A1(apbi[24]), .A2(n31840), .B(n26517), .Y(
        n2272) );
  NAND2xp5_ASAP7_75t_SL U28851 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[62]), .B(n24583), .Y(n25249) );
  AOI21xp33_ASAP7_75t_SL U28852 ( .A1(n31117), .A2(uart1_r_RHOLD__15__6_), .B(
        n31116), .Y(n2089) );
  AOI22xp33_ASAP7_75t_SL U28853 ( .A1(n31242), .A2(uart1_r_RHOLD__0__1_), .B1(
        uart1_r_RHOLD__24__1_), .B2(n31241), .Y(n27486) );
  AOI21xp33_ASAP7_75t_SL U28854 ( .A1(n31105), .A2(uart1_r_RHOLD__3__5_), .B(
        n30042), .Y(n2108) );
  AOI21xp33_ASAP7_75t_SL U28855 ( .A1(n31097), .A2(uart1_r_RHOLD__14__6_), .B(
        n31096), .Y(n2088) );
  INVxp33_ASAP7_75t_SL U28856 ( .A(n32165), .Y(n26851) );
  AOI21xp33_ASAP7_75t_SL U28857 ( .A1(n31113), .A2(uart1_r_RHOLD__1__1_), .B(
        n26109), .Y(n2390) );
  AOI21xp33_ASAP7_75t_SL U28858 ( .A1(n31089), .A2(uart1_r_RHOLD__13__6_), .B(
        n31088), .Y(n2087) );
  AOI21xp33_ASAP7_75t_SL U28859 ( .A1(n31113), .A2(uart1_r_RHOLD__1__0_), .B(
        n26024), .Y(n2391) );
  AOI21xp33_ASAP7_75t_SL U28860 ( .A1(n31121), .A2(uart1_r_RHOLD__12__6_), .B(
        n31120), .Y(n2086) );
  AOI21xp33_ASAP7_75t_SL U28861 ( .A1(n31093), .A2(uart1_r_RHOLD__11__6_), .B(
        n31092), .Y(n2085) );
  INVx1_ASAP7_75t_SL U28862 ( .A(mult_x_1196_n873), .Y(mult_x_1196_n861) );
  AOI21xp33_ASAP7_75t_SL U28863 ( .A1(n31105), .A2(uart1_r_RHOLD__3__1_), .B(
        n26107), .Y(n2394) );
  AOI22xp33_ASAP7_75t_SL U28864 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__30_), .B1(u0_0_leon3x0_p0_ici[58]), 
        .B2(n29059), .Y(n25889) );
  AOI21xp33_ASAP7_75t_SL U28865 ( .A1(n31105), .A2(uart1_r_RHOLD__3__0_), .B(
        n26020), .Y(n2395) );
  AOI21xp33_ASAP7_75t_SL U28866 ( .A1(n31133), .A2(uart1_r_RHOLD__6__5_), .B(
        n30049), .Y(n2111) );
  AOI21xp33_ASAP7_75t_SL U28867 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__22_), 
        .A2(n30655), .B(n29133), .Y(n1788) );
  OAI22xp33_ASAP7_75t_SL U28868 ( .A1(n26842), .A2(n32166), .B1(
        u0_0_leon3x0_p0_iu_v_M__CTRL__RD__5_), .B2(n32165), .Y(n24767) );
  AOI21xp33_ASAP7_75t_SL U28869 ( .A1(n31133), .A2(uart1_r_RHOLD__6__1_), .B(
        n26113), .Y(n2400) );
  AOI21xp33_ASAP7_75t_SL U28870 ( .A1(n31133), .A2(uart1_r_RHOLD__6__0_), .B(
        n26028), .Y(n2401) );
  AOI21xp33_ASAP7_75t_SL U28871 ( .A1(n31133), .A2(uart1_r_RHOLD__6__6_), .B(
        n31132), .Y(n2080) );
  INVx1_ASAP7_75t_SL U28872 ( .A(n26202), .Y(n31889) );
  AOI21xp33_ASAP7_75t_SL U28873 ( .A1(n31101), .A2(uart1_r_RHOLD__29__6_), .B(
        n31100), .Y(n2103) );
  OAI21xp33_ASAP7_75t_SL U28874 ( .A1(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .A2(
        n27246), .B(n27489), .Y(n28406) );
  AOI22xp33_ASAP7_75t_SL U28875 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__6_), .B1(u0_0_leon3x0_p0_ici[34]), 
        .B2(n29059), .Y(n29056) );
  AOI21xp33_ASAP7_75t_SL U28876 ( .A1(n31125), .A2(uart1_r_RHOLD__26__6_), .B(
        n31124), .Y(n2100) );
  NAND2xp33_ASAP7_75t_SL U28877 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[52]), .B(
        n24583), .Y(n30831) );
  AOI22xp33_ASAP7_75t_SL U28878 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__7_), .B1(u0_0_leon3x0_p0_ici[35]), 
        .B2(n29059), .Y(n29055) );
  AOI22xp33_ASAP7_75t_SL U28879 ( .A1(apbi[6]), .A2(n28060), .B1(uart1_r_FLOW_), .B2(n28059), .Y(n4710) );
  AOI22xp33_ASAP7_75t_SL U28880 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__8_), .B1(u0_0_leon3x0_p0_ici[36]), 
        .B2(n29059), .Y(n29054) );
  NAND2xp33_ASAP7_75t_SL U28881 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[56]), .B(
        n24583), .Y(n25247) );
  NAND2xp5_ASAP7_75t_SL U28882 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[58]), .B(n24583), .Y(n25248) );
  AOI21xp33_ASAP7_75t_SL U28883 ( .A1(n31065), .A2(uart1_r_RHOLD__24__6_), .B(
        n31064), .Y(n2098) );
  AOI22xp33_ASAP7_75t_SL U28884 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__4_), .B1(u0_0_leon3x0_p0_ici[32]), 
        .B2(n29059), .Y(n29058) );
  AOI22xp33_ASAP7_75t_SL U28885 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__5_), .B1(u0_0_leon3x0_p0_ici[33]), 
        .B2(n29059), .Y(n29057) );
  OAI21xp33_ASAP7_75t_SL U28886 ( .A1(n30304), .A2(n30625), .B(n25779), .Y(
        n25780) );
  AOI21xp33_ASAP7_75t_SL U28887 ( .A1(n31085), .A2(uart1_r_RHOLD__23__6_), .B(
        n31084), .Y(n2097) );
  OAI21xp33_ASAP7_75t_SL U28888 ( .A1(n18876), .A2(n32669), .B(n28908), .Y(
        u0_0_leon3x0_p0_iu_fe_pc_2_) );
  AOI22xp33_ASAP7_75t_SL U28889 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__3_), .B1(u0_0_leon3x0_p0_ici[31]), 
        .B2(n29059), .Y(n29061) );
  AOI21xp33_ASAP7_75t_SL U28890 ( .A1(n31081), .A2(uart1_r_RHOLD__22__6_), .B(
        n31080), .Y(n2096) );
  NAND2xp33_ASAP7_75t_SL U28891 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[53]), .B(
        n24583), .Y(n25254) );
  NAND2xp33_ASAP7_75t_SL U28892 ( .A(n24327), .B(n24406), .Y(n24328) );
  NOR2xp33_ASAP7_75t_SRAM U28893 ( .A(n31658), .B(n29115), .Y(n29116) );
  NAND2xp33_ASAP7_75t_SL U28894 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[59]), .B(
        n24583), .Y(n25255) );
  INVxp67_ASAP7_75t_SL U28895 ( .A(n26199), .Y(n26197) );
  OAI21xp33_ASAP7_75t_SL U28896 ( .A1(apbi[14]), .A2(n29383), .B(n25637), .Y(
        n2324) );
  AOI21xp33_ASAP7_75t_SL U28897 ( .A1(n31129), .A2(uart1_r_RHOLD__21__6_), .B(
        n31128), .Y(n2095) );
  NAND2xp33_ASAP7_75t_SL U28898 ( .A(n22556), .B(n28402), .Y(n26229) );
  AOI22xp33_ASAP7_75t_SL U28899 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__10_), .B1(u0_0_leon3x0_p0_ici[38]), 
        .B2(n29059), .Y(n29053) );
  AOI22xp33_ASAP7_75t_SL U28900 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__11_), .B1(u0_0_leon3x0_p0_ici[39]), 
        .B2(n29059), .Y(n29052) );
  AOI22xp33_ASAP7_75t_SL U28901 ( .A1(u0_0_leon3x0_p0_c0mmu_mcii[19]), .A2(
        n31877), .B1(u0_0_leon3x0_p0_c0mmu_mcdi[55]), .B2(n24583), .Y(n33033)
         );
  INVxp33_ASAP7_75t_SL U28902 ( .A(n30250), .Y(n29134) );
  NOR2x1_ASAP7_75t_SL U28903 ( .A(n23259), .B(n23258), .Y(n23257) );
  INVxp33_ASAP7_75t_SL U28904 ( .A(n28825), .Y(n28840) );
  AOI22xp33_ASAP7_75t_SL U28905 ( .A1(u0_0_leon3x0_p0_c0mmu_mcii[21]), .A2(
        n31877), .B1(u0_0_leon3x0_p0_c0mmu_mcdi[57]), .B2(n24583), .Y(n33040)
         );
  AOI22xp33_ASAP7_75t_SL U28906 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__28_), .B1(u0_0_leon3x0_p0_ici[56]), 
        .B2(n29059), .Y(n29031) );
  OAI21xp33_ASAP7_75t_SL U28907 ( .A1(apbi[9]), .A2(n29383), .B(n29248), .Y(
        n1796) );
  AOI21xp33_ASAP7_75t_SL U28908 ( .A1(n31073), .A2(uart1_r_RHOLD__18__6_), .B(
        n31072), .Y(n2092) );
  AOI22xp33_ASAP7_75t_SL U28909 ( .A1(it_q[15]), .A2(n24636), .B1(n32635), 
        .B2(n30130), .Y(n25742) );
  AOI22xp33_ASAP7_75t_SL U28910 ( .A1(apbi[8]), .A2(n28060), .B1(
        uart1_r_EXTCLKEN_), .B2(n28059), .Y(n4684) );
  AOI21xp33_ASAP7_75t_SL U28911 ( .A1(n31065), .A2(uart1_r_RHOLD__24__1_), .B(
        n26096), .Y(n2432) );
  AOI21xp33_ASAP7_75t_SL U28912 ( .A1(n31109), .A2(uart1_r_RHOLD__28__2_), .B(
        n29536), .Y(n2226) );
  AOI21xp33_ASAP7_75t_SL U28913 ( .A1(n31065), .A2(uart1_r_RHOLD__24__0_), .B(
        n26000), .Y(n2433) );
  NAND2xp33_ASAP7_75t_SL U28914 ( .A(n24576), .B(n27092), .Y(n26156) );
  AOI21xp33_ASAP7_75t_SL U28915 ( .A1(n31073), .A2(uart1_r_RHOLD__18__5_), .B(
        n30034), .Y(n2123) );
  AOI22xp33_ASAP7_75t_SL U28916 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__26_), .B1(u0_0_leon3x0_p0_ici[54]), 
        .B2(n29059), .Y(n29033) );
  AOI21xp33_ASAP7_75t_SL U28917 ( .A1(n31125), .A2(uart1_r_RHOLD__26__2_), .B(
        n29540), .Y(n2224) );
  AOI21xp33_ASAP7_75t_SL U28918 ( .A1(n31125), .A2(uart1_r_RHOLD__26__7_), .B(
        n30850), .Y(n2069) );
  AOI21xp33_ASAP7_75t_SL U28919 ( .A1(n31125), .A2(uart1_r_RHOLD__26__1_), .B(
        n26111), .Y(n2436) );
  INVxp33_ASAP7_75t_SL U28920 ( .A(n28964), .Y(n29143) );
  AOI21xp33_ASAP7_75t_SL U28921 ( .A1(n31065), .A2(uart1_r_RHOLD__24__2_), .B(
        n29525), .Y(n2222) );
  AOI21xp33_ASAP7_75t_SL U28922 ( .A1(n31125), .A2(uart1_r_RHOLD__26__0_), .B(
        n26026), .Y(n2437) );
  INVx1_ASAP7_75t_SL U28923 ( .A(n25790), .Y(n26152) );
  AOI21xp33_ASAP7_75t_SL U28924 ( .A1(n31085), .A2(uart1_r_RHOLD__23__2_), .B(
        n29530), .Y(n2221) );
  AOI21xp33_ASAP7_75t_SL U28925 ( .A1(n31081), .A2(uart1_r_RHOLD__22__2_), .B(
        n29529), .Y(n2220) );
  OAI22xp33_ASAP7_75t_SL U28926 ( .A1(n28869), .A2(n27109), .B1(n27108), .B2(
        n27106), .Y(n26154) );
  AOI21xp33_ASAP7_75t_SL U28927 ( .A1(n31129), .A2(uart1_r_RHOLD__21__2_), .B(
        n29541), .Y(n2219) );
  AOI21xp33_ASAP7_75t_SL U28928 ( .A1(n31109), .A2(uart1_r_RHOLD__28__1_), .B(
        n26108), .Y(n2440) );
  AOI21xp33_ASAP7_75t_SL U28929 ( .A1(n31065), .A2(uart1_r_RHOLD__24__7_), .B(
        n30835), .Y(n2067) );
  AOI21xp33_ASAP7_75t_SL U28930 ( .A1(n31109), .A2(uart1_r_RHOLD__28__0_), .B(
        n26022), .Y(n2441) );
  AOI21xp33_ASAP7_75t_SL U28931 ( .A1(n31073), .A2(uart1_r_RHOLD__18__2_), .B(
        n29527), .Y(n2216) );
  NAND2xp33_ASAP7_75t_SL U28932 ( .A(n30394), .B(n30226), .Y(n30229) );
  INVxp67_ASAP7_75t_SL U28933 ( .A(n30225), .Y(n30233) );
  AOI21xp33_ASAP7_75t_SL U28934 ( .A1(n31085), .A2(uart1_r_RHOLD__23__7_), .B(
        n30840), .Y(n2066) );
  AOI21xp33_ASAP7_75t_SL U28935 ( .A1(n31117), .A2(uart1_r_RHOLD__15__2_), .B(
        n29538), .Y(n2213) );
  AOI21xp33_ASAP7_75t_SL U28936 ( .A1(n31097), .A2(uart1_r_RHOLD__14__2_), .B(
        n29533), .Y(n2212) );
  AOI21xp33_ASAP7_75t_SL U28937 ( .A1(n31129), .A2(uart1_r_RHOLD__21__5_), .B(
        n30048), .Y(n2126) );
  AOI21xp33_ASAP7_75t_SL U28938 ( .A1(n31089), .A2(uart1_r_RHOLD__13__2_), .B(
        n29531), .Y(n2211) );
  AOI21xp33_ASAP7_75t_SL U28939 ( .A1(n31081), .A2(uart1_r_RHOLD__22__7_), .B(
        n30839), .Y(n2065) );
  NAND2xp33_ASAP7_75t_SL U28940 ( .A(n27098), .B(n26555), .Y(n26556) );
  AOI21xp33_ASAP7_75t_SL U28941 ( .A1(n31121), .A2(uart1_r_RHOLD__12__2_), .B(
        n29539), .Y(n2210) );
  AOI21xp33_ASAP7_75t_SL U28942 ( .A1(n31093), .A2(uart1_r_RHOLD__11__2_), .B(
        n29532), .Y(n2209) );
  AOI21xp33_ASAP7_75t_SL U28943 ( .A1(n31129), .A2(uart1_r_RHOLD__21__7_), .B(
        n30851), .Y(n2064) );
  NAND2xp33_ASAP7_75t_SL U28944 ( .A(n24576), .B(n26552), .Y(n26553) );
  NAND2xp33_ASAP7_75t_SL U28945 ( .A(n28967), .B(n26551), .Y(n26554) );
  AOI21xp33_ASAP7_75t_SL U28946 ( .A1(n31081), .A2(uart1_r_RHOLD__22__5_), .B(
        n30036), .Y(n2127) );
  AOI22xp33_ASAP7_75t_SL U28947 ( .A1(n28967), .A2(n27097), .B1(n24576), .B2(
        n27100), .Y(n26149) );
  AOI21xp33_ASAP7_75t_SL U28948 ( .A1(n31133), .A2(uart1_r_RHOLD__6__2_), .B(
        n29542), .Y(n2204) );
  AOI21xp33_ASAP7_75t_SL U28949 ( .A1(n31085), .A2(uart1_r_RHOLD__23__5_), .B(
        n30037), .Y(n2128) );
  AOI21xp33_ASAP7_75t_SL U28950 ( .A1(n31073), .A2(uart1_r_RHOLD__18__7_), .B(
        n30837), .Y(n2061) );
  NAND2xp5_ASAP7_75t_SL U28951 ( .A(n30110), .B(n30109), .Y(n30111) );
  INVxp67_ASAP7_75t_SL U28952 ( .A(n32184), .Y(n24782) );
  INVxp67_ASAP7_75t_SL U28953 ( .A(n27100), .Y(n26279) );
  AOI21xp33_ASAP7_75t_SL U28954 ( .A1(n31093), .A2(uart1_r_RHOLD__11__1_), .B(
        n26105), .Y(n2408) );
  NAND2xp33_ASAP7_75t_SL U28955 ( .A(n32627), .B(n30130), .Y(n25042) );
  OAI22xp33_ASAP7_75t_SL U28956 ( .A1(n27108), .A2(n28916), .B1(n28850), .B2(
        n27106), .Y(n26252) );
  AOI21xp33_ASAP7_75t_SL U28957 ( .A1(n31093), .A2(uart1_r_RHOLD__11__5_), .B(
        n30039), .Y(n2116) );
  AOI21xp33_ASAP7_75t_SL U28958 ( .A1(n31093), .A2(uart1_r_RHOLD__11__0_), .B(
        n26018), .Y(n2409) );
  AOI22xp33_ASAP7_75t_SL U28959 ( .A1(n30995), .A2(n25040), .B1(ic_q[15]), 
        .B2(n22387), .Y(n25043) );
  AOI21xp33_ASAP7_75t_SL U28960 ( .A1(n31121), .A2(uart1_r_RHOLD__12__1_), .B(
        n26110), .Y(n2410) );
  AND2x2_ASAP7_75t_SL U28961 ( .A(u0_0_leon3x0_p0_iu_r_X__LADDR__1_), .B(
        n30017), .Y(n25038) );
  AOI21xp33_ASAP7_75t_SL U28962 ( .A1(n31105), .A2(uart1_r_RHOLD__3__6_), .B(
        n31104), .Y(n2077) );
  AOI21xp33_ASAP7_75t_SL U28963 ( .A1(n31121), .A2(uart1_r_RHOLD__12__5_), .B(
        n30046), .Y(n2117) );
  AOI21xp33_ASAP7_75t_SL U28964 ( .A1(n31121), .A2(uart1_r_RHOLD__12__0_), .B(
        n26025), .Y(n2411) );
  AOI21xp33_ASAP7_75t_SL U28965 ( .A1(n31089), .A2(uart1_r_RHOLD__13__1_), .B(
        n26104), .Y(n2412) );
  INVxp67_ASAP7_75t_SL U28966 ( .A(mult_x_1196_n2396), .Y(n22824) );
  AOI21xp33_ASAP7_75t_SL U28967 ( .A1(n31089), .A2(uart1_r_RHOLD__13__0_), .B(
        n26017), .Y(n2413) );
  AOI22xp33_ASAP7_75t_SL U28968 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__31_), .A2(n30207), .B1(
        ic_q[31]), .B2(n22387), .Y(n25035) );
  AOI21xp33_ASAP7_75t_SL U28969 ( .A1(n31097), .A2(uart1_r_RHOLD__14__1_), .B(
        n26106), .Y(n2414) );
  AOI21xp33_ASAP7_75t_SL U28970 ( .A1(n31097), .A2(uart1_r_RHOLD__14__0_), .B(
        n26019), .Y(n2415) );
  AOI21xp33_ASAP7_75t_SL U28971 ( .A1(n31089), .A2(uart1_r_RHOLD__13__5_), .B(
        n30038), .Y(n2118) );
  AOI22xp33_ASAP7_75t_SL U28972 ( .A1(ic_q[23]), .A2(n22387), .B1(n32643), 
        .B2(n30130), .Y(n25061) );
  AOI21xp33_ASAP7_75t_SL U28973 ( .A1(n31113), .A2(uart1_r_RHOLD__1__6_), .B(
        n31112), .Y(n2075) );
  AOI22xp33_ASAP7_75t_SL U28974 ( .A1(it_q[7]), .A2(n24636), .B1(n32611), .B2(
        n30130), .Y(n25056) );
  INVx1_ASAP7_75t_SL U28975 ( .A(mult_x_1196_n2631), .Y(n23256) );
  AOI21xp33_ASAP7_75t_SL U28976 ( .A1(n22387), .A2(ic_q[7]), .B(n30559), .Y(
        n25057) );
  AOI21xp33_ASAP7_75t_SL U28977 ( .A1(n31073), .A2(uart1_r_RHOLD__18__1_), .B(
        n26100), .Y(n2420) );
  AOI21xp33_ASAP7_75t_SL U28978 ( .A1(n31097), .A2(uart1_r_RHOLD__14__5_), .B(
        n30040), .Y(n2119) );
  AOI21xp33_ASAP7_75t_SL U28979 ( .A1(n31073), .A2(uart1_r_RHOLD__18__0_), .B(
        n26007), .Y(n2421) );
  AOI21xp33_ASAP7_75t_SL U28980 ( .A1(n22387), .A2(ic_q[21]), .B(n27249), .Y(
        n26333) );
  AOI22xp33_ASAP7_75t_SL U28981 ( .A1(it_q[25]), .A2(n24636), .B1(n32655), 
        .B2(n30130), .Y(n25414) );
  AOI22xp33_ASAP7_75t_SL U28982 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__29_), .A2(n30207), .B1(
        ic_q[29]), .B2(n22387), .Y(n25415) );
  AOI21xp33_ASAP7_75t_SL U28983 ( .A1(n31117), .A2(uart1_r_RHOLD__15__5_), .B(
        n30045), .Y(n2120) );
  AOI21xp33_ASAP7_75t_SL U28984 ( .A1(n31129), .A2(uart1_r_RHOLD__21__1_), .B(
        n26112), .Y(n2426) );
  AOI21xp33_ASAP7_75t_SL U28985 ( .A1(n31129), .A2(uart1_r_RHOLD__21__0_), .B(
        n26027), .Y(n2427) );
  AOI21xp33_ASAP7_75t_SL U28986 ( .A1(n31101), .A2(uart1_r_RHOLD__29__7_), .B(
        n30844), .Y(n2072) );
  AOI22xp33_ASAP7_75t_SL U28987 ( .A1(it_q[9]), .A2(n24636), .B1(n32623), .B2(
        n30130), .Y(n29989) );
  AOI21xp33_ASAP7_75t_SL U28988 ( .A1(n31081), .A2(uart1_r_RHOLD__22__1_), .B(
        n26102), .Y(n2428) );
  AOI21xp33_ASAP7_75t_SL U28989 ( .A1(n31081), .A2(uart1_r_RHOLD__22__0_), .B(
        n26010), .Y(n2429) );
  AOI21xp33_ASAP7_75t_SL U28990 ( .A1(n31109), .A2(uart1_r_RHOLD__28__7_), .B(
        n30846), .Y(n2071) );
  AOI21xp33_ASAP7_75t_SL U28991 ( .A1(n31085), .A2(uart1_r_RHOLD__23__1_), .B(
        n26103), .Y(n2430) );
  AOI21xp33_ASAP7_75t_SL U28992 ( .A1(n31101), .A2(uart1_r_RHOLD__29__2_), .B(
        n29534), .Y(n2227) );
  AOI21xp33_ASAP7_75t_SL U28993 ( .A1(n31085), .A2(uart1_r_RHOLD__23__0_), .B(
        n26011), .Y(n2431) );
  NOR2x1_ASAP7_75t_SL U28994 ( .A(n24680), .B(n27241), .Y(n31054) );
  OAI21xp33_ASAP7_75t_SL U28995 ( .A1(n32986), .A2(n32719), .B(n32988), .Y(
        n31321) );
  AOI22xp33_ASAP7_75t_SL U28996 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__28_), .A2(n30207), .B1(
        ic_q[28]), .B2(n22387), .Y(n25443) );
  AOI22xp33_ASAP7_75t_SL U28997 ( .A1(n27065), .A2(n27064), .B1(n28521), .B2(
        n29598), .Y(n27074) );
  OAI21xp33_ASAP7_75t_SL U28998 ( .A1(apbi[6]), .A2(n29383), .B(n29303), .Y(
        n1731) );
  AOI22xp33_ASAP7_75t_SL U28999 ( .A1(n28967), .A2(n26389), .B1(n28847), .B2(
        n26555), .Y(n25459) );
  NAND2xp33_ASAP7_75t_SL U29000 ( .A(n23665), .B(n28402), .Y(n26446) );
  OAI21xp33_ASAP7_75t_SL U29001 ( .A1(n4520), .A2(n24633), .B(n25944), .Y(
        n17804) );
  NOR2x1_ASAP7_75t_SL U29002 ( .A(n23663), .B(n23662), .Y(n23661) );
  AOI22xp33_ASAP7_75t_SL U29003 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__19_), .B1(u0_0_leon3x0_p0_ici[47]), 
        .B2(n29059), .Y(n29044) );
  AOI22xp33_ASAP7_75t_SL U29004 ( .A1(ic_q[27]), .A2(n22387), .B1(n32651), 
        .B2(n30130), .Y(n26344) );
  OAI21xp33_ASAP7_75t_SL U29005 ( .A1(apbi[20]), .A2(n31840), .B(n31525), .Y(
        n2833) );
  INVxp67_ASAP7_75t_SL U29006 ( .A(mult_x_1196_n2335), .Y(n23065) );
  AOI22xp33_ASAP7_75t_SL U29007 ( .A1(n30995), .A2(n31451), .B1(ic_q[2]), .B2(
        n22387), .Y(n30996) );
  OAI21xp33_ASAP7_75t_SL U29008 ( .A1(apbi[21]), .A2(n31840), .B(n31839), .Y(
        n2832) );
  AOI22xp33_ASAP7_75t_SL U29009 ( .A1(it_q[14]), .A2(n24636), .B1(n32633), 
        .B2(n30130), .Y(n25715) );
  AOI22xp33_ASAP7_75t_SL U29010 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__18_), .B1(u0_0_leon3x0_p0_ici[46]), 
        .B2(n29059), .Y(n29045) );
  INVxp67_ASAP7_75t_SL U29011 ( .A(n24168), .Y(n24207) );
  AOI22xp33_ASAP7_75t_SL U29012 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__25_), .B1(u0_0_leon3x0_p0_ici[53]), 
        .B2(n29059), .Y(n29035) );
  AOI22xp33_ASAP7_75t_SL U29013 ( .A1(it_q[16]), .A2(n24636), .B1(n32637), 
        .B2(n30130), .Y(n26964) );
  AOI22xp33_ASAP7_75t_SL U29014 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__24_), .A2(n30207), .B1(
        ic_q[24]), .B2(n22387), .Y(n26512) );
  NAND2xp33_ASAP7_75t_SL U29015 ( .A(n24576), .B(n27101), .Y(n27102) );
  NAND2xp5_ASAP7_75t_SL U29016 ( .A(n27507), .B(n27512), .Y(n29981) );
  AOI22xp33_ASAP7_75t_SL U29017 ( .A1(it_q[20]), .A2(n24636), .B1(n32645), 
        .B2(n30130), .Y(n26511) );
  AOI22xp33_ASAP7_75t_SL U29018 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__25_), .A2(n30207), .B1(
        ic_q[25]), .B2(n22387), .Y(n28409) );
  OAI21xp33_ASAP7_75t_SL U29019 ( .A1(n30426), .A2(n30304), .B(n30303), .Y(
        n30305) );
  AOI22xp33_ASAP7_75t_SL U29020 ( .A1(it_q[21]), .A2(n24636), .B1(n32647), 
        .B2(n30130), .Y(n28408) );
  NAND2xp33_ASAP7_75t_SL U29021 ( .A(n28967), .B(n27100), .Y(n27103) );
  NAND2xp33_ASAP7_75t_SL U29022 ( .A(n27098), .B(n27097), .Y(n27099) );
  AOI22xp33_ASAP7_75t_SL U29023 ( .A1(ic_q[12]), .A2(n22387), .B1(n32621), 
        .B2(n30130), .Y(n25435) );
  INVxp67_ASAP7_75t_SL U29024 ( .A(add_x_735_n47), .Y(add_x_735_n274) );
  AOI22xp33_ASAP7_75t_SL U29025 ( .A1(n28980), .A2(n22939), .B1(n24571), .B2(
        n28979), .Y(n28915) );
  OAI21xp33_ASAP7_75t_SL U29026 ( .A1(n32719), .A2(n25328), .B(n25327), .Y(
        n32984) );
  AOI22xp33_ASAP7_75t_SL U29027 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__23_), .B1(u0_0_leon3x0_p0_ici[51]), 
        .B2(n29059), .Y(n29039) );
  AOI22xp33_ASAP7_75t_SL U29028 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__20_), .B1(u0_0_leon3x0_p0_ici[48]), 
        .B2(n29059), .Y(n29042) );
  XOR2xp5_ASAP7_75t_SL U29029 ( .A(n22878), .B(mult_x_1196_n2158), .Y(n22877)
         );
  NAND2xp5_ASAP7_75t_SL U29030 ( .A(n29136), .B(n29154), .Y(n30672) );
  AOI22xp33_ASAP7_75t_SL U29031 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__21_), .B1(u0_0_leon3x0_p0_ici[49]), 
        .B2(n29059), .Y(n29041) );
  AOI22xp33_ASAP7_75t_SL U29032 ( .A1(ahb0_r_HADDR__3_), .A2(n22393), .B1(
        n32705), .B2(n32985), .Y(n2928) );
  AOI22xp33_ASAP7_75t_SL U29033 ( .A1(it_q[18]), .A2(n24636), .B1(n32641), 
        .B2(n30130), .Y(n26221) );
  AOI22xp33_ASAP7_75t_SL U29034 ( .A1(it_q[24]), .A2(n24636), .B1(n32653), 
        .B2(n30130), .Y(n25442) );
  OAI21xp33_ASAP7_75t_SL U29035 ( .A1(apbi[5]), .A2(n29383), .B(n29288), .Y(
        n2852) );
  OAI21xp33_ASAP7_75t_SL U29036 ( .A1(n29587), .A2(n24427), .B(n29586), .Y(
        n29601) );
  INVxp33_ASAP7_75t_SL U29037 ( .A(mult_x_1196_n2440), .Y(n24119) );
  AOI22xp33_ASAP7_75t_SL U29038 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__14_), .B1(u0_0_leon3x0_p0_ici[42]), 
        .B2(n29059), .Y(n29048) );
  INVxp67_ASAP7_75t_SL U29039 ( .A(n29638), .Y(n30159) );
  OAI21xp33_ASAP7_75t_SL U29040 ( .A1(uart1_r_LOOPB_), .A2(n24633), .B(n29943), 
        .Y(n2869) );
  NAND2xp33_ASAP7_75t_SL U29041 ( .A(n28967), .B(n26376), .Y(n25788) );
  INVxp67_ASAP7_75t_SL U29042 ( .A(n32998), .Y(n32999) );
  INVxp67_ASAP7_75t_SL U29043 ( .A(n32996), .Y(n32997) );
  AOI21xp33_ASAP7_75t_SL U29044 ( .A1(n26298), .A2(n25782), .B(n25191), .Y(
        n25464) );
  NAND2xp5_ASAP7_75t_SL U29045 ( .A(n29137), .B(n29155), .Y(n30295) );
  OAI21xp33_ASAP7_75t_SL U29046 ( .A1(n27503), .A2(n31503), .B(n27511), .Y(
        n27515) );
  AOI22xp33_ASAP7_75t_SL U29047 ( .A1(apbi[0]), .A2(n28060), .B1(
        uart1_uarto_RXEN_), .B2(n28059), .Y(n4545) );
  INVxp67_ASAP7_75t_SL U29048 ( .A(n28142), .Y(n28141) );
  AOI22xp33_ASAP7_75t_SL U29049 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__17_), .B1(u0_0_leon3x0_p0_ici[45]), 
        .B2(n29059), .Y(n29046) );
  XOR2xp5_ASAP7_75t_SL U29050 ( .A(mult_x_1196_n2194), .B(mult_x_1196_n2255), 
        .Y(n24128) );
  AOI22xp33_ASAP7_75t_SL U29051 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__12_), .B1(u0_0_leon3x0_p0_ici[40]), 
        .B2(n29059), .Y(n29051) );
  NAND2xp33_ASAP7_75t_SL U29052 ( .A(n23965), .B(n28402), .Y(n27247) );
  AOI22xp33_ASAP7_75t_SL U29053 ( .A1(n27098), .A2(n26390), .B1(n24576), .B2(
        n26551), .Y(n25799) );
  INVxp67_ASAP7_75t_SL U29054 ( .A(add_x_735_n75), .Y(add_x_735_n73) );
  OAI211xp5_ASAP7_75t_SRAM U29055 ( .A1(n29639), .A2(n29638), .B(
        u0_0_leon3x0_p0_iu_r_M__CTRL__TT__2_), .C(n30707), .Y(n29641) );
  INVxp67_ASAP7_75t_SL U29056 ( .A(add_x_735_n115), .Y(add_x_735_n117) );
  OAI21xp33_ASAP7_75t_SL U29057 ( .A1(n32004), .A2(n30151), .B(n30150), .Y(
        n30152) );
  NAND2xp33_ASAP7_75t_SL U29058 ( .A(n24634), .B(n28825), .Y(n26998) );
  XOR2xp5_ASAP7_75t_SL U29059 ( .A(n24117), .B(mult_x_1196_n2440), .Y(n24118)
         );
  INVxp67_ASAP7_75t_SL U29060 ( .A(add_x_735_n116), .Y(add_x_735_n118) );
  OAI21xp33_ASAP7_75t_SL U29061 ( .A1(n31412), .A2(n31411), .B(n31410), .Y(
        n31414) );
  AOI22xp33_ASAP7_75t_SL U29062 ( .A1(n29585), .A2(n27064), .B1(n29579), .B2(
        n29598), .Y(n25904) );
  AOI22xp33_ASAP7_75t_SL U29063 ( .A1(n28967), .A2(n26555), .B1(n28847), .B2(
        n26552), .Y(n25798) );
  NAND2xp33_ASAP7_75t_SL U29064 ( .A(n24571), .B(n28402), .Y(n25713) );
  AOI22xp33_ASAP7_75t_SL U29065 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__16_), .B1(u0_0_leon3x0_p0_ici[44]), 
        .B2(n29059), .Y(n29047) );
  AOI22xp33_ASAP7_75t_SL U29066 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__26_), .A2(n30207), .B1(
        ic_q[26]), .B2(n22387), .Y(n26234) );
  INVxp67_ASAP7_75t_SL U29067 ( .A(n33002), .Y(n33003) );
  NAND2xp33_ASAP7_75t_SL U29068 ( .A(n27098), .B(n26377), .Y(n26378) );
  AOI22xp33_ASAP7_75t_SL U29069 ( .A1(n27098), .A2(n26423), .B1(n28847), .B2(
        n27097), .Y(n26428) );
  OAI21xp33_ASAP7_75t_SL U29070 ( .A1(n26298), .A2(n26297), .B(n26296), .Y(
        n28974) );
  NAND2xp33_ASAP7_75t_SL U29071 ( .A(n28967), .B(n26424), .Y(n26427) );
  OAI21xp33_ASAP7_75t_SL U29072 ( .A1(apbi[25]), .A2(n31840), .B(n31367), .Y(
        n2829) );
  INVxp67_ASAP7_75t_SL U29073 ( .A(n33000), .Y(n33001) );
  AOI22xp33_ASAP7_75t_SL U29074 ( .A1(apbi[1]), .A2(n28060), .B1(
        uart1_uarto_TXEN_), .B2(n28059), .Y(n2894) );
  NAND2xp33_ASAP7_75t_SL U29075 ( .A(n23161), .B(n28402), .Y(n26960) );
  AOI22xp5_ASAP7_75t_SL U29076 ( .A1(n26926), .A2(n26925), .B1(n26924), .B2(
        n26923), .Y(n30237) );
  AOI22xp33_ASAP7_75t_SL U29077 ( .A1(it_q[22]), .A2(n24636), .B1(n32649), 
        .B2(n30130), .Y(n26233) );
  INVxp33_ASAP7_75t_SL U29078 ( .A(n25133), .Y(n25135) );
  OAI22xp33_ASAP7_75t_SL U29079 ( .A1(n31155), .A2(n31184), .B1(n31154), .B2(
        n31182), .Y(n31156) );
  OAI21xp33_ASAP7_75t_SL U29080 ( .A1(uart1_r_THOLD__25__2_), .A2(n27920), .B(
        n27852), .Y(n1860) );
  OAI22xp33_ASAP7_75t_SL U29081 ( .A1(n31107), .A2(n30063), .B1(n31106), .B2(
        n30062), .Y(n30043) );
  OAI21xp33_ASAP7_75t_SL U29082 ( .A1(uart1_r_THOLD__24__3_), .A2(n27947), .B(
        n27795), .Y(n1993) );
  OAI21xp33_ASAP7_75t_SL U29083 ( .A1(n30446), .A2(n30312), .B(n30311), .Y(
        n30315) );
  OAI22xp33_ASAP7_75t_SL U29084 ( .A1(n31163), .A2(n30866), .B1(n31162), .B2(
        n30865), .Y(n30860) );
  OAI21xp33_ASAP7_75t_SL U29085 ( .A1(uart1_r_THOLD__9__1_), .A2(n27929), .B(
        n27352), .Y(n2023) );
  OAI21xp33_ASAP7_75t_SL U29086 ( .A1(uart1_r_THOLD__25__0_), .A2(n27920), .B(
        n27919), .Y(n1862) );
  OAI22xp33_ASAP7_75t_SL U29087 ( .A1(n31171), .A2(n30772), .B1(n31170), .B2(
        n30771), .Y(n30768) );
  OAI21xp33_ASAP7_75t_SL U29088 ( .A1(uart1_r_THOLD__11__7_), .A2(n27977), .B(
        n27579), .Y(n1905) );
  OAI21xp33_ASAP7_75t_SL U29089 ( .A1(uart1_r_THOLD__30__3_), .A2(n27950), .B(
        n27807), .Y(n1994) );
  OAI21xp33_ASAP7_75t_SL U29090 ( .A1(uart1_r_THOLD__13__5_), .A2(n27931), .B(
        n27669), .Y(n1947) );
  OAI21xp33_ASAP7_75t_SL U29091 ( .A1(uart1_r_THOLD__20__4_), .A2(n27939), .B(
        n27727), .Y(n1842) );
  OAI22xp33_ASAP7_75t_SL U29092 ( .A1(n31167), .A2(n30063), .B1(n31166), .B2(
        n30062), .Y(n30058) );
  OAI22xp33_ASAP7_75t_SL U29093 ( .A1(n31127), .A2(n31184), .B1(n31126), .B2(
        n31182), .Y(n31128) );
  OAI22xp33_ASAP7_75t_SL U29094 ( .A1(n31179), .A2(n30063), .B1(n31178), .B2(
        n30062), .Y(n30061) );
  OAI21xp33_ASAP7_75t_SL U29095 ( .A1(uart1_r_THOLD__28__3_), .A2(n27935), .B(
        n27787), .Y(n1883) );
  OAI22xp33_ASAP7_75t_SL U29096 ( .A1(n31127), .A2(n30866), .B1(n31126), .B2(
        n30865), .Y(n30851) );
  OAI21xp33_ASAP7_75t_SL U29097 ( .A1(uart1_r_THOLD__31__1_), .A2(n27975), .B(
        n27384), .Y(n2042) );
  OAI21xp33_ASAP7_75t_SL U29098 ( .A1(uart1_r_THOLD__30__0_), .A2(n27950), .B(
        n27949), .Y(n2035) );
  OAI22xp33_ASAP7_75t_SL U29099 ( .A1(n31151), .A2(n30063), .B1(n31150), .B2(
        n30062), .Y(n30054) );
  OAI22xp33_ASAP7_75t_SL U29100 ( .A1(n31115), .A2(n31184), .B1(n31114), .B2(
        n31182), .Y(n31116) );
  OAI21xp33_ASAP7_75t_SL U29101 ( .A1(uart1_r_THOLD__22__4_), .A2(n27952), .B(
        n27737), .Y(n1972) );
  OAI22xp33_ASAP7_75t_SL U29102 ( .A1(n31087), .A2(n30063), .B1(n31086), .B2(
        n30062), .Y(n30038) );
  OAI22xp33_ASAP7_75t_SL U29103 ( .A1(n31147), .A2(n30063), .B1(n31146), .B2(
        n30062), .Y(n30053) );
  OAI21xp33_ASAP7_75t_SL U29104 ( .A1(uart1_r_THOLD__10__1_), .A2(n27948), .B(
        n27356), .Y(n2024) );
  OAI21xp33_ASAP7_75t_SL U29105 ( .A1(uart1_r_THOLD__20__6_), .A2(n27939), .B(
        n27595), .Y(n1840) );
  OAI21xp33_ASAP7_75t_SL U29106 ( .A1(uart1_r_THOLD__16__6_), .A2(n27946), .B(
        n27600), .Y(n1929) );
  OAI21xp33_ASAP7_75t_SL U29107 ( .A1(uart1_r_THOLD__22__3_), .A2(n27952), .B(
        n27809), .Y(n1992) );
  OAI21xp33_ASAP7_75t_SL U29108 ( .A1(uart1_r_THOLD__28__1_), .A2(n27935), .B(
        n27323), .Y(n1885) );
  OAI22xp33_ASAP7_75t_SL U29109 ( .A1(n31095), .A2(n30063), .B1(n31094), .B2(
        n30062), .Y(n30040) );
  OAI21xp33_ASAP7_75t_SL U29110 ( .A1(uart1_r_THOLD__12__5_), .A2(n27937), .B(
        n27652), .Y(n1946) );
  OAI22xp33_ASAP7_75t_SL U29111 ( .A1(n31079), .A2(n30866), .B1(n31078), .B2(
        n30865), .Y(n30839) );
  OAI21xp33_ASAP7_75t_SL U29112 ( .A1(n30645), .A2(n27030), .B(n27011), .Y(
        n27012) );
  OAI22xp33_ASAP7_75t_SL U29113 ( .A1(n31099), .A2(n30063), .B1(n31098), .B2(
        n30062), .Y(n30041) );
  OAI22xp33_ASAP7_75t_SL U29114 ( .A1(n31139), .A2(n31184), .B1(n31138), .B2(
        n31182), .Y(n31140) );
  OAI21xp33_ASAP7_75t_SL U29115 ( .A1(uart1_r_THOLD__31__0_), .A2(n27975), .B(
        n27974), .Y(n2043) );
  OAI22xp33_ASAP7_75t_SL U29116 ( .A1(n31095), .A2(n31184), .B1(n31094), .B2(
        n31182), .Y(n31096) );
  OAI21xp33_ASAP7_75t_SL U29117 ( .A1(uart1_r_THOLD__25__3_), .A2(n27920), .B(
        n27798), .Y(n1859) );
  OAI21xp33_ASAP7_75t_SL U29118 ( .A1(uart1_r_THOLD__28__0_), .A2(n27935), .B(
        n27934), .Y(n1886) );
  OAI21xp33_ASAP7_75t_SL U29119 ( .A1(n31412), .A2(n30366), .B(n30365), .Y(
        n30368) );
  OAI21xp33_ASAP7_75t_SL U29120 ( .A1(uart1_r_THOLD__29__6_), .A2(n27928), .B(
        n27589), .Y(n1888) );
  OAI21xp33_ASAP7_75t_SL U29121 ( .A1(uart1_r_THOLD__19__6_), .A2(n27968), .B(
        n27615), .Y(n1930) );
  OAI22xp33_ASAP7_75t_SL U29122 ( .A1(n31127), .A2(n30063), .B1(n31126), .B2(
        n30062), .Y(n30048) );
  OAI21xp33_ASAP7_75t_SL U29123 ( .A1(uart1_r_THOLD__28__2_), .A2(n27935), .B(
        n27861), .Y(n1884) );
  OAI21xp33_ASAP7_75t_SL U29124 ( .A1(uart1_r_THOLD__24__1_), .A2(n27947), .B(
        n27339), .Y(n2033) );
  OAI22xp33_ASAP7_75t_SL U29125 ( .A1(n31119), .A2(n31184), .B1(n31118), .B2(
        n31182), .Y(n31120) );
  OAI21xp33_ASAP7_75t_SL U29126 ( .A1(n30645), .A2(n29907), .B(n28797), .Y(
        n28798) );
  OAI21xp33_ASAP7_75t_SL U29127 ( .A1(uart1_r_THOLD__23__6_), .A2(n27973), .B(
        n27618), .Y(n1848) );
  OAI21xp33_ASAP7_75t_SL U29128 ( .A1(uart1_r_THOLD__31__5_), .A2(n27975), .B(
        n27687), .Y(n2038) );
  OAI21xp33_ASAP7_75t_SL U29129 ( .A1(uart1_r_THOLD__27__6_), .A2(n27967), .B(
        n27614), .Y(n1872) );
  OAI21xp33_ASAP7_75t_SL U29130 ( .A1(uart1_r_THOLD__16__1_), .A2(n27946), .B(
        n27337), .Y(n2029) );
  OAI21xp33_ASAP7_75t_SL U29131 ( .A1(uart1_r_THOLD__9__5_), .A2(n27929), .B(
        n27668), .Y(n1943) );
  OAI21xp33_ASAP7_75t_SL U29132 ( .A1(uart1_r_THOLD__19__1_), .A2(n27968), .B(
        n27375), .Y(n2030) );
  OAI21xp33_ASAP7_75t_SL U29133 ( .A1(uart1_r_THOLD__8__7_), .A2(n27933), .B(
        n27551), .Y(n1902) );
  OAI21xp33_ASAP7_75t_SL U29134 ( .A1(uart1_r_THOLD__30__4_), .A2(n27950), .B(
        n27735), .Y(n1974) );
  OAI21xp33_ASAP7_75t_SL U29135 ( .A1(uart1_r_THOLD__31__4_), .A2(n27975), .B(
        n27751), .Y(n2039) );
  OAI22xp33_ASAP7_75t_SL U29136 ( .A1(n31111), .A2(n30772), .B1(n31110), .B2(
        n30771), .Y(n30753) );
  OAI22xp33_ASAP7_75t_SL U29137 ( .A1(n31175), .A2(n30063), .B1(n31174), .B2(
        n30062), .Y(n30060) );
  OAI21xp33_ASAP7_75t_SL U29138 ( .A1(uart1_r_THOLD__31__6_), .A2(n27975), .B(
        n27619), .Y(n2037) );
  OAI21xp33_ASAP7_75t_SL U29139 ( .A1(uart1_r_THOLD__19__4_), .A2(n27968), .B(
        n27747), .Y(n1970) );
  OAI21xp33_ASAP7_75t_SL U29140 ( .A1(uart1_r_THOLD__22__6_), .A2(n27952), .B(
        n27605), .Y(n1932) );
  OAI22xp33_ASAP7_75t_SL U29141 ( .A1(n31163), .A2(n31184), .B1(n31162), .B2(
        n31182), .Y(n31164) );
  OAI22xp33_ASAP7_75t_SL U29142 ( .A1(n31185), .A2(n31184), .B1(n31183), .B2(
        n31182), .Y(n31186) );
  OAI22xp33_ASAP7_75t_SL U29143 ( .A1(n31091), .A2(n31184), .B1(n31090), .B2(
        n31182), .Y(n31092) );
  OAI22xp33_ASAP7_75t_SL U29144 ( .A1(n31143), .A2(n30866), .B1(n31142), .B2(
        n30865), .Y(n30855) );
  OAI21xp33_ASAP7_75t_SL U29145 ( .A1(uart1_r_THOLD__24__6_), .A2(n27947), .B(
        n27601), .Y(n1933) );
  OAI21xp33_ASAP7_75t_SL U29146 ( .A1(uart1_r_THOLD__14__1_), .A2(n27951), .B(
        n27359), .Y(n2028) );
  OAI22xp33_ASAP7_75t_SL U29147 ( .A1(n31063), .A2(n30866), .B1(n31062), .B2(
        n30865), .Y(n30835) );
  OAI21xp33_ASAP7_75t_SL U29148 ( .A1(uart1_r_THOLD__29__7_), .A2(n27928), .B(
        n27548), .Y(n1887) );
  OAI21xp33_ASAP7_75t_SL U29149 ( .A1(uart1_r_THOLD__16__4_), .A2(n27946), .B(
        n27732), .Y(n1969) );
  OAI22xp33_ASAP7_75t_SL U29150 ( .A1(n31155), .A2(n30063), .B1(n31154), .B2(
        n30062), .Y(n30055) );
  OAI21xp33_ASAP7_75t_SL U29151 ( .A1(uart1_r_THOLD__8__5_), .A2(n27933), .B(
        n27650), .Y(n1942) );
  OAI21xp33_ASAP7_75t_SL U29152 ( .A1(uart1_r_THOLD__27__5_), .A2(n27967), .B(
        n27682), .Y(n1873) );
  OAI21xp33_ASAP7_75t_SL U29153 ( .A1(uart1_r_THOLD__26__7_), .A2(n27962), .B(
        n27570), .Y(n1863) );
  OAI22xp33_ASAP7_75t_SL U29154 ( .A1(n31091), .A2(n30063), .B1(n31090), .B2(
        n30062), .Y(n30039) );
  OAI21xp33_ASAP7_75t_SL U29155 ( .A1(uart1_r_THOLD__10__5_), .A2(n27948), .B(
        n27670), .Y(n1944) );
  OAI21xp33_ASAP7_75t_SL U29156 ( .A1(uart1_r_THOLD__13__1_), .A2(n27931), .B(
        n27354), .Y(n2027) );
  OAI22xp33_ASAP7_75t_SL U29157 ( .A1(n31147), .A2(n31184), .B1(n31146), .B2(
        n31182), .Y(n31148) );
  NAND2xp33_ASAP7_75t_SL U29158 ( .A(n30435), .B(n28835), .Y(n28836) );
  OAI22xp33_ASAP7_75t_SL U29159 ( .A1(n31075), .A2(n30063), .B1(n31074), .B2(
        n30062), .Y(n30035) );
  OAI21xp33_ASAP7_75t_SL U29160 ( .A1(uart1_r_THOLD__25__1_), .A2(n27920), .B(
        n27344), .Y(n1861) );
  OAI21xp33_ASAP7_75t_SL U29161 ( .A1(n30645), .A2(n30464), .B(n28954), .Y(
        n28955) );
  OAI21xp33_ASAP7_75t_SL U29162 ( .A1(uart1_r_THOLD__31__3_), .A2(n27975), .B(
        n27823), .Y(n2040) );
  OAI22xp33_ASAP7_75t_SL U29163 ( .A1(n31071), .A2(n31184), .B1(n31070), .B2(
        n31182), .Y(n31072) );
  OAI21xp33_ASAP7_75t_SL U29164 ( .A1(uart1_r_THOLD__9__7_), .A2(n27929), .B(
        n27549), .Y(n1903) );
  OAI21xp33_ASAP7_75t_SL U29165 ( .A1(uart1_r_THOLD__21__1_), .A2(n27926), .B(
        n27349), .Y(n2031) );
  INVxp67_ASAP7_75t_SL U29166 ( .A(n28774), .Y(n28777) );
  OAI22xp33_ASAP7_75t_SL U29167 ( .A1(n31087), .A2(n31184), .B1(n31086), .B2(
        n31182), .Y(n31088) );
  INVxp33_ASAP7_75t_SL U29168 ( .A(n31617), .Y(n31619) );
  OAI21xp33_ASAP7_75t_SL U29169 ( .A1(uart1_r_THOLD__12__1_), .A2(n27937), .B(
        n27324), .Y(n2026) );
  OAI21xp33_ASAP7_75t_SL U29170 ( .A1(uart1_r_THOLD__22__1_), .A2(n27952), .B(
        n27360), .Y(n2032) );
  OAI22xp33_ASAP7_75t_SL U29171 ( .A1(n31119), .A2(n30063), .B1(n31118), .B2(
        n30062), .Y(n30046) );
  OAI22xp33_ASAP7_75t_SL U29172 ( .A1(n31143), .A2(n31184), .B1(n31142), .B2(
        n31182), .Y(n31144) );
  OAI22xp33_ASAP7_75t_SL U29173 ( .A1(n31179), .A2(n31184), .B1(n31178), .B2(
        n31182), .Y(n31180) );
  OAI22xp33_ASAP7_75t_SL U29174 ( .A1(n31083), .A2(n30866), .B1(n31082), .B2(
        n30865), .Y(n30840) );
  OAI21xp33_ASAP7_75t_SL U29175 ( .A1(uart1_r_THOLD__21__6_), .A2(n27926), .B(
        n27588), .Y(n1931) );
  OAI21xp33_ASAP7_75t_SL U29176 ( .A1(uart1_r_THOLD__14__4_), .A2(n27951), .B(
        n27736), .Y(n1968) );
  OAI21xp33_ASAP7_75t_SL U29177 ( .A1(uart1_r_THOLD__11__5_), .A2(n27977), .B(
        n27688), .Y(n1945) );
  OAI22xp33_ASAP7_75t_SL U29178 ( .A1(n31135), .A2(n30866), .B1(n31134), .B2(
        n30865), .Y(n30853) );
  OAI21xp33_ASAP7_75t_SL U29179 ( .A1(uart1_r_THOLD__10__7_), .A2(n27948), .B(
        n27561), .Y(n1904) );
  OAI21xp33_ASAP7_75t_SL U29180 ( .A1(uart1_r_THOLD__20__5_), .A2(n27939), .B(
        n27653), .Y(n1841) );
  OAI22xp33_ASAP7_75t_SL U29181 ( .A1(n31131), .A2(n30063), .B1(n31130), .B2(
        n30062), .Y(n30049) );
  OAI21xp33_ASAP7_75t_SL U29182 ( .A1(uart1_r_THOLD__11__1_), .A2(n27977), .B(
        n27386), .Y(n2025) );
  OAI21xp33_ASAP7_75t_SL U29183 ( .A1(uart1_r_THOLD__27__7_), .A2(n27967), .B(
        n27573), .Y(n1871) );
  OAI22xp33_ASAP7_75t_SL U29184 ( .A1(n31159), .A2(n30063), .B1(n31158), .B2(
        n30062), .Y(n30056) );
  OAI21xp33_ASAP7_75t_SL U29185 ( .A1(uart1_r_THOLD__23__5_), .A2(n27973), .B(
        n27686), .Y(n1849) );
  OAI21xp33_ASAP7_75t_SL U29186 ( .A1(uart1_r_THOLD__30__6_), .A2(n27950), .B(
        n27603), .Y(n1934) );
  OAI21xp33_ASAP7_75t_SL U29187 ( .A1(uart1_r_THOLD__31__7_), .A2(n27975), .B(
        n27578), .Y(n2036) );
  OAI22xp33_ASAP7_75t_SL U29188 ( .A1(n31175), .A2(n31184), .B1(n31174), .B2(
        n31182), .Y(n31176) );
  OAI21xp33_ASAP7_75t_SL U29189 ( .A1(uart1_r_THOLD__24__4_), .A2(n27947), .B(
        n27733), .Y(n1973) );
  OAI22xp33_ASAP7_75t_SL U29190 ( .A1(n31071), .A2(n30866), .B1(n31070), .B2(
        n30865), .Y(n30837) );
  OAI21xp33_ASAP7_75t_SL U29191 ( .A1(uart1_r_THOLD__31__2_), .A2(n27975), .B(
        n27887), .Y(n2041) );
  OAI21xp33_ASAP7_75t_SL U29192 ( .A1(uart1_r_THOLD__27__4_), .A2(n27967), .B(
        n27746), .Y(n1874) );
  OAI21xp33_ASAP7_75t_SL U29193 ( .A1(uart1_r_THOLD__26__6_), .A2(n27962), .B(
        n27611), .Y(n1864) );
  OAI22xp33_ASAP7_75t_SL U29194 ( .A1(n31139), .A2(n30866), .B1(n31138), .B2(
        n30865), .Y(n30854) );
  OAI21xp33_ASAP7_75t_SL U29195 ( .A1(uart1_r_THOLD__21__4_), .A2(n27926), .B(
        n27720), .Y(n1971) );
  AOI21xp33_ASAP7_75t_SL U29196 ( .A1(n28774), .A2(n28830), .B(n28773), .Y(
        n28775) );
  OAI21xp33_ASAP7_75t_SL U29197 ( .A1(uart1_r_THOLD__22__5_), .A2(n27952), .B(
        n27673), .Y(n1952) );
  OAI21xp33_ASAP7_75t_SL U29198 ( .A1(uart1_r_THOLD__22__7_), .A2(n27952), .B(
        n27564), .Y(n1912) );
  OAI21xp33_ASAP7_75t_SL U29199 ( .A1(uart1_r_THOLD__26__2_), .A2(n27962), .B(
        n27879), .Y(n1868) );
  OAI21xp33_ASAP7_75t_SL U29200 ( .A1(uart1_r_THOLD__10__3_), .A2(n27948), .B(
        n27806), .Y(n1984) );
  OAI21xp33_ASAP7_75t_SL U29201 ( .A1(uart1_r_THOLD__29__0_), .A2(n27928), .B(
        n27927), .Y(n1894) );
  OAI22xp33_ASAP7_75t_SL U29202 ( .A1(n31071), .A2(n30063), .B1(n31070), .B2(
        n30062), .Y(n30034) );
  OAI21xp33_ASAP7_75t_SL U29203 ( .A1(uart1_r_THOLD__20__1_), .A2(n27939), .B(
        n27326), .Y(n1845) );
  NOR2xp33_ASAP7_75t_SRAM U29204 ( .A(n3068), .B(n32193), .Y(n32201) );
  OAI22xp33_ASAP7_75t_SL U29205 ( .A1(n31123), .A2(n31184), .B1(n31122), .B2(
        n31182), .Y(n31124) );
  OAI21xp33_ASAP7_75t_SL U29206 ( .A1(uart1_r_THOLD__9__4_), .A2(n27929), .B(
        n27722), .Y(n1963) );
  OAI22xp33_ASAP7_75t_SL U29207 ( .A1(n31107), .A2(n30866), .B1(n31106), .B2(
        n30865), .Y(n30846) );
  OAI22xp33_ASAP7_75t_SL U29208 ( .A1(n31131), .A2(n30866), .B1(n31130), .B2(
        n30865), .Y(n30852) );
  OAI22xp33_ASAP7_75t_SL U29209 ( .A1(n31063), .A2(n30063), .B1(n31062), .B2(
        n30062), .Y(n30032) );
  OAI21xp33_ASAP7_75t_SL U29210 ( .A1(uart1_r_THOLD__24__5_), .A2(n27947), .B(
        n27659), .Y(n1953) );
  INVxp67_ASAP7_75t_SL U29211 ( .A(n24173), .Y(n22650) );
  OAI21xp33_ASAP7_75t_SL U29212 ( .A1(uart1_r_THOLD__12__2_), .A2(n27937), .B(
        n27862), .Y(n2006) );
  OAI21xp33_ASAP7_75t_SL U29213 ( .A1(uart1_r_THOLD__30__2_), .A2(n27950), .B(
        n27871), .Y(n2014) );
  OAI21xp33_ASAP7_75t_SL U29214 ( .A1(uart1_r_THOLD__24__2_), .A2(n27947), .B(
        n27869), .Y(n2013) );
  OAI21xp33_ASAP7_75t_SL U29215 ( .A1(uart1_r_THOLD__27__0_), .A2(n27967), .B(
        n27966), .Y(n1878) );
  OAI22xp33_ASAP7_75t_SL U29216 ( .A1(n31067), .A2(n31184), .B1(n31066), .B2(
        n31182), .Y(n31068) );
  OAI22xp33_ASAP7_75t_SL U29217 ( .A1(n31155), .A2(n30866), .B1(n31154), .B2(
        n30865), .Y(n30858) );
  OAI21xp33_ASAP7_75t_SL U29218 ( .A1(uart1_r_THOLD__24__7_), .A2(n27947), .B(
        n27560), .Y(n1913) );
  OAI22xp33_ASAP7_75t_SL U29219 ( .A1(n31087), .A2(n30866), .B1(n31086), .B2(
        n30865), .Y(n30841) );
  OAI22xp33_ASAP7_75t_SL U29220 ( .A1(n31171), .A2(n31184), .B1(n31170), .B2(
        n31182), .Y(n31172) );
  OAI21xp33_ASAP7_75t_SL U29221 ( .A1(n30446), .A2(n30291), .B(n30290), .Y(
        n30294) );
  OAI21xp33_ASAP7_75t_SL U29222 ( .A1(uart1_r_THOLD__26__1_), .A2(n27962), .B(
        n27370), .Y(n1869) );
  OAI21xp33_ASAP7_75t_SL U29223 ( .A1(uart1_r_THOLD__8__4_), .A2(n27933), .B(
        n27724), .Y(n1962) );
  OAI21xp33_ASAP7_75t_SL U29224 ( .A1(uart1_r_THOLD__22__2_), .A2(n27952), .B(
        n27873), .Y(n2012) );
  OAI21xp33_ASAP7_75t_SL U29225 ( .A1(uart1_r_THOLD__30__5_), .A2(n27950), .B(
        n27671), .Y(n1954) );
  OAI21xp33_ASAP7_75t_SL U29226 ( .A1(uart1_r_THOLD__11__6_), .A2(n27977), .B(
        n27620), .Y(n1925) );
  OAI22xp33_ASAP7_75t_SL U29227 ( .A1(n31099), .A2(n30866), .B1(n31098), .B2(
        n30865), .Y(n30844) );
  OAI22xp33_ASAP7_75t_SL U29228 ( .A1(n31075), .A2(n31184), .B1(n31074), .B2(
        n31182), .Y(n31076) );
  OAI21xp33_ASAP7_75t_SL U29229 ( .A1(uart1_r_THOLD__30__7_), .A2(n27950), .B(
        n27562), .Y(n1914) );
  OAI21xp33_ASAP7_75t_SL U29230 ( .A1(uart1_r_THOLD__29__1_), .A2(n27928), .B(
        n27350), .Y(n1893) );
  OAI22xp33_ASAP7_75t_SL U29231 ( .A1(n31107), .A2(n31184), .B1(n31106), .B2(
        n31182), .Y(n31108) );
  OAI22xp33_ASAP7_75t_SL U29232 ( .A1(n31143), .A2(n30063), .B1(n31142), .B2(
        n30062), .Y(n30052) );
  OAI21xp33_ASAP7_75t_SL U29233 ( .A1(uart1_r_THOLD__23__0_), .A2(n27973), .B(
        n27972), .Y(n1854) );
  OAI21xp33_ASAP7_75t_SL U29234 ( .A1(uart1_r_THOLD__13__2_), .A2(n27931), .B(
        n27859), .Y(n2007) );
  OAI22xp33_ASAP7_75t_SL U29235 ( .A1(n31083), .A2(n30063), .B1(n31082), .B2(
        n30062), .Y(n30037) );
  OAI21xp33_ASAP7_75t_SL U29236 ( .A1(n30645), .A2(n28576), .B(n28575), .Y(
        n28577) );
  OAI22xp33_ASAP7_75t_SL U29237 ( .A1(n31119), .A2(n30866), .B1(n31118), .B2(
        n30865), .Y(n30849) );
  OAI21xp33_ASAP7_75t_SL U29238 ( .A1(uart1_r_THOLD__11__3_), .A2(n27977), .B(
        n27824), .Y(n1985) );
  OAI21xp33_ASAP7_75t_SL U29239 ( .A1(uart1_r_THOLD__26__0_), .A2(n27962), .B(
        n27961), .Y(n1870) );
  OAI21xp33_ASAP7_75t_SL U29240 ( .A1(uart1_r_THOLD__16__3_), .A2(n27946), .B(
        n27794), .Y(n1989) );
  OAI22xp33_ASAP7_75t_SL U29241 ( .A1(n31111), .A2(n31184), .B1(n31110), .B2(
        n31182), .Y(n31112) );
  OAI21xp33_ASAP7_75t_SL U29242 ( .A1(uart1_r_THOLD__21__2_), .A2(n27926), .B(
        n27856), .Y(n2011) );
  OAI21xp33_ASAP7_75t_SL U29243 ( .A1(uart1_r_THOLD__27__1_), .A2(n27967), .B(
        n27374), .Y(n1877) );
  OAI21xp33_ASAP7_75t_SL U29244 ( .A1(uart1_r_THOLD__29__2_), .A2(n27928), .B(
        n27857), .Y(n1892) );
  INVxp33_ASAP7_75t_SL U29245 ( .A(n31572), .Y(n31618) );
  OAI21xp33_ASAP7_75t_SL U29246 ( .A1(uart1_r_THOLD__14__3_), .A2(n27951), .B(
        n27808), .Y(n1988) );
  OAI22xp33_ASAP7_75t_SL U29247 ( .A1(n31175), .A2(n30866), .B1(n31174), .B2(
        n30865), .Y(n30863) );
  OAI21xp33_ASAP7_75t_SL U29248 ( .A1(uart1_r_THOLD__10__6_), .A2(n27948), .B(
        n27602), .Y(n1924) );
  OAI21xp33_ASAP7_75t_SL U29249 ( .A1(uart1_r_THOLD__19__2_), .A2(n27968), .B(
        n27883), .Y(n2010) );
  OAI22xp33_ASAP7_75t_SL U29250 ( .A1(n31099), .A2(n31184), .B1(n31098), .B2(
        n31182), .Y(n31100) );
  OAI22xp33_ASAP7_75t_SL U29251 ( .A1(n31079), .A2(n30063), .B1(n31078), .B2(
        n30062), .Y(n30036) );
  OAI21xp33_ASAP7_75t_SL U29252 ( .A1(uart1_r_THOLD__23__1_), .A2(n27973), .B(
        n27382), .Y(n1853) );
  OAI21xp33_ASAP7_75t_SL U29253 ( .A1(uart1_r_THOLD__29__3_), .A2(n27928), .B(
        n27803), .Y(n1891) );
  OAI22xp33_ASAP7_75t_SL U29254 ( .A1(n31139), .A2(n30063), .B1(n31138), .B2(
        n30062), .Y(n30051) );
  NAND2xp5_ASAP7_75t_SL U29255 ( .A(n23358), .B(n22706), .Y(n22705) );
  OAI22xp33_ASAP7_75t_SL U29256 ( .A1(n31159), .A2(n30866), .B1(n31158), .B2(
        n30865), .Y(n30859) );
  OAI21xp33_ASAP7_75t_SL U29257 ( .A1(uart1_r_THOLD__23__7_), .A2(n27973), .B(
        n27577), .Y(n1847) );
  OAI21xp33_ASAP7_75t_SL U29258 ( .A1(uart1_r_THOLD__12__3_), .A2(n27937), .B(
        n27788), .Y(n1986) );
  OAI21xp33_ASAP7_75t_SL U29259 ( .A1(uart1_r_THOLD__20__0_), .A2(n27939), .B(
        n27938), .Y(n1846) );
  OAI22xp33_ASAP7_75t_SL U29260 ( .A1(n31179), .A2(n30866), .B1(n31178), .B2(
        n30865), .Y(n30864) );
  INVxp67_ASAP7_75t_SL U29261 ( .A(n29584), .Y(n26216) );
  OAI21xp33_ASAP7_75t_SL U29262 ( .A1(uart1_r_THOLD__14__2_), .A2(n27951), .B(
        n27872), .Y(n2008) );
  OAI21xp33_ASAP7_75t_SL U29263 ( .A1(uart1_r_THOLD__27__2_), .A2(n27967), .B(
        n27882), .Y(n1876) );
  OAI21xp33_ASAP7_75t_SL U29264 ( .A1(uart1_r_THOLD__13__3_), .A2(n27931), .B(
        n27805), .Y(n1987) );
  OAI22xp33_ASAP7_75t_SL U29265 ( .A1(n31147), .A2(n30866), .B1(n31146), .B2(
        n30865), .Y(n30856) );
  OAI21xp33_ASAP7_75t_SL U29266 ( .A1(n30445), .A2(n29595), .B(n28891), .Y(
        n28892) );
  OAI22xp33_ASAP7_75t_SL U29267 ( .A1(n31091), .A2(n30866), .B1(n31090), .B2(
        n30865), .Y(n30842) );
  OAI21xp33_ASAP7_75t_SL U29268 ( .A1(uart1_r_THOLD__8__6_), .A2(n27933), .B(
        n27592), .Y(n1922) );
  OAI21xp33_ASAP7_75t_SL U29269 ( .A1(uart1_r_THOLD__23__2_), .A2(n27973), .B(
        n27886), .Y(n1852) );
  OAI22xp33_ASAP7_75t_SL U29270 ( .A1(n31075), .A2(n30866), .B1(n31074), .B2(
        n30865), .Y(n30838) );
  OAI22xp33_ASAP7_75t_SL U29271 ( .A1(n31159), .A2(n31184), .B1(n31158), .B2(
        n31182), .Y(n31160) );
  OAI21xp33_ASAP7_75t_SL U29272 ( .A1(uart1_r_THOLD__16__2_), .A2(n27946), .B(
        n27868), .Y(n2009) );
  OAI21xp33_ASAP7_75t_SL U29273 ( .A1(uart1_r_THOLD__9__6_), .A2(n27929), .B(
        n27590), .Y(n1923) );
  OAI22xp33_ASAP7_75t_SL U29274 ( .A1(n31185), .A2(n30866), .B1(n31183), .B2(
        n30865), .Y(n30867) );
  OAI21xp33_ASAP7_75t_SL U29275 ( .A1(uart1_r_THOLD__13__4_), .A2(n27931), .B(
        n27723), .Y(n1967) );
  OAI21xp33_ASAP7_75t_SL U29276 ( .A1(uart1_r_THOLD__8__2_), .A2(n27933), .B(
        n27860), .Y(n2002) );
  OAI21xp33_ASAP7_75t_SL U29277 ( .A1(uart1_r_THOLD__14__5_), .A2(n27951), .B(
        n27672), .Y(n1948) );
  OAI21xp33_ASAP7_75t_SL U29278 ( .A1(uart1_r_THOLD__8__1_), .A2(n27933), .B(
        n27311), .Y(n2022) );
  OAI22xp33_ASAP7_75t_SL U29279 ( .A1(n31115), .A2(n30063), .B1(n31114), .B2(
        n30062), .Y(n30045) );
  OAI22xp33_ASAP7_75t_SL U29280 ( .A1(n31131), .A2(n31184), .B1(n31130), .B2(
        n31182), .Y(n31132) );
  OAI22xp33_ASAP7_75t_SL U29281 ( .A1(n31111), .A2(n30866), .B1(n31110), .B2(
        n30865), .Y(n30847) );
  NAND2xp33_ASAP7_75t_SL U29282 ( .A(n30453), .B(n30452), .Y(n30457) );
  OAI21xp33_ASAP7_75t_SL U29283 ( .A1(uart1_r_THOLD__23__4_), .A2(n27973), .B(
        n27750), .Y(n1850) );
  OAI21xp33_ASAP7_75t_SL U29284 ( .A1(uart1_r_THOLD__16__5_), .A2(n27946), .B(
        n27658), .Y(n1949) );
  OAI21xp33_ASAP7_75t_SL U29285 ( .A1(uart1_r_THOLD__14__6_), .A2(n27951), .B(
        n27604), .Y(n1928) );
  OAI21xp33_ASAP7_75t_SL U29286 ( .A1(uart1_r_THOLD__25__4_), .A2(n27920), .B(
        n27716), .Y(n1858) );
  OAI21xp33_ASAP7_75t_SL U29287 ( .A1(uart1_r_THOLD__29__5_), .A2(n27928), .B(
        n27667), .Y(n1889) );
  OAI21xp33_ASAP7_75t_SL U29288 ( .A1(uart1_r_THOLD__20__3_), .A2(n27939), .B(
        n27789), .Y(n1843) );
  OAI22xp33_ASAP7_75t_SL U29289 ( .A1(n31115), .A2(n30866), .B1(n31114), .B2(
        n30865), .Y(n30848) );
  OAI22xp33_ASAP7_75t_SL U29290 ( .A1(n31067), .A2(n30063), .B1(n31066), .B2(
        n30062), .Y(n30033) );
  OAI22xp33_ASAP7_75t_SL U29291 ( .A1(n31123), .A2(n30866), .B1(n31122), .B2(
        n30865), .Y(n30850) );
  OAI21xp33_ASAP7_75t_SL U29292 ( .A1(uart1_r_THOLD__12__7_), .A2(n27937), .B(
        n27553), .Y(n1906) );
  OAI21xp33_ASAP7_75t_SL U29293 ( .A1(uart1_r_THOLD__29__4_), .A2(n27928), .B(
        n27721), .Y(n1890) );
  OAI21xp33_ASAP7_75t_SL U29294 ( .A1(uart1_r_THOLD__28__5_), .A2(n27935), .B(
        n27651), .Y(n1881) );
  OAI22xp33_ASAP7_75t_SL U29295 ( .A1(n31171), .A2(n30866), .B1(n31170), .B2(
        n30865), .Y(n30862) );
  OAI22xp33_ASAP7_75t_SL U29296 ( .A1(n31079), .A2(n31184), .B1(n31078), .B2(
        n31182), .Y(n31080) );
  OAI22xp33_ASAP7_75t_SL U29297 ( .A1(n31103), .A2(n30063), .B1(n31102), .B2(
        n30062), .Y(n30042) );
  NOR2x1_ASAP7_75t_SL U29298 ( .A(n24240), .B(n24239), .Y(n24241) );
  OAI21xp33_ASAP7_75t_SL U29299 ( .A1(uart1_r_THOLD__12__4_), .A2(n27937), .B(
        n27726), .Y(n1966) );
  OAI21xp33_ASAP7_75t_SL U29300 ( .A1(uart1_r_THOLD__9__2_), .A2(n27929), .B(
        n27858), .Y(n2003) );
  OAI21xp33_ASAP7_75t_SL U29301 ( .A1(n30446), .A2(n30376), .B(n30375), .Y(
        n30379) );
  OAI22xp33_ASAP7_75t_SL U29302 ( .A1(n31167), .A2(n31184), .B1(n31166), .B2(
        n31182), .Y(n31168) );
  OAI22xp33_ASAP7_75t_SL U29303 ( .A1(n31123), .A2(n30063), .B1(n31122), .B2(
        n30062), .Y(n30047) );
  OAI21xp33_ASAP7_75t_SL U29304 ( .A1(uart1_r_THOLD__26__5_), .A2(n27962), .B(
        n27679), .Y(n1865) );
  OAI21xp33_ASAP7_75t_SL U29305 ( .A1(uart1_r_THOLD__13__6_), .A2(n27931), .B(
        n27591), .Y(n1927) );
  OAI22xp33_ASAP7_75t_SL U29306 ( .A1(n31103), .A2(n30866), .B1(n31102), .B2(
        n30865), .Y(n30845) );
  OAI22xp33_ASAP7_75t_SL U29307 ( .A1(n31083), .A2(n31184), .B1(n31082), .B2(
        n31182), .Y(n31084) );
  OAI22xp33_ASAP7_75t_SL U29308 ( .A1(n31185), .A2(n30063), .B1(n31183), .B2(
        n30062), .Y(n30064) );
  OAI21xp33_ASAP7_75t_SL U29309 ( .A1(uart1_r_THOLD__13__7_), .A2(n27931), .B(
        n27550), .Y(n1907) );
  OAI21xp33_ASAP7_75t_SL U29310 ( .A1(uart1_r_THOLD__28__6_), .A2(n27935), .B(
        n27593), .Y(n1880) );
  OAI21xp33_ASAP7_75t_SL U29311 ( .A1(uart1_r_THOLD__25__5_), .A2(n27920), .B(
        n27662), .Y(n1857) );
  INVxp67_ASAP7_75t_SL U29312 ( .A(n30451), .Y(n30462) );
  OAI21xp33_ASAP7_75t_SL U29313 ( .A1(uart1_r_THOLD__28__4_), .A2(n27935), .B(
        n27725), .Y(n1882) );
  OAI22xp33_ASAP7_75t_SL U29314 ( .A1(n31171), .A2(n30063), .B1(n31170), .B2(
        n30062), .Y(n30059) );
  OAI21xp33_ASAP7_75t_SL U29315 ( .A1(uart1_r_THOLD__19__5_), .A2(n27968), .B(
        n27683), .Y(n1950) );
  OAI21xp33_ASAP7_75t_SL U29316 ( .A1(uart1_r_THOLD__20__2_), .A2(n27939), .B(
        n27863), .Y(n1844) );
  OAI21xp33_ASAP7_75t_SL U29317 ( .A1(uart1_r_THOLD__8__3_), .A2(n27933), .B(
        n27786), .Y(n1982) );
  OAI21xp33_ASAP7_75t_SL U29318 ( .A1(uart1_r_THOLD__11__4_), .A2(n27977), .B(
        n27752), .Y(n1965) );
  OAI21xp33_ASAP7_75t_SL U29319 ( .A1(uart1_r_THOLD__21__3_), .A2(n27926), .B(
        n27802), .Y(n1991) );
  OAI21xp33_ASAP7_75t_SL U29320 ( .A1(uart1_r_THOLD__26__4_), .A2(n27962), .B(
        n27743), .Y(n1866) );
  OAI21xp33_ASAP7_75t_SL U29321 ( .A1(uart1_r_THOLD__21__5_), .A2(n27926), .B(
        n27666), .Y(n1951) );
  OAI22xp33_ASAP7_75t_SL U29322 ( .A1(n31151), .A2(n31184), .B1(n31150), .B2(
        n31182), .Y(n31152) );
  OAI22xp33_ASAP7_75t_SL U29323 ( .A1(n31151), .A2(n30866), .B1(n31150), .B2(
        n30865), .Y(n30857) );
  OAI22xp33_ASAP7_75t_SL U29324 ( .A1(n31063), .A2(n31184), .B1(n31062), .B2(
        n31182), .Y(n31064) );
  OAI21xp33_ASAP7_75t_SL U29325 ( .A1(uart1_r_THOLD__25__6_), .A2(n27920), .B(
        n27584), .Y(n1856) );
  OAI21xp33_ASAP7_75t_SL U29326 ( .A1(uart1_r_THOLD__14__7_), .A2(n27951), .B(
        n27563), .Y(n1908) );
  OAI22xp33_ASAP7_75t_SL U29327 ( .A1(n31163), .A2(n30063), .B1(n31162), .B2(
        n30062), .Y(n30057) );
  OAI21xp33_ASAP7_75t_SL U29328 ( .A1(uart1_r_THOLD__10__2_), .A2(n27948), .B(
        n27870), .Y(n2004) );
  OAI21xp33_ASAP7_75t_SL U29329 ( .A1(uart1_r_THOLD__16__7_), .A2(n27946), .B(
        n27559), .Y(n1909) );
  OAI21xp33_ASAP7_75t_SL U29330 ( .A1(uart1_r_THOLD__28__7_), .A2(n27935), .B(
        n27552), .Y(n1879) );
  OAI21xp33_ASAP7_75t_SL U29331 ( .A1(uart1_r_THOLD__10__4_), .A2(n27948), .B(
        n27734), .Y(n1964) );
  OAI22xp33_ASAP7_75t_SL U29332 ( .A1(n31067), .A2(n30866), .B1(n31066), .B2(
        n30865), .Y(n30836) );
  OAI21xp33_ASAP7_75t_SL U29333 ( .A1(uart1_r_THOLD__19__7_), .A2(n27968), .B(
        n27574), .Y(n1910) );
  OAI21xp33_ASAP7_75t_SL U29334 ( .A1(uart1_r_THOLD__12__6_), .A2(n27937), .B(
        n27594), .Y(n1926) );
  OAI21xp33_ASAP7_75t_SL U29335 ( .A1(uart1_r_THOLD__27__3_), .A2(n27967), .B(
        n27818), .Y(n1875) );
  OAI21xp33_ASAP7_75t_SL U29336 ( .A1(uart1_r_THOLD__9__3_), .A2(n27929), .B(
        n27804), .Y(n1983) );
  OAI21xp33_ASAP7_75t_SL U29337 ( .A1(uart1_r_THOLD__19__3_), .A2(n27968), .B(
        n27819), .Y(n1990) );
  OAI22xp33_ASAP7_75t_SL U29338 ( .A1(n31135), .A2(n30063), .B1(n31134), .B2(
        n30062), .Y(n30050) );
  OAI21xp33_ASAP7_75t_SL U29339 ( .A1(uart1_r_THOLD__11__2_), .A2(n27977), .B(
        n27888), .Y(n2005) );
  OAI22xp33_ASAP7_75t_SL U29340 ( .A1(n31111), .A2(n30063), .B1(n31110), .B2(
        n30062), .Y(n30044) );
  OAI22xp33_ASAP7_75t_SL U29341 ( .A1(n31167), .A2(n30866), .B1(n31166), .B2(
        n30865), .Y(n30861) );
  OAI22xp33_ASAP7_75t_SL U29342 ( .A1(n31135), .A2(n31184), .B1(n31134), .B2(
        n31182), .Y(n31136) );
  OAI21xp33_ASAP7_75t_SL U29343 ( .A1(uart1_r_THOLD__25__7_), .A2(n27920), .B(
        n27543), .Y(n1855) );
  OAI21xp33_ASAP7_75t_SL U29344 ( .A1(uart1_r_THOLD__26__3_), .A2(n27962), .B(
        n27815), .Y(n1867) );
  OAI22xp33_ASAP7_75t_SL U29345 ( .A1(n31103), .A2(n31184), .B1(n31102), .B2(
        n31182), .Y(n31104) );
  INVx1_ASAP7_75t_SL U29346 ( .A(n30783), .Y(n31241) );
  OAI21xp33_ASAP7_75t_SL U29347 ( .A1(uart1_r_THOLD__23__3_), .A2(n27973), .B(
        n27822), .Y(n1851) );
  OAI22xp33_ASAP7_75t_SL U29348 ( .A1(n31095), .A2(n30866), .B1(n31094), .B2(
        n30865), .Y(n30843) );
  OAI21xp33_ASAP7_75t_SL U29349 ( .A1(uart1_r_THOLD__21__7_), .A2(n27926), .B(
        n27547), .Y(n1911) );
  OAI21xp33_ASAP7_75t_SL U29350 ( .A1(uart1_r_THOLD__30__1_), .A2(n27950), .B(
        n27358), .Y(n2034) );
  NAND2xp33_ASAP7_75t_SL U29351 ( .A(n25901), .B(n25627), .Y(n29587) );
  AOI22xp33_ASAP7_75t_SL U29352 ( .A1(n28835), .A2(n30340), .B1(
        u0_0_leon3x0_p0_divi[46]), .B2(n28782), .Y(n26577) );
  INVxp33_ASAP7_75t_SL U29353 ( .A(n26567), .Y(n26569) );
  NAND2xp33_ASAP7_75t_SL U29354 ( .A(n28132), .B(n26585), .Y(n26586) );
  OAI21xp33_ASAP7_75t_SL U29355 ( .A1(n30645), .A2(n28556), .B(n28555), .Y(
        n28557) );
  AOI22xp33_ASAP7_75t_SL U29356 ( .A1(n28554), .A2(n29598), .B1(n23665), .B2(
        n29583), .Y(n26689) );
  NAND2xp33_ASAP7_75t_SL U29357 ( .A(n28830), .B(n26684), .Y(n26685) );
  INVxp33_ASAP7_75t_SL U29358 ( .A(n26684), .Y(n26688) );
  INVxp33_ASAP7_75t_SL U29359 ( .A(n29003), .Y(n26674) );
  INVx1_ASAP7_75t_SL U29360 ( .A(n28855), .Y(n28920) );
  NAND2xp5_ASAP7_75t_SL U29361 ( .A(n25097), .B(n25096), .Y(n26424) );
  NAND2xp33_ASAP7_75t_SL U29362 ( .A(n29426), .B(n29383), .Y(n29233) );
  OAI22xp33_ASAP7_75t_SL U29363 ( .A1(n30376), .A2(n29595), .B1(n28633), .B2(
        n28632), .Y(n28639) );
  NAND2xp33_ASAP7_75t_SL U29364 ( .A(n29988), .B(n31840), .Y(n26491) );
  OAI21xp33_ASAP7_75t_SL U29365 ( .A1(n30407), .A2(n30701), .B(n29210), .Y(
        n29222) );
  NAND2xp33_ASAP7_75t_SL U29366 ( .A(n29270), .B(n29383), .Y(n29271) );
  INVxp33_ASAP7_75t_SL U29367 ( .A(n28668), .Y(n28672) );
  AOI22xp33_ASAP7_75t_SL U29368 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__2_), 
        .A2(n24648), .B1(n31442), .B2(n29699), .Y(n3354) );
  NAND2xp33_ASAP7_75t_SL U29369 ( .A(n26626), .B(n31840), .Y(n26623) );
  NAND2xp33_ASAP7_75t_SL U29370 ( .A(n25907), .B(n25476), .Y(n25794) );
  OAI21xp33_ASAP7_75t_SL U29371 ( .A1(n30645), .A2(n29693), .B(n28813), .Y(
        n28814) );
  OAI22xp33_ASAP7_75t_SL U29372 ( .A1(n31059), .A2(n30772), .B1(n31058), .B2(
        n30771), .Y(n30740) );
  OAI21xp33_ASAP7_75t_SL U29373 ( .A1(n30701), .A2(n30699), .B(n30698), .Y(
        n18089) );
  OAI22xp33_ASAP7_75t_SL U29374 ( .A1(n31059), .A2(n30063), .B1(n31058), .B2(
        n30062), .Y(n30031) );
  OAI21xp33_ASAP7_75t_SL U29375 ( .A1(n30701), .A2(n30696), .B(n30695), .Y(
        n18090) );
  OAI21xp33_ASAP7_75t_SL U29376 ( .A1(n18614), .A2(n25198), .B(n25189), .Y(
        n25782) );
  INVxp67_ASAP7_75t_SL U29377 ( .A(n28966), .Y(n26299) );
  OAI22xp33_ASAP7_75t_SL U29378 ( .A1(n31059), .A2(n31184), .B1(n31058), .B2(
        n31182), .Y(n31060) );
  OAI22xp33_ASAP7_75t_SL U29379 ( .A1(n31059), .A2(n30866), .B1(n31058), .B2(
        n30865), .Y(n30834) );
  INVxp33_ASAP7_75t_SL U29380 ( .A(n26293), .Y(n26297) );
  NOR2xp33_ASAP7_75t_SL U29381 ( .A(n23162), .B(u0_0_leon3x0_p0_divi[25]), .Y(
        n25493) );
  AND2x2_ASAP7_75t_SL U29382 ( .A(n22556), .B(n29583), .Y(n23163) );
  NAND2xp33_ASAP7_75t_SL U29383 ( .A(n29420), .B(n29383), .Y(n29303) );
  NAND2xp33_ASAP7_75t_SL U29384 ( .A(n31941), .B(n31840), .Y(n26478) );
  NAND2xp33_ASAP7_75t_SL U29385 ( .A(n31244), .B(n31840), .Y(n26630) );
  INVxp67_ASAP7_75t_SL U29386 ( .A(mult_x_1196_n2151), .Y(n22796) );
  INVx1_ASAP7_75t_SL U29387 ( .A(n28970), .Y(n28979) );
  AOI22xp33_ASAP7_75t_SL U29388 ( .A1(dc_q[25]), .A2(n31004), .B1(dt_q[21]), 
        .B2(n29991), .Y(n28410) );
  OAI21xp33_ASAP7_75t_SL U29389 ( .A1(n30446), .A2(n30445), .B(n30444), .Y(
        n30448) );
  NAND2xp33_ASAP7_75t_SL U29390 ( .A(n25626), .B(n29584), .Y(n28488) );
  AOI22xp33_ASAP7_75t_SL U29391 ( .A1(dc_q[29]), .A2(n31004), .B1(dt_q[25]), 
        .B2(n24573), .Y(n25416) );
  OAI22xp33_ASAP7_75t_SL U29392 ( .A1(n31139), .A2(n26127), .B1(n31138), .B2(
        n26126), .Y(n26115) );
  AOI22xp33_ASAP7_75t_SL U29393 ( .A1(it_q[17]), .A2(n24636), .B1(dc_q[21]), 
        .B2(n31473), .Y(n26332) );
  OAI22xp33_ASAP7_75t_SL U29394 ( .A1(n31139), .A2(n26069), .B1(n29956), .B2(
        n31138), .Y(n26030) );
  INVxp33_ASAP7_75t_SL U29395 ( .A(n31873), .Y(n30819) );
  OAI22xp33_ASAP7_75t_SL U29396 ( .A1(n31127), .A2(n26127), .B1(n31126), .B2(
        n26126), .Y(n26112) );
  OAI22xp33_ASAP7_75t_SL U29397 ( .A1(n31127), .A2(n26069), .B1(n29956), .B2(
        n31126), .Y(n26027) );
  OAI22xp33_ASAP7_75t_SL U29398 ( .A1(n31079), .A2(n26127), .B1(n31078), .B2(
        n26126), .Y(n26102) );
  OAI22xp33_ASAP7_75t_SL U29399 ( .A1(n31079), .A2(n26069), .B1(n29956), .B2(
        n31078), .Y(n26010) );
  OAI22xp33_ASAP7_75t_SL U29400 ( .A1(n31083), .A2(n26127), .B1(n31082), .B2(
        n26126), .Y(n26103) );
  OAI22xp33_ASAP7_75t_SL U29401 ( .A1(n31083), .A2(n26069), .B1(n29956), .B2(
        n31082), .Y(n26011) );
  OAI22xp33_ASAP7_75t_SL U29402 ( .A1(n31063), .A2(n26127), .B1(n31062), .B2(
        n26126), .Y(n26096) );
  OAI22xp33_ASAP7_75t_SL U29403 ( .A1(n31063), .A2(n26069), .B1(n29956), .B2(
        n31062), .Y(n26000) );
  OAI22xp33_ASAP7_75t_SL U29404 ( .A1(n31135), .A2(n26127), .B1(n31134), .B2(
        n26126), .Y(n26114) );
  AOI211xp5_ASAP7_75t_SL U29405 ( .A1(n24578), .A2(n23665), .B(n26155), .C(
        n24473), .Y(n28849) );
  OAI22xp33_ASAP7_75t_SL U29406 ( .A1(n31135), .A2(n26069), .B1(n29956), .B2(
        n31134), .Y(n26029) );
  OAI22xp33_ASAP7_75t_SL U29407 ( .A1(n31123), .A2(n26127), .B1(n31122), .B2(
        n26126), .Y(n26111) );
  OAI22xp33_ASAP7_75t_SL U29408 ( .A1(n31123), .A2(n26069), .B1(n29956), .B2(
        n31122), .Y(n26026) );
  OAI22xp33_ASAP7_75t_SL U29409 ( .A1(n31067), .A2(n26127), .B1(n31066), .B2(
        n26126), .Y(n26099) );
  OAI22xp33_ASAP7_75t_SL U29410 ( .A1(n31067), .A2(n26069), .B1(n29956), .B2(
        n31066), .Y(n26002) );
  NAND2xp33_ASAP7_75t_SL U29411 ( .A(n30356), .B(n28835), .Y(n27204) );
  OAI22xp33_ASAP7_75t_SL U29412 ( .A1(n31107), .A2(n26127), .B1(n31106), .B2(
        n26126), .Y(n26108) );
  AOI22xp33_ASAP7_75t_SL U29413 ( .A1(u0_0_leon3x0_p0_divi[13]), .A2(n27200), 
        .B1(n28830), .B2(n27199), .Y(n27201) );
  OAI22xp33_ASAP7_75t_SL U29414 ( .A1(n31107), .A2(n26069), .B1(n29956), .B2(
        n31106), .Y(n26022) );
  INVxp33_ASAP7_75t_SL U29415 ( .A(n27199), .Y(n27202) );
  OAI22xp33_ASAP7_75t_SL U29416 ( .A1(n31159), .A2(n26127), .B1(n31158), .B2(
        n26126), .Y(n26120) );
  NAND2xp5_ASAP7_75t_SL U29417 ( .A(n24477), .B(n25797), .Y(n26552) );
  OAI22xp33_ASAP7_75t_SL U29418 ( .A1(n31159), .A2(n26069), .B1(n29956), .B2(
        n31158), .Y(n26046) );
  NAND2xp5_ASAP7_75t_SL U29419 ( .A(n25796), .B(n25795), .Y(n26551) );
  OAI22xp33_ASAP7_75t_SL U29420 ( .A1(n31075), .A2(n26127), .B1(n31074), .B2(
        n26126), .Y(n26101) );
  OAI22xp33_ASAP7_75t_SL U29421 ( .A1(n31075), .A2(n26069), .B1(n29956), .B2(
        n31074), .Y(n26008) );
  OAI22xp33_ASAP7_75t_SL U29422 ( .A1(n31059), .A2(n26069), .B1(n31058), .B2(
        n29956), .Y(n25982) );
  OAI22xp33_ASAP7_75t_SL U29423 ( .A1(n31155), .A2(n26127), .B1(n31154), .B2(
        n26126), .Y(n26119) );
  OAI22xp33_ASAP7_75t_SL U29424 ( .A1(n31155), .A2(n26069), .B1(n29956), .B2(
        n31154), .Y(n26040) );
  OAI22xp33_ASAP7_75t_SL U29425 ( .A1(n31143), .A2(n26069), .B1(n29956), .B2(
        n31142), .Y(n26033) );
  NAND2xp5_ASAP7_75t_SL U29426 ( .A(n24967), .B(n26736), .Y(n27241) );
  INVxp33_ASAP7_75t_SL U29427 ( .A(n30009), .Y(n27064) );
  AOI21xp33_ASAP7_75t_SL U29428 ( .A1(n24631), .A2(n26168), .B(n26164), .Y(
        n26165) );
  AOI21xp33_ASAP7_75t_SL U29429 ( .A1(n26168), .A2(n29150), .B(n23164), .Y(
        n26162) );
  AOI22xp33_ASAP7_75t_SL U29430 ( .A1(u0_0_leon3x0_p0_c0mmu_dcache0_r_NOFLUSH_), .A2(n30995), .B1(it_q[26]), .B2(n24636), .Y(n25617) );
  OAI21xp33_ASAP7_75t_SL U29431 ( .A1(n30645), .A2(n29768), .B(n28465), .Y(
        n28466) );
  OAI21xp33_ASAP7_75t_SL U29432 ( .A1(n29864), .A2(n26522), .B(n26484), .Y(
        n26485) );
  OAI21xp33_ASAP7_75t_SL U29433 ( .A1(n30645), .A2(n29081), .B(n28511), .Y(
        n28512) );
  OAI21xp33_ASAP7_75t_SL U29434 ( .A1(n30645), .A2(n30821), .B(n28530), .Y(
        n28531) );
  NAND2xp33_ASAP7_75t_SL U29435 ( .A(n30874), .B(n31840), .Y(n26627) );
  NAND2xp33_ASAP7_75t_SL U29436 ( .A(apbi[13]), .B(n24633), .Y(n29333) );
  INVxp67_ASAP7_75t_SL U29437 ( .A(mult_x_1196_n2364), .Y(n22473) );
  INVxp33_ASAP7_75t_SL U29438 ( .A(n25627), .Y(n25623) );
  OAI21xp33_ASAP7_75t_SL U29439 ( .A1(n25336), .A2(n32719), .B(n25335), .Y(
        n32985) );
  INVxp67_ASAP7_75t_SL U29440 ( .A(n29583), .Y(n27075) );
  INVx1_ASAP7_75t_SL U29441 ( .A(mult_x_1196_n2185), .Y(mult_x_1196_n953) );
  INVxp33_ASAP7_75t_SL U29442 ( .A(add_x_735_n135), .Y(add_x_735_n133) );
  INVxp33_ASAP7_75t_SL U29443 ( .A(add_x_735_n100), .Y(add_x_735_n102) );
  NAND2xp5_ASAP7_75t_SL U29444 ( .A(n29700), .B(n29699), .Y(n29875) );
  BUFx4f_ASAP7_75t_SL U29445 ( .A(n24039), .Y(n22412) );
  INVxp67_ASAP7_75t_SL U29446 ( .A(mult_x_1196_n2279), .Y(n23148) );
  OAI21xp33_ASAP7_75t_SL U29447 ( .A1(n30149), .A2(n30148), .B(n31954), .Y(
        n30150) );
  OAI21xp33_ASAP7_75t_SL U29448 ( .A1(n1792), .A2(n30141), .B(n30979), .Y(
        n30153) );
  INVxp33_ASAP7_75t_SL U29449 ( .A(n31004), .Y(n30126) );
  OAI21xp33_ASAP7_75t_SL U29450 ( .A1(n2962), .A2(n31312), .B(n32445), .Y(
        n31317) );
  OAI21xp33_ASAP7_75t_SL U29451 ( .A1(add_x_735_n199), .A2(add_x_735_n191), 
        .B(add_x_735_n192), .Y(add_x_735_n190) );
  OAI21xp33_ASAP7_75t_SL U29452 ( .A1(u0_0_leon3x0_p0_c0mmu_dcache0_r_BMEXC_), 
        .A2(n32199), .B(n32198), .Y(n2999) );
  INVxp33_ASAP7_75t_SL U29453 ( .A(n26385), .Y(n26387) );
  AOI22xp33_ASAP7_75t_SL U29454 ( .A1(u0_0_leon3x0_p0_divi[23]), .A2(n27200), 
        .B1(n28830), .B2(n26385), .Y(n26386) );
  INVxp67_ASAP7_75t_SL U29455 ( .A(mult_x_1196_n2360), .Y(n23432) );
  AOI22xp33_ASAP7_75t_SL U29456 ( .A1(dc_q[24]), .A2(n31004), .B1(dt_q[20]), 
        .B2(n29991), .Y(n26513) );
  INVx1_ASAP7_75t_SL U29457 ( .A(n28051), .Y(n28052) );
  INVxp33_ASAP7_75t_SL U29458 ( .A(n28044), .Y(n28048) );
  AOI22xp33_ASAP7_75t_SL U29459 ( .A1(it_q[3]), .A2(n24636), .B1(dc_q[3]), 
        .B2(n31473), .Y(n30880) );
  NAND2xp5_ASAP7_75t_SL U29460 ( .A(n29356), .B(n29357), .Y(n28042) );
  AOI22xp33_ASAP7_75t_SL U29461 ( .A1(dc_q[27]), .A2(n31004), .B1(dt_q[23]), 
        .B2(n24573), .Y(n26346) );
  NAND2xp33_ASAP7_75t_SL U29462 ( .A(apbi[11]), .B(n24633), .Y(n25944) );
  AOI22xp33_ASAP7_75t_SL U29463 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__27_), .A2(n30207), .B1(
        it_q[23]), .B2(n24636), .Y(n26345) );
  AOI22xp5_ASAP7_75t_SL U29464 ( .A1(n27146), .A2(n27145), .B1(n27144), .B2(
        n27154), .Y(n30386) );
  OAI21xp33_ASAP7_75t_SL U29465 ( .A1(n28121), .A2(n32004), .B(n28120), .Y(
        n28130) );
  OAI21xp33_ASAP7_75t_SL U29466 ( .A1(n30446), .A2(n30219), .B(n30218), .Y(
        n30222) );
  NAND2xp33_ASAP7_75t_SL U29467 ( .A(n30614), .B(n30609), .Y(n28998) );
  AOI21xp33_ASAP7_75t_SL U29468 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__5_), 
        .A2(n22378), .B(n26814), .Y(n2796) );
  AOI22xp33_ASAP7_75t_SL U29469 ( .A1(dc_q[26]), .A2(n31004), .B1(dt_q[22]), 
        .B2(n24573), .Y(n26235) );
  NAND2xp5_ASAP7_75t_SL U29470 ( .A(n26774), .B(n26773), .Y(n31431) );
  INVxp33_ASAP7_75t_SL U29471 ( .A(add_x_735_n191), .Y(add_x_735_n290) );
  NAND2xp33_ASAP7_75t_SL U29472 ( .A(n31328), .B(n31840), .Y(n26497) );
  INVxp67_ASAP7_75t_SL U29473 ( .A(mult_x_1196_n2252), .Y(n22971) );
  NAND2xp33_ASAP7_75t_SL U29474 ( .A(n30106), .B(n31840), .Y(n26633) );
  NAND2xp33_ASAP7_75t_SL U29475 ( .A(n28254), .B(n31840), .Y(n26640) );
  NAND2xp33_ASAP7_75t_SL U29476 ( .A(n26646), .B(n31840), .Y(n26643) );
  INVxp33_ASAP7_75t_SL U29477 ( .A(add_x_735_n203), .Y(add_x_735_n201) );
  INVxp67_ASAP7_75t_SL U29478 ( .A(add_x_735_n204), .Y(add_x_735_n202) );
  NAND2xp33_ASAP7_75t_SL U29479 ( .A(n29287), .B(n29383), .Y(n29288) );
  AOI22xp33_ASAP7_75t_SL U29480 ( .A1(dc_q[28]), .A2(n31004), .B1(dt_q[24]), 
        .B2(n24573), .Y(n25444) );
  AOI22xp33_ASAP7_75t_SL U29481 ( .A1(n28272), .A2(n29598), .B1(n22906), .B2(
        n29583), .Y(n26933) );
  NAND2xp33_ASAP7_75t_SL U29482 ( .A(n30833), .B(n24633), .Y(n29943) );
  OAI21xp33_ASAP7_75t_SL U29483 ( .A1(n25393), .A2(n30212), .B(n32074), .Y(
        n25394) );
  AOI21xp33_ASAP7_75t_SL U29484 ( .A1(n29598), .A2(n27027), .B(n26996), .Y(
        n27001) );
  NAND2xp33_ASAP7_75t_SL U29485 ( .A(n23161), .B(n29583), .Y(n26999) );
  INVxp33_ASAP7_75t_SL U29486 ( .A(uart1_scaler_11_), .Y(n28140) );
  INVxp33_ASAP7_75t_SL U29487 ( .A(u0_0_leon3x0_p0_divi[29]), .Y(n29149) );
  AND2x2_ASAP7_75t_SL U29488 ( .A(n24579), .B(u0_0_leon3x0_p0_divi[29]), .Y(
        n29145) );
  AOI22xp33_ASAP7_75t_SL U29489 ( .A1(n29583), .A2(n23365), .B1(n29584), .B2(
        n29585), .Y(n29586) );
  O2A1O1Ixp33_ASAP7_75t_SL U29490 ( .A1(n27196), .A2(n25198), .B(n25116), .C(
        n28850), .Y(n25117) );
  AOI21xp33_ASAP7_75t_SL U29491 ( .A1(n30272), .A2(n28835), .B(n28493), .Y(
        n28494) );
  AOI22xp33_ASAP7_75t_SL U29492 ( .A1(apbi[8]), .A2(n31736), .B1(
        sr1_r_MCFG1__ROMWIDTH__0_), .B2(n31735), .Y(n2916) );
  AOI22xp33_ASAP7_75t_SL U29493 ( .A1(apbi[11]), .A2(n31736), .B1(
        sr1_r_MCFG1__ROMWRITE_), .B2(n31735), .Y(n2917) );
  AOI22xp33_ASAP7_75t_SL U29494 ( .A1(apbi[23]), .A2(n31736), .B1(
        sr1_r_MCFG1__IOWS__3_), .B2(n31735), .Y(n2918) );
  AOI22xp33_ASAP7_75t_SL U29495 ( .A1(apbi[22]), .A2(n31736), .B1(
        sr1_r_MCFG1__IOWS__2_), .B2(n31735), .Y(n2919) );
  AOI22xp33_ASAP7_75t_SL U29496 ( .A1(apbi[21]), .A2(n31736), .B1(
        sr1_r_MCFG1__IOWS__1_), .B2(n31735), .Y(n2920) );
  AOI22xp33_ASAP7_75t_SL U29497 ( .A1(apbi[20]), .A2(n31736), .B1(
        sr1_r_MCFG1__IOWS__0_), .B2(n31735), .Y(n2921) );
  AOI22xp33_ASAP7_75t_SL U29498 ( .A1(apbi[25]), .A2(n31736), .B1(
        sr1_r_MCFG1__BEXCEN_), .B2(n31735), .Y(n2922) );
  OAI22xp33_ASAP7_75t_SL U29499 ( .A1(n25175), .A2(n29592), .B1(n31418), .B2(
        n28941), .Y(n25181) );
  AOI22xp33_ASAP7_75t_SL U29500 ( .A1(apbi[26]), .A2(n31736), .B1(
        sr1_r_MCFG1__BRDYEN_), .B2(n31735), .Y(n2923) );
  AOI22xp33_ASAP7_75t_SL U29501 ( .A1(u0_0_leon3x0_p0_divi[22]), .A2(n27200), 
        .B1(n28830), .B2(n26430), .Y(n26431) );
  OAI21xp33_ASAP7_75t_SL U29502 ( .A1(apbi[1]), .A2(n30030), .B(n26098), .Y(
        n4532) );
  OAI22xp33_ASAP7_75t_SL U29503 ( .A1(n31063), .A2(n29556), .B1(n31062), .B2(
        n29555), .Y(n29525) );
  OAI21xp33_ASAP7_75t_SL U29504 ( .A1(n30800), .A2(n32719), .B(n25261), .Y(
        n32995) );
  OAI22xp33_ASAP7_75t_SL U29505 ( .A1(n31135), .A2(n29556), .B1(n31134), .B2(
        n29555), .Y(n29543) );
  OAI22xp33_ASAP7_75t_SL U29506 ( .A1(n31123), .A2(n29556), .B1(n31122), .B2(
        n29555), .Y(n29540) );
  OAI22xp33_ASAP7_75t_SL U29507 ( .A1(n31067), .A2(n29556), .B1(n31066), .B2(
        n29555), .Y(n29526) );
  OAI21xp33_ASAP7_75t_SL U29508 ( .A1(uart1_r_THOLD__17__6_), .A2(n27922), .B(
        n27585), .Y(n1824) );
  OAI22xp33_ASAP7_75t_SL U29509 ( .A1(n31107), .A2(n29556), .B1(n31106), .B2(
        n29555), .Y(n29536) );
  OAI22xp33_ASAP7_75t_SL U29510 ( .A1(n31099), .A2(n29556), .B1(n31098), .B2(
        n29555), .Y(n29534) );
  OAI21xp33_ASAP7_75t_SL U29511 ( .A1(uart1_r_THOLD__17__7_), .A2(n27922), .B(
        n27544), .Y(n1823) );
  OAI22xp33_ASAP7_75t_SL U29512 ( .A1(n31159), .A2(n29556), .B1(n31158), .B2(
        n29555), .Y(n29549) );
  OAI22xp33_ASAP7_75t_SL U29513 ( .A1(n31075), .A2(n29556), .B1(n31074), .B2(
        n29555), .Y(n29528) );
  OAI21xp33_ASAP7_75t_SL U29514 ( .A1(uart1_r_THOLD__15__0_), .A2(n27979), .B(
        n27978), .Y(n1822) );
  OAI21xp33_ASAP7_75t_SL U29515 ( .A1(uart1_r_THOLD__15__1_), .A2(n27979), .B(
        n27389), .Y(n1821) );
  INVxp67_ASAP7_75t_SL U29516 ( .A(n29218), .Y(n29217) );
  OAI21xp33_ASAP7_75t_SL U29517 ( .A1(uart1_r_THOLD__15__2_), .A2(n27979), .B(
        n27889), .Y(n1820) );
  AOI22xp33_ASAP7_75t_SL U29518 ( .A1(uart1_r_TRADDR__2_), .A2(n27315), .B1(
        n27312), .B2(n27314), .Y(n2240) );
  OAI21xp33_ASAP7_75t_SL U29519 ( .A1(uart1_r_THOLD__15__3_), .A2(n27979), .B(
        n27825), .Y(n1819) );
  NAND2xp33_ASAP7_75t_SL U29520 ( .A(n24694), .B(n27319), .Y(n2242) );
  OAI21xp33_ASAP7_75t_SL U29521 ( .A1(uart1_r_THOLD__15__4_), .A2(n27979), .B(
        n27753), .Y(n1818) );
  OAI21xp33_ASAP7_75t_SL U29522 ( .A1(uart1_r_THOLD__15__5_), .A2(n27979), .B(
        n27689), .Y(n1817) );
  OAI21xp33_ASAP7_75t_SL U29523 ( .A1(uart1_r_THOLD__15__6_), .A2(n27979), .B(
        n27621), .Y(n1816) );
  OAI21xp33_ASAP7_75t_SL U29524 ( .A1(uart1_r_THOLD__15__7_), .A2(n27979), .B(
        n27580), .Y(n1815) );
  AOI21xp33_ASAP7_75t_SL U29525 ( .A1(n29003), .A2(n26534), .B(n30006), .Y(
        n26447) );
  NAND2xp33_ASAP7_75t_SL U29526 ( .A(n24950), .B(n31873), .Y(n24951) );
  OAI21xp33_ASAP7_75t_SL U29527 ( .A1(uart1_r_THOLD__8__0_), .A2(n27933), .B(
        n27932), .Y(n2254) );
  OAI21xp33_ASAP7_75t_SL U29528 ( .A1(uart1_r_THOLD__11__0_), .A2(n27977), .B(
        n27976), .Y(n2257) );
  OAI21xp33_ASAP7_75t_SL U29529 ( .A1(uart1_r_THOLD__12__0_), .A2(n27937), .B(
        n27936), .Y(n2258) );
  OAI21xp33_ASAP7_75t_SL U29530 ( .A1(uart1_r_THOLD__13__0_), .A2(n27931), .B(
        n27930), .Y(n2259) );
  OAI21xp5_ASAP7_75t_SL U29531 ( .A1(n31982), .A2(n29810), .B(n29809), .Y(
        n29818) );
  NAND2xp33_ASAP7_75t_SL U29532 ( .A(n26520), .B(n31840), .Y(n26517) );
  OAI21xp33_ASAP7_75t_SL U29533 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_r_E__CTRL__ANNUL_), .B(n32067), .Y(n3709) );
  OAI21xp33_ASAP7_75t_SL U29534 ( .A1(n30446), .A2(n30282), .B(n30281), .Y(
        n30284) );
  NAND2xp5_ASAP7_75t_SL U29535 ( .A(n28286), .B(n28288), .Y(n28287) );
  NAND2xp5_ASAP7_75t_SL U29536 ( .A(n26534), .B(n30619), .Y(n27246) );
  OAI21xp33_ASAP7_75t_SL U29537 ( .A1(n30645), .A2(n27172), .B(n27131), .Y(
        n27132) );
  OAI21xp33_ASAP7_75t_SL U29538 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__9_), 
        .A2(n30701), .B(n27137), .Y(n2312) );
  OAI21xp33_ASAP7_75t_SL U29539 ( .A1(n30645), .A2(n29932), .B(n28752), .Y(
        n28753) );
  OAI21xp33_ASAP7_75t_SL U29540 ( .A1(n31412), .A2(n30412), .B(n30411), .Y(
        n30415) );
  OAI22xp33_ASAP7_75t_SL U29541 ( .A1(n31151), .A2(n30772), .B1(n31150), .B2(
        n30771), .Y(n30763) );
  OAI22xp33_ASAP7_75t_SL U29542 ( .A1(n31167), .A2(n30772), .B1(n31166), .B2(
        n30771), .Y(n30767) );
  OAI21xp33_ASAP7_75t_SL U29543 ( .A1(uart1_r_THOLD__20__7_), .A2(n27939), .B(
        n27554), .Y(n1839) );
  OAI22xp33_ASAP7_75t_SL U29544 ( .A1(n31131), .A2(n30772), .B1(n31130), .B2(
        n30771), .Y(n30758) );
  OAI22xp33_ASAP7_75t_SL U29545 ( .A1(n31155), .A2(n30772), .B1(n31154), .B2(
        n30771), .Y(n30764) );
  OAI22xp33_ASAP7_75t_SL U29546 ( .A1(n31175), .A2(n30772), .B1(n31174), .B2(
        n30771), .Y(n30769) );
  OAI22xp33_ASAP7_75t_SL U29547 ( .A1(n31179), .A2(n30772), .B1(n31178), .B2(
        n30771), .Y(n30770) );
  OAI22xp33_ASAP7_75t_SL U29548 ( .A1(n31147), .A2(n30772), .B1(n31146), .B2(
        n30771), .Y(n30762) );
  OAI21xp33_ASAP7_75t_SL U29549 ( .A1(uart1_r_THOLD__18__0_), .A2(n27960), .B(
        n27959), .Y(n1838) );
  OAI22xp33_ASAP7_75t_SL U29550 ( .A1(n31091), .A2(n30772), .B1(n31090), .B2(
        n30771), .Y(n30748) );
  OAI22xp33_ASAP7_75t_SL U29551 ( .A1(n31119), .A2(n30772), .B1(n31118), .B2(
        n30771), .Y(n30755) );
  NAND2xp5_ASAP7_75t_SL U29552 ( .A(n31574), .B(n31572), .Y(n32022) );
  OAI22xp33_ASAP7_75t_SL U29553 ( .A1(n31087), .A2(n30772), .B1(n31086), .B2(
        n30771), .Y(n30747) );
  OAI21xp33_ASAP7_75t_SL U29554 ( .A1(uart1_r_THOLD__18__1_), .A2(n27960), .B(
        n27368), .Y(n1837) );
  OAI22xp33_ASAP7_75t_SL U29555 ( .A1(n31095), .A2(n30772), .B1(n31094), .B2(
        n30771), .Y(n30749) );
  OAI22xp33_ASAP7_75t_SL U29556 ( .A1(n31115), .A2(n30772), .B1(n31114), .B2(
        n30771), .Y(n30754) );
  OAI22xp33_ASAP7_75t_SL U29557 ( .A1(n31185), .A2(n30772), .B1(n31183), .B2(
        n30771), .Y(n30773) );
  OAI21xp33_ASAP7_75t_SL U29558 ( .A1(uart1_r_THOLD__18__2_), .A2(n27960), .B(
        n27878), .Y(n1836) );
  OAI22xp33_ASAP7_75t_SL U29559 ( .A1(n31163), .A2(n30772), .B1(n31162), .B2(
        n30771), .Y(n30766) );
  OAI22xp33_ASAP7_75t_SL U29560 ( .A1(n31071), .A2(n30772), .B1(n31070), .B2(
        n30771), .Y(n30743) );
  OAI22xp33_ASAP7_75t_SL U29561 ( .A1(n31143), .A2(n30772), .B1(n31142), .B2(
        n30771), .Y(n30761) );
  OAI22xp33_ASAP7_75t_SL U29562 ( .A1(n31139), .A2(n30772), .B1(n31138), .B2(
        n30771), .Y(n30760) );
  OAI22xp33_ASAP7_75t_SL U29563 ( .A1(n31127), .A2(n30772), .B1(n31126), .B2(
        n30771), .Y(n30757) );
  OAI22xp33_ASAP7_75t_SL U29564 ( .A1(n31079), .A2(n30772), .B1(n31078), .B2(
        n30771), .Y(n30745) );
  OAI21xp33_ASAP7_75t_SL U29565 ( .A1(uart1_r_THOLD__18__3_), .A2(n27960), .B(
        n27814), .Y(n1835) );
  OAI22xp33_ASAP7_75t_SL U29566 ( .A1(n31083), .A2(n30772), .B1(n31082), .B2(
        n30771), .Y(n30746) );
  OAI22xp33_ASAP7_75t_SL U29567 ( .A1(n31063), .A2(n30772), .B1(n31062), .B2(
        n30771), .Y(n30741) );
  OAI21xp33_ASAP7_75t_SL U29568 ( .A1(uart1_r_THOLD__18__4_), .A2(n27960), .B(
        n27742), .Y(n1834) );
  OAI22xp33_ASAP7_75t_SL U29569 ( .A1(n31135), .A2(n30772), .B1(n31134), .B2(
        n30771), .Y(n30759) );
  OAI22xp33_ASAP7_75t_SL U29570 ( .A1(n31123), .A2(n30772), .B1(n31122), .B2(
        n30771), .Y(n30756) );
  AOI21xp33_ASAP7_75t_SL U29571 ( .A1(n32719), .A2(n31602), .B(n4076), .Y(
        n32035) );
  OAI22xp33_ASAP7_75t_SL U29572 ( .A1(n31067), .A2(n30772), .B1(n31066), .B2(
        n30771), .Y(n30742) );
  OAI21xp33_ASAP7_75t_SL U29573 ( .A1(uart1_r_THOLD__18__5_), .A2(n27960), .B(
        n27678), .Y(n1833) );
  OAI22xp33_ASAP7_75t_SL U29574 ( .A1(n31107), .A2(n30772), .B1(n31106), .B2(
        n30771), .Y(n30752) );
  OAI22xp33_ASAP7_75t_SL U29575 ( .A1(n31099), .A2(n30772), .B1(n31098), .B2(
        n30771), .Y(n30750) );
  OAI22xp33_ASAP7_75t_SL U29576 ( .A1(n31159), .A2(n30772), .B1(n31158), .B2(
        n30771), .Y(n30765) );
  OAI22xp33_ASAP7_75t_SL U29577 ( .A1(n31075), .A2(n30772), .B1(n31074), .B2(
        n30771), .Y(n30744) );
  OAI22xp33_ASAP7_75t_SL U29578 ( .A1(n31111), .A2(n28225), .B1(n31110), .B2(
        n28224), .Y(n28206) );
  OAI22xp33_ASAP7_75t_SL U29579 ( .A1(n31171), .A2(n28225), .B1(n31170), .B2(
        n28224), .Y(n28221) );
  OAI22xp33_ASAP7_75t_SL U29580 ( .A1(n31103), .A2(n28225), .B1(n31102), .B2(
        n28224), .Y(n28204) );
  OAI22xp33_ASAP7_75t_SL U29581 ( .A1(n31151), .A2(n28225), .B1(n31150), .B2(
        n28224), .Y(n28216) );
  OAI22xp33_ASAP7_75t_SL U29582 ( .A1(n31167), .A2(n28225), .B1(n31166), .B2(
        n28224), .Y(n28220) );
  OAI22xp33_ASAP7_75t_SL U29583 ( .A1(n31131), .A2(n28225), .B1(n31130), .B2(
        n28224), .Y(n28211) );
  OAI22xp33_ASAP7_75t_SL U29584 ( .A1(n31155), .A2(n28225), .B1(n31154), .B2(
        n28224), .Y(n28217) );
  OAI22xp33_ASAP7_75t_SL U29585 ( .A1(n31175), .A2(n28225), .B1(n31174), .B2(
        n28224), .Y(n28222) );
  OAI21xp33_ASAP7_75t_SL U29586 ( .A1(uart1_r_THOLD__18__6_), .A2(n27960), .B(
        n27610), .Y(n1832) );
  OAI22xp33_ASAP7_75t_SL U29587 ( .A1(n31179), .A2(n28225), .B1(n31178), .B2(
        n28224), .Y(n28223) );
  OAI22xp33_ASAP7_75t_SL U29588 ( .A1(n31147), .A2(n28225), .B1(n31146), .B2(
        n28224), .Y(n28215) );
  OAI22xp33_ASAP7_75t_SL U29589 ( .A1(n31091), .A2(n28225), .B1(n31090), .B2(
        n28224), .Y(n28201) );
  OAI21xp33_ASAP7_75t_SL U29590 ( .A1(uart1_r_THOLD__18__7_), .A2(n27960), .B(
        n27569), .Y(n1831) );
  OAI22xp33_ASAP7_75t_SL U29591 ( .A1(n31119), .A2(n28225), .B1(n31118), .B2(
        n28224), .Y(n28208) );
  OAI22xp33_ASAP7_75t_SL U29592 ( .A1(n31087), .A2(n28225), .B1(n31086), .B2(
        n28224), .Y(n28200) );
  OAI22xp33_ASAP7_75t_SL U29593 ( .A1(n31095), .A2(n28225), .B1(n31094), .B2(
        n28224), .Y(n28202) );
  OAI21xp33_ASAP7_75t_SL U29594 ( .A1(uart1_r_THOLD__17__0_), .A2(n27922), .B(
        n27921), .Y(n1830) );
  OAI22xp33_ASAP7_75t_SL U29595 ( .A1(n31103), .A2(n30772), .B1(n31102), .B2(
        n30771), .Y(n30751) );
  OAI22xp33_ASAP7_75t_SL U29596 ( .A1(n31115), .A2(n28225), .B1(n31114), .B2(
        n28224), .Y(n28207) );
  OAI22xp33_ASAP7_75t_SL U29597 ( .A1(n31185), .A2(n28225), .B1(n31183), .B2(
        n28224), .Y(n28226) );
  OAI22xp33_ASAP7_75t_SL U29598 ( .A1(n31163), .A2(n28225), .B1(n31162), .B2(
        n28224), .Y(n28219) );
  OAI22xp33_ASAP7_75t_SL U29599 ( .A1(n31071), .A2(n28225), .B1(n31070), .B2(
        n28224), .Y(n28196) );
  OAI21xp33_ASAP7_75t_SL U29600 ( .A1(uart1_r_THOLD__17__1_), .A2(n27922), .B(
        n27345), .Y(n1829) );
  INVxp67_ASAP7_75t_SL U29601 ( .A(n27303), .Y(n27304) );
  OAI22xp33_ASAP7_75t_SL U29602 ( .A1(n31143), .A2(n28225), .B1(n31142), .B2(
        n28224), .Y(n28214) );
  OAI22xp33_ASAP7_75t_SL U29603 ( .A1(n31139), .A2(n28225), .B1(n31138), .B2(
        n28224), .Y(n28213) );
  OAI22xp33_ASAP7_75t_SL U29604 ( .A1(n31127), .A2(n28225), .B1(n31126), .B2(
        n28224), .Y(n28210) );
  OAI22xp33_ASAP7_75t_SL U29605 ( .A1(n31079), .A2(n28225), .B1(n31078), .B2(
        n28224), .Y(n28198) );
  OAI22xp33_ASAP7_75t_SL U29606 ( .A1(n31083), .A2(n28225), .B1(n31082), .B2(
        n28224), .Y(n28199) );
  OAI22xp33_ASAP7_75t_SL U29607 ( .A1(n31063), .A2(n28225), .B1(n31062), .B2(
        n28224), .Y(n28194) );
  NAND2xp5_ASAP7_75t_SL U29608 ( .A(n23195), .B(n23194), .Y(n23193) );
  OAI22xp33_ASAP7_75t_SL U29609 ( .A1(n31135), .A2(n28225), .B1(n31134), .B2(
        n28224), .Y(n28212) );
  OAI22xp33_ASAP7_75t_SL U29610 ( .A1(n31123), .A2(n28225), .B1(n31122), .B2(
        n28224), .Y(n28209) );
  OAI22xp33_ASAP7_75t_SL U29611 ( .A1(n31067), .A2(n28225), .B1(n31066), .B2(
        n28224), .Y(n28195) );
  OAI22xp33_ASAP7_75t_SL U29612 ( .A1(n31107), .A2(n28225), .B1(n31106), .B2(
        n28224), .Y(n28205) );
  OAI22xp33_ASAP7_75t_SL U29613 ( .A1(n31099), .A2(n28225), .B1(n31098), .B2(
        n28224), .Y(n28203) );
  OAI22xp33_ASAP7_75t_SL U29614 ( .A1(n31159), .A2(n28225), .B1(n31158), .B2(
        n28224), .Y(n28218) );
  OAI22xp33_ASAP7_75t_SL U29615 ( .A1(n31075), .A2(n28225), .B1(n31074), .B2(
        n28224), .Y(n28197) );
  OAI21xp33_ASAP7_75t_SL U29616 ( .A1(uart1_r_THOLD__17__2_), .A2(n27922), .B(
        n27853), .Y(n1828) );
  OAI22xp33_ASAP7_75t_SL U29617 ( .A1(n31111), .A2(n29556), .B1(n31110), .B2(
        n29555), .Y(n29537) );
  OAI22xp33_ASAP7_75t_SL U29618 ( .A1(n31171), .A2(n29556), .B1(n31170), .B2(
        n29555), .Y(n29552) );
  OAI21xp33_ASAP7_75t_SL U29619 ( .A1(uart1_r_THOLD__17__3_), .A2(n27922), .B(
        n27799), .Y(n1827) );
  OAI22xp33_ASAP7_75t_SL U29620 ( .A1(n31103), .A2(n29556), .B1(n31102), .B2(
        n29555), .Y(n29535) );
  OAI22xp33_ASAP7_75t_SL U29621 ( .A1(n31151), .A2(n29556), .B1(n31150), .B2(
        n29555), .Y(n29547) );
  OAI22xp33_ASAP7_75t_SL U29622 ( .A1(n31167), .A2(n29556), .B1(n31166), .B2(
        n29555), .Y(n29551) );
  OAI21xp33_ASAP7_75t_SL U29623 ( .A1(uart1_r_THOLD__17__4_), .A2(n27922), .B(
        n27717), .Y(n1826) );
  OAI22xp33_ASAP7_75t_SL U29624 ( .A1(n31131), .A2(n29556), .B1(n31130), .B2(
        n29555), .Y(n29542) );
  OAI22xp33_ASAP7_75t_SL U29625 ( .A1(n31155), .A2(n29556), .B1(n31154), .B2(
        n29555), .Y(n29548) );
  OAI22xp33_ASAP7_75t_SL U29626 ( .A1(n31175), .A2(n29556), .B1(n31174), .B2(
        n29555), .Y(n29553) );
  OAI22xp33_ASAP7_75t_SL U29627 ( .A1(n31179), .A2(n29556), .B1(n31178), .B2(
        n29555), .Y(n29554) );
  AOI21xp33_ASAP7_75t_SL U29628 ( .A1(n31242), .A2(uart1_r_RHOLD__0__5_), .B(
        n30108), .Y(n30109) );
  OAI22xp33_ASAP7_75t_SL U29629 ( .A1(n31147), .A2(n29556), .B1(n31146), .B2(
        n29555), .Y(n29546) );
  OAI22xp33_ASAP7_75t_SL U29630 ( .A1(n31091), .A2(n29556), .B1(n31090), .B2(
        n29555), .Y(n29532) );
  OAI22xp33_ASAP7_75t_SL U29631 ( .A1(n31119), .A2(n29556), .B1(n31118), .B2(
        n29555), .Y(n29539) );
  OAI22xp33_ASAP7_75t_SL U29632 ( .A1(n31087), .A2(n29556), .B1(n31086), .B2(
        n29555), .Y(n29531) );
  OAI22xp33_ASAP7_75t_SL U29633 ( .A1(n31095), .A2(n29556), .B1(n31094), .B2(
        n29555), .Y(n29533) );
  OAI22xp33_ASAP7_75t_SL U29634 ( .A1(n31115), .A2(n29556), .B1(n31114), .B2(
        n29555), .Y(n29538) );
  OAI22xp33_ASAP7_75t_SL U29635 ( .A1(n31185), .A2(n29556), .B1(n31183), .B2(
        n29555), .Y(n29557) );
  OAI22xp33_ASAP7_75t_SL U29636 ( .A1(n31163), .A2(n29556), .B1(n31162), .B2(
        n29555), .Y(n29550) );
  OAI22xp33_ASAP7_75t_SL U29637 ( .A1(n31071), .A2(n29556), .B1(n31070), .B2(
        n29555), .Y(n29527) );
  OAI22xp33_ASAP7_75t_SL U29638 ( .A1(n31143), .A2(n29556), .B1(n31142), .B2(
        n29555), .Y(n29545) );
  OAI22xp33_ASAP7_75t_SL U29639 ( .A1(n31139), .A2(n29556), .B1(n31138), .B2(
        n29555), .Y(n29544) );
  OAI21xp33_ASAP7_75t_SL U29640 ( .A1(uart1_r_THOLD__17__5_), .A2(n27922), .B(
        n27663), .Y(n1825) );
  OAI22xp33_ASAP7_75t_SL U29641 ( .A1(n31127), .A2(n29556), .B1(n31126), .B2(
        n29555), .Y(n29541) );
  OAI22xp33_ASAP7_75t_SL U29642 ( .A1(n31079), .A2(n29556), .B1(n31078), .B2(
        n29555), .Y(n29529) );
  OAI22xp33_ASAP7_75t_SL U29643 ( .A1(n31083), .A2(n29556), .B1(n31082), .B2(
        n29555), .Y(n29530) );
  OAI22xp33_ASAP7_75t_SL U29644 ( .A1(n31087), .A2(n26069), .B1(n29956), .B2(
        n31086), .Y(n26017) );
  OAI21xp33_ASAP7_75t_SL U29645 ( .A1(n31340), .A2(n29693), .B(n26323), .Y(
        n26324) );
  NAND2xp5_ASAP7_75t_SL U29646 ( .A(n29131), .B(n29130), .Y(n29171) );
  OAI22xp33_ASAP7_75t_SL U29647 ( .A1(n31087), .A2(n26127), .B1(n31086), .B2(
        n26126), .Y(n26104) );
  OAI22xp33_ASAP7_75t_SL U29648 ( .A1(n31103), .A2(n26127), .B1(n31102), .B2(
        n26126), .Y(n26107) );
  OAI22xp33_ASAP7_75t_SL U29649 ( .A1(n31119), .A2(n26069), .B1(n29956), .B2(
        n31118), .Y(n26025) );
  NAND2xp33_ASAP7_75t_SL U29650 ( .A(n28405), .B(n27155), .Y(n26227) );
  AOI21xp33_ASAP7_75t_SL U29651 ( .A1(n29564), .A2(n26534), .B(n30006), .Y(
        n26230) );
  INVxp67_ASAP7_75t_SL U29652 ( .A(n29255), .Y(n29256) );
  NAND2xp33_ASAP7_75t_SL U29653 ( .A(n32005), .B(n31840), .Y(n26543) );
  OAI21xp5_ASAP7_75t_SL U29654 ( .A1(n29146), .A2(n26304), .B(n26303), .Y(
        n26305) );
  OAI22xp33_ASAP7_75t_SL U29655 ( .A1(n31103), .A2(n26069), .B1(n29956), .B2(
        n31102), .Y(n26020) );
  AOI21xp5_ASAP7_75t_SL U29656 ( .A1(n29564), .A2(n29563), .B(n29562), .Y(
        n32302) );
  INVxp33_ASAP7_75t_SL U29657 ( .A(add_x_735_n230), .Y(add_x_735_n232) );
  NAND2xp5_ASAP7_75t_SL U29658 ( .A(n2883), .B(uart1_scaler_11_), .Y(n28142)
         );
  OAI22xp33_ASAP7_75t_SL U29659 ( .A1(n29166), .A2(n30654), .B1(n29132), .B2(
        n30653), .Y(n29133) );
  OAI22xp33_ASAP7_75t_SL U29660 ( .A1(n31119), .A2(n26127), .B1(n31118), .B2(
        n26126), .Y(n26110) );
  OAI22xp33_ASAP7_75t_SL U29661 ( .A1(n31151), .A2(n26127), .B1(n31150), .B2(
        n26126), .Y(n26118) );
  OAI22xp33_ASAP7_75t_SL U29662 ( .A1(n31091), .A2(n26069), .B1(n29956), .B2(
        n31090), .Y(n26018) );
  OAI22xp33_ASAP7_75t_SL U29663 ( .A1(n31091), .A2(n26127), .B1(n31090), .B2(
        n26126), .Y(n26105) );
  OAI22xp33_ASAP7_75t_SL U29664 ( .A1(n31151), .A2(n26069), .B1(n29956), .B2(
        n31150), .Y(n26037) );
  NAND2xp33_ASAP7_75t_SL U29665 ( .A(n30151), .B(n31840), .Y(n26620) );
  OAI22xp33_ASAP7_75t_SL U29666 ( .A1(n31167), .A2(n26127), .B1(n31166), .B2(
        n26126), .Y(n26122) );
  NAND2xp5_ASAP7_75t_SL U29667 ( .A(it_q[11]), .B(n24636), .Y(n25041) );
  OAI22xp33_ASAP7_75t_SL U29668 ( .A1(n31147), .A2(n26069), .B1(n29956), .B2(
        n31146), .Y(n26034) );
  NAND2xp33_ASAP7_75t_SL U29669 ( .A(n28540), .B(n29598), .Y(n25830) );
  OAI22xp33_ASAP7_75t_SL U29670 ( .A1(n31167), .A2(n26069), .B1(n29956), .B2(
        n31166), .Y(n26050) );
  AOI22xp33_ASAP7_75t_SL U29671 ( .A1(apbi[19]), .A2(n31736), .B1(
        sr1_r_MCFG1__IOEN_), .B2(n31735), .Y(n2350) );
  OAI22xp33_ASAP7_75t_SL U29672 ( .A1(n31147), .A2(n26127), .B1(n31146), .B2(
        n26126), .Y(n26117) );
  OAI22xp33_ASAP7_75t_SL U29673 ( .A1(n31131), .A2(n26127), .B1(n31130), .B2(
        n26126), .Y(n26113) );
  OAI22xp33_ASAP7_75t_SL U29674 ( .A1(n31131), .A2(n26069), .B1(n29956), .B2(
        n31130), .Y(n26028) );
  OAI22xp33_ASAP7_75t_SL U29675 ( .A1(n31179), .A2(n26069), .B1(n29956), .B2(
        n31178), .Y(n26063) );
  OAI22xp33_ASAP7_75t_SL U29676 ( .A1(n31179), .A2(n26127), .B1(n31178), .B2(
        n26126), .Y(n26125) );
  OAI22xp33_ASAP7_75t_SL U29677 ( .A1(n31175), .A2(n26069), .B1(n29956), .B2(
        n31174), .Y(n26057) );
  INVxp33_ASAP7_75t_SL U29678 ( .A(n26262), .Y(n26264) );
  OAI22xp33_ASAP7_75t_SL U29679 ( .A1(n31175), .A2(n26127), .B1(n31174), .B2(
        n26126), .Y(n26124) );
  AOI22xp33_ASAP7_75t_SL U29680 ( .A1(dc_q[19]), .A2(n31004), .B1(dt_q[15]), 
        .B2(n24573), .Y(n25744) );
  NAND2xp33_ASAP7_75t_SL U29681 ( .A(n29430), .B(n29383), .Y(n29248) );
  AOI22xp33_ASAP7_75t_SL U29682 ( .A1(u0_0_leon3x0_p0_divi[5]), .A2(n27200), 
        .B1(n28830), .B2(n26262), .Y(n26263) );
  INVx1_ASAP7_75t_SL U29683 ( .A(n32004), .Y(n30993) );
  NAND2xp33_ASAP7_75t_SL U29684 ( .A(n28405), .B(n28668), .Y(n26887) );
  OAI22xp33_ASAP7_75t_SL U29685 ( .A1(n31163), .A2(n26069), .B1(n29956), .B2(
        n31162), .Y(n26047) );
  NAND2xp5_ASAP7_75t_SL U29686 ( .A(n28879), .B(n28878), .Y(n29505) );
  INVx1_ASAP7_75t_SL U29687 ( .A(n30562), .Y(n22413) );
  AOI21xp33_ASAP7_75t_SL U29688 ( .A1(n31950), .A2(uart1_r_EXTCLKEN_), .B(
        n29751), .Y(n29755) );
  OAI22xp33_ASAP7_75t_SL U29689 ( .A1(n31163), .A2(n26127), .B1(n31162), .B2(
        n26126), .Y(n26121) );
  AOI22xp33_ASAP7_75t_SL U29690 ( .A1(dc_q[23]), .A2(n31004), .B1(dt_q[19]), 
        .B2(n29991), .Y(n25063) );
  OAI22xp33_ASAP7_75t_SL U29691 ( .A1(n31185), .A2(n26069), .B1(n29956), .B2(
        n31183), .Y(n26070) );
  OAI22xp33_ASAP7_75t_SL U29692 ( .A1(n31071), .A2(n26127), .B1(n31070), .B2(
        n26126), .Y(n26100) );
  OAI22xp33_ASAP7_75t_SL U29693 ( .A1(n31111), .A2(n26127), .B1(n31110), .B2(
        n26126), .Y(n26109) );
  OAI22xp33_ASAP7_75t_SL U29694 ( .A1(n31185), .A2(n26127), .B1(n31183), .B2(
        n26126), .Y(n26128) );
  AOI22xp33_ASAP7_75t_SL U29695 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__23_), .A2(n30207), .B1(
        it_q[19]), .B2(n24636), .Y(n25062) );
  NAND2xp33_ASAP7_75t_SL U29696 ( .A(n30549), .B(n31840), .Y(n26594) );
  OAI22xp33_ASAP7_75t_SL U29697 ( .A1(n31171), .A2(n26127), .B1(n31170), .B2(
        n26126), .Y(n26123) );
  OAI21xp33_ASAP7_75t_SL U29698 ( .A1(n31017), .A2(n32719), .B(n25263), .Y(
        n32994) );
  OAI22xp33_ASAP7_75t_SL U29699 ( .A1(n31095), .A2(n26069), .B1(n29956), .B2(
        n31094), .Y(n26019) );
  OAI22xp33_ASAP7_75t_SL U29700 ( .A1(n31071), .A2(n26069), .B1(n29956), .B2(
        n31070), .Y(n26007) );
  NAND2xp33_ASAP7_75t_SL U29701 ( .A(n30552), .B(n29383), .Y(n25637) );
  OAI21xp33_ASAP7_75t_SL U29702 ( .A1(n30446), .A2(n30402), .B(n30401), .Y(
        n30405) );
  OAI22xp33_ASAP7_75t_SL U29703 ( .A1(n28095), .A2(n28094), .B1(n30783), .B2(
        n28093), .Y(n28098) );
  OAI22xp33_ASAP7_75t_SL U29704 ( .A1(n31111), .A2(n26069), .B1(n29956), .B2(
        n31110), .Y(n26024) );
  AOI21xp33_ASAP7_75t_SL U29705 ( .A1(n31240), .A2(n28084), .B(n28083), .Y(
        n28092) );
  OAI22xp33_ASAP7_75t_SL U29706 ( .A1(n31143), .A2(n26127), .B1(n31142), .B2(
        n26126), .Y(n26116) );
  OAI22xp33_ASAP7_75t_SL U29707 ( .A1(n31095), .A2(n26127), .B1(n31094), .B2(
        n26126), .Y(n26106) );
  OAI22xp33_ASAP7_75t_SL U29708 ( .A1(n31171), .A2(n26069), .B1(n29956), .B2(
        n31170), .Y(n26056) );
  NAND2xp33_ASAP7_75t_SL U29709 ( .A(apbi[2]), .B(n30738), .Y(n4670) );
  AOI22xp33_ASAP7_75t_SL U29710 ( .A1(n29060), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PC__2_), .B1(u0_0_leon3x0_p0_ici[30]), 
        .B2(n29059), .Y(n28908) );
  OAI21xp33_ASAP7_75t_SL U29711 ( .A1(n24690), .A2(n26147), .B(n26141), .Y(
        n26293) );
  AOI22xp33_ASAP7_75t_SL U29712 ( .A1(dc_q[16]), .A2(n31473), .B1(dt_q[12]), 
        .B2(n24573), .Y(n26668) );
  NAND2xp33_ASAP7_75t_SL U29713 ( .A(n28108), .B(n27979), .Y(n27978) );
  OAI21xp33_ASAP7_75t_SL U29714 ( .A1(n28941), .A2(n26429), .B(n26417), .Y(
        n26418) );
  INVxp33_ASAP7_75t_SL U29715 ( .A(add_x_735_n199), .Y(add_x_735_n197) );
  NAND2xp33_ASAP7_75t_SL U29716 ( .A(n29568), .B(n27967), .Y(n27882) );
  NAND2xp5_ASAP7_75t_SL U29717 ( .A(n32194), .B(n30198), .Y(n30205) );
  NAND2xp33_ASAP7_75t_SL U29718 ( .A(n29510), .B(n27922), .Y(n27799) );
  NAND2xp33_ASAP7_75t_SL U29719 ( .A(n27493), .B(n27935), .Y(n27323) );
  NAND2xp33_ASAP7_75t_SL U29720 ( .A(n28108), .B(n27922), .Y(n27921) );
  NAND2xp33_ASAP7_75t_SL U29721 ( .A(n29568), .B(n27979), .Y(n27889) );
  NAND2xp33_ASAP7_75t_SL U29722 ( .A(n30780), .B(n27979), .Y(n27753) );
  NAND2xp33_ASAP7_75t_SL U29723 ( .A(n30833), .B(n27935), .Y(n27552) );
  NAND2xp33_ASAP7_75t_SL U29724 ( .A(n30833), .B(n27979), .Y(n27580) );
  NAND2xp33_ASAP7_75t_SL U29725 ( .A(n31197), .B(n27922), .Y(n27585) );
  INVxp33_ASAP7_75t_SL U29726 ( .A(n32008), .Y(n30141) );
  NAND2xp33_ASAP7_75t_SL U29727 ( .A(n27493), .B(n27979), .Y(n27389) );
  NAND2xp33_ASAP7_75t_SL U29728 ( .A(n31197), .B(n27935), .Y(n27593) );
  OAI21xp33_ASAP7_75t_SL U29729 ( .A1(apbi[3]), .A2(n27965), .B(n27817), .Y(
        n1811) );
  NAND2xp33_ASAP7_75t_SL U29730 ( .A(n30780), .B(n27935), .Y(n27725) );
  INVxp33_ASAP7_75t_SL U29731 ( .A(n29883), .Y(n30707) );
  INVx1_ASAP7_75t_SL U29732 ( .A(n28924), .Y(n28618) );
  NAND2xp33_ASAP7_75t_SL U29733 ( .A(n29568), .B(n27922), .Y(n27853) );
  NAND2xp33_ASAP7_75t_SL U29734 ( .A(n29510), .B(n27979), .Y(n27825) );
  NAND2xp33_ASAP7_75t_SL U29735 ( .A(n28108), .B(n27967), .Y(n27966) );
  NAND2xp33_ASAP7_75t_SL U29736 ( .A(n30780), .B(n27922), .Y(n27717) );
  NAND2xp33_ASAP7_75t_SL U29737 ( .A(n27136), .B(n30701), .Y(n27137) );
  NAND2xp33_ASAP7_75t_SL U29738 ( .A(n27493), .B(n27922), .Y(n27345) );
  NAND2xp33_ASAP7_75t_SL U29739 ( .A(n30833), .B(n27922), .Y(n27544) );
  NAND2xp5_ASAP7_75t_SL U29740 ( .A(n28847), .B(n28844), .Y(n27094) );
  OAI21xp33_ASAP7_75t_SL U29741 ( .A1(n31645), .A2(n31973), .B(n31644), .Y(
        n31648) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U29742 ( .A1(n31438), .A2(n29195), .B(n29184), 
        .C(n29202), .Y(n29188) );
  NAND2xp33_ASAP7_75t_SL U29743 ( .A(n30073), .B(n27935), .Y(n27651) );
  NAND2xp33_ASAP7_75t_SL U29744 ( .A(n29510), .B(n27935), .Y(n27787) );
  NAND2xp5_ASAP7_75t_SL U29745 ( .A(n32673), .B(n32674), .Y(n32682) );
  OAI21xp33_ASAP7_75t_SL U29746 ( .A1(apbi[2]), .A2(n27965), .B(n27881), .Y(
        n1812) );
  OAI22xp33_ASAP7_75t_SL U29747 ( .A1(apbi[6]), .A2(n29515), .B1(
        timer0_r_RELOAD__6_), .B2(n29514), .Y(n1727) );
  NAND2xp33_ASAP7_75t_SL U29748 ( .A(n27493), .B(n27967), .Y(n27374) );
  OAI21xp33_ASAP7_75t_SL U29749 ( .A1(apbi[0]), .A2(n27965), .B(n27964), .Y(
        n1814) );
  NAND2xp33_ASAP7_75t_SL U29750 ( .A(n30073), .B(n27922), .Y(n27663) );
  OAI21xp33_ASAP7_75t_SL U29751 ( .A1(apbi[1]), .A2(n27965), .B(n27372), .Y(
        n1813) );
  NAND2xp33_ASAP7_75t_SL U29752 ( .A(n31197), .B(n27979), .Y(n27621) );
  NAND2xp33_ASAP7_75t_SL U29753 ( .A(n30073), .B(n27979), .Y(n27689) );
  NAND2xp33_ASAP7_75t_SL U29754 ( .A(n29568), .B(n27935), .Y(n27861) );
  INVx1_ASAP7_75t_SL U29755 ( .A(n28762), .Y(n28914) );
  NAND2xp33_ASAP7_75t_SL U29756 ( .A(dc_q[7]), .B(n31473), .Y(n25055) );
  INVxp67_ASAP7_75t_SL U29757 ( .A(n25142), .Y(n25110) );
  OAI22xp33_ASAP7_75t_SL U29758 ( .A1(n30812), .A2(n28257), .B1(n23229), .B2(
        u0_0_leon3x0_p0_iu_r_A__RSEL2__2_), .Y(n2820) );
  INVx1_ASAP7_75t_SL U29759 ( .A(n26155), .Y(n25785) );
  NAND2xp33_ASAP7_75t_SL U29760 ( .A(n30780), .B(n27920), .Y(n27716) );
  INVxp67_ASAP7_75t_SL U29761 ( .A(n29300), .Y(n29295) );
  NAND2xp33_ASAP7_75t_SL U29762 ( .A(n28108), .B(n27939), .Y(n27938) );
  OAI21xp33_ASAP7_75t_SL U29763 ( .A1(n27196), .A2(n22392), .B(n25622), .Y(
        n25627) );
  NAND2xp33_ASAP7_75t_SL U29764 ( .A(n24694), .B(n25995), .Y(n25993) );
  NAND2xp33_ASAP7_75t_SL U29765 ( .A(n27493), .B(n27939), .Y(n27326) );
  INVxp67_ASAP7_75t_SL U29766 ( .A(mult_x_1196_n2786), .Y(n23410) );
  INVx1_ASAP7_75t_SL U29767 ( .A(n29745), .Y(n29325) );
  NAND2xp33_ASAP7_75t_SL U29768 ( .A(n29568), .B(n27939), .Y(n27863) );
  INVxp67_ASAP7_75t_SL U29769 ( .A(n29267), .Y(n29262) );
  NAND2xp33_ASAP7_75t_SL U29770 ( .A(n29510), .B(n27920), .Y(n27798) );
  NAND2xp33_ASAP7_75t_SL U29771 ( .A(n30073), .B(n27920), .Y(n27662) );
  NAND2xp33_ASAP7_75t_SL U29772 ( .A(n29568), .B(n27920), .Y(n27852) );
  NAND2xp33_ASAP7_75t_SL U29773 ( .A(n29510), .B(n27939), .Y(n27789) );
  NAND2xp33_ASAP7_75t_SL U29774 ( .A(n27493), .B(n27920), .Y(n27344) );
  NAND2xp33_ASAP7_75t_SL U29775 ( .A(n28108), .B(n27920), .Y(n27919) );
  OAI21xp33_ASAP7_75t_SL U29776 ( .A1(n31503), .A2(n31973), .B(n31502), .Y(
        n31506) );
  NAND2xp33_ASAP7_75t_SL U29777 ( .A(n30780), .B(n27939), .Y(n27727) );
  NAND2xp33_ASAP7_75t_SL U29778 ( .A(n30833), .B(n27962), .Y(n27570) );
  NOR2xp33_ASAP7_75t_SL U29779 ( .A(n23651), .B(n22392), .Y(n25168) );
  NAND2xp33_ASAP7_75t_SL U29780 ( .A(n30073), .B(n27939), .Y(n27653) );
  INVx1_ASAP7_75t_SL U29781 ( .A(n29605), .Y(n28502) );
  OAI22xp33_ASAP7_75t_SL U29782 ( .A1(irqctrl0_r_IPEND__9_), .A2(n29745), .B1(
        irqctrl0_r_IFORCE__0__9_), .B2(n29254), .Y(n29255) );
  OAI21xp33_ASAP7_75t_SL U29783 ( .A1(irqctrl0_r_IFORCE__0__15_), .A2(n29394), 
        .B(n24694), .Y(n29396) );
  NAND2xp33_ASAP7_75t_SL U29784 ( .A(n31197), .B(n27939), .Y(n27595) );
  AOI21xp33_ASAP7_75t_SL U29785 ( .A1(n27197), .A2(n29150), .B(n27196), .Y(
        n27199) );
  NAND2xp33_ASAP7_75t_SL U29786 ( .A(n30780), .B(n27973), .Y(n27750) );
  NOR2x1_ASAP7_75t_SL U29787 ( .A(n25023), .B(n25044), .Y(n31004) );
  AOI21xp33_ASAP7_75t_SL U29788 ( .A1(n24575), .A2(n23160), .B(n28987), .Y(
        n28983) );
  NAND2xp33_ASAP7_75t_SL U29789 ( .A(n29510), .B(n27973), .Y(n27822) );
  AOI21xp33_ASAP7_75t_SL U29790 ( .A1(n31424), .A2(n31398), .B(n31397), .Y(
        n31399) );
  NAND2xp33_ASAP7_75t_SL U29791 ( .A(n29568), .B(n27973), .Y(n27886) );
  NAND2xp33_ASAP7_75t_SL U29792 ( .A(n27493), .B(n27973), .Y(n27382) );
  NAND2xp33_ASAP7_75t_SL U29793 ( .A(n30073), .B(n27973), .Y(n27686) );
  AOI22xp33_ASAP7_75t_SL U29794 ( .A1(dc_q[15]), .A2(n31473), .B1(dt_q[11]), 
        .B2(n24573), .Y(n25047) );
  NAND2xp33_ASAP7_75t_SL U29795 ( .A(n28108), .B(n27973), .Y(n27972) );
  NAND2xp33_ASAP7_75t_SL U29796 ( .A(n25901), .B(n28620), .Y(n26918) );
  INVx1_ASAP7_75t_SL U29797 ( .A(n23396), .Y(n23164) );
  OAI21xp33_ASAP7_75t_SL U29798 ( .A1(n31327), .A2(n31973), .B(n31326), .Y(
        n31330) );
  NAND2xp33_ASAP7_75t_SL U29799 ( .A(n31197), .B(n27973), .Y(n27618) );
  NAND2xp33_ASAP7_75t_SL U29800 ( .A(n30833), .B(n27920), .Y(n27543) );
  OAI21xp33_ASAP7_75t_SL U29801 ( .A1(n31372), .A2(n31973), .B(n31371), .Y(
        n31375) );
  NAND2xp33_ASAP7_75t_SL U29802 ( .A(n28132), .B(n28620), .Y(n25425) );
  AOI22xp33_ASAP7_75t_SL U29803 ( .A1(u0_0_leon3x0_p0_iu_r_E__CTRL__WREG_), 
        .A2(n24648), .B1(u0_0_leon3x0_p0_iu_r_A__CTRL__WREG_), .B2(n32065), 
        .Y(n2712) );
  AOI21xp33_ASAP7_75t_SL U29804 ( .A1(n24578), .A2(n23002), .B(n26155), .Y(
        n25787) );
  NAND2xp33_ASAP7_75t_SL U29805 ( .A(n31197), .B(n27920), .Y(n27584) );
  AOI21xp33_ASAP7_75t_SL U29806 ( .A1(n29787), .A2(n31398), .B(n29786), .Y(
        n29788) );
  OR2x2_ASAP7_75t_SL U29807 ( .A(n22578), .B(n24469), .Y(n23642) );
  NAND2xp5_ASAP7_75t_SL U29808 ( .A(n24478), .B(n25625), .Y(n29584) );
  NAND2xp33_ASAP7_75t_SL U29809 ( .A(n30833), .B(n27973), .Y(n27577) );
  NAND2xp33_ASAP7_75t_SL U29810 ( .A(n29568), .B(n27960), .Y(n27878) );
  OR2x2_ASAP7_75t_SL U29811 ( .A(n22578), .B(n22392), .Y(n23641) );
  NAND2xp33_ASAP7_75t_SL U29812 ( .A(n29510), .B(n27960), .Y(n27814) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U29813 ( .A1(n31027), .A2(n31848), .B(n31323), 
        .C(n31026), .Y(n31028) );
  OAI22xp33_ASAP7_75t_SL U29814 ( .A1(n28193), .A2(n28192), .B1(
        uart1_r_RWADDR__0_), .B2(n28191), .Y(n2453) );
  NAND2xp33_ASAP7_75t_SL U29815 ( .A(n27493), .B(n27962), .Y(n27370) );
  NAND2xp33_ASAP7_75t_SL U29816 ( .A(n31868), .B(n28601), .Y(n28606) );
  OA21x2_ASAP7_75t_SRAM U29817 ( .A1(n26001), .A2(n28192), .B(n26021), .Y(
        n25973) );
  NAND2xp33_ASAP7_75t_SL U29818 ( .A(n30780), .B(n27960), .Y(n27742) );
  NAND2xp5_ASAP7_75t_SL U29819 ( .A(n27425), .B(n27424), .Y(n27915) );
  AOI22xp33_ASAP7_75t_SL U29820 ( .A1(n25974), .A2(n28191), .B1(
        uart1_r_RWADDR__2_), .B2(n28192), .Y(n2455) );
  OAI21xp33_ASAP7_75t_SL U29821 ( .A1(n32027), .A2(n31452), .B(n32243), .Y(
        n25518) );
  OAI22xp33_ASAP7_75t_SL U29822 ( .A1(sr1_r_MCFG1__ROMRWS__2_), .A2(n29522), 
        .B1(apbi[2]), .B2(n30779), .Y(n2899) );
  NAND2xp33_ASAP7_75t_SL U29823 ( .A(n28108), .B(n27962), .Y(n27961) );
  NAND2xp33_ASAP7_75t_SL U29824 ( .A(n30833), .B(n27967), .Y(n27573) );
  INVxp33_ASAP7_75t_SL U29825 ( .A(n28191), .Y(n25976) );
  OAI21xp33_ASAP7_75t_SL U29826 ( .A1(apbi[7]), .A2(n27965), .B(n27572), .Y(
        n1807) );
  NAND2xp33_ASAP7_75t_SL U29827 ( .A(n30073), .B(n27960), .Y(n27678) );
  AOI22xp33_ASAP7_75t_SL U29828 ( .A1(apbi[1]), .A2(n29524), .B1(
        sr1_r_MCFG2__RAMRWS__1_), .B2(n29523), .Y(n2907) );
  AOI22xp33_ASAP7_75t_SL U29829 ( .A1(apbi[0]), .A2(n29524), .B1(
        sr1_r_MCFG2__RAMRWS__0_), .B2(n29523), .Y(n2908) );
  AOI22xp33_ASAP7_75t_SL U29830 ( .A1(apbi[3]), .A2(n29524), .B1(
        sr1_r_MCFG2__RAMWWS__1_), .B2(n29523), .Y(n2909) );
  OAI21xp33_ASAP7_75t_SL U29831 ( .A1(apbi[6]), .A2(n27965), .B(n27613), .Y(
        n1808) );
  NAND2xp33_ASAP7_75t_SL U29832 ( .A(n31197), .B(n27967), .Y(n27614) );
  AOI22xp33_ASAP7_75t_SL U29833 ( .A1(apbi[2]), .A2(n29524), .B1(
        sr1_r_MCFG2__RAMWWS__0_), .B2(n29523), .Y(n2910) );
  NAND2xp33_ASAP7_75t_SL U29834 ( .A(n30073), .B(n27967), .Y(n27682) );
  NAND2xp33_ASAP7_75t_SL U29835 ( .A(n31197), .B(n27960), .Y(n27610) );
  AOI21xp33_ASAP7_75t_SL U29836 ( .A1(n26682), .A2(n29150), .B(n23666), .Y(
        n26684) );
  AOI22xp5_ASAP7_75t_SL U29837 ( .A1(n27895), .A2(n27849), .B1(n27848), .B2(
        n27847), .Y(n28249) );
  NAND2xp33_ASAP7_75t_SL U29838 ( .A(n30780), .B(n27967), .Y(n27746) );
  OAI22xp33_ASAP7_75t_SL U29839 ( .A1(apbi[3]), .A2(n29515), .B1(
        timer0_r_RELOAD__3_), .B2(n29514), .Y(n1740) );
  NAND2xp33_ASAP7_75t_SL U29840 ( .A(n29510), .B(n27967), .Y(n27818) );
  OAI21xp33_ASAP7_75t_SL U29841 ( .A1(apbi[5]), .A2(n27965), .B(n27681), .Y(
        n1809) );
  OAI21xp33_ASAP7_75t_SL U29842 ( .A1(apbi[4]), .A2(n27965), .B(n27745), .Y(
        n1810) );
  NAND2xp33_ASAP7_75t_SL U29843 ( .A(n30833), .B(n27960), .Y(n27569) );
  INVx1_ASAP7_75t_SL U29844 ( .A(n30779), .Y(n31736) );
  OAI21xp33_ASAP7_75t_SL U29845 ( .A1(n29748), .A2(n31973), .B(n29747), .Y(
        n29757) );
  NAND2xp33_ASAP7_75t_SL U29846 ( .A(n31197), .B(n27962), .Y(n27611) );
  NAND2xp33_ASAP7_75t_SL U29847 ( .A(n29750), .B(n29749), .Y(n29751) );
  AOI21xp33_ASAP7_75t_SL U29848 ( .A1(n28403), .A2(n29796), .B(n26226), .Y(
        n26228) );
  NAND2xp33_ASAP7_75t_SL U29849 ( .A(n30073), .B(n27962), .Y(n27679) );
  NAND2xp33_ASAP7_75t_SL U29850 ( .A(n29752), .B(n32008), .Y(n29753) );
  INVxp67_ASAP7_75t_SL U29851 ( .A(n28243), .Y(n28238) );
  INVx1_ASAP7_75t_SL U29852 ( .A(n28403), .Y(n26522) );
  NAND2xp33_ASAP7_75t_SL U29853 ( .A(n30833), .B(n27939), .Y(n27554) );
  AOI21xp33_ASAP7_75t_SL U29854 ( .A1(uart1_r_BRATE__0_), .A2(n28056), .B(
        n28178), .Y(n2873) );
  NOR2xp33_ASAP7_75t_SL U29855 ( .A(n23980), .B(mult_x_1196_n3255), .Y(n23663)
         );
  INVxp67_ASAP7_75t_SL U29856 ( .A(n29245), .Y(n29240) );
  NAND2xp33_ASAP7_75t_SL U29857 ( .A(n30780), .B(n27962), .Y(n27743) );
  AOI21xp33_ASAP7_75t_SL U29858 ( .A1(u0_0_leon3x0_p0_divi[24]), .A2(n24579), 
        .B(n28433), .Y(n28434) );
  NAND2xp33_ASAP7_75t_SL U29859 ( .A(n28108), .B(n27960), .Y(n27959) );
  AOI21xp33_ASAP7_75t_SL U29860 ( .A1(n29846), .A2(n31868), .B(n28651), .Y(
        n28652) );
  NAND2xp33_ASAP7_75t_SL U29861 ( .A(n29510), .B(n27962), .Y(n27815) );
  NAND2xp33_ASAP7_75t_SL U29862 ( .A(n29568), .B(n27962), .Y(n27879) );
  OAI22xp33_ASAP7_75t_SL U29863 ( .A1(apbi[2]), .A2(n29515), .B1(
        timer0_r_RELOAD__2_), .B2(n29514), .Y(n1750) );
  NAND2xp33_ASAP7_75t_SL U29864 ( .A(n27493), .B(n27960), .Y(n27368) );
  OAI21xp33_ASAP7_75t_SL U29865 ( .A1(n31974), .A2(n31973), .B(n31972), .Y(
        n31977) );
  NAND2xp33_ASAP7_75t_SL U29866 ( .A(n31197), .B(n27929), .Y(n27590) );
  NAND2xp33_ASAP7_75t_SL U29867 ( .A(n31197), .B(n27948), .Y(n27602) );
  NAND2xp33_ASAP7_75t_SL U29868 ( .A(n31197), .B(n27977), .Y(n27620) );
  OAI21xp33_ASAP7_75t_SL U29869 ( .A1(n31851), .A2(n31973), .B(n31850), .Y(
        n31854) );
  NAND2xp33_ASAP7_75t_SL U29870 ( .A(n31197), .B(n27937), .Y(n27594) );
  NAND2xp33_ASAP7_75t_SL U29871 ( .A(n31197), .B(n27931), .Y(n27591) );
  NAND2xp33_ASAP7_75t_SL U29872 ( .A(n31197), .B(n27951), .Y(n27604) );
  NAND2xp33_ASAP7_75t_SL U29873 ( .A(n31197), .B(n27946), .Y(n27600) );
  OAI22xp33_ASAP7_75t_SL U29874 ( .A1(apbi[5]), .A2(n29515), .B1(
        timer0_r_RELOAD__5_), .B2(n29514), .Y(n1639) );
  NAND2xp33_ASAP7_75t_SL U29875 ( .A(n31197), .B(n27968), .Y(n27615) );
  NAND2xp33_ASAP7_75t_SL U29876 ( .A(n31197), .B(n27926), .Y(n27588) );
  AOI21xp33_ASAP7_75t_SL U29877 ( .A1(n28806), .A2(n31398), .B(n26288), .Y(
        n26289) );
  NAND2xp33_ASAP7_75t_SL U29878 ( .A(n31197), .B(n27952), .Y(n27605) );
  AOI21xp33_ASAP7_75t_SL U29879 ( .A1(uart1_r_BREAKIRQEN_), .A2(n31950), .B(
        n29853), .Y(n29855) );
  NAND2xp33_ASAP7_75t_SL U29880 ( .A(n31197), .B(n27947), .Y(n27601) );
  OAI22xp33_ASAP7_75t_SL U29881 ( .A1(apbi[4]), .A2(n29515), .B1(
        timer0_r_RELOAD__4_), .B2(n29514), .Y(n1629) );
  NAND2xp33_ASAP7_75t_SL U29882 ( .A(n31197), .B(n27950), .Y(n27603) );
  OAI21xp33_ASAP7_75t_SL U29883 ( .A1(apbi[5]), .A2(n27942), .B(n27655), .Y(
        n1935) );
  OAI22xp33_ASAP7_75t_SL U29884 ( .A1(apbi[0]), .A2(n29515), .B1(
        timer0_r_RELOAD__0_), .B2(n29514), .Y(n4370) );
  OAI21xp33_ASAP7_75t_SL U29885 ( .A1(apbi[5]), .A2(n27925), .B(n27665), .Y(
        n1936) );
  INVxp33_ASAP7_75t_SL U29886 ( .A(n31242), .Y(n28094) );
  OAI22xp33_ASAP7_75t_SL U29887 ( .A1(apbi[7]), .A2(n29515), .B1(
        timer0_r_RELOAD__7_), .B2(n29514), .Y(n1625) );
  INVx1_ASAP7_75t_SL U29888 ( .A(mult_x_1196_n855), .Y(mult_x_1196_n856) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U29889 ( .A1(n28082), .A2(n28081), .B(n31238), 
        .C(n28080), .Y(n28083) );
  OAI21xp33_ASAP7_75t_SL U29890 ( .A1(apbi[5]), .A2(n27955), .B(n27675), .Y(
        n1937) );
  OAI21xp33_ASAP7_75t_SL U29891 ( .A1(apbi[5]), .A2(n27971), .B(n27685), .Y(
        n1938) );
  INVxp33_ASAP7_75t_SL U29892 ( .A(add_x_735_n250), .Y(add_x_735_n299) );
  AOI21xp33_ASAP7_75t_SL U29893 ( .A1(u0_0_leon3x0_p0_divi[17]), .A2(n24580), 
        .B(n25824), .Y(n25825) );
  OAI21xp33_ASAP7_75t_SL U29894 ( .A1(apbi[5]), .A2(n27945), .B(n27657), .Y(
        n1939) );
  AOI21xp33_ASAP7_75t_SL U29895 ( .A1(u0_0_leon3x0_p0_divi[18]), .A2(n24579), 
        .B(n25775), .Y(n25776) );
  OAI21xp33_ASAP7_75t_SL U29896 ( .A1(apbi[5]), .A2(n27918), .B(n27661), .Y(
        n1940) );
  INVxp33_ASAP7_75t_SL U29897 ( .A(add_x_735_n236), .Y(add_x_735_n296) );
  OAI21xp33_ASAP7_75t_SL U29898 ( .A1(apbi[5]), .A2(n27958), .B(n27677), .Y(
        n1941) );
  NAND2xp33_ASAP7_75t_SL U29899 ( .A(n32066), .B(n32065), .Y(n32067) );
  AOI22xp33_ASAP7_75t_SL U29900 ( .A1(u0_0_leon3x0_p0_iu_r_E__CTRL__WICC_), 
        .A2(n24649), .B1(u0_0_leon3x0_p0_iu_r_A__CTRL__WICC_), .B2(n32065), 
        .Y(n3715) );
  INVxp33_ASAP7_75t_SL U29901 ( .A(n18895), .Y(add_x_735_n240) );
  NAND2xp5_ASAP7_75t_SL U29902 ( .A(n30653), .B(n30701), .Y(n30654) );
  NAND2xp33_ASAP7_75t_SL U29903 ( .A(n30833), .B(n27951), .Y(n27563) );
  INVx1_ASAP7_75t_SL U29904 ( .A(mult_x_1196_n3059), .Y(n22459) );
  NAND2xp33_ASAP7_75t_SL U29905 ( .A(n30833), .B(n27946), .Y(n27559) );
  NAND2xp33_ASAP7_75t_SL U29906 ( .A(n30833), .B(n27968), .Y(n27574) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U29907 ( .A1(n24997), .A2(n25230), .B(n31946), 
        .C(n24996), .Y(n3308) );
  INVx1_ASAP7_75t_SL U29908 ( .A(n30030), .Y(n30738) );
  AOI22xp33_ASAP7_75t_SL U29909 ( .A1(n28846), .A2(u0_0_leon3x0_p0_muli[41]), 
        .B1(n28845), .B2(n28844), .Y(n28976) );
  OAI22xp33_ASAP7_75t_SL U29910 ( .A1(n23651), .A2(n28843), .B1(n22493), .B2(
        n26294), .Y(n26277) );
  INVxp67_ASAP7_75t_SL U29911 ( .A(n26295), .Y(n26296) );
  NAND2xp33_ASAP7_75t_SL U29912 ( .A(n30833), .B(n27926), .Y(n27547) );
  INVxp33_ASAP7_75t_SL U29913 ( .A(add_x_735_n144), .Y(add_x_735_n285) );
  INVx1_ASAP7_75t_SL U29914 ( .A(n26469), .Y(n31841) );
  NAND2xp5_ASAP7_75t_SL U29915 ( .A(n28933), .B(n28932), .Y(n30451) );
  NAND2xp33_ASAP7_75t_SL U29916 ( .A(n30833), .B(n27952), .Y(n27564) );
  NAND2xp33_ASAP7_75t_SL U29917 ( .A(n30694), .B(n30701), .Y(n30695) );
  NAND2xp33_ASAP7_75t_SL U29918 ( .A(n30697), .B(n30701), .Y(n30698) );
  NAND2xp33_ASAP7_75t_SL U29919 ( .A(n30833), .B(n27947), .Y(n27560) );
  NAND2xp33_ASAP7_75t_SL U29920 ( .A(n30833), .B(n27950), .Y(n27562) );
  AOI21xp33_ASAP7_75t_SL U29921 ( .A1(u0_0_leon3x0_p0_divi[10]), .A2(n28680), 
        .B(n28679), .Y(n28681) );
  OR2x2_ASAP7_75t_SL U29922 ( .A(n23651), .B(n30008), .Y(n23650) );
  OAI21xp33_ASAP7_75t_SL U29923 ( .A1(apbi[6]), .A2(n27942), .B(n27597), .Y(
        n1915) );
  NAND2xp33_ASAP7_75t_SL U29924 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_STPEND_), 
        .B(n31452), .Y(n32024) );
  NAND2xp5_ASAP7_75t_SL U29925 ( .A(n25409), .B(n30203), .Y(n25401) );
  OAI21xp33_ASAP7_75t_SL U29926 ( .A1(apbi[6]), .A2(n27925), .B(n27587), .Y(
        n1916) );
  NAND2xp33_ASAP7_75t_SL U29927 ( .A(n31398), .B(n29846), .Y(n29836) );
  NAND2xp33_ASAP7_75t_SL U29928 ( .A(n30987), .B(n32008), .Y(n30988) );
  OAI21xp33_ASAP7_75t_SL U29929 ( .A1(apbi[6]), .A2(n27955), .B(n27607), .Y(
        n1917) );
  OAI21xp33_ASAP7_75t_SL U29930 ( .A1(apbi[6]), .A2(n27971), .B(n27617), .Y(
        n1918) );
  OAI21xp33_ASAP7_75t_SL U29931 ( .A1(apbi[6]), .A2(n27945), .B(n27599), .Y(
        n1919) );
  OAI21xp33_ASAP7_75t_SL U29932 ( .A1(apbi[6]), .A2(n27918), .B(n27583), .Y(
        n1920) );
  OAI21xp33_ASAP7_75t_SL U29933 ( .A1(n30700), .A2(n28727), .B(n28726), .Y(
        n28728) );
  AOI22xp33_ASAP7_75t_SL U29934 ( .A1(n28981), .A2(n28844), .B1(n28847), .B2(
        n28978), .Y(n26257) );
  OAI21xp33_ASAP7_75t_SL U29935 ( .A1(apbi[6]), .A2(n27958), .B(n27609), .Y(
        n1921) );
  INVx1_ASAP7_75t_SL U29936 ( .A(n32512), .Y(n32458) );
  NAND2xp33_ASAP7_75t_SL U29937 ( .A(n31197), .B(n27933), .Y(n27592) );
  INVxp67_ASAP7_75t_SL U29938 ( .A(mult_x_1196_n3174), .Y(n22801) );
  NAND2xp33_ASAP7_75t_SL U29939 ( .A(n29568), .B(n27933), .Y(n27860) );
  NAND2xp33_ASAP7_75t_SL U29940 ( .A(n31398), .B(n29623), .Y(n29687) );
  INVxp67_ASAP7_75t_SL U29941 ( .A(n24779), .Y(n24781) );
  NAND2xp33_ASAP7_75t_SL U29942 ( .A(n30073), .B(n27946), .Y(n27658) );
  OAI21xp33_ASAP7_75t_SL U29943 ( .A1(apbi[2]), .A2(n27958), .B(n27877), .Y(
        n2001) );
  NOR2xp33_ASAP7_75t_SL U29944 ( .A(n23980), .B(mult_x_1196_n3270), .Y(n23259)
         );
  OAI22xp33_ASAP7_75t_SL U29945 ( .A1(n30549), .A2(n31243), .B1(n2322), .B2(
        n31953), .Y(n30554) );
  OAI21xp33_ASAP7_75t_SL U29946 ( .A1(apbi[2]), .A2(n27918), .B(n27851), .Y(
        n2000) );
  OAI21xp33_ASAP7_75t_SL U29947 ( .A1(apbi[2]), .A2(n27945), .B(n27867), .Y(
        n1999) );
  NAND2xp33_ASAP7_75t_SL U29948 ( .A(n30073), .B(n27968), .Y(n27683) );
  OAI21xp33_ASAP7_75t_SL U29949 ( .A1(apbi[2]), .A2(n27971), .B(n27885), .Y(
        n1998) );
  OAI21xp33_ASAP7_75t_SL U29950 ( .A1(apbi[2]), .A2(n27955), .B(n27875), .Y(
        n1997) );
  OAI21xp33_ASAP7_75t_SL U29951 ( .A1(apbi[2]), .A2(n27925), .B(n27855), .Y(
        n1996) );
  NAND2xp33_ASAP7_75t_SL U29952 ( .A(n30073), .B(n27926), .Y(n27666) );
  OAI21xp33_ASAP7_75t_SL U29953 ( .A1(apbi[2]), .A2(n27942), .B(n27865), .Y(
        n1995) );
  NAND2xp33_ASAP7_75t_SL U29954 ( .A(n29510), .B(n27950), .Y(n27807) );
  NAND2xp33_ASAP7_75t_SL U29955 ( .A(n29510), .B(n27947), .Y(n27795) );
  NAND2xp33_ASAP7_75t_SL U29956 ( .A(n29510), .B(n27952), .Y(n27809) );
  NAND2xp33_ASAP7_75t_SL U29957 ( .A(n29510), .B(n27926), .Y(n27802) );
  NAND2xp33_ASAP7_75t_SL U29958 ( .A(n29510), .B(n27968), .Y(n27819) );
  NAND2xp33_ASAP7_75t_SL U29959 ( .A(n29510), .B(n27946), .Y(n27794) );
  NAND2xp33_ASAP7_75t_SL U29960 ( .A(n32197), .B(n31897), .Y(n31603) );
  NAND2xp33_ASAP7_75t_SL U29961 ( .A(n29510), .B(n27951), .Y(n27808) );
  BUFx6f_ASAP7_75t_SL U29962 ( .A(n24003), .Y(n22756) );
  NAND2xp33_ASAP7_75t_SL U29963 ( .A(n29510), .B(n27931), .Y(n27805) );
  NAND2xp33_ASAP7_75t_SL U29964 ( .A(n29510), .B(n27937), .Y(n27788) );
  INVxp33_ASAP7_75t_SL U29965 ( .A(add_x_735_n212), .Y(add_x_735_n293) );
  NAND2xp33_ASAP7_75t_SL U29966 ( .A(n29510), .B(n27977), .Y(n27824) );
  NAND2xp33_ASAP7_75t_SL U29967 ( .A(n29510), .B(n27948), .Y(n27806) );
  NAND2xp33_ASAP7_75t_SL U29968 ( .A(n29510), .B(n27929), .Y(n27804) );
  NAND2xp33_ASAP7_75t_SL U29969 ( .A(n29510), .B(n27933), .Y(n27786) );
  OAI21xp33_ASAP7_75t_SL U29970 ( .A1(apbi[3]), .A2(n27958), .B(n27813), .Y(
        n1981) );
  NAND2xp33_ASAP7_75t_SL U29971 ( .A(n30073), .B(n27952), .Y(n27673) );
  OAI21xp33_ASAP7_75t_SL U29972 ( .A1(apbi[3]), .A2(n27918), .B(n27797), .Y(
        n1980) );
  NAND2xp33_ASAP7_75t_SL U29973 ( .A(n30073), .B(n27947), .Y(n27659) );
  OAI21xp33_ASAP7_75t_SL U29974 ( .A1(apbi[3]), .A2(n27945), .B(n27793), .Y(
        n1979) );
  NAND2xp33_ASAP7_75t_SL U29975 ( .A(n29568), .B(n27929), .Y(n27858) );
  OAI21xp33_ASAP7_75t_SL U29976 ( .A1(apbi[3]), .A2(n27971), .B(n27821), .Y(
        n1978) );
  OAI21xp33_ASAP7_75t_SL U29977 ( .A1(apbi[3]), .A2(n27955), .B(n27811), .Y(
        n1977) );
  OAI21xp33_ASAP7_75t_SL U29978 ( .A1(apbi[3]), .A2(n27925), .B(n27801), .Y(
        n1976) );
  OAI21xp33_ASAP7_75t_SL U29979 ( .A1(apbi[3]), .A2(n27942), .B(n27791), .Y(
        n1975) );
  NAND2xp33_ASAP7_75t_SL U29980 ( .A(n30780), .B(n27950), .Y(n27735) );
  NAND2xp33_ASAP7_75t_SL U29981 ( .A(n30780), .B(n27947), .Y(n27733) );
  NAND2xp33_ASAP7_75t_SL U29982 ( .A(n30780), .B(n27952), .Y(n27737) );
  NAND2xp33_ASAP7_75t_SL U29983 ( .A(n30780), .B(n27926), .Y(n27720) );
  NAND2xp5_ASAP7_75t_SL U29984 ( .A(uart1_r_RCNT__1_), .B(n27506), .Y(n27505)
         );
  NAND2xp33_ASAP7_75t_SL U29985 ( .A(n30780), .B(n27968), .Y(n27747) );
  INVxp67_ASAP7_75t_SL U29986 ( .A(n27507), .Y(n27500) );
  INVxp67_ASAP7_75t_SL U29987 ( .A(mult_x_1196_n3157), .Y(n22454) );
  NAND2xp33_ASAP7_75t_SL U29988 ( .A(n30780), .B(n27946), .Y(n27732) );
  NAND2xp33_ASAP7_75t_SL U29989 ( .A(n30780), .B(n27951), .Y(n27736) );
  NAND2xp33_ASAP7_75t_SL U29990 ( .A(n30073), .B(n27950), .Y(n27671) );
  NAND2xp33_ASAP7_75t_SL U29991 ( .A(n30780), .B(n27931), .Y(n27723) );
  NAND2xp33_ASAP7_75t_SL U29992 ( .A(n30780), .B(n27937), .Y(n27726) );
  INVxp67_ASAP7_75t_SL U29993 ( .A(mult_x_1196_n3235), .Y(n24172) );
  NAND2xp33_ASAP7_75t_SL U29994 ( .A(n30780), .B(n27977), .Y(n27752) );
  OAI21xp33_ASAP7_75t_SL U29995 ( .A1(apbi[4]), .A2(n27942), .B(n27729), .Y(
        n1955) );
  NAND2xp33_ASAP7_75t_SL U29996 ( .A(n30780), .B(n27948), .Y(n27734) );
  NAND2xp33_ASAP7_75t_SL U29997 ( .A(n30780), .B(n27929), .Y(n27722) );
  INVxp33_ASAP7_75t_SL U29998 ( .A(n27506), .Y(n27497) );
  NAND2xp33_ASAP7_75t_SL U29999 ( .A(n30780), .B(n27933), .Y(n27724) );
  OAI21xp33_ASAP7_75t_SL U30000 ( .A1(apbi[4]), .A2(n27925), .B(n27719), .Y(
        n1956) );
  OAI21xp33_ASAP7_75t_SL U30001 ( .A1(apbi[4]), .A2(n27958), .B(n27741), .Y(
        n1961) );
  INVx3_ASAP7_75t_SL U30002 ( .A(n23443), .Y(n24008) );
  OAI21xp33_ASAP7_75t_SL U30003 ( .A1(apbi[4]), .A2(n27918), .B(n27715), .Y(
        n1960) );
  OAI21xp33_ASAP7_75t_SL U30004 ( .A1(apbi[4]), .A2(n27945), .B(n27731), .Y(
        n1959) );
  OAI21xp33_ASAP7_75t_SL U30005 ( .A1(apbi[4]), .A2(n27955), .B(n27739), .Y(
        n1957) );
  OAI21xp33_ASAP7_75t_SL U30006 ( .A1(apbi[4]), .A2(n27971), .B(n27749), .Y(
        n1958) );
  INVxp67_ASAP7_75t_SL U30007 ( .A(mult_x_1196_n3160), .Y(n22508) );
  NAND2xp5_ASAP7_75t_SL U30008 ( .A(n30922), .B(n30921), .Y(n30926) );
  NAND2xp33_ASAP7_75t_SL U30009 ( .A(n30073), .B(n27933), .Y(n27650) );
  NAND2xp33_ASAP7_75t_SL U30010 ( .A(n30073), .B(n27929), .Y(n27668) );
  NAND2xp33_ASAP7_75t_SL U30011 ( .A(n30073), .B(n27948), .Y(n27670) );
  NAND2xp33_ASAP7_75t_SL U30012 ( .A(n28108), .B(n27975), .Y(n27974) );
  NAND2xp33_ASAP7_75t_SL U30013 ( .A(n27493), .B(n27975), .Y(n27384) );
  NAND2xp33_ASAP7_75t_SL U30014 ( .A(n29568), .B(n27975), .Y(n27887) );
  INVxp33_ASAP7_75t_SL U30015 ( .A(add_x_735_n220), .Y(add_x_735_n294) );
  NAND2xp33_ASAP7_75t_SL U30016 ( .A(n29510), .B(n27975), .Y(n27823) );
  NAND2xp33_ASAP7_75t_SL U30017 ( .A(n30780), .B(n27975), .Y(n27751) );
  NAND2xp33_ASAP7_75t_SL U30018 ( .A(n30073), .B(n27975), .Y(n27687) );
  OAI21xp33_ASAP7_75t_SL U30019 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_r_X__ICC__1_), .B(n30678), .Y(n3856) );
  NAND2xp33_ASAP7_75t_SL U30020 ( .A(n31197), .B(n27975), .Y(n27619) );
  NAND2xp33_ASAP7_75t_SL U30021 ( .A(n30833), .B(n27975), .Y(n27578) );
  NAND2xp33_ASAP7_75t_SL U30022 ( .A(n28108), .B(n27950), .Y(n27949) );
  NAND2xp33_ASAP7_75t_SL U30023 ( .A(n27493), .B(n27950), .Y(n27358) );
  NAND2xp33_ASAP7_75t_SL U30024 ( .A(n27493), .B(n27947), .Y(n27339) );
  NAND2xp33_ASAP7_75t_SL U30025 ( .A(n27493), .B(n27952), .Y(n27360) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30026 ( .A1(n27316), .A2(uart1_r_TRADDR__0_), 
        .B(uart1_r_TRADDR__1_), .C(n27302), .Y(n27303) );
  NAND2xp33_ASAP7_75t_SL U30027 ( .A(n27493), .B(n27926), .Y(n27349) );
  NAND2xp33_ASAP7_75t_SL U30028 ( .A(n27493), .B(n27968), .Y(n27375) );
  NAND2xp33_ASAP7_75t_SL U30029 ( .A(n27493), .B(n27946), .Y(n27337) );
  NAND2xp33_ASAP7_75t_SL U30030 ( .A(n27493), .B(n27951), .Y(n27359) );
  NAND2xp33_ASAP7_75t_SL U30031 ( .A(n27493), .B(n27931), .Y(n27354) );
  NAND2xp33_ASAP7_75t_SL U30032 ( .A(n27493), .B(n27937), .Y(n27324) );
  NAND2xp33_ASAP7_75t_SL U30033 ( .A(n27493), .B(n27977), .Y(n27386) );
  NAND2xp33_ASAP7_75t_SL U30034 ( .A(n27493), .B(n27948), .Y(n27356) );
  NAND2xp33_ASAP7_75t_SL U30035 ( .A(n27493), .B(n27929), .Y(n27352) );
  NAND2xp33_ASAP7_75t_SL U30036 ( .A(n27493), .B(n27933), .Y(n27311) );
  OAI21xp33_ASAP7_75t_SL U30037 ( .A1(apbi[1]), .A2(n27958), .B(n27367), .Y(
        n2021) );
  OAI21xp33_ASAP7_75t_SL U30038 ( .A1(apbi[1]), .A2(n27918), .B(n27342), .Y(
        n2020) );
  NAND2xp33_ASAP7_75t_SL U30039 ( .A(n30073), .B(n27977), .Y(n27688) );
  OAI21xp33_ASAP7_75t_SL U30040 ( .A1(apbi[1]), .A2(n27945), .B(n27336), .Y(
        n2019) );
  INVx1_ASAP7_75t_SL U30041 ( .A(n24832), .Y(n32173) );
  INVxp67_ASAP7_75t_SL U30042 ( .A(n24748), .Y(n24762) );
  NAND2xp33_ASAP7_75t_SL U30043 ( .A(n30073), .B(n27937), .Y(n27652) );
  OAI21xp33_ASAP7_75t_SL U30044 ( .A1(n26855), .A2(n24748), .B(n25005), .Y(
        n24760) );
  OAI21xp33_ASAP7_75t_SL U30045 ( .A1(apbi[1]), .A2(n27971), .B(n27379), .Y(
        n2018) );
  NAND2xp33_ASAP7_75t_SL U30046 ( .A(n30073), .B(n27931), .Y(n27669) );
  OAI21xp33_ASAP7_75t_SL U30047 ( .A1(apbi[1]), .A2(n27955), .B(n27363), .Y(
        n2017) );
  OAI22xp33_ASAP7_75t_SL U30048 ( .A1(n24935), .A2(n24934), .B1(n23229), .B2(
        u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .Y(n3558) );
  NAND2xp5_ASAP7_75t_SL U30049 ( .A(n24793), .B(n24792), .Y(n24802) );
  OAI21xp33_ASAP7_75t_SL U30050 ( .A1(apbi[1]), .A2(n27925), .B(n27348), .Y(
        n2016) );
  OAI21xp33_ASAP7_75t_SL U30051 ( .A1(apbi[1]), .A2(n27942), .B(n27332), .Y(
        n2015) );
  NAND2xp33_ASAP7_75t_SL U30052 ( .A(n29568), .B(n27950), .Y(n27871) );
  INVxp67_ASAP7_75t_SL U30053 ( .A(mult_x_1196_n3224), .Y(n23359) );
  NAND2xp33_ASAP7_75t_SL U30054 ( .A(n30073), .B(n27951), .Y(n27672) );
  NAND2xp33_ASAP7_75t_SL U30055 ( .A(n29568), .B(n27947), .Y(n27869) );
  NAND2xp33_ASAP7_75t_SL U30056 ( .A(n29568), .B(n27952), .Y(n27873) );
  NAND2xp33_ASAP7_75t_SL U30057 ( .A(n29568), .B(n27926), .Y(n27856) );
  NAND2xp33_ASAP7_75t_SL U30058 ( .A(n29568), .B(n27968), .Y(n27883) );
  NAND2xp33_ASAP7_75t_SL U30059 ( .A(n29568), .B(n27946), .Y(n27868) );
  OAI22xp33_ASAP7_75t_SL U30060 ( .A1(n4742), .A2(n30107), .B1(n30106), .B2(
        n31243), .Y(n30108) );
  AOI21xp33_ASAP7_75t_SL U30061 ( .A1(n28770), .A2(n29150), .B(n23651), .Y(
        n28774) );
  NAND2xp33_ASAP7_75t_SL U30062 ( .A(n29568), .B(n27951), .Y(n27872) );
  NAND2xp33_ASAP7_75t_SL U30063 ( .A(n29568), .B(n27931), .Y(n27859) );
  NAND2xp33_ASAP7_75t_SL U30064 ( .A(n29568), .B(n27937), .Y(n27862) );
  NAND2xp33_ASAP7_75t_SL U30065 ( .A(n29568), .B(n27977), .Y(n27888) );
  AOI21xp33_ASAP7_75t_SL U30066 ( .A1(n29887), .A2(n31398), .B(n29496), .Y(
        n29497) );
  NAND2xp33_ASAP7_75t_SL U30067 ( .A(n29568), .B(n27948), .Y(n27870) );
  OAI21xp33_ASAP7_75t_SL U30068 ( .A1(n24631), .A2(u0_0_leon3x0_p0_divi[20]), 
        .B(n27058), .Y(n29136) );
  AOI21xp33_ASAP7_75t_SL U30069 ( .A1(n32972), .A2(n32982), .B(n32907), .Y(
        n1695) );
  NAND2xp33_ASAP7_75t_SL U30070 ( .A(n30833), .B(n27977), .Y(n27579) );
  OAI21xp33_ASAP7_75t_SL U30071 ( .A1(apbi[7]), .A2(n27942), .B(n27556), .Y(
        n1895) );
  NAND2xp33_ASAP7_75t_SL U30072 ( .A(n29150), .B(n27059), .Y(n27063) );
  NAND2xp33_ASAP7_75t_SL U30073 ( .A(n28108), .B(n27977), .Y(n27976) );
  AOI21xp33_ASAP7_75t_SL U30074 ( .A1(n32972), .A2(n32970), .B(n32902), .Y(
        n1696) );
  OAI21xp33_ASAP7_75t_SL U30075 ( .A1(apbi[0]), .A2(n27918), .B(n27917), .Y(
        n2252) );
  INVxp67_ASAP7_75t_SL U30076 ( .A(add_x_735_n141), .Y(add_x_735_n284) );
  INVxp67_ASAP7_75t_SL U30077 ( .A(add_x_735_n131), .Y(add_x_735_n129) );
  NAND2xp33_ASAP7_75t_SL U30078 ( .A(n30073), .B(n27928), .Y(n27667) );
  NAND2xp33_ASAP7_75t_SL U30079 ( .A(n28108), .B(n27937), .Y(n27936) );
  NAND2xp33_ASAP7_75t_SL U30080 ( .A(n26465), .B(n30030), .Y(n26098) );
  NAND2xp33_ASAP7_75t_SL U30081 ( .A(n30833), .B(n27948), .Y(n27561) );
  AOI21xp33_ASAP7_75t_SL U30082 ( .A1(n32972), .A2(n32962), .B(n32900), .Y(
        n1697) );
  NAND2xp33_ASAP7_75t_SL U30083 ( .A(n31895), .B(n31892), .Y(n31878) );
  OAI21xp33_ASAP7_75t_SL U30084 ( .A1(n30898), .A2(n31973), .B(n30897), .Y(
        n30901) );
  OAI21xp33_ASAP7_75t_SL U30085 ( .A1(apbi[7]), .A2(n27918), .B(n27542), .Y(
        n1900) );
  OAI21xp33_ASAP7_75t_SL U30086 ( .A1(apbi[0]), .A2(n27945), .B(n27944), .Y(
        n2251) );
  NAND2xp33_ASAP7_75t_SL U30087 ( .A(n28108), .B(n27931), .Y(n27930) );
  NAND2xp33_ASAP7_75t_SL U30088 ( .A(n30780), .B(n27928), .Y(n27721) );
  INVxp33_ASAP7_75t_SL U30089 ( .A(add_x_735_n209), .Y(add_x_735_n292) );
  OAI22xp33_ASAP7_75t_SL U30090 ( .A1(apbi[1]), .A2(n29515), .B1(
        timer0_r_RELOAD__1_), .B2(n29514), .Y(n2231) );
  AOI21xp33_ASAP7_75t_SL U30091 ( .A1(n28403), .A2(n27275), .B(n27244), .Y(
        n27245) );
  NAND2xp33_ASAP7_75t_SL U30092 ( .A(n28108), .B(n27928), .Y(n27927) );
  NAND2xp33_ASAP7_75t_SL U30093 ( .A(n30833), .B(n27929), .Y(n27549) );
  NAND2xp33_ASAP7_75t_SL U30094 ( .A(n29510), .B(n27928), .Y(n27803) );
  AOI21xp33_ASAP7_75t_SL U30095 ( .A1(n32972), .A2(n32954), .B(n32898), .Y(
        n1698) );
  OAI21xp33_ASAP7_75t_SL U30096 ( .A1(apbi[0]), .A2(n27971), .B(n27970), .Y(
        n2250) );
  NAND2xp33_ASAP7_75t_SL U30097 ( .A(n24387), .B(n24409), .Y(n24320) );
  INVxp67_ASAP7_75t_SL U30098 ( .A(add_x_735_n54), .Y(add_x_735_n275) );
  NAND2xp33_ASAP7_75t_SL U30099 ( .A(n28125), .B(n32008), .Y(n28126) );
  OAI21xp33_ASAP7_75t_SL U30100 ( .A1(apbi[0]), .A2(n27955), .B(n27954), .Y(
        n2249) );
  AOI21xp33_ASAP7_75t_SL U30101 ( .A1(n32972), .A2(n32946), .B(n32896), .Y(
        n1699) );
  AOI21xp33_ASAP7_75t_SL U30102 ( .A1(u0_0_leon3x0_p0_divi[19]), .A2(n24579), 
        .B(n26990), .Y(n26993) );
  OAI21xp33_ASAP7_75t_SL U30103 ( .A1(apbi[0]), .A2(n27925), .B(n27924), .Y(
        n2248) );
  AOI21xp33_ASAP7_75t_SL U30104 ( .A1(n32972), .A2(n32938), .B(n32894), .Y(
        n1700) );
  OAI21xp33_ASAP7_75t_SL U30105 ( .A1(apbi[7]), .A2(n27958), .B(n27568), .Y(
        n1901) );
  NAND2xp33_ASAP7_75t_SL U30106 ( .A(n30833), .B(n27933), .Y(n27551) );
  NAND2xp33_ASAP7_75t_SL U30107 ( .A(n24694), .B(n27301), .Y(n2238) );
  OAI21xp33_ASAP7_75t_SL U30108 ( .A1(apbi[0]), .A2(n27942), .B(n27941), .Y(
        n2247) );
  NAND2xp33_ASAP7_75t_SL U30109 ( .A(n29568), .B(n27928), .Y(n27857) );
  NAND2xp33_ASAP7_75t_SL U30110 ( .A(n28821), .B(u0_0_leon3x0_p0_divi[30]), 
        .Y(n25131) );
  NAND2xp33_ASAP7_75t_SL U30111 ( .A(n24694), .B(n26083), .Y(n2246) );
  AOI21xp33_ASAP7_75t_SL U30112 ( .A1(n32972), .A2(n32930), .B(n32892), .Y(
        n1701) );
  NAND2xp33_ASAP7_75t_SL U30113 ( .A(n27493), .B(n27928), .Y(n27350) );
  INVxp67_ASAP7_75t_SL U30114 ( .A(add_x_735_n85), .Y(add_x_735_n278) );
  AOI21xp33_ASAP7_75t_SL U30115 ( .A1(n32972), .A2(n32922), .B(n32890), .Y(
        n1702) );
  OAI21xp33_ASAP7_75t_SL U30116 ( .A1(n27316), .A2(n31531), .B(n26080), .Y(
        n29357) );
  AOI21xp33_ASAP7_75t_SL U30117 ( .A1(n28403), .A2(n28529), .B(n26533), .Y(
        n26536) );
  OAI21xp33_ASAP7_75t_SL U30118 ( .A1(apbi[7]), .A2(n27945), .B(n27558), .Y(
        n1899) );
  NAND2xp33_ASAP7_75t_SL U30119 ( .A(n30833), .B(n27928), .Y(n27548) );
  INVxp67_ASAP7_75t_SL U30120 ( .A(n30198), .Y(n30210) );
  INVxp33_ASAP7_75t_SL U30121 ( .A(add_x_735_n153), .Y(add_x_735_n286) );
  INVxp33_ASAP7_75t_SL U30122 ( .A(n31608), .Y(n31312) );
  OAI21xp33_ASAP7_75t_SL U30123 ( .A1(apbi[7]), .A2(n27955), .B(n27566), .Y(
        n1897) );
  NAND2xp33_ASAP7_75t_SL U30124 ( .A(n30833), .B(n27937), .Y(n27553) );
  INVxp67_ASAP7_75t_SL U30125 ( .A(add_x_735_n123), .Y(add_x_735_n282) );
  OAI21xp33_ASAP7_75t_SL U30126 ( .A1(apbi[0]), .A2(n27958), .B(n27957), .Y(
        n2253) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30127 ( .A1(n22919), .A2(n18908), .B(n30662), 
        .C(n30661), .Y(n30665) );
  INVxp33_ASAP7_75t_SL U30128 ( .A(add_x_735_n113), .Y(add_x_735_n111) );
  NAND2xp33_ASAP7_75t_SL U30129 ( .A(n30833), .B(n27931), .Y(n27550) );
  NAND2xp33_ASAP7_75t_SL U30130 ( .A(n28108), .B(n27933), .Y(n27932) );
  NAND2xp33_ASAP7_75t_SL U30131 ( .A(n28108), .B(n27935), .Y(n27934) );
  OAI21xp33_ASAP7_75t_SL U30132 ( .A1(add_x_735_n113), .A2(add_x_735_n105), 
        .B(add_x_735_n106), .Y(add_x_735_n100) );
  OAI21xp33_ASAP7_75t_SL U30133 ( .A1(apbi[7]), .A2(n27971), .B(n27576), .Y(
        n1898) );
  OAI21xp33_ASAP7_75t_SL U30134 ( .A1(n31531), .A2(n31973), .B(n31530), .Y(
        n31534) );
  OAI21xp33_ASAP7_75t_SL U30135 ( .A1(apbi[7]), .A2(n27925), .B(n27546), .Y(
        n1896) );
  NAND2xp33_ASAP7_75t_SL U30136 ( .A(n31197), .B(n27928), .Y(n27589) );
  INVxp67_ASAP7_75t_SL U30137 ( .A(mult_x_1196_n3154), .Y(n22567) );
  NAND2xp33_ASAP7_75t_SL U30138 ( .A(n30502), .B(n24875), .Y(n24892) );
  INVxp33_ASAP7_75t_SL U30139 ( .A(n26080), .Y(n26079) );
  NAND2xp33_ASAP7_75t_SL U30140 ( .A(n27085), .B(n27489), .Y(n26327) );
  INVx1_ASAP7_75t_SL U30141 ( .A(n18610), .Y(n27196) );
  NAND2xp33_ASAP7_75t_SL U30142 ( .A(n27557), .B(n27945), .Y(n27558) );
  NOR2xp33_ASAP7_75t_SRAM U30143 ( .A(n2844), .B(n31953), .Y(n27482) );
  NAND2xp33_ASAP7_75t_SL U30144 ( .A(n27481), .B(n27480), .Y(n27483) );
  INVxp67_ASAP7_75t_SL U30145 ( .A(mult_x_1196_n3095), .Y(n23098) );
  NAND2xp33_ASAP7_75t_SL U30146 ( .A(n29012), .B(n22392), .Y(n25520) );
  NAND2xp33_ASAP7_75t_SL U30147 ( .A(n27880), .B(n27965), .Y(n27881) );
  OAI21xp5_ASAP7_75t_SL U30148 ( .A1(n32847), .A2(n32856), .B(n32846), .Y(
        n32946) );
  NAND2xp33_ASAP7_75t_SL U30149 ( .A(n27816), .B(n27965), .Y(n27817) );
  OAI21xp5_ASAP7_75t_SL U30150 ( .A1(n32845), .A2(n32856), .B(n32844), .Y(
        n32938) );
  NAND2xp33_ASAP7_75t_SL U30151 ( .A(n27744), .B(n27965), .Y(n27745) );
  OAI22xp33_ASAP7_75t_SL U30152 ( .A1(n29274), .A2(n29649), .B1(n29744), .B2(
        n29651), .Y(n29276) );
  NAND2xp33_ASAP7_75t_SL U30153 ( .A(n28805), .B(n22392), .Y(n25625) );
  NAND2xp33_ASAP7_75t_SL U30154 ( .A(n27616), .B(n27971), .Y(n27617) );
  NAND2xp33_ASAP7_75t_SL U30155 ( .A(n27680), .B(n27965), .Y(n27681) );
  NAND2xp33_ASAP7_75t_SL U30156 ( .A(n27541), .B(n27918), .Y(n27542) );
  OAI21xp5_ASAP7_75t_SL U30157 ( .A1(n32843), .A2(n32856), .B(n32842), .Y(
        n32930) );
  NAND2xp33_ASAP7_75t_SL U30158 ( .A(n27612), .B(n27965), .Y(n27613) );
  NAND2xp33_ASAP7_75t_SL U30159 ( .A(n29490), .B(n22392), .Y(n25763) );
  NAND2xp33_ASAP7_75t_SL U30160 ( .A(n27571), .B(n27965), .Y(n27572) );
  INVxp67_ASAP7_75t_SL U30161 ( .A(mult_x_1196_n3089), .Y(n24246) );
  NAND2xp33_ASAP7_75t_SL U30162 ( .A(n27608), .B(n27958), .Y(n27609) );
  NOR2x1_ASAP7_75t_SL U30163 ( .A(n25390), .B(n32071), .Y(n29883) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U30164 ( .A1(n32245), .A2(n32244), .B(n32243), .C(
        n32242), .Y(n32247) );
  NAND2xp33_ASAP7_75t_SL U30165 ( .A(n27676), .B(n27958), .Y(n27677) );
  OAI21xp33_ASAP7_75t_SL U30166 ( .A1(n24527), .A2(dataout[10]), .B(n32931), 
        .Y(n1708) );
  OAI21xp33_ASAP7_75t_SL U30167 ( .A1(n23980), .A2(n29909), .B(n28102), .Y(
        n28100) );
  NAND2xp33_ASAP7_75t_SL U30168 ( .A(n27718), .B(n27925), .Y(n27719) );
  OAI21xp33_ASAP7_75t_SL U30169 ( .A1(n29831), .A2(n26338), .B(n25424), .Y(
        n28620) );
  OAI21xp5_ASAP7_75t_SL U30170 ( .A1(n32857), .A2(n32856), .B(n32855), .Y(
        n32982) );
  OAI22xp33_ASAP7_75t_SL U30171 ( .A1(n29744), .A2(n29652), .B1(n29274), .B2(
        n29650), .Y(n29278) );
  OAI21xp5_ASAP7_75t_SL U30172 ( .A1(n32853), .A2(n32856), .B(n32852), .Y(
        n32970) );
  NAND2xp33_ASAP7_75t_SL U30173 ( .A(n27555), .B(n27942), .Y(n27556) );
  NAND2xp33_ASAP7_75t_SL U30174 ( .A(n27728), .B(n27942), .Y(n27729) );
  NAND2xp33_ASAP7_75t_SL U30175 ( .A(n27582), .B(n27918), .Y(n27583) );
  NAND2xp33_ASAP7_75t_SL U30176 ( .A(n27545), .B(n27925), .Y(n27546) );
  OAI21xp5_ASAP7_75t_SL U30177 ( .A1(n32851), .A2(n32856), .B(n32850), .Y(
        n32962) );
  OAI21xp33_ASAP7_75t_SL U30178 ( .A1(apbi[28]), .A2(n31501), .B(n31500), .Y(
        n1780) );
  NAND2xp33_ASAP7_75t_SL U30179 ( .A(n27565), .B(n27955), .Y(n27566) );
  NAND2xp33_ASAP7_75t_SL U30180 ( .A(n27963), .B(n27965), .Y(n27964) );
  NAND2xp33_ASAP7_75t_SL U30181 ( .A(n27598), .B(n27945), .Y(n27599) );
  NAND2xp33_ASAP7_75t_SL U30182 ( .A(n28586), .B(n22392), .Y(n25622) );
  NAND2xp33_ASAP7_75t_SL U30183 ( .A(n27575), .B(n27971), .Y(n27576) );
  NAND2xp33_ASAP7_75t_SL U30184 ( .A(n27371), .B(n27965), .Y(n27372) );
  OAI21xp5_ASAP7_75t_SL U30185 ( .A1(n32849), .A2(n32856), .B(n32848), .Y(
        n32954) );
  OAI22xp5_ASAP7_75t_SL U30186 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_), 
        .A2(n24770), .B1(n24753), .B2(n24744), .Y(n24832) );
  NAND2xp33_ASAP7_75t_SL U30187 ( .A(uart1_r_OVF_), .B(n31190), .Y(n30775) );
  OAI21xp33_ASAP7_75t_SL U30188 ( .A1(n2924), .A2(n31198), .B(n25943), .Y(
        n17805) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U30189 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), .A2(n24983), .B(n24933), .C(
        n25668), .Y(n24934) );
  NAND2xp33_ASAP7_75t_SL U30190 ( .A(n29275), .B(n29390), .Y(n29254) );
  NAND2xp5_ASAP7_75t_SL U30191 ( .A(n30197), .B(n31458), .Y(n30198) );
  AOI22xp33_ASAP7_75t_SL U30192 ( .A1(uart1_r_TSEMPTYIRQEN_), .A2(n31950), 
        .B1(irqctrl0_r_IPEND__14_), .B2(n31247), .Y(n30551) );
  NAND2xp33_ASAP7_75t_SL U30193 ( .A(n27674), .B(n27955), .Y(n27675) );
  NAND2xp33_ASAP7_75t_SL U30194 ( .A(timer0_r_RELOAD__5_), .B(n31237), .Y(
        n30080) );
  OAI21xp33_ASAP7_75t_SL U30195 ( .A1(apbi[25]), .A2(n29650), .B(n29649), .Y(
        n29253) );
  NAND2xp33_ASAP7_75t_SL U30196 ( .A(uart1_r_FRAME_), .B(n31190), .Y(n31189)
         );
  NAND2xp33_ASAP7_75t_SL U30197 ( .A(n27684), .B(n27971), .Y(n27685) );
  INVxp67_ASAP7_75t_SL U30198 ( .A(mult_x_1196_n2835), .Y(n22716) );
  AOI22xp33_ASAP7_75t_SL U30199 ( .A1(uart1_r_TSEMPTY_), .A2(n31951), .B1(
        timer0_r_RELOAD__1_), .B2(n31237), .Y(n27465) );
  OAI21xp33_ASAP7_75t_SL U30200 ( .A1(apbi[28]), .A2(n29650), .B(n29649), .Y(
        n29242) );
  OAI21xp33_ASAP7_75t_SL U30201 ( .A1(n29561), .A2(n30008), .B(n29560), .Y(
        n29562) );
  NAND2xp33_ASAP7_75t_SL U30202 ( .A(n27895), .B(n27316), .Y(n27302) );
  INVxp67_ASAP7_75t_SL U30203 ( .A(n29313), .Y(n29308) );
  INVxp67_ASAP7_75t_SL U30204 ( .A(n25882), .Y(n25884) );
  NAND2xp33_ASAP7_75t_SL U30205 ( .A(n30465), .B(n22392), .Y(n25495) );
  OAI22xp33_ASAP7_75t_SL U30206 ( .A1(n29312), .A2(n29649), .B1(n31197), .B2(
        n29651), .Y(n29309) );
  NAND2xp33_ASAP7_75t_SL U30207 ( .A(n28714), .B(n22392), .Y(n25496) );
  NAND2xp33_ASAP7_75t_SL U30208 ( .A(uart1_r_PARERR_), .B(n31190), .Y(n30067)
         );
  NAND2xp33_ASAP7_75t_SL U30209 ( .A(n27656), .B(n27945), .Y(n27657) );
  OAI21xp33_ASAP7_75t_SL U30210 ( .A1(n27144), .A2(n30008), .B(n27164), .Y(
        n26611) );
  NAND2xp33_ASAP7_75t_SL U30211 ( .A(n27567), .B(n27958), .Y(n27568) );
  XNOR2xp5_ASAP7_75t_SL U30212 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__1_), .B(
        n30938), .Y(n24834) );
  XNOR2xp5_ASAP7_75t_SL U30213 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__2_), .B(
        n32178), .Y(n24835) );
  NAND2xp33_ASAP7_75t_SL U30214 ( .A(n27606), .B(n27955), .Y(n27607) );
  XNOR2xp5_ASAP7_75t_SL U30215 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__3_), .B(
        n32179), .Y(n24836) );
  NAND2xp33_ASAP7_75t_SL U30216 ( .A(n27660), .B(n27918), .Y(n27661) );
  NAND2xp33_ASAP7_75t_SL U30217 ( .A(n18610), .B(n28131), .Y(n25629) );
  OAI21xp33_ASAP7_75t_SL U30218 ( .A1(n32762), .A2(n30982), .B(n29852), .Y(
        n29853) );
  NAND2xp33_ASAP7_75t_SL U30219 ( .A(n27586), .B(n27925), .Y(n27587) );
  OAI21xp5_ASAP7_75t_SL U30220 ( .A1(n32841), .A2(n32856), .B(n32840), .Y(
        n32922) );
  NAND2xp33_ASAP7_75t_SL U30221 ( .A(n27169), .B(n22392), .Y(n25404) );
  OAI21xp33_ASAP7_75t_SL U30222 ( .A1(sr1_r_MCFG2__RAMBANKSZ__0_), .A2(n31198), 
        .B(n30140), .Y(n1803) );
  OAI21xp5_ASAP7_75t_SL U30223 ( .A1(n24771), .A2(n24876), .B(n24770), .Y(
        n32187) );
  NAND2xp33_ASAP7_75t_SL U30224 ( .A(n27596), .B(n27942), .Y(n27597) );
  NAND2xp33_ASAP7_75t_SL U30225 ( .A(n27654), .B(n27942), .Y(n27655) );
  NAND2xp33_ASAP7_75t_SL U30226 ( .A(uart1_r_BREAK_), .B(n31190), .Y(n28233)
         );
  NAND2xp33_ASAP7_75t_SL U30227 ( .A(n27664), .B(n27925), .Y(n27665) );
  NAND2xp33_ASAP7_75t_SL U30228 ( .A(n31335), .B(n22392), .Y(n25407) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30229 ( .A1(irqctrl0_r_ILEVEL__15_), .A2(n31248), 
        .B(n31025), .C(n31954), .Y(n31026) );
  AOI22xp33_ASAP7_75t_SL U30230 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__13_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__1_), .B2(n24584), .Y(
        n2655) );
  AOI22xp33_ASAP7_75t_SL U30231 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__14_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__2_), .B2(n31986), .Y(
        n3599) );
  AOI22xp33_ASAP7_75t_SL U30232 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__15_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__3_), .B2(n31986), .Y(
        n3598) );
  AOI22xp33_ASAP7_75t_SL U30233 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__21_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__9_), .B2(n24584), .Y(
        n3597) );
  AOI22xp33_ASAP7_75t_SL U30234 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__23_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__11_), .B2(n31986), 
        .Y(n3596) );
  AOI22xp33_ASAP7_75t_SL U30235 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__26_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__14_), .B2(n24584), 
        .Y(n3595) );
  AOI22xp33_ASAP7_75t_SL U30236 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__28_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__16_), .B2(n31986), 
        .Y(n3594) );
  AOI22xp33_ASAP7_75t_SL U30237 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__29_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__17_), .B2(n31986), 
        .Y(n3593) );
  AOI22xp33_ASAP7_75t_SL U30238 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__31_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__19_), .B2(n31986), 
        .Y(n3592) );
  AOI22xp33_ASAP7_75t_SL U30239 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__12_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__0_), .B2(n24584), .Y(
        n2679) );
  OAI21xp33_ASAP7_75t_SL U30240 ( .A1(n28725), .A2(n25198), .B(n25476), .Y(
        n25470) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30241 ( .A1(u0_0_leon3x0_p0_iu_v_X__DCI__LOCK_), 
        .A2(n24648), .B(n32020), .C(n32019), .Y(n3586) );
  OAI21xp33_ASAP7_75t_SL U30242 ( .A1(apbi[31]), .A2(n29650), .B(n29649), .Y(
        n29393) );
  NAND2xp33_ASAP7_75t_SL U30243 ( .A(n29391), .B(n29390), .Y(n29394) );
  OAI21xp33_ASAP7_75t_SL U30244 ( .A1(apbi[20]), .A2(n29650), .B(n29649), .Y(
        n29319) );
  INVx1_ASAP7_75t_SL U30245 ( .A(n28802), .Y(n28808) );
  INVxp67_ASAP7_75t_SL U30246 ( .A(n29322), .Y(n29317) );
  OAI21xp33_ASAP7_75t_SL U30247 ( .A1(apbi[18]), .A2(n29650), .B(n29649), .Y(
        n29332) );
  INVxp67_ASAP7_75t_SL U30248 ( .A(n29379), .Y(n29330) );
  AOI22xp33_ASAP7_75t_SL U30249 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__16_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__4_), .B2(n31986), .Y(
        n2631) );
  AO21x1_ASAP7_75t_SL U30250 ( .A1(n28928), .A2(n22556), .B(n24631), .Y(n23162) );
  OAI21xp33_ASAP7_75t_SL U30251 ( .A1(apbi[23]), .A2(n29650), .B(n29649), .Y(
        n29281) );
  OAI21xp33_ASAP7_75t_SL U30252 ( .A1(n24495), .A2(DP_OP_1196_128_7433_n456), 
        .B(n28584), .Y(n3554) );
  OAI21xp33_ASAP7_75t_SL U30253 ( .A1(apbi[21]), .A2(n29650), .B(n29649), .Y(
        n29297) );
  OAI21xp33_ASAP7_75t_SL U30254 ( .A1(apbi[17]), .A2(n29650), .B(n29649), .Y(
        n27296) );
  OAI21xp33_ASAP7_75t_SL U30255 ( .A1(n24495), .A2(DP_OP_1196_128_7433_n455), 
        .B(n28589), .Y(n3548) );
  OAI21xp33_ASAP7_75t_SL U30256 ( .A1(n24495), .A2(DP_OP_1196_128_7433_n454), 
        .B(n28614), .Y(n3534) );
  AOI22xp33_ASAP7_75t_SL U30257 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__27_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__15_), .B2(n24584), 
        .Y(n4396) );
  NAND2xp33_ASAP7_75t_SL U30258 ( .A(n24681), .B(n29624), .Y(n29625) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30259 ( .A1(n25564), .A2(n26356), .B(n25563), 
        .C(n25562), .Y(n18252) );
  AOI21xp33_ASAP7_75t_SL U30260 ( .A1(n28995), .A2(
        u0_0_leon3x0_p0_iu_r_E__CWP__0_), .B(n28994), .Y(n28997) );
  INVx1_ASAP7_75t_SL U30261 ( .A(n27208), .Y(n30632) );
  INVxp67_ASAP7_75t_SL U30262 ( .A(n31463), .Y(n31591) );
  AOI22xp33_ASAP7_75t_SL U30263 ( .A1(n18610), .A2(n26278), .B1(n23365), .B2(
        n28982), .Y(n27109) );
  AOI22xp33_ASAP7_75t_SL U30264 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__14_), 
        .A2(n28888), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__2_), .B2(n28779), .Y(
        n27205) );
  INVxp33_ASAP7_75t_SL U30265 ( .A(u0_0_leon3x0_p0_divi[13]), .Y(n27197) );
  OA21x2_ASAP7_75t_SL U30266 ( .A1(n18610), .A2(n28827), .B(
        u0_0_leon3x0_p0_divi[13]), .Y(n27198) );
  AOI22xp33_ASAP7_75t_SL U30267 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__30_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__18_), .B2(n31986), 
        .Y(n4321) );
  NAND2xp5_ASAP7_75t_SL U30268 ( .A(n29669), .B(n29667), .Y(n31442) );
  NAND2xp5_ASAP7_75t_SL U30269 ( .A(u0_0_leon3x0_p0_div0_r_CNT__0_), .B(n24909), .Y(n24901) );
  NAND2xp33_ASAP7_75t_SL U30270 ( .A(n28821), .B(u0_0_leon3x0_p0_divi[12]), 
        .Y(n26163) );
  OAI21xp33_ASAP7_75t_SL U30271 ( .A1(n31188), .A2(n31057), .B(n27524), .Y(
        n28191) );
  NOR2x1_ASAP7_75t_SL U30272 ( .A(n22375), .B(n27208), .Y(n28762) );
  NAND2xp5_ASAP7_75t_SL U30273 ( .A(n24681), .B(n29211), .Y(n30701) );
  OAI21xp33_ASAP7_75t_SL U30274 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_M__CTRL__ANNUL_), .B(n32070), .Y(n3707) );
  OAI21xp33_ASAP7_75t_SL U30275 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_r_X__CTRL__ANNUL_), .B(n32071), .Y(n3705) );
  AOI22xp33_ASAP7_75t_SL U30276 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__24_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__12_), .B2(n24584), 
        .Y(n2481) );
  AOI22xp33_ASAP7_75t_SL U30277 ( .A1(u0_0_leon3x0_p0_divo[24]), .A2(n31421), 
        .B1(u0_0_leon3x0_p0_divi[55]), .B2(n31662), .Y(n28307) );
  AOI22xp33_ASAP7_75t_SL U30278 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__22_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__10_), .B2(n24584), 
        .Y(n2508) );
  AOI22xp33_ASAP7_75t_SL U30279 ( .A1(u0_0_leon3x0_p0_divo[22]), .A2(n31421), 
        .B1(u0_0_leon3x0_p0_divi[53]), .B2(n31662), .Y(n28311) );
  AOI22xp33_ASAP7_75t_SL U30280 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__20_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__8_), .B2(n31986), .Y(
        n2535) );
  AOI22xp33_ASAP7_75t_SL U30281 ( .A1(u0_0_leon3x0_p0_divo[20]), .A2(n31421), 
        .B1(u0_0_leon3x0_p0_divi[51]), .B2(n31662), .Y(n27023) );
  NAND2xp33_ASAP7_75t_SL U30282 ( .A(n23980), .B(n29144), .Y(n26742) );
  INVxp67_ASAP7_75t_SL U30283 ( .A(DP_OP_1196_128_7433_n179), .Y(
        DP_OP_1196_128_7433_n177) );
  AOI22xp33_ASAP7_75t_SL U30284 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__19_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__7_), .B2(n24584), .Y(
        n2558) );
  INVxp67_ASAP7_75t_SL U30285 ( .A(n32043), .Y(n25600) );
  NAND2xp33_ASAP7_75t_SL U30286 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[5]), .B(n31877), .Y(n25267) );
  OAI21xp33_ASAP7_75t_SL U30287 ( .A1(n23980), .A2(n30008), .B(n28102), .Y(
        n28104) );
  NAND2xp33_ASAP7_75t_SL U30288 ( .A(n31001), .B(n31465), .Y(n27249) );
  AOI22xp33_ASAP7_75t_SL U30289 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__18_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__6_), .B2(n24584), .Y(
        n2586) );
  AOI22xp33_ASAP7_75t_SL U30290 ( .A1(uart1_r_BRATE__0_), .A2(n31246), .B1(
        timer0_r_RELOAD__0_), .B2(n31237), .Y(n28080) );
  AOI21xp33_ASAP7_75t_SL U30291 ( .A1(n30622), .A2(u0_0_leon3x0_p0_divi[14]), 
        .B(n26573), .Y(n26578) );
  INVxp67_ASAP7_75t_SL U30292 ( .A(DP_OP_1196_128_7433_n207), .Y(
        DP_OP_1196_128_7433_n205) );
  NAND2xp5_ASAP7_75t_SL U30293 ( .A(n27256), .B(n28562), .Y(n3636) );
  OAI21xp33_ASAP7_75t_SL U30294 ( .A1(n28096), .A2(n31973), .B(n30979), .Y(
        n28097) );
  AOI22xp33_ASAP7_75t_SL U30295 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__17_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__5_), .B2(n24584), .Y(
        n2607) );
  NAND2xp5_ASAP7_75t_SL U30296 ( .A(n25849), .B(n25848), .Y(n29515) );
  NAND2xp33_ASAP7_75t_SL U30297 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__4_), .B(
        n28779), .Y(n26677) );
  NAND2xp5_ASAP7_75t_SL U30298 ( .A(n29225), .B(n29230), .Y(n31443) );
  NAND2xp33_ASAP7_75t_SL U30299 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[6]), .B(n31877), .Y(n24980) );
  AOI22xp33_ASAP7_75t_SL U30300 ( .A1(uart1_r_TCNT__5_), .A2(n31951), .B1(
        irqctrl0_r_IPEND__9_), .B2(n31247), .Y(n30146) );
  NAND3xp33_ASAP7_75t_SRAM U30301 ( .A(n24988), .B(n24987), .C(n24986), .Y(
        n24997) );
  OAI21xp5_ASAP7_75t_SL U30302 ( .A1(n28725), .A2(n28868), .B(n26254), .Y(
        n28978) );
  NAND2xp33_ASAP7_75t_SL U30303 ( .A(n18614), .B(n26358), .Y(n26364) );
  AOI22xp33_ASAP7_75t_SL U30304 ( .A1(n22837), .A2(n24577), .B1(n22556), .B2(
        n28982), .Y(n28916) );
  INVxp67_ASAP7_75t_SL U30305 ( .A(mult_x_1196_n2782), .Y(n22997) );
  OAI21xp5_ASAP7_75t_SL U30306 ( .A1(n28621), .A2(n28868), .B(n26253), .Y(
        n28844) );
  OAI22xp33_ASAP7_75t_SL U30307 ( .A1(n22902), .A2(n28843), .B1(n28490), .B2(
        n26294), .Y(n26250) );
  OAI21xp33_ASAP7_75t_SL U30308 ( .A1(n31001), .A2(n30881), .B(n31465), .Y(
        n30882) );
  NAND2xp33_ASAP7_75t_SL U30309 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[8]), .B(n31877), .Y(n25270) );
  NAND2xp33_ASAP7_75t_SL U30310 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[7]), .B(n31877), .Y(n25269) );
  INVxp33_ASAP7_75t_SL U30311 ( .A(n30682), .Y(n24875) );
  NAND2xp33_ASAP7_75t_SL U30312 ( .A(sr1_r_MCFG1__IOWIDTH__0_), .B(n32003), 
        .Y(n30897) );
  INVxp33_ASAP7_75t_SL U30313 ( .A(n31589), .Y(n31592) );
  AOI22xp33_ASAP7_75t_SL U30314 ( .A1(uart1_r_BRATE__11_), .A2(n31246), .B1(
        irqctrl0_r_IPEND__11_), .B2(n31247), .Y(n28127) );
  OAI21xp33_ASAP7_75t_SL U30315 ( .A1(n2924), .A2(n30982), .B(n28122), .Y(
        n28124) );
  AOI21xp33_ASAP7_75t_SL U30316 ( .A1(n32003), .A2(sr1_r_MCFG1__ROMWRITE_), 
        .B(n31849), .Y(n28120) );
  OAI21xp33_ASAP7_75t_SL U30317 ( .A1(n22396), .A2(n31301), .B(n31300), .Y(
        n2968) );
  NAND2xp33_ASAP7_75t_SL U30318 ( .A(n24579), .B(u0_0_leon3x0_p0_divi[20]), 
        .Y(n27058) );
  OAI22xp33_ASAP7_75t_SL U30319 ( .A1(n29352), .A2(n31973), .B1(n26502), .B2(
        n31323), .Y(n26504) );
  INVxp33_ASAP7_75t_SL U30320 ( .A(u0_0_leon3x0_p0_divi[23]), .Y(n26383) );
  OA21x2_ASAP7_75t_SL U30321 ( .A1(n23002), .A2(n28827), .B(
        u0_0_leon3x0_p0_divi[23]), .Y(n26384) );
  NAND2xp33_ASAP7_75t_SL U30322 ( .A(n31567), .B(n31566), .Y(n31569) );
  INVxp33_ASAP7_75t_SL U30323 ( .A(n26788), .Y(n26772) );
  AOI22xp33_ASAP7_75t_SL U30324 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__25_), 
        .A2(n31987), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__13_), .B2(n31986), 
        .Y(n4601) );
  INVxp67_ASAP7_75t_SL U30325 ( .A(mult_x_1196_n2879), .Y(n23085) );
  INVxp67_ASAP7_75t_SL U30326 ( .A(mult_x_1196_n3228), .Y(n23309) );
  NAND2xp33_ASAP7_75t_SL U30327 ( .A(sr1_r_MCFG1__IOWIDTH__1_), .B(n32003), 
        .Y(n31502) );
  OAI21xp33_ASAP7_75t_SL U30328 ( .A1(n30980), .A2(n31973), .B(n30979), .Y(
        n30992) );
  OAI21xp33_ASAP7_75t_SL U30329 ( .A1(n32774), .A2(n30982), .B(n30981), .Y(
        n30986) );
  AOI22xp33_ASAP7_75t_SL U30330 ( .A1(uart1_r_BRATE__10_), .A2(n31246), .B1(
        irqctrl0_r_IPEND__10_), .B2(n31247), .Y(n30989) );
  NAND2xp5_ASAP7_75t_SL U30331 ( .A(n26097), .B(n31248), .Y(n29383) );
  NAND2xp33_ASAP7_75t_SL U30332 ( .A(n24580), .B(u0_0_leon3x0_p0_divi[11]), 
        .Y(n28625) );
  INVxp33_ASAP7_75t_SL U30333 ( .A(n26923), .Y(n26919) );
  INVxp67_ASAP7_75t_SL U30334 ( .A(n28190), .Y(n2864) );
  AOI21xp33_ASAP7_75t_SL U30335 ( .A1(n29214), .A2(n30118), .B(n29213), .Y(
        n29215) );
  AOI21xp33_ASAP7_75t_SL U30336 ( .A1(n28779), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__0_), .B(n28634), .Y(n28635) );
  INVxp33_ASAP7_75t_SL U30337 ( .A(n29667), .Y(n29668) );
  AOI22xp33_ASAP7_75t_SL U30338 ( .A1(n30694), .A2(n30621), .B1(
        u0_0_leon3x0_p0_iu_r_W__S__TT__7_), .B2(n28779), .Y(n28686) );
  AO21x1_ASAP7_75t_SL U30339 ( .A1(n29150), .A2(n23365), .B(n23361), .Y(n23360) );
  OAI21xp33_ASAP7_75t_SL U30340 ( .A1(n29144), .A2(n23365), .B(n23364), .Y(
        n23363) );
  INVx1_ASAP7_75t_SL U30341 ( .A(n31735), .Y(n29522) );
  AOI21xp33_ASAP7_75t_SL U30342 ( .A1(n29226), .A2(n29225), .B(n24510), .Y(
        n29229) );
  OAI21xp33_ASAP7_75t_SL U30343 ( .A1(n30273), .A2(n29594), .B(n28492), .Y(
        n28493) );
  OAI21xp33_ASAP7_75t_SL U30344 ( .A1(n3325), .A2(n29738), .B(n25949), .Y(
        n18049) );
  OAI21xp33_ASAP7_75t_SL U30345 ( .A1(sr1_r_MCFG2__RAMWIDTH__1_), .A2(n31198), 
        .B(n30074), .Y(n2911) );
  OAI21xp33_ASAP7_75t_SL U30346 ( .A1(sr1_r_MCFG2__RAMWIDTH__0_), .A2(n31198), 
        .B(n30781), .Y(n2912) );
  INVxp33_ASAP7_75t_SL U30347 ( .A(u0_0_leon3x0_p0_divi[22]), .Y(n26429) );
  OAI21xp33_ASAP7_75t_SL U30348 ( .A1(n30965), .A2(n29199), .B(n29186), .Y(
        n29187) );
  INVxp33_ASAP7_75t_SL U30349 ( .A(n28843), .Y(n28846) );
  NAND2xp33_ASAP7_75t_SL U30350 ( .A(n28830), .B(u0_0_leon3x0_p0_divi[19]), 
        .Y(n26991) );
  NAND2xp33_ASAP7_75t_SL U30351 ( .A(n27738), .B(n27955), .Y(n27739) );
  NAND2xp5_ASAP7_75t_SL U30352 ( .A(n25400), .B(n31566), .Y(n30203) );
  OAI22xp33_ASAP7_75t_SL U30353 ( .A1(n4775), .A2(n29385), .B1(n30833), .B2(
        n29384), .Y(n17853) );
  NAND2xp5_ASAP7_75t_SL U30354 ( .A(n26097), .B(n30790), .Y(n30030) );
  OAI21xp33_ASAP7_75t_SL U30355 ( .A1(n28829), .A2(n30008), .B(n25871), .Y(
        n25873) );
  AOI22xp33_ASAP7_75t_SL U30356 ( .A1(n30622), .A2(u0_0_leon3x0_p0_divi[6]), 
        .B1(u0_0_leon3x0_p0_iu_r_W__S__WIM__7_), .B2(n28890), .Y(n28783) );
  OAI22xp33_ASAP7_75t_SL U30357 ( .A1(n2235), .A2(n29385), .B1(n28116), .B2(
        n29384), .Y(n17857) );
  NAND2xp33_ASAP7_75t_SL U30358 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[2]), .B(n31877), .Y(n25265) );
  NAND2xp33_ASAP7_75t_SL U30359 ( .A(n27317), .B(n27316), .Y(n27318) );
  INVxp33_ASAP7_75t_SL U30360 ( .A(n30790), .Y(n30107) );
  NAND2xp33_ASAP7_75t_SL U30361 ( .A(n27940), .B(n27942), .Y(n27941) );
  NAND2xp33_ASAP7_75t_SL U30362 ( .A(n27923), .B(n27925), .Y(n27924) );
  NAND2xp33_ASAP7_75t_SL U30363 ( .A(n27953), .B(n27955), .Y(n27954) );
  NAND2xp33_ASAP7_75t_SL U30364 ( .A(n27969), .B(n27971), .Y(n27970) );
  NAND2xp33_ASAP7_75t_SL U30365 ( .A(n27943), .B(n27945), .Y(n27944) );
  INVxp67_ASAP7_75t_SL U30366 ( .A(n29376), .Y(n29657) );
  NAND2xp33_ASAP7_75t_SL U30367 ( .A(n27916), .B(n27918), .Y(n27917) );
  XNOR2xp5_ASAP7_75t_SL U30368 ( .A(n24063), .B(n23971), .Y(mult_x_1196_n2858)
         );
  NAND2xp33_ASAP7_75t_SL U30369 ( .A(n27956), .B(n27958), .Y(n27957) );
  INVxp67_ASAP7_75t_SL U30370 ( .A(n32662), .Y(n31892) );
  AO21x1_ASAP7_75t_SRAM U30371 ( .A1(n27305), .A2(n29356), .B(
        uart1_r_TWADDR__2_), .Y(n27306) );
  NAND2xp33_ASAP7_75t_SL U30372 ( .A(n27380), .B(n29356), .Y(n27307) );
  OAI22xp33_ASAP7_75t_SL U30373 ( .A1(n18801), .A2(n31628), .B1(n32033), .B2(
        n31628), .Y(n31630) );
  NAND2xp33_ASAP7_75t_SL U30374 ( .A(n28821), .B(u0_0_leon3x0_p0_divi[6]), .Y(
        n28772) );
  NAND2xp5_ASAP7_75t_SL U30375 ( .A(n25992), .B(n27496), .Y(n25995) );
  NAND2xp5_ASAP7_75t_SL U30376 ( .A(n31954), .B(n31956), .Y(n32004) );
  NAND2xp33_ASAP7_75t_SL U30377 ( .A(n27730), .B(n27945), .Y(n27731) );
  NAND2xp33_ASAP7_75t_SL U30378 ( .A(n27714), .B(n27918), .Y(n27715) );
  NAND2xp33_ASAP7_75t_SL U30379 ( .A(n27740), .B(n27958), .Y(n27741) );
  NAND2xp33_ASAP7_75t_SL U30380 ( .A(n27790), .B(n27942), .Y(n27791) );
  NAND2xp33_ASAP7_75t_SL U30381 ( .A(n27800), .B(n27925), .Y(n27801) );
  NAND2xp33_ASAP7_75t_SL U30382 ( .A(n27810), .B(n27955), .Y(n27811) );
  NAND2xp33_ASAP7_75t_SL U30383 ( .A(n27820), .B(n27971), .Y(n27821) );
  NAND2xp33_ASAP7_75t_SL U30384 ( .A(n27792), .B(n27945), .Y(n27793) );
  NAND2xp33_ASAP7_75t_SL U30385 ( .A(n27796), .B(n27918), .Y(n27797) );
  NAND2xp33_ASAP7_75t_SL U30386 ( .A(n27812), .B(n27958), .Y(n27813) );
  NAND2xp33_ASAP7_75t_SL U30387 ( .A(n27864), .B(n27942), .Y(n27865) );
  NAND2xp33_ASAP7_75t_SL U30388 ( .A(n27854), .B(n27925), .Y(n27855) );
  NAND2xp33_ASAP7_75t_SL U30389 ( .A(n27874), .B(n27955), .Y(n27875) );
  NAND2xp33_ASAP7_75t_SL U30390 ( .A(n27884), .B(n27971), .Y(n27885) );
  NAND2xp33_ASAP7_75t_SL U30391 ( .A(n27866), .B(n27945), .Y(n27867) );
  NAND2xp33_ASAP7_75t_SL U30392 ( .A(n27850), .B(n27918), .Y(n27851) );
  NAND2xp33_ASAP7_75t_SL U30393 ( .A(n27876), .B(n27958), .Y(n27877) );
  NAND2xp33_ASAP7_75t_SL U30394 ( .A(n27331), .B(n27942), .Y(n27332) );
  NAND2xp33_ASAP7_75t_SL U30395 ( .A(n27347), .B(n27925), .Y(n27348) );
  NAND2xp33_ASAP7_75t_SL U30396 ( .A(n27362), .B(n27955), .Y(n27363) );
  NAND2xp33_ASAP7_75t_SL U30397 ( .A(n27378), .B(n27971), .Y(n27379) );
  NAND2xp33_ASAP7_75t_SL U30398 ( .A(n27335), .B(n27945), .Y(n27336) );
  NAND2xp33_ASAP7_75t_SL U30399 ( .A(n27341), .B(n27918), .Y(n27342) );
  NAND2xp33_ASAP7_75t_SL U30400 ( .A(n27366), .B(n27958), .Y(n27367) );
  NAND2xp33_ASAP7_75t_SL U30401 ( .A(n24681), .B(n30938), .Y(n32177) );
  NAND2xp33_ASAP7_75t_SL U30402 ( .A(n27748), .B(n27971), .Y(n27749) );
  INVxp67_ASAP7_75t_SL U30403 ( .A(mult_x_1196_n3192), .Y(n23158) );
  OAI21xp33_ASAP7_75t_SL U30404 ( .A1(n32159), .A2(n26788), .B(n26800), .Y(
        n26799) );
  NAND2xp5_ASAP7_75t_SL U30405 ( .A(n31327), .B(n27496), .Y(n27506) );
  NAND2xp5_ASAP7_75t_SL U30406 ( .A(n29516), .B(timer0_v_TICK_), .Y(n29517) );
  INVxp67_ASAP7_75t_SL U30407 ( .A(n29516), .Y(n25851) );
  INVxp67_ASAP7_75t_SL U30408 ( .A(n29390), .Y(n29237) );
  INVxp33_ASAP7_75t_SL U30409 ( .A(n27496), .Y(n25994) );
  OAI21xp33_ASAP7_75t_SL U30410 ( .A1(apbi[26]), .A2(n29650), .B(n29649), .Y(
        n29264) );
  NAND2xp5_ASAP7_75t_SL U30411 ( .A(n27914), .B(n27913), .Y(n29559) );
  OR2x2_ASAP7_75t_SL U30412 ( .A(n25025), .B(n25024), .Y(n31469) );
  INVx1_ASAP7_75t_SL U30413 ( .A(n31466), .Y(n30995) );
  NOR2x1_ASAP7_75t_SL U30414 ( .A(n25476), .B(n25092), .Y(n26155) );
  OAI21xp33_ASAP7_75t_SL U30415 ( .A1(n22902), .A2(n30008), .B(n25857), .Y(
        n25859) );
  AOI22xp33_ASAP7_75t_SL U30416 ( .A1(uart1_r_BRATE__8_), .A2(n31246), .B1(
        irqctrl0_r_IPEND__8_), .B2(n31247), .Y(n29754) );
  INVxp67_ASAP7_75t_SL U30417 ( .A(n31465), .Y(n30559) );
  OAI21xp33_ASAP7_75t_SL U30418 ( .A1(apbi[19]), .A2(n29650), .B(n29649), .Y(
        n28240) );
  INVxp67_ASAP7_75t_SL U30419 ( .A(mult_x_1196_n3112), .Y(n22718) );
  INVxp33_ASAP7_75t_SL U30420 ( .A(DP_OP_1196_128_7433_n354), .Y(
        DP_OP_1196_128_7433_n386) );
  INVxp33_ASAP7_75t_SL U30421 ( .A(n32391), .Y(n32645) );
  OAI21xp33_ASAP7_75t_SL U30422 ( .A1(n31261), .A2(n25402), .B(n24684), .Y(
        n31566) );
  AOI21xp33_ASAP7_75t_SL U30423 ( .A1(n30644), .A2(n28540), .B(n28539), .Y(
        n28541) );
  OAI22xp33_ASAP7_75t_SL U30424 ( .A1(n32814), .A2(n32820), .B1(n32813), .B2(
        n32812), .Y(n32819) );
  INVxp33_ASAP7_75t_SL U30425 ( .A(DP_OP_1196_128_7433_n350), .Y(
        DP_OP_1196_128_7433_n385) );
  NAND2xp33_ASAP7_75t_SL U30426 ( .A(n26770), .B(n29214), .Y(n26788) );
  NAND2xp33_ASAP7_75t_SL U30427 ( .A(n24874), .B(n29177), .Y(n24895) );
  NAND2xp33_ASAP7_75t_SL U30428 ( .A(n32244), .B(n22396), .Y(n31300) );
  INVx1_ASAP7_75t_SL U30429 ( .A(n24511), .Y(n22414) );
  INVxp67_ASAP7_75t_SL U30430 ( .A(n30872), .Y(n31240) );
  XNOR2xp5_ASAP7_75t_SL U30431 ( .A(n24063), .B(n23969), .Y(mult_x_1196_n2926)
         );
  AOI22xp33_ASAP7_75t_SL U30432 ( .A1(uart1_uarto_TXEN_), .A2(n31950), .B1(
        n31245), .B2(timer0_r_SCALER__1_), .Y(n27467) );
  AOI21xp33_ASAP7_75t_SL U30433 ( .A1(n30644), .A2(n27169), .B(n27130), .Y(
        n27131) );
  NAND2xp33_ASAP7_75t_SL U30434 ( .A(n27459), .B(n28231), .Y(n30548) );
  NAND2xp5_ASAP7_75t_SL U30435 ( .A(n28032), .B(n27581), .Y(n29954) );
  AOI21xp33_ASAP7_75t_SL U30436 ( .A1(n30644), .A2(n30721), .B(n28751), .Y(
        n28752) );
  OAI21xp33_ASAP7_75t_SL U30437 ( .A1(n3916), .A2(n29592), .B(n27113), .Y(
        n27117) );
  NAND2xp33_ASAP7_75t_SL U30438 ( .A(n22721), .B(n29146), .Y(n28626) );
  NAND2xp5_ASAP7_75t_SL U30439 ( .A(n27895), .B(n27894), .Y(n27914) );
  OAI31xp33_ASAP7_75t_SRAM U30440 ( .A1(n29214), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__PS_), .A3(n29212), .B(n24681), .Y(n29213)
         );
  NAND2xp33_ASAP7_75t_SL U30441 ( .A(u0_0_leon3x0_p0_divi[43]), .B(n28782), 
        .Y(n28636) );
  NOR3xp33_ASAP7_75t_SRAM U30442 ( .A(n31657), .B(n24912), .C(n26817), .Y(
        n24913) );
  INVx1_ASAP7_75t_SL U30443 ( .A(DP_OP_1196_128_7433_n338), .Y(
        DP_OP_1196_128_7433_n6) );
  INVxp33_ASAP7_75t_SL U30444 ( .A(n31440), .Y(n29227) );
  INVxp33_ASAP7_75t_SL U30445 ( .A(n31672), .Y(n29108) );
  NAND2xp5_ASAP7_75t_SL U30446 ( .A(n24881), .B(n25216), .Y(n31817) );
  NAND2xp5_ASAP7_75t_SL U30447 ( .A(n29738), .B(n29676), .Y(n25949) );
  AOI22xp5_ASAP7_75t_SL U30448 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TT__6_), .A2(
        n29740), .B1(n29739), .B2(n29738), .Y(n3324) );
  OAI21xp33_ASAP7_75t_SL U30449 ( .A1(n22939), .A2(n29144), .B(n28925), .Y(
        n28927) );
  OAI21xp33_ASAP7_75t_SL U30450 ( .A1(n32075), .A2(n29648), .B(n29647), .Y(
        n3322) );
  AOI22xp33_ASAP7_75t_SL U30451 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), 
        .A2(n24649), .B1(u0_0_leon3x0_p0_iu_r_M__CTRL__WICC_), .B2(n32068), 
        .Y(n3711) );
  NAND2xp33_ASAP7_75t_SL U30452 ( .A(n22449), .B(n29146), .Y(n28882) );
  NAND2xp33_ASAP7_75t_SL U30453 ( .A(n24579), .B(u0_0_leon3x0_p0_divi[2]), .Y(
        n28881) );
  NAND2xp5_ASAP7_75t_SL U30454 ( .A(n24750), .B(n24749), .Y(n24751) );
  NAND2xp33_ASAP7_75t_SL U30455 ( .A(uart1_r_BRATE__9_), .B(n31246), .Y(n30145) );
  OAI21xp33_ASAP7_75t_SL U30456 ( .A1(n29206), .A2(n29202), .B(n26806), .Y(
        n26808) );
  NAND2xp5_ASAP7_75t_SL U30457 ( .A(n25561), .B(n25560), .Y(n25562) );
  NAND2xp33_ASAP7_75t_SL U30458 ( .A(n27194), .B(n25610), .Y(n25563) );
  OAI22xp33_ASAP7_75t_SL U30459 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__27_), 
        .A2(n27143), .B1(n22426), .B2(n27141), .Y(n26902) );
  OAI21xp33_ASAP7_75t_SL U30460 ( .A1(n26896), .A2(n29592), .B(n26895), .Y(
        n26897) );
  AOI22xp33_ASAP7_75t_SL U30461 ( .A1(uart1_r_BRATE__5_), .A2(n31246), .B1(
        n31951), .B2(uart1_r_PARERR_), .Y(n30100) );
  OAI21xp33_ASAP7_75t_SL U30462 ( .A1(n32075), .A2(n29476), .B(n25950), .Y(
        n2766) );
  AOI22xp33_ASAP7_75t_SL U30463 ( .A1(uart1_r_PAREN_), .A2(n31950), .B1(n31245), .B2(timer0_r_SCALER__5_), .Y(n30075) );
  NAND2xp33_ASAP7_75t_SL U30464 ( .A(uart1_r_TXCLK__0_), .B(n29949), .Y(n26082) );
  NAND2xp5_ASAP7_75t_SL U30465 ( .A(n27330), .B(n27376), .Y(n27942) );
  NAND2xp5_ASAP7_75t_SL U30466 ( .A(n27346), .B(n27376), .Y(n27925) );
  NAND2xp5_ASAP7_75t_SL U30467 ( .A(n27361), .B(n27376), .Y(n27955) );
  NAND2xp5_ASAP7_75t_SL U30468 ( .A(n27377), .B(n27376), .Y(n27971) );
  NAND2xp33_ASAP7_75t_SL U30469 ( .A(u0_0_leon3x0_p0_divi[48]), .B(n28782), 
        .Y(n26701) );
  NOR2x1_ASAP7_75t_SL U30470 ( .A(n31529), .B(n29743), .Y(n29745) );
  AOI22xp33_ASAP7_75t_SL U30471 ( .A1(n30612), .A2(u0_0_leon3x0_p0_divi[31]), 
        .B1(u0_0_leon3x0_p0_iu_r_W__S__WIM__0_), .B2(n30611), .Y(n28999) );
  NAND2xp5_ASAP7_75t_SL U30472 ( .A(n27334), .B(n27376), .Y(n27945) );
  NAND2xp5_ASAP7_75t_SL U30473 ( .A(n27340), .B(n27376), .Y(n27918) );
  NAND2xp5_ASAP7_75t_SL U30474 ( .A(n27365), .B(n27376), .Y(n27958) );
  INVxp33_ASAP7_75t_SL U30475 ( .A(n29474), .Y(n29475) );
  AND2x2_ASAP7_75t_SL U30476 ( .A(n23161), .B(n28982), .Y(n23160) );
  INVxp33_ASAP7_75t_SL U30477 ( .A(n30621), .Y(n28727) );
  OAI22xp5_ASAP7_75t_SL U30478 ( .A1(n4701), .A2(n29948), .B1(n28028), .B2(
        n28027), .Y(n28029) );
  NAND2xp5_ASAP7_75t_SL U30479 ( .A(n2267), .B(n27325), .Y(n27381) );
  XNOR2xp5_ASAP7_75t_SL U30480 ( .A(n24064), .B(n23969), .Y(mult_x_1196_n2927)
         );
  OAI21xp33_ASAP7_75t_SL U30481 ( .A1(n31396), .A2(n29930), .B(n29929), .Y(
        n29931) );
  INVx1_ASAP7_75t_SL U30482 ( .A(n26278), .Y(n28868) );
  AOI21xp33_ASAP7_75t_SL U30483 ( .A1(n30644), .A2(n27027), .B(n27010), .Y(
        n27011) );
  NAND2xp33_ASAP7_75t_SL U30484 ( .A(n24694), .B(n32705), .Y(n32040) );
  INVxp67_ASAP7_75t_SL U30485 ( .A(n33061), .Y(n32822) );
  INVxp33_ASAP7_75t_SL U30486 ( .A(n32704), .Y(n32706) );
  OAI22xp33_ASAP7_75t_SL U30487 ( .A1(n32912), .A2(n32943), .B1(n32906), .B2(
        n32895), .Y(n32896) );
  NAND2xp33_ASAP7_75t_SL U30488 ( .A(n31195), .B(n31501), .Y(n31196) );
  OAI22xp33_ASAP7_75t_SL U30489 ( .A1(n32912), .A2(n32951), .B1(n32906), .B2(
        n32897), .Y(n32898) );
  NAND2xp33_ASAP7_75t_SL U30490 ( .A(n30137), .B(n31501), .Y(n30138) );
  NAND2xp33_ASAP7_75t_SL U30491 ( .A(n30139), .B(n31198), .Y(n30140) );
  OAI22xp33_ASAP7_75t_SL U30492 ( .A1(n32912), .A2(n32959), .B1(n32906), .B2(
        n32899), .Y(n32900) );
  AOI22xp33_ASAP7_75t_SL U30493 ( .A1(u0_0_leon3x0_p0_iu_r_M__CTRL__WICC_), 
        .A2(n24649), .B1(u0_0_leon3x0_p0_iu_r_E__CTRL__WICC_), .B2(n32068), 
        .Y(n3713) );
  NAND2xp33_ASAP7_75t_SL U30494 ( .A(n32069), .B(n32068), .Y(n32070) );
  NAND2xp33_ASAP7_75t_SL U30495 ( .A(n30868), .B(n31501), .Y(n30869) );
  OAI22xp33_ASAP7_75t_SL U30496 ( .A1(n32912), .A2(n32967), .B1(n32906), .B2(
        n32901), .Y(n32902) );
  NOR2x1_ASAP7_75t_SL U30497 ( .A(n24464), .B(n27057), .Y(
        u0_0_leon3x0_p0_divi[20]) );
  NAND2xp33_ASAP7_75t_SL U30498 ( .A(n28057), .B(n31501), .Y(n28058) );
  NAND2xp5_ASAP7_75t_SL U30499 ( .A(n27380), .B(n27376), .Y(n27965) );
  NOR2x1_ASAP7_75t_SL U30500 ( .A(n24466), .B(n28479), .Y(
        u0_0_leon3x0_p0_divi[21]) );
  OAI22xp33_ASAP7_75t_SL U30501 ( .A1(n32912), .A2(n32978), .B1(n32906), .B2(
        n32905), .Y(n32907) );
  NAND2xp33_ASAP7_75t_SL U30502 ( .A(n28236), .B(n31501), .Y(n28237) );
  NOR2x1_ASAP7_75t_SL U30503 ( .A(n26382), .B(n26381), .Y(
        u0_0_leon3x0_p0_divi[23]) );
  OAI21xp33_ASAP7_75t_SL U30504 ( .A1(n25765), .A2(n29592), .B(n25764), .Y(
        n25767) );
  NAND2xp33_ASAP7_75t_SL U30505 ( .A(ahbso_0__HRDATA__24_), .B(n32973), .Y(
        n32914) );
  NAND2xp5_ASAP7_75t_SL U30506 ( .A(n29738), .B(n29729), .Y(n29730) );
  NAND2xp33_ASAP7_75t_SL U30507 ( .A(n23365), .B(n29146), .Y(n23364) );
  OAI22xp33_ASAP7_75t_SL U30508 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__6_), 
        .A2(n31256), .B1(n22421), .B2(u0_0_leon3x0_p0_dci[38]), .Y(n3680) );
  NAND2xp33_ASAP7_75t_SL U30509 ( .A(ahbso_0__HRDATA__25_), .B(n32973), .Y(
        n32924) );
  OAI21xp33_ASAP7_75t_SL U30510 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__7_), .B(n30877), .Y(n3675) );
  INVxp67_ASAP7_75t_SL U30511 ( .A(n30814), .Y(n28760) );
  NAND2xp33_ASAP7_75t_SL U30512 ( .A(ahbso_0__HRDATA__26_), .B(n32973), .Y(
        n32932) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30513 ( .A1(n32522), .A2(n32521), .B(n32565), 
        .C(n32520), .Y(it_data[7]) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30514 ( .A1(n32509), .A2(n32508), .B(n32565), 
        .C(n32507), .Y(it_data[6]) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30515 ( .A1(n32502), .A2(n32501), .B(n32565), 
        .C(n32500), .Y(it_data[5]) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30516 ( .A1(n32488), .A2(n32487), .B(n32565), 
        .C(n32486), .Y(it_data[3]) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30517 ( .A1(n32480), .A2(n32479), .B(n32565), 
        .C(n32478), .Y(it_data[2]) );
  NAND2xp33_ASAP7_75t_SL U30518 ( .A(n24382), .B(n24412), .Y(n24383) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30519 ( .A1(n32473), .A2(n32472), .B(n32565), 
        .C(n32471), .Y(it_data[1]) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30520 ( .A1(n32466), .A2(n32465), .B(n32565), 
        .C(n32464), .Y(it_data[0]) );
  NAND2xp33_ASAP7_75t_SL U30521 ( .A(n28232), .B(n28231), .Y(n31190) );
  NAND2xp33_ASAP7_75t_SL U30522 ( .A(n30780), .B(n31198), .Y(n30781) );
  NAND2xp33_ASAP7_75t_SL U30523 ( .A(n30073), .B(n31198), .Y(n30074) );
  NAND2xp33_ASAP7_75t_SL U30524 ( .A(ahbso_0__HRDATA__0_), .B(n32854), .Y(
        n32840) );
  INVx1_ASAP7_75t_SL U30525 ( .A(n30006), .Y(n27489) );
  INVxp67_ASAP7_75t_SL U30526 ( .A(n28131), .Y(n29909) );
  NAND2xp33_ASAP7_75t_SL U30527 ( .A(ahbso_0__HRDATA__1_), .B(n32854), .Y(
        n32842) );
  NAND2xp33_ASAP7_75t_SL U30528 ( .A(ahbso_0__HRDATA__2_), .B(n32854), .Y(
        n32844) );
  NAND2xp33_ASAP7_75t_SL U30529 ( .A(ahbso_0__HRDATA__3_), .B(n32854), .Y(
        n32846) );
  NAND2xp33_ASAP7_75t_SL U30530 ( .A(ahbso_0__HRDATA__4_), .B(n32854), .Y(
        n32848) );
  INVx1_ASAP7_75t_SL U30531 ( .A(n31501), .Y(n28119) );
  NAND2xp33_ASAP7_75t_SL U30532 ( .A(ahbso_0__HRDATA__5_), .B(n32854), .Y(
        n32850) );
  NAND2xp33_ASAP7_75t_SL U30533 ( .A(ahbso_0__HRDATA__6_), .B(n32854), .Y(
        n32852) );
  NAND2xp33_ASAP7_75t_SL U30534 ( .A(ahbso_0__HRDATA__7_), .B(n32854), .Y(
        n32855) );
  OAI21xp33_ASAP7_75t_SL U30535 ( .A1(n32874), .A2(n32859), .B(n32858), .Y(
        n32923) );
  INVxp67_ASAP7_75t_SL U30536 ( .A(n22436), .Y(n28490) );
  INVxp67_ASAP7_75t_SL U30537 ( .A(n31198), .Y(n26136) );
  NAND2xp5_ASAP7_75t_SL U30538 ( .A(n32862), .B(n32861), .Y(n32931) );
  AOI21xp33_ASAP7_75t_SL U30539 ( .A1(n30652), .A2(
        u0_0_leon3x0_p0_iu_de_icc_3_), .B(n24680), .Y(n29809) );
  OAI21xp33_ASAP7_75t_SL U30540 ( .A1(n32874), .A2(n32864), .B(n32863), .Y(
        n32939) );
  NAND2xp33_ASAP7_75t_SL U30541 ( .A(n31499), .B(n31501), .Y(n31500) );
  OAI21xp33_ASAP7_75t_SL U30542 ( .A1(n32874), .A2(n32866), .B(n32865), .Y(
        n32947) );
  OAI21xp33_ASAP7_75t_SL U30543 ( .A1(n32874), .A2(n32868), .B(n32867), .Y(
        n32955) );
  AOI22xp33_ASAP7_75t_SL U30544 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__12_), .A2(
        n22375), .B1(n22721), .B2(n28131), .Y(n25426) );
  OAI21xp33_ASAP7_75t_SL U30545 ( .A1(n32874), .A2(n32870), .B(n32869), .Y(
        n32963) );
  OAI21xp33_ASAP7_75t_SL U30546 ( .A1(n32874), .A2(n32873), .B(n32872), .Y(
        n32971) );
  INVx1_ASAP7_75t_SL U30547 ( .A(n24907), .Y(n24909) );
  OAI22xp33_ASAP7_75t_SL U30548 ( .A1(n32912), .A2(n32919), .B1(n32906), .B2(
        n32889), .Y(n32890) );
  INVx1_ASAP7_75t_SL U30549 ( .A(n26454), .Y(n26534) );
  OAI22xp33_ASAP7_75t_SL U30550 ( .A1(n32912), .A2(n32927), .B1(n32906), .B2(
        n32891), .Y(n32892) );
  OAI22xp33_ASAP7_75t_SL U30551 ( .A1(n32912), .A2(n32935), .B1(n32906), .B2(
        n32893), .Y(n32894) );
  OAI21xp33_ASAP7_75t_SL U30552 ( .A1(n30397), .A2(n29198), .B(n29183), .Y(
        n30796) );
  INVx1_ASAP7_75t_SL U30553 ( .A(n30134), .Y(n25848) );
  AOI21xp33_ASAP7_75t_SL U30554 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__WIM__5_), 
        .A2(n29198), .B(n29182), .Y(n31438) );
  NAND2xp33_ASAP7_75t_SL U30555 ( .A(u0_0_leon3x0_p0_divi[38]), .B(n28782), 
        .Y(n28784) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30556 ( .A1(n28189), .A2(n29964), .B(n29974), 
        .C(n28188), .Y(n28190) );
  AOI21xp33_ASAP7_75t_SL U30557 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__WIM__1_), 
        .A2(n29198), .B(n29181), .Y(n31347) );
  NOR2xp33_ASAP7_75t_SL U30558 ( .A(n23375), .B(n28827), .Y(n23447) );
  OAI22xp33_ASAP7_75t_SL U30559 ( .A1(n32794), .A2(n32820), .B1(n32813), .B2(
        n32793), .Y(n32795) );
  OAI22xp33_ASAP7_75t_SL U30560 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__28_), 
        .A2(n27143), .B1(n26917), .B2(n27141), .Y(n26923) );
  INVxp33_ASAP7_75t_SL U30561 ( .A(n29861), .Y(n32621) );
  OAI22xp33_ASAP7_75t_SL U30562 ( .A1(n32798), .A2(n32820), .B1(n32813), .B2(
        n32797), .Y(n32800) );
  INVxp33_ASAP7_75t_SL U30563 ( .A(n30808), .Y(n32623) );
  NAND2xp5_ASAP7_75t_SL U30564 ( .A(n31954), .B(n31951), .Y(n31973) );
  OAI21xp33_ASAP7_75t_SL U30565 ( .A1(n23229), .A2(n32730), .B(n32134), .Y(
        n32136) );
  AOI21xp33_ASAP7_75t_SL U30566 ( .A1(n30644), .A2(n28574), .B(n28573), .Y(
        n28575) );
  INVx1_ASAP7_75t_SL U30567 ( .A(n31023), .Y(n31247) );
  INVx1_ASAP7_75t_SL U30568 ( .A(n22721), .Y(n28621) );
  AND3x1_ASAP7_75t_SRAM U30569 ( .A(n25077), .B(n25680), .C(n25230), .Y(n25078) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30570 ( .A1(n25077), .A2(n25230), .B(n24924), 
        .C(n24923), .Y(n3570) );
  OAI22xp33_ASAP7_75t_SL U30571 ( .A1(n32805), .A2(n32820), .B1(n32813), .B2(
        n32804), .Y(n32806) );
  NAND2xp5_ASAP7_75t_SL U30572 ( .A(n25604), .B(n32068), .Y(n32071) );
  AOI21xp33_ASAP7_75t_SL U30573 ( .A1(n30644), .A2(n29899), .B(n28796), .Y(
        n28797) );
  OAI22xp33_ASAP7_75t_SL U30574 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__8_), 
        .A2(n31256), .B1(n23229), .B2(u0_0_leon3x0_p0_dci[40]), .Y(n3662) );
  NAND2xp33_ASAP7_75t_SL U30575 ( .A(ahbso_0__HRDATA__27_), .B(n32973), .Y(
        n32940) );
  NAND2xp33_ASAP7_75t_SL U30576 ( .A(ahbso_0__HRDATA__28_), .B(n32973), .Y(
        n32948) );
  OAI22xp33_ASAP7_75t_SL U30577 ( .A1(n25892), .A2(n27141), .B1(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__29_), .B2(n27143), .Y(n25900) );
  NAND2xp33_ASAP7_75t_SL U30578 ( .A(ahbso_0__HRDATA__29_), .B(n32973), .Y(
        n32956) );
  NAND2xp33_ASAP7_75t_SL U30579 ( .A(ahbso_0__HRDATA__30_), .B(n32973), .Y(
        n32964) );
  INVxp67_ASAP7_75t_SL U30580 ( .A(n30580), .Y(n28562) );
  NAND2xp33_ASAP7_75t_SL U30581 ( .A(ahbso_0__HRDATA__31_), .B(n32973), .Y(
        n32974) );
  AOI21xp33_ASAP7_75t_SL U30582 ( .A1(n30644), .A2(n30465), .B(n28953), .Y(
        n28954) );
  INVxp67_ASAP7_75t_SL U30583 ( .A(n32986), .Y(n32990) );
  XNOR2xp5_ASAP7_75t_SL U30584 ( .A(n24063), .B(n23965), .Y(mult_x_1196_n2994)
         );
  OAI21xp33_ASAP7_75t_SL U30585 ( .A1(n30407), .A2(n29198), .B(n29193), .Y(
        n31014) );
  AOI21xp33_ASAP7_75t_SL U30586 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__WIM__4_), 
        .A2(n29198), .B(n29192), .Y(n29624) );
  OAI21xp33_ASAP7_75t_SL U30587 ( .A1(n30454), .A2(n29594), .B(n28889), .Y(
        n28893) );
  AOI22xp33_ASAP7_75t_SL U30588 ( .A1(n30622), .A2(u0_0_leon3x0_p0_divi[2]), 
        .B1(u0_0_leon3x0_p0_iu_r_W__S__WIM__3_), .B2(n28890), .Y(n28891) );
  AOI21xp33_ASAP7_75t_SL U30589 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__WIM__0_), 
        .A2(n29198), .B(n29190), .Y(n31437) );
  INVxp67_ASAP7_75t_SL U30590 ( .A(n29195), .Y(n29191) );
  NAND2xp5_ASAP7_75t_SL U30591 ( .A(n25369), .B(n29474), .Y(n29674) );
  AOI21xp33_ASAP7_75t_SL U30592 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__WIM__3_), 
        .A2(n29198), .B(n29185), .Y(n30965) );
  NAND2xp33_ASAP7_75t_SL U30593 ( .A(n25392), .B(n31960), .Y(n25393) );
  NAND2xp33_ASAP7_75t_SL U30594 ( .A(n26049), .B(n26060), .Y(n31087) );
  NAND2xp33_ASAP7_75t_SL U30595 ( .A(n26068), .B(n26043), .Y(n31063) );
  NAND2xp33_ASAP7_75t_SL U30596 ( .A(n23161), .B(n24577), .Y(n25786) );
  OAI21xp33_ASAP7_75t_SL U30597 ( .A1(n27069), .A2(n29592), .B(n27068), .Y(
        n27072) );
  NAND2xp33_ASAP7_75t_SL U30598 ( .A(n26045), .B(n26043), .Y(n31159) );
  NAND2xp5_ASAP7_75t_SL U30599 ( .A(n29275), .B(n29279), .Y(n27297) );
  XNOR2xp5_ASAP7_75t_SL U30600 ( .A(n23969), .B(n24051), .Y(mult_x_1196_n2914)
         );
  NAND2xp33_ASAP7_75t_SL U30601 ( .A(n26036), .B(n26060), .Y(n31119) );
  NAND3xp33_ASAP7_75t_SRAM U30602 ( .A(n31575), .B(n31574), .C(n31573), .Y(
        n31576) );
  INVx1_ASAP7_75t_SL U30603 ( .A(n25200), .Y(n25198) );
  NAND2xp33_ASAP7_75t_SL U30604 ( .A(n26032), .B(n26060), .Y(n31091) );
  NOR2x1_ASAP7_75t_SL U30605 ( .A(n32171), .B(n24763), .Y(n26854) );
  XNOR2xp5_ASAP7_75t_SL U30606 ( .A(n24054), .B(n22968), .Y(mult_x_1196_n2781)
         );
  INVx1_ASAP7_75t_SL U30607 ( .A(n29279), .Y(n29294) );
  NAND2xp33_ASAP7_75t_SL U30608 ( .A(n32457), .B(n31582), .Y(n25024) );
  BUFx6f_ASAP7_75t_SL U30609 ( .A(n23966), .Y(n23050) );
  INVxp67_ASAP7_75t_SL U30610 ( .A(DP_OP_1196_128_7433_n138), .Y(
        DP_OP_1196_128_7433_n140) );
  OAI21xp33_ASAP7_75t_SL U30611 ( .A1(n26572), .A2(n29592), .B(n26571), .Y(
        n26573) );
  NAND2xp33_ASAP7_75t_SL U30612 ( .A(n26055), .B(n26060), .Y(n31147) );
  INVxp67_ASAP7_75t_SL U30613 ( .A(n25045), .Y(n25030) );
  NAND2xp5_ASAP7_75t_SL U30614 ( .A(n29391), .B(n29279), .Y(n29282) );
  NAND2xp33_ASAP7_75t_SL U30615 ( .A(n25028), .B(n31582), .Y(n25029) );
  INVx1_ASAP7_75t_SL U30616 ( .A(n28424), .Y(n28637) );
  NAND2xp33_ASAP7_75t_SL U30617 ( .A(n26298), .B(n28982), .Y(n26294) );
  NAND2xp33_ASAP7_75t_SL U30618 ( .A(n26298), .B(n24578), .Y(n28843) );
  OAI21xp33_ASAP7_75t_SL U30619 ( .A1(n32075), .A2(n30709), .B(n29735), .Y(
        n2724) );
  AOI21xp33_ASAP7_75t_SL U30620 ( .A1(n30644), .A2(n29680), .B(n28812), .Y(
        n28813) );
  NAND2xp5_ASAP7_75t_SL U30621 ( .A(n26039), .B(n26043), .Y(n31075) );
  OAI21xp5_ASAP7_75t_SL U30622 ( .A1(n24791), .A2(n18838), .B(n24790), .Y(
        n30939) );
  NAND2xp5_ASAP7_75t_SL U30623 ( .A(n26039), .B(n26053), .Y(n31155) );
  AOI21xp33_ASAP7_75t_SL U30624 ( .A1(n30644), .A2(n29074), .B(n28510), .Y(
        n28511) );
  NAND2xp33_ASAP7_75t_SL U30625 ( .A(n26055), .B(n26066), .Y(n31071) );
  INVxp33_ASAP7_75t_SL U30626 ( .A(n29955), .Y(n26094) );
  INVxp67_ASAP7_75t_SL U30627 ( .A(n24786), .Y(n24787) );
  NAND2xp33_ASAP7_75t_SL U30628 ( .A(n3067), .B(n22396), .Y(n31304) );
  NAND2xp5_ASAP7_75t_SL U30629 ( .A(n26039), .B(n26066), .Y(n31083) );
  INVxp67_ASAP7_75t_SL U30630 ( .A(n28982), .Y(n26147) );
  NAND2xp33_ASAP7_75t_SL U30631 ( .A(n24684), .B(n32705), .Y(n32043) );
  NAND2xp33_ASAP7_75t_SL U30632 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[3]), .B(
        n31259), .Y(n31465) );
  NAND2xp33_ASAP7_75t_SL U30633 ( .A(n26068), .B(n26066), .Y(n31185) );
  OAI21xp33_ASAP7_75t_SL U30634 ( .A1(n31024), .A2(n31023), .B(n31022), .Y(
        n31025) );
  NAND2xp5_ASAP7_75t_SL U30635 ( .A(n25230), .B(n24987), .Y(n24984) );
  AOI22xp33_ASAP7_75t_SL U30636 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__WREG_), 
        .A2(n24648), .B1(u0_0_leon3x0_p0_iu_r_E__CTRL__WREG_), .B2(n32068), 
        .Y(n2710) );
  NAND2xp33_ASAP7_75t_SL U30637 ( .A(n26045), .B(n26060), .Y(n31095) );
  NAND2xp5_ASAP7_75t_SL U30638 ( .A(n26039), .B(n26060), .Y(n31115) );
  NAND2xp33_ASAP7_75t_SL U30639 ( .A(n26062), .B(n26043), .Y(n31135) );
  NAND2xp33_ASAP7_75t_SL U30640 ( .A(n26045), .B(n26066), .Y(n31079) );
  OAI22xp33_ASAP7_75t_SL U30641 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__10_), 
        .A2(n27143), .B1(n27142), .B2(n27141), .Y(n27154) );
  NAND2xp33_ASAP7_75t_SL U30642 ( .A(n26055), .B(n26043), .Y(n31123) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U30643 ( .A1(n32055), .A2(n32054), .B(n32053), 
        .C(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), .Y(n32056) );
  NAND2xp33_ASAP7_75t_SL U30644 ( .A(n26036), .B(n26043), .Y(n31107) );
  AOI21xp33_ASAP7_75t_SL U30645 ( .A1(n30644), .A2(n28529), .B(n28528), .Y(
        n28530) );
  NAND2xp33_ASAP7_75t_SL U30646 ( .A(apbi[11]), .B(n31198), .Y(n25943) );
  AOI21xp33_ASAP7_75t_SL U30647 ( .A1(n30644), .A2(n28554), .B(n28553), .Y(
        n28555) );
  NAND2xp33_ASAP7_75t_SL U30648 ( .A(add_x_735_A_2_), .B(n29146), .Y(n26363)
         );
  NAND2xp33_ASAP7_75t_SL U30649 ( .A(n23002), .B(n28982), .Y(n26254) );
  AOI21xp33_ASAP7_75t_SL U30650 ( .A1(n30644), .A2(n29778), .B(n28464), .Y(
        n28465) );
  OAI21xp33_ASAP7_75t_SL U30651 ( .A1(n29889), .A2(n32075), .B(n26138), .Y(
        n18051) );
  OAI21xp33_ASAP7_75t_SL U30652 ( .A1(n31396), .A2(n27166), .B(n27165), .Y(
        n27167) );
  INVx1_ASAP7_75t_SL U30653 ( .A(n28968), .Y(n28987) );
  NAND2xp33_ASAP7_75t_SL U30654 ( .A(n26032), .B(n26043), .Y(n31067) );
  INVx1_ASAP7_75t_SL U30655 ( .A(n31605), .Y(n31447) );
  NAND2xp33_ASAP7_75t_SL U30656 ( .A(n24634), .B(n28132), .Y(n28671) );
  NAND2xp33_ASAP7_75t_SL U30657 ( .A(n22968), .B(n24577), .Y(n25458) );
  NAND2xp33_ASAP7_75t_SL U30658 ( .A(n26062), .B(n26060), .Y(n31179) );
  NAND2xp33_ASAP7_75t_SL U30659 ( .A(n28425), .B(n28424), .Y(n28427) );
  NAND2xp33_ASAP7_75t_SL U30660 ( .A(n26068), .B(n26060), .Y(n31175) );
  AND2x2_ASAP7_75t_SL U30661 ( .A(n23365), .B(n24577), .Y(n23362) );
  INVxp67_ASAP7_75t_SL U30662 ( .A(n29985), .Y(n27499) );
  XNOR2xp5_ASAP7_75t_SL U30663 ( .A(n24055), .B(n23976), .Y(n23534) );
  NAND2xp33_ASAP7_75t_SL U30664 ( .A(n26049), .B(n26043), .Y(n31099) );
  NAND2xp5_ASAP7_75t_SL U30665 ( .A(n30204), .B(n25033), .Y(n25022) );
  OAI21xp33_ASAP7_75t_SL U30666 ( .A1(n24638), .A2(n30342), .B(n30341), .Y(
        n30343) );
  OAI22xp33_ASAP7_75t_SL U30667 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__16_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__26_), .Y(
        n28384) );
  INVx1_ASAP7_75t_SL U30668 ( .A(n32132), .Y(n32014) );
  OAI22xp33_ASAP7_75t_SL U30669 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__14_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__24_), .Y(
        n28462) );
  OAI21xp33_ASAP7_75t_SL U30670 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__10_), 
        .A2(n24651), .B(n28709), .Y(n3168) );
  OAI21xp33_ASAP7_75t_SL U30671 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__9_), 
        .A2(n22377), .B(n26215), .Y(n3420) );
  OAI21xp33_ASAP7_75t_SL U30672 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__WY_), .A2(
        n24654), .B(n25276), .Y(n3152) );
  NAND2xp5_ASAP7_75t_SL U30673 ( .A(n26097), .B(n27463), .Y(n30134) );
  NAND2xp33_ASAP7_75t_SL U30674 ( .A(n26062), .B(n26067), .Y(n31162) );
  INVxp33_ASAP7_75t_SL U30675 ( .A(timer0_v_TICK_), .Y(n33064) );
  OAI21xp33_ASAP7_75t_SL U30676 ( .A1(n24638), .A2(n30363), .B(n30362), .Y(
        n30364) );
  OAI21xp33_ASAP7_75t_SL U30677 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__WY_), .A2(
        n24655), .B(n25275), .Y(n3154) );
  OAI22xp33_ASAP7_75t_SL U30678 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__28_), .Y(
        n25939) );
  OAI21xp33_ASAP7_75t_SL U30679 ( .A1(n28509), .A2(n30642), .B(n28508), .Y(
        n28510) );
  INVxp33_ASAP7_75t_SL U30680 ( .A(n29499), .Y(n29482) );
  OAI21xp33_ASAP7_75t_SL U30681 ( .A1(u0_0_leon3x0_p0_ici[48]), .A2(n24649), 
        .B(n26976), .Y(n2529) );
  INVxp33_ASAP7_75t_SL U30682 ( .A(n28805), .Y(n26287) );
  INVxp67_ASAP7_75t_SL U30683 ( .A(n29012), .Y(n31395) );
  OAI21xp33_ASAP7_75t_SL U30684 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__20_), 
        .A2(n24649), .B(n26978), .Y(n2527) );
  OAI21xp5_ASAP7_75t_SL U30685 ( .A1(ahb0_r_HADDR__3_), .A2(n17288), .B(n25413), .Y(n31019) );
  OAI21xp33_ASAP7_75t_SL U30686 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__20_), 
        .A2(n24650), .B(n26980), .Y(n2525) );
  OAI21xp33_ASAP7_75t_SL U30687 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__19_), 
        .A2(n24658), .B(n24702), .Y(n3600) );
  OAI21xp33_ASAP7_75t_SL U30688 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__20_), 
        .A2(n24650), .B(n26982), .Y(n2523) );
  OAI21xp33_ASAP7_75t_SL U30689 ( .A1(n27009), .A2(n30642), .B(n27008), .Y(
        n27010) );
  OAI21xp33_ASAP7_75t_SL U30690 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__WY_), .A2(
        n24657), .B(n31390), .Y(n3156) );
  NAND2xp5_ASAP7_75t_SL U30691 ( .A(n28373), .B(n23102), .Y(n28375) );
  OAI21xp33_ASAP7_75t_SL U30692 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), 
        .A2(n24654), .B(n31538), .Y(n4179) );
  OAI21xp33_ASAP7_75t_SL U30693 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__0_), 
        .A2(n24649), .B(n29232), .Y(n3340) );
  AOI21xp33_ASAP7_75t_SL U30694 ( .A1(n28018), .A2(uart1_r_THOLD__30__1_), .B(
        n27416), .Y(n27420) );
  NAND2xp33_ASAP7_75t_SL U30695 ( .A(n31336), .B(n29899), .Y(n29900) );
  OAI22xp33_ASAP7_75t_SL U30696 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__27_), .Y(
        n26348) );
  OAI21xp33_ASAP7_75t_SL U30697 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__18_), 
        .A2(n24656), .B(n25730), .Y(n2574) );
  INVx1_ASAP7_75t_SL U30698 ( .A(n29987), .Y(n27524) );
  OAI21xp33_ASAP7_75t_SL U30699 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__18_), 
        .A2(n24656), .B(n25728), .Y(n2576) );
  OAI21xp33_ASAP7_75t_SL U30700 ( .A1(u0_0_leon3x0_p0_ici[55]), .A2(n22377), 
        .B(n26880), .Y(n3396) );
  AND4x1_ASAP7_75t_SL U30701 ( .A(n27432), .B(n27431), .C(n27430), .D(n27429), 
        .Y(n27433) );
  NAND2xp5_ASAP7_75t_SL U30702 ( .A(n25243), .B(n31020), .Y(n4643) );
  OAI21xp33_ASAP7_75t_SL U30703 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__18_), 
        .A2(n24656), .B(n25726), .Y(n2578) );
  OAI21xp33_ASAP7_75t_SL U30704 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__27_), 
        .A2(n22377), .B(n26882), .Y(n3394) );
  OAI21xp33_ASAP7_75t_SL U30705 ( .A1(u0_0_leon3x0_p0_ici[46]), .A2(n24656), 
        .B(n25720), .Y(n2580) );
  OAI21xp33_ASAP7_75t_SL U30706 ( .A1(n27129), .A2(n30642), .B(n27128), .Y(
        n27130) );
  OAI21xp33_ASAP7_75t_SL U30707 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__27_), 
        .A2(n22377), .B(n26884), .Y(n3392) );
  NAND2xp33_ASAP7_75t_SL U30708 ( .A(n30120), .B(n30878), .Y(n30121) );
  OAI21xp33_ASAP7_75t_SL U30709 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__27_), 
        .A2(n22377), .B(n26886), .Y(n3390) );
  NAND2xp33_ASAP7_75t_SL U30710 ( .A(n25731), .B(n32075), .Y(n25710) );
  NAND2xp5_ASAP7_75t_SL U30711 ( .A(u0_0_leon3x0_p0_iu_r_M__NALIGN_), .B(
        n29721), .Y(n29474) );
  NAND2xp5_ASAP7_75t_SL U30712 ( .A(n31336), .B(n28574), .Y(n30491) );
  OAI21xp33_ASAP7_75t_SL U30713 ( .A1(n30730), .A2(n30642), .B(n28750), .Y(
        n28751) );
  AOI22xp33_ASAP7_75t_SL U30714 ( .A1(u0_0_leon3x0_p0_iu_r_X__NERROR_), .A2(
        n24648), .B1(n33057), .B2(n33056), .Y(n3376) );
  OAI21xp33_ASAP7_75t_SL U30715 ( .A1(u0_0_leon3x0_p0_iu_v_M__IRQEN2_), .A2(
        n24658), .B(n30693), .Y(n3383) );
  OAI21xp33_ASAP7_75t_SL U30716 ( .A1(n31584), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DCS__1_), .B(n30915), .Y(n31600) );
  NAND2xp33_ASAP7_75t_SL U30717 ( .A(n28830), .B(u0_0_leon3x0_p0_divi[0]), .Y(
        n26743) );
  NAND2xp33_ASAP7_75t_SL U30718 ( .A(n31336), .B(n29837), .Y(n29838) );
  OAI21xp33_ASAP7_75t_SL U30719 ( .A1(n28527), .A2(n30642), .B(n28526), .Y(
        n28528) );
  OAI22xp33_ASAP7_75t_SL U30720 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__23_), .Y(
        n28471) );
  OAI21xp33_ASAP7_75t_SL U30721 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__19_), 
        .A2(n24657), .B(n25752), .Y(n2546) );
  OAI21xp33_ASAP7_75t_SL U30722 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__19_), 
        .A2(n24657), .B(n25750), .Y(n2548) );
  OAI21xp33_ASAP7_75t_SL U30723 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__19_), 
        .A2(n24657), .B(n25748), .Y(n2550) );
  OAI21xp33_ASAP7_75t_SL U30724 ( .A1(u0_0_leon3x0_p0_ici[47]), .A2(n24656), 
        .B(n25746), .Y(n2552) );
  INVxp67_ASAP7_75t_SL U30725 ( .A(n26014), .Y(n25979) );
  NAND2xp33_ASAP7_75t_SL U30726 ( .A(n26068), .B(n26054), .Y(n31058) );
  INVxp33_ASAP7_75t_SL U30727 ( .A(n29831), .Y(n29832) );
  OAI21xp33_ASAP7_75t_SL U30728 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__2_), 
        .A2(n24656), .B(n25708), .Y(n3352) );
  NAND2xp5_ASAP7_75t_SL U30729 ( .A(n27641), .B(n27640), .Y(n27646) );
  OAI22xp33_ASAP7_75t_SL U30730 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__10_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__20_), .Y(
        n26970) );
  OAI22xp33_ASAP7_75t_SL U30731 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__9_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__19_), .Y(
        n28525) );
  OAI21xp33_ASAP7_75t_SL U30732 ( .A1(u0_0_leon3x0_p0_iu_v_E__SU_), .A2(n22377), .B(n30798), .Y(n3360) );
  OAI21xp33_ASAP7_75t_SL U30733 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__25_), 
        .A2(n24652), .B(n28418), .Y(n3404) );
  NAND2xp5_ASAP7_75t_SL U30734 ( .A(n25004), .B(n25003), .Y(n26812) );
  AOI21xp33_ASAP7_75t_SL U30735 ( .A1(n28018), .A2(uart1_r_THOLD__28__1_), .B(
        n27406), .Y(n27415) );
  OAI21xp33_ASAP7_75t_SL U30736 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__25_), 
        .A2(n24652), .B(n28454), .Y(n3402) );
  OAI21xp33_ASAP7_75t_SL U30737 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__25_), 
        .A2(n24652), .B(n28456), .Y(n3400) );
  NAND2xp33_ASAP7_75t_SL U30738 ( .A(n26055), .B(n26044), .Y(n31122) );
  OAI21xp33_ASAP7_75t_SL U30739 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__LD_), .A2(
        n24654), .B(n31867), .Y(n3514) );
  NAND2xp33_ASAP7_75t_SL U30740 ( .A(n31336), .B(n31335), .Y(n31337) );
  NAND2xp33_ASAP7_75t_SL U30741 ( .A(n26055), .B(n26061), .Y(n31146) );
  OAI21xp33_ASAP7_75t_SL U30742 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__LD_), .A2(
        n24654), .B(n31865), .Y(n3516) );
  OAI21xp33_ASAP7_75t_SL U30743 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__3_), 
        .A2(n22377), .B(n26839), .Y(n3478) );
  OAI21xp33_ASAP7_75t_SL U30744 ( .A1(u0_0_leon3x0_p0_ici[51]), .A2(n24652), 
        .B(n29038), .Y(n3248) );
  OAI21xp33_ASAP7_75t_SL U30745 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__3_), 
        .A2(n24655), .B(n31521), .Y(n3476) );
  NAND2xp33_ASAP7_75t_SL U30746 ( .A(n26032), .B(n26044), .Y(n31066) );
  O2A1O1Ixp33_ASAP7_75t_SL U30747 ( .A1(n25575), .A2(n30196), .B(n25027), .C(
        n25026), .Y(n25045) );
  NAND2xp33_ASAP7_75t_SL U30748 ( .A(n26062), .B(n26061), .Y(n31178) );
  OAI21xp33_ASAP7_75t_SL U30749 ( .A1(irqctrl0_r_ILEVEL__3_), .A2(n29415), .B(
        n29636), .Y(n29406) );
  OAI21xp33_ASAP7_75t_SL U30750 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__LD_), .B(n31863), .Y(n3518) );
  NAND2xp33_ASAP7_75t_SL U30751 ( .A(n26036), .B(n26044), .Y(n31106) );
  NAND2xp33_ASAP7_75t_SL U30752 ( .A(n26049), .B(n26044), .Y(n31098) );
  NAND2xp33_ASAP7_75t_SL U30753 ( .A(n26062), .B(n26044), .Y(n31134) );
  OAI21xp33_ASAP7_75t_SL U30754 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__6_), 
        .A2(n24655), .B(n31519), .Y(n4006) );
  NAND2xp33_ASAP7_75t_SL U30755 ( .A(n26068), .B(n26061), .Y(n31174) );
  OAI22xp33_ASAP7_75t_SL U30756 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), 
        .A2(n24495), .B1(n23229), .B2(u0_0_leon3x0_p0_iu_r_A__IMM__29_), .Y(
        n29862) );
  NAND2xp33_ASAP7_75t_SL U30757 ( .A(n26045), .B(n26054), .Y(n31130) );
  OAI21xp33_ASAP7_75t_SL U30758 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_), 
        .A2(n22377), .B(n24700), .Y(n4107) );
  AOI22xp33_ASAP7_75t_SL U30759 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__4_), .A2(
        n24648), .B1(n30813), .B2(DP_OP_1196_128_7433_n456), .Y(n3522) );
  INVx1_ASAP7_75t_SL U30760 ( .A(DP_OP_1196_128_7433_n233), .Y(
        DP_OP_1196_128_7433_n235) );
  OAI21xp33_ASAP7_75t_SL U30761 ( .A1(n28538), .A2(n30642), .B(n28537), .Y(
        n28539) );
  NAND2xp33_ASAP7_75t_SL U30762 ( .A(n26045), .B(n26044), .Y(n31158) );
  INVx1_ASAP7_75t_SL U30763 ( .A(n26308), .Y(n30611) );
  INVx1_ASAP7_75t_SL U30764 ( .A(DP_OP_1196_128_7433_n232), .Y(
        DP_OP_1196_128_7433_n234) );
  INVxp33_ASAP7_75t_SL U30765 ( .A(n24753), .Y(n24754) );
  NAND2xp5_ASAP7_75t_SL U30766 ( .A(n26039), .B(n26044), .Y(n31074) );
  NAND2xp33_ASAP7_75t_SL U30767 ( .A(n26049), .B(n26054), .Y(n31166) );
  OAI21xp33_ASAP7_75t_SL U30768 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__23_), 
        .A2(n24654), .B(n31983), .Y(n4103) );
  INVx4_ASAP7_75t_SL U30769 ( .A(n22216), .Y(n23966) );
  AND2x2_ASAP7_75t_SL U30770 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WY_), .B(
        n32161), .Y(n31402) );
  NAND2xp5_ASAP7_75t_SL U30771 ( .A(n26039), .B(n26054), .Y(n31154) );
  INVx1_ASAP7_75t_SL U30772 ( .A(n29637), .Y(n29880) );
  OAI21xp33_ASAP7_75t_SL U30773 ( .A1(u0_0_leon3x0_p0_ici[49]), .A2(n24649), 
        .B(n27046), .Y(n3236) );
  OAI21xp33_ASAP7_75t_SL U30774 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__21_), 
        .A2(n24649), .B(n27050), .Y(n3232) );
  OAI21xp33_ASAP7_75t_SL U30775 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__0_), 
        .A2(n24658), .B(n26830), .Y(n3530) );
  OAI21xp33_ASAP7_75t_SL U30776 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__21_), 
        .A2(n24649), .B(n27052), .Y(n3230) );
  INVxp33_ASAP7_75t_SL U30777 ( .A(n24783), .Y(n24784) );
  NAND2xp33_ASAP7_75t_SL U30778 ( .A(n26055), .B(n26067), .Y(n31070) );
  AOI21xp33_ASAP7_75t_SL U30779 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__28_), 
        .A2(n24647), .B(n26809), .Y(n3490) );
  OAI21xp33_ASAP7_75t_SL U30780 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__31_), 
        .A2(n22377), .B(n26722), .Y(n4151) );
  NAND2xp33_ASAP7_75t_SL U30781 ( .A(n26032), .B(n26067), .Y(n31142) );
  OAI21xp33_ASAP7_75t_SL U30782 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__2_), 
        .A2(n24655), .B(n31520), .Y(n3493) );
  NAND2xp33_ASAP7_75t_SL U30783 ( .A(n26036), .B(n26067), .Y(n31138) );
  OAI21xp33_ASAP7_75t_SL U30784 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__28_), 
        .A2(n24655), .B(n25546), .Y(n3486) );
  AOI22xp33_ASAP7_75t_SL U30785 ( .A1(irqctrl0_r_IMASK__0__14_), .A2(n31249), 
        .B1(irqctrl0_r_IFORCE__0__14_), .B2(n31251), .Y(n30550) );
  NAND2xp33_ASAP7_75t_SL U30786 ( .A(n26068), .B(n26067), .Y(n31183) );
  NAND2xp33_ASAP7_75t_SL U30787 ( .A(n26049), .B(n26067), .Y(n31126) );
  OAI21xp33_ASAP7_75t_SL U30788 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__28_), 
        .A2(n24655), .B(n25548), .Y(n3484) );
  OAI21xp33_ASAP7_75t_SL U30789 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__2_), 
        .A2(n24658), .B(n26836), .Y(n3495) );
  NOR4xp25_ASAP7_75t_SRAM U30790 ( .A(n25559), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__26_), .C(n30351), .D(n25558), .Y(
        n25560) );
  OAI21xp33_ASAP7_75t_SL U30791 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), 
        .A2(n22377), .B(n24954), .Y(n4155) );
  NAND2xp33_ASAP7_75t_SL U30792 ( .A(n31336), .B(n28586), .Y(n27219) );
  OAI21xp33_ASAP7_75t_SL U30793 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__2_), 
        .A2(n24658), .B(n26834), .Y(n3497) );
  NAND2xp33_ASAP7_75t_SL U30794 ( .A(n26045), .B(n26061), .Y(n31094) );
  NAND2xp33_ASAP7_75t_SL U30795 ( .A(n26049), .B(n26061), .Y(n31086) );
  NAND2xp33_ASAP7_75t_SL U30796 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__16_), 
        .B(n24796), .Y(n24795) );
  NAND2xp33_ASAP7_75t_SL U30797 ( .A(n26045), .B(n26067), .Y(n31078) );
  OAI21xp33_ASAP7_75t_SL U30798 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__27_), 
        .A2(n24655), .B(n25552), .Y(n3503) );
  INVxp33_ASAP7_75t_SL U30799 ( .A(DP_OP_1196_128_7433_n84), .Y(
        DP_OP_1196_128_7433_n86) );
  NOR2x1_ASAP7_75t_SL U30800 ( .A(n25086), .B(n28880), .Y(n26298) );
  NAND2xp5_ASAP7_75t_SL U30801 ( .A(n26039), .B(n26067), .Y(n31082) );
  INVxp33_ASAP7_75t_SL U30802 ( .A(DP_OP_1196_128_7433_n85), .Y(
        DP_OP_1196_128_7433_n87) );
  INVxp67_ASAP7_75t_SL U30803 ( .A(n24808), .Y(n24773) );
  NAND2xp33_ASAP7_75t_SL U30804 ( .A(n26036), .B(n26061), .Y(n31118) );
  OAI21xp33_ASAP7_75t_SL U30805 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__29_), 
        .A2(n24650), .B(n29578), .Y(n3282) );
  OAI21xp33_ASAP7_75t_SL U30806 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__0_), 
        .A2(n22377), .B(n24955), .Y(n4163) );
  OAI21xp33_ASAP7_75t_SL U30807 ( .A1(n31396), .A2(n26734), .B(n25211), .Y(
        n25212) );
  OAI21xp33_ASAP7_75t_SL U30808 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__27_), 
        .A2(n24655), .B(n25550), .Y(n3507) );
  NAND2xp33_ASAP7_75t_SL U30809 ( .A(n26068), .B(n26044), .Y(n31062) );
  NAND2xp33_ASAP7_75t_SL U30810 ( .A(n26032), .B(n26061), .Y(n31090) );
  OAI21xp33_ASAP7_75t_SL U30811 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), 
        .A2(n24654), .B(n31820), .Y(n4165) );
  OAI21xp33_ASAP7_75t_SL U30812 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__3_), 
        .A2(n24658), .B(n26838), .Y(n3480) );
  AOI21xp33_ASAP7_75t_SL U30813 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__27_), 
        .A2(n24647), .B(n26825), .Y(n3509) );
  INVx1_ASAP7_75t_SL U30814 ( .A(n32075), .Y(n29738) );
  OAI21xp33_ASAP7_75t_SL U30815 ( .A1(u0_0_leon3x0_p0_ici[58]), .A2(n24657), 
        .B(n25888), .Y(n2380) );
  NAND2xp33_ASAP7_75t_SL U30816 ( .A(n31336), .B(n27027), .Y(n27028) );
  OAI21xp33_ASAP7_75t_SL U30817 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), 
        .A2(n24655), .B(n32011), .Y(n3606) );
  OAI21xp33_ASAP7_75t_SL U30818 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__8_), 
        .A2(n22377), .B(n30716), .Y(n3434) );
  NAND2xp33_ASAP7_75t_SL U30819 ( .A(n28946), .B(n22375), .Y(n28947) );
  OAI21xp33_ASAP7_75t_SL U30820 ( .A1(n29782), .A2(n30642), .B(n28463), .Y(
        n28464) );
  INVxp33_ASAP7_75t_SL U30821 ( .A(u0_0_leon3x0_p0_divi[1]), .Y(n28940) );
  OAI21xp33_ASAP7_75t_SL U30822 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__8_), 
        .A2(n24658), .B(n30718), .Y(n3432) );
  NAND2xp33_ASAP7_75t_SL U30823 ( .A(n31336), .B(n29680), .Y(n29685) );
  NAND2xp5_ASAP7_75t_SL U30824 ( .A(n31751), .B(n32790), .Y(n32749) );
  INVxp67_ASAP7_75t_SL U30825 ( .A(n27462), .Y(n25636) );
  INVxp33_ASAP7_75t_SL U30826 ( .A(n30465), .Y(n30467) );
  OAI21xp33_ASAP7_75t_SL U30827 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__8_), 
        .A2(n24658), .B(n30720), .Y(n3430) );
  OAI21xp33_ASAP7_75t_SL U30828 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__3_), 
        .A2(n24651), .B(n29487), .Y(n3182) );
  OAI21xp33_ASAP7_75t_SL U30829 ( .A1(n28572), .A2(n30642), .B(n28571), .Y(
        n28573) );
  OAI21xp33_ASAP7_75t_SL U30830 ( .A1(u0_0_leon3x0_p0_dci[4]), .A2(n24657), 
        .B(n24969), .Y(n3582) );
  OAI21xp33_ASAP7_75t_SL U30831 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__30_), 
        .A2(n24650), .B(n30582), .Y(n2378) );
  OAI21xp33_ASAP7_75t_SL U30832 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__3_), 
        .A2(n24650), .B(n29489), .Y(n3180) );
  OAI21xp33_ASAP7_75t_SL U30833 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_), 
        .A2(n22377), .B(n24959), .Y(n4105) );
  NAND2xp33_ASAP7_75t_SL U30834 ( .A(n22939), .B(n29146), .Y(n28925) );
  NAND2xp33_ASAP7_75t_SL U30835 ( .A(n28232), .B(n27462), .Y(n31023) );
  NAND2xp33_ASAP7_75t_SL U30836 ( .A(n29646), .B(n32075), .Y(n29647) );
  OAI21xp33_ASAP7_75t_SL U30837 ( .A1(u0_0_leon3x0_p0_ici[37]), .A2(n22377), 
        .B(n26209), .Y(n3426) );
  NAND2xp33_ASAP7_75t_SL U30838 ( .A(n32133), .B(n32132), .Y(n32134) );
  INVx1_ASAP7_75t_SL U30839 ( .A(n32050), .Y(n24912) );
  OAI21xp33_ASAP7_75t_SL U30840 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__9_), 
        .A2(n22377), .B(n26211), .Y(n3424) );
  OAI21xp33_ASAP7_75t_SL U30841 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__30_), 
        .A2(n24650), .B(n30584), .Y(n2376) );
  INVxp33_ASAP7_75t_SL U30842 ( .A(n29737), .Y(n29740) );
  NAND2xp5_ASAP7_75t_SL U30843 ( .A(n25846), .B(n27463), .Y(n26467) );
  NAND2xp33_ASAP7_75t_SL U30844 ( .A(n32018), .B(n32017), .Y(n32019) );
  OAI21xp33_ASAP7_75t_SL U30845 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__9_), 
        .A2(n22377), .B(n26213), .Y(n3422) );
  OAI21xp33_ASAP7_75t_SL U30846 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__10_), 
        .A2(n24653), .B(n28707), .Y(n3170) );
  OAI21xp33_ASAP7_75t_SL U30847 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__30_), 
        .A2(n24650), .B(n30586), .Y(n2374) );
  OAI21xp33_ASAP7_75t_SL U30848 ( .A1(u0_0_leon3x0_p0_dci[5]), .A2(n24657), 
        .B(n24973), .Y(n3588) );
  NAND2xp33_ASAP7_75t_SL U30849 ( .A(n26036), .B(n26054), .Y(n31150) );
  OAI21xp33_ASAP7_75t_SL U30850 ( .A1(n24995), .A2(n24928), .B(n24927), .Y(
        n24935) );
  NAND2xp5_ASAP7_75t_SL U30851 ( .A(n26039), .B(n26061), .Y(n31114) );
  INVxp67_ASAP7_75t_SL U30852 ( .A(n28602), .Y(n27189) );
  NAND2xp33_ASAP7_75t_SL U30853 ( .A(n25955), .B(n25963), .Y(n27292) );
  INVxp67_ASAP7_75t_SL U30854 ( .A(n29635), .Y(n29877) );
  NAND2xp33_ASAP7_75t_SL U30855 ( .A(n31336), .B(n27275), .Y(n26716) );
  NAND2xp5_ASAP7_75t_SL U30856 ( .A(n28769), .B(n29144), .Y(n27143) );
  NAND2xp33_ASAP7_75t_SL U30857 ( .A(n26032), .B(n26054), .Y(n31102) );
  NAND2xp33_ASAP7_75t_SL U30858 ( .A(n26097), .B(n31251), .Y(n27291) );
  NAND2xp5_ASAP7_75t_SL U30859 ( .A(n25639), .B(n31249), .Y(n29384) );
  NAND2xp5_ASAP7_75t_SL U30860 ( .A(n25962), .B(n25963), .Y(n29743) );
  INVxp67_ASAP7_75t_SL U30861 ( .A(n28521), .Y(n27086) );
  NAND2xp33_ASAP7_75t_SL U30862 ( .A(n26055), .B(n26054), .Y(n31170) );
  OAI21xp33_ASAP7_75t_SL U30863 ( .A1(n24638), .A2(n30309), .B(n30308), .Y(
        n30310) );
  OAI21xp33_ASAP7_75t_SL U30864 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__24_), 
        .A2(n24653), .B(n29777), .Y(n2469) );
  OAI21xp33_ASAP7_75t_SL U30865 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__28_), 
        .A2(n24654), .B(n25456), .Y(n3488) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U30866 ( .A1(n30955), .A2(n24940), .B(n24986), .C(
        n25668), .Y(n24941) );
  OAI21xp33_ASAP7_75t_SL U30867 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__31_), 
        .A2(n22377), .B(n26724), .Y(n4095) );
  OAI21xp33_ASAP7_75t_SL U30868 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__24_), 
        .A2(n24653), .B(n29775), .Y(n2471) );
  NAND2xp33_ASAP7_75t_SL U30869 ( .A(n26062), .B(n26054), .Y(n31110) );
  OAI21xp33_ASAP7_75t_SL U30870 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__24_), 
        .A2(n24653), .B(n29766), .Y(n2473) );
  OAI21xp33_ASAP7_75t_SL U30871 ( .A1(u0_0_leon3x0_p0_ici[42]), .A2(n24649), 
        .B(n27180), .Y(n3212) );
  NAND2xp5_ASAP7_75t_SL U30872 ( .A(n31667), .B(n31674), .Y(n31422) );
  NAND2xp33_ASAP7_75t_SL U30873 ( .A(n30677), .B(n29884), .Y(n29727) );
  OAI21xp33_ASAP7_75t_SL U30874 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), 
        .A2(n24656), .B(n32013), .Y(n3604) );
  OAI21xp33_ASAP7_75t_SL U30875 ( .A1(n24638), .A2(n30399), .B(n30398), .Y(
        n30400) );
  NAND2xp33_ASAP7_75t_SL U30876 ( .A(u0_0_leon3x0_p0_iu_r_W__S__WIM__6_), .B(
        n29198), .Y(n29193) );
  OAI21xp33_ASAP7_75t_SL U30877 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_), 
        .A2(n24658), .B(n24704), .Y(n3862) );
  NAND2xp5_ASAP7_75t_SL U30878 ( .A(n26803), .B(n26782), .Y(n29195) );
  OAI21xp33_ASAP7_75t_SL U30879 ( .A1(n29898), .A2(n30642), .B(n28795), .Y(
        n28796) );
  AOI21xp33_ASAP7_75t_SL U30880 ( .A1(n29359), .A2(n29344), .B(n29342), .Y(
        n29343) );
  OAI21xp33_ASAP7_75t_SL U30881 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__31_), 
        .A2(n22377), .B(n26374), .Y(n4328) );
  NAND2xp5_ASAP7_75t_SL U30882 ( .A(n32909), .B(n32839), .Y(n32856) );
  OAI21xp33_ASAP7_75t_SL U30883 ( .A1(u0_0_leon3x0_p0_muli[8]), .A2(n22377), 
        .B(n24960), .Y(n3860) );
  INVx1_ASAP7_75t_SL U30884 ( .A(n32044), .Y(n32122) );
  OAI21xp33_ASAP7_75t_SL U30885 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_), 
        .A2(n24654), .B(n31985), .Y(n3858) );
  AOI22xp33_ASAP7_75t_SL U30886 ( .A1(ahbso_0__HRDATA__23_), .A2(n32904), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[27]), .B2(n32903), .Y(n32978) );
  NAND2xp33_ASAP7_75t_SL U30887 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[16]), .B(
        n32871), .Y(n32865) );
  OAI21xp33_ASAP7_75t_SL U30888 ( .A1(u0_0_leon3x0_p0_ici[40]), .A2(n24652), 
        .B(n29050), .Y(n2673) );
  INVx1_ASAP7_75t_SL U30889 ( .A(n32839), .Y(n32854) );
  NAND2xp33_ASAP7_75t_SL U30890 ( .A(n29196), .B(n29198), .Y(n29197) );
  INVxp67_ASAP7_75t_SL U30891 ( .A(n28714), .Y(n27166) );
  OAI21xp33_ASAP7_75t_SL U30892 ( .A1(n28482), .A2(n28995), .B(n24634), .Y(
        n29591) );
  NAND2xp33_ASAP7_75t_SL U30893 ( .A(n29307), .B(n32075), .Y(n26138) );
  OAI21xp33_ASAP7_75t_SL U30894 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__12_), 
        .A2(n24653), .B(n29826), .Y(n2671) );
  OAI21xp33_ASAP7_75t_SL U30895 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__6_), 
        .A2(n22377), .B(n26248), .Y(n3934) );
  NAND2xp5_ASAP7_75t_SL U30896 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__19_), .B(
        n28769), .Y(n25772) );
  OR3x1_ASAP7_75t_SRAM U30897 ( .A(n25608), .B(n33054), .C(n33055), .Y(n25609)
         );
  OAI21xp33_ASAP7_75t_SL U30898 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__12_), 
        .A2(n24653), .B(n29828), .Y(n2669) );
  OAI21xp33_ASAP7_75t_SL U30899 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__6_), 
        .A2(n22377), .B(n26246), .Y(n3936) );
  OAI21xp33_ASAP7_75t_SL U30900 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__12_), 
        .A2(n24653), .B(n29830), .Y(n2667) );
  AOI22xp33_ASAP7_75t_SL U30901 ( .A1(u0_0_leon3x0_p0_dci[41]), .A2(n24648), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__9_), .B2(n30878), .Y(n3653) );
  OAI21xp33_ASAP7_75t_SL U30902 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__6_), 
        .A2(n22377), .B(n26244), .Y(n3938) );
  OAI21xp33_ASAP7_75t_SL U30903 ( .A1(u0_0_leon3x0_p0_ici[34]), .A2(n22377), 
        .B(n26242), .Y(n3940) );
  NAND2xp33_ASAP7_75t_SL U30904 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[17]), .B(
        n32871), .Y(n32867) );
  AOI21xp5_ASAP7_75t_SL U30905 ( .A1(n31560), .A2(n32591), .B(n31562), .Y(
        n31561) );
  INVx1_ASAP7_75t_SL U30906 ( .A(add_x_735_A_9_), .Y(n28725) );
  INVx1_ASAP7_75t_SL U30907 ( .A(n31412), .Y(n30394) );
  NAND2xp33_ASAP7_75t_SL U30908 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[18]), .B(
        n32871), .Y(n32869) );
  INVxp67_ASAP7_75t_SL U30909 ( .A(DP_OP_1196_128_7433_n263), .Y(
        DP_OP_1196_128_7433_n261) );
  INVxp67_ASAP7_75t_SL U30910 ( .A(DP_OP_1196_128_7433_n262), .Y(
        DP_OP_1196_128_7433_n260) );
  OAI21xp33_ASAP7_75t_SL U30911 ( .A1(n24638), .A2(n30279), .B(n30278), .Y(
        n30280) );
  INVxp33_ASAP7_75t_SL U30912 ( .A(n30813), .Y(n28701) );
  OAI21xp33_ASAP7_75t_SL U30913 ( .A1(n29684), .A2(n30642), .B(n28811), .Y(
        n28812) );
  AOI21xp33_ASAP7_75t_SL U30914 ( .A1(n18867), .A2(n32094), .B(n32093), .Y(
        n32096) );
  AOI22xp33_ASAP7_75t_SL U30915 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__5_), .A2(
        n24648), .B1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__5_), .B2(n30813), .Y(
        n3687) );
  AOI21xp33_ASAP7_75t_SL U30916 ( .A1(uart1_r_DPAR_), .A2(n27533), .B(n27532), 
        .Y(n2859) );
  OAI21xp33_ASAP7_75t_SL U30917 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__WREG_), 
        .A2(n24658), .B(n24953), .Y(n2708) );
  OAI21xp33_ASAP7_75t_SL U30918 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__6_), 
        .A2(n22377), .B(n31255), .Y(n3684) );
  NAND2xp5_ASAP7_75t_SL U30919 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__1_), 
        .B(n30163), .Y(n30169) );
  OAI21xp33_ASAP7_75t_SL U30920 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__7_), 
        .A2(n24656), .B(n31513), .Y(n2716) );
  INVxp67_ASAP7_75t_SL U30921 ( .A(n26226), .Y(n25509) );
  OAI21xp33_ASAP7_75t_SL U30922 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__29_), 
        .A2(n24655), .B(n25544), .Y(n3743) );
  NOR2xp33_ASAP7_75t_SL U30923 ( .A(n22906), .B(n29148), .Y(n26922) );
  OAI21xp33_ASAP7_75t_SL U30924 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__7_), 
        .A2(n24658), .B(n26841), .Y(n2718) );
  OAI21xp33_ASAP7_75t_SL U30925 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__7_), 
        .A2(n24656), .B(n31512), .Y(n2720) );
  INVx1_ASAP7_75t_SL U30926 ( .A(n29342), .Y(n29350) );
  INVxp67_ASAP7_75t_SL U30927 ( .A(n30878), .Y(n31256) );
  OAI21xp33_ASAP7_75t_SL U30928 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__29_), 
        .A2(n24657), .B(n32064), .Y(n3745) );
  NAND2xp33_ASAP7_75t_SL U30929 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[13]), .B(
        n32871), .Y(n32858) );
  OAI21xp33_ASAP7_75t_SL U30930 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_), 
        .A2(n24655), .B(n25235), .Y(n3871) );
  OAI21xp33_ASAP7_75t_SL U30931 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__7_), .B(n31510), .Y(n2722) );
  NAND2xp33_ASAP7_75t_SL U30932 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[14]), .B(
        n32871), .Y(n32861) );
  NAND2xp33_ASAP7_75t_SL U30933 ( .A(n31336), .B(n28529), .Y(n25806) );
  NAND2xp33_ASAP7_75t_SL U30934 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__6_), .B(
        n28769), .Y(n26261) );
  OAI21xp33_ASAP7_75t_SL U30935 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__1_), 
        .A2(n24656), .B(n31517), .Y(n3750) );
  OAI211xp5_ASAP7_75t_SRAM U30936 ( .A1(n3055), .A2(n30185), .B(n24684), .C(
        n30184), .Y(n30188) );
  INVxp67_ASAP7_75t_SL U30937 ( .A(n28540), .Y(n25809) );
  NAND2xp33_ASAP7_75t_SL U30938 ( .A(u0_0_leon3x0_p0_iu_r_W__S__WIM__7_), .B(
        n29198), .Y(n29183) );
  INVx1_ASAP7_75t_SL U30939 ( .A(n23002), .Y(n22418) );
  OAI21xp33_ASAP7_75t_SL U30940 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__1_), 
        .A2(n24658), .B(n26832), .Y(n3752) );
  INVx1_ASAP7_75t_SL U30941 ( .A(n28759), .Y(n30877) );
  INVxp67_ASAP7_75t_SL U30942 ( .A(n29796), .Y(n29798) );
  NAND2xp5_ASAP7_75t_SL U30943 ( .A(n31296), .B(n31301), .Y(n32284) );
  OAI21xp33_ASAP7_75t_SL U30944 ( .A1(n24638), .A2(n30409), .B(n30408), .Y(
        n30410) );
  INVx1_ASAP7_75t_SL U30945 ( .A(u0_0_leon3x0_p0_muli[41]), .Y(n28829) );
  AOI22xp33_ASAP7_75t_SL U30946 ( .A1(u0_0_leon3x0_p0_dci[39]), .A2(n24648), 
        .B1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__7_), .B2(n30878), .Y(n3671) );
  INVxp33_ASAP7_75t_SL U30947 ( .A(n32076), .Y(n25610) );
  OAI21xp33_ASAP7_75t_SL U30948 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), 
        .A2(n24658), .B(n24703), .Y(n3864) );
  AND2x2_ASAP7_75t_SL U30949 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__28_), .B(
        n28769), .Y(n26920) );
  NAND2xp33_ASAP7_75t_SL U30950 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[15]), .B(
        n32871), .Y(n32863) );
  AOI22xp33_ASAP7_75t_SL U30951 ( .A1(ahbso_0__HRDATA__16_), .A2(n32904), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[20]), .B2(n32903), .Y(n32919) );
  OAI21xp33_ASAP7_75t_SL U30952 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__5_), 
        .A2(n22377), .B(n26843), .Y(n2794) );
  OAI21xp33_ASAP7_75t_SL U30953 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__30_), 
        .A2(n22377), .B(n24958), .Y(n3889) );
  AOI22xp33_ASAP7_75t_SL U30954 ( .A1(ahbso_0__HRDATA__21_), .A2(n32904), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[25]), .B2(n32903), .Y(n32959) );
  AOI22xp33_ASAP7_75t_SL U30955 ( .A1(ahbso_0__HRDATA__19_), .A2(n32904), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[23]), .B2(n32903), .Y(n32943) );
  NAND2xp33_ASAP7_75t_SL U30956 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__12_), 
        .B(n28769), .Y(n28624) );
  AOI21xp33_ASAP7_75t_SL U30957 ( .A1(n24582), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__23_), .B(n28887), .Y(n26417) );
  OAI21xp33_ASAP7_75t_SL U30958 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__5_), 
        .A2(n24658), .B(n26844), .Y(n2792) );
  OAI21xp33_ASAP7_75t_SL U30959 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__5_), 
        .A2(n24656), .B(n31515), .Y(n2790) );
  OAI21xp33_ASAP7_75t_SL U30960 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__25_), 
        .A2(n24654), .B(n25542), .Y(n3769) );
  NAND2xp33_ASAP7_75t_SL U30961 ( .A(n22379), .B(DP_OP_1196_128_7433_n454), 
        .Y(n32163) );
  INVxp33_ASAP7_75t_SL U30962 ( .A(n31427), .Y(n31432) );
  INVxp33_ASAP7_75t_SL U30963 ( .A(n26734), .Y(n26725) );
  NAND2xp33_ASAP7_75t_SL U30964 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__13_), 
        .B(n28769), .Y(n26161) );
  NAND2xp33_ASAP7_75t_SL U30965 ( .A(n31336), .B(n29074), .Y(n29075) );
  NAND2xp5_ASAP7_75t_SL U30966 ( .A(n3704), .B(n25608), .Y(n29214) );
  OAI21xp33_ASAP7_75t_SL U30967 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__25_), 
        .A2(n24654), .B(n25540), .Y(n3771) );
  AOI22xp33_ASAP7_75t_SL U30968 ( .A1(ahbso_0__HRDATA__17_), .A2(n32904), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[21]), .B2(n32903), .Y(n32927) );
  NAND2xp33_ASAP7_75t_SL U30969 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), .B(
        n32161), .Y(n30653) );
  OAI21xp33_ASAP7_75t_SL U30970 ( .A1(n28552), .A2(n30642), .B(n28551), .Y(
        n28553) );
  OAI21xp33_ASAP7_75t_SL U30971 ( .A1(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .A2(
        n24657), .B(n32116), .Y(n2786) );
  BUFx12f_ASAP7_75t_SL U30972 ( .A(u0_0_leon3x0_p0_muli[37]), .Y(n24044) );
  AOI22xp33_ASAP7_75t_SL U30973 ( .A1(ahbso_0__HRDATA__20_), .A2(n32904), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[24]), .B2(n32903), .Y(n32951) );
  NOR2xp33_ASAP7_75t_SRAM U30974 ( .A(n32160), .B(n24641), .Y(rf_addr_w[7]) );
  OAI21xp33_ASAP7_75t_SL U30975 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__25_), 
        .A2(n24654), .B(n25538), .Y(n3773) );
  NOR2xp33_ASAP7_75t_SRAM U30976 ( .A(n32155), .B(n24641), .Y(rf_addr_w[2]) );
  OAI21xp33_ASAP7_75t_SL U30977 ( .A1(u0_0_leon3x0_p0_iu_v_E__CWP__0_), .A2(
        n24657), .B(n32118), .Y(n2784) );
  NOR2xp33_ASAP7_75t_SRAM U30978 ( .A(n32156), .B(n24641), .Y(rf_addr_w[3]) );
  NAND2xp5_ASAP7_75t_SL U30979 ( .A(n28013), .B(n28012), .Y(n28023) );
  AOI21xp33_ASAP7_75t_SL U30980 ( .A1(n28888), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__3_), .B(n28887), .Y(n28889) );
  INVxp33_ASAP7_75t_SL U30981 ( .A(DP_OP_1196_128_7433_n452), .Y(n26845) );
  OAI21xp33_ASAP7_75t_SL U30982 ( .A1(u0_0_leon3x0_p0_iu_v_A__CTRL__TRAP_), 
        .A2(n24654), .B(n31808), .Y(n3700) );
  INVxp33_ASAP7_75t_SL U30983 ( .A(DP_OP_1196_128_7433_n454), .Y(n26846) );
  INVxp67_ASAP7_75t_SL U30984 ( .A(DP_OP_1196_128_7433_n453), .Y(n26847) );
  AOI22xp33_ASAP7_75t_SL U30985 ( .A1(ahbso_0__HRDATA__22_), .A2(n32904), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[26]), .B2(n32903), .Y(n32967) );
  OAI21xp33_ASAP7_75t_SL U30986 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__13_), 
        .A2(n24653), .B(n28595), .Y(n2645) );
  NAND2xp33_ASAP7_75t_SL U30987 ( .A(n31336), .B(n26950), .Y(n26951) );
  NAND2xp33_ASAP7_75t_SL U30988 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[19]), .B(
        n32871), .Y(n32872) );
  INVx4_ASAP7_75t_SL U30989 ( .A(n23974), .Y(n23975) );
  NAND2xp5_ASAP7_75t_SL U30990 ( .A(n31579), .B(n31457), .Y(n31263) );
  OAI21xp33_ASAP7_75t_SL U30991 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__13_), 
        .A2(n24653), .B(n28597), .Y(n2643) );
  INVx1_ASAP7_75t_SL U30992 ( .A(n22939), .Y(n29561) );
  OAI21xp33_ASAP7_75t_SL U30993 ( .A1(n18839), .A2(n24654), .B(n31944), .Y(
        n3891) );
  NAND2xp33_ASAP7_75t_SL U30994 ( .A(n31336), .B(n27169), .Y(n27170) );
  OAI21xp5_ASAP7_75t_SL U30995 ( .A1(n28952), .A2(n30642), .B(n28951), .Y(
        n28953) );
  NAND2xp33_ASAP7_75t_SL U30996 ( .A(n30644), .B(n28602), .Y(n28604) );
  AOI22xp33_ASAP7_75t_SL U30997 ( .A1(ahbso_0__HRDATA__18_), .A2(n32904), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[22]), .B2(n32903), .Y(n32935) );
  NAND2xp33_ASAP7_75t_SL U30998 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__30_), .B(
        n22375), .Y(n29612) );
  NAND2xp33_ASAP7_75t_SL U30999 ( .A(n28833), .B(n32075), .Y(n25950) );
  AOI21xp33_ASAP7_75t_SL U31000 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__26_), 
        .A2(n22378), .B(n26822), .Y(n3766) );
  NAND2xp33_ASAP7_75t_SL U31001 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__16_), 
        .B(n28769), .Y(n26681) );
  INVxp67_ASAP7_75t_SL U31002 ( .A(n29613), .Y(n30591) );
  NAND2xp33_ASAP7_75t_SL U31003 ( .A(n29144), .B(u0_0_leon3x0_p0_divi[0]), .Y(
        n28996) );
  OAI21xp33_ASAP7_75t_SL U31004 ( .A1(n25331), .A2(n31607), .B(n25330), .Y(
        n25336) );
  INVx1_ASAP7_75t_SL U31005 ( .A(n24531), .Y(n22419) );
  NAND2xp33_ASAP7_75t_SL U31006 ( .A(n31264), .B(n32243), .Y(n25338) );
  OAI21xp33_ASAP7_75t_SL U31007 ( .A1(u0_0_leon3x0_p0_iu_v_E__CWP__1_), .A2(
        n24657), .B(n31349), .Y(n2798) );
  NAND2xp33_ASAP7_75t_SL U31008 ( .A(n25745), .B(n24670), .Y(n25746) );
  NAND2xp33_ASAP7_75t_SL U31009 ( .A(n27235), .B(n22378), .Y(n27236) );
  NAND2xp33_ASAP7_75t_SL U31010 ( .A(n26979), .B(n24667), .Y(n26980) );
  NAND2xp33_ASAP7_75t_SL U31011 ( .A(n30372), .B(n24664), .Y(n30367) );
  AND2x2_ASAP7_75t_SL U31012 ( .A(n25319), .B(n24671), .Y(n25318) );
  NAND2xp33_ASAP7_75t_SL U31013 ( .A(u0_0_leon3x0_p0_div0_r_X__31_), .B(n28371), .Y(n28376) );
  NAND2xp33_ASAP7_75t_SL U31014 ( .A(n25729), .B(n24670), .Y(n25730) );
  NAND2xp33_ASAP7_75t_SL U31015 ( .A(n28877), .B(n30007), .Y(n28898) );
  NAND2xp5_ASAP7_75t_SL U31016 ( .A(n24533), .B(n32455), .Y(n32456) );
  AOI21xp33_ASAP7_75t_SL U31017 ( .A1(n31824), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__7_), .B(n24679), .Y(n30822) );
  NAND2xp33_ASAP7_75t_SL U31018 ( .A(n25288), .B(n24673), .Y(n25287) );
  NAND2xp33_ASAP7_75t_SL U31019 ( .A(n25300), .B(n24672), .Y(n25299) );
  NAND2xp33_ASAP7_75t_SL U31020 ( .A(n23845), .B(n24678), .Y(n28532) );
  BUFx3_ASAP7_75t_SL U31021 ( .A(u0_0_leon3x0_p0_muli[40]), .Y(n22939) );
  NAND2xp33_ASAP7_75t_SL U31022 ( .A(n31834), .B(n24667), .Y(n31831) );
  NAND2xp33_ASAP7_75t_SL U31023 ( .A(n25747), .B(n24670), .Y(n25748) );
  NAND2xp33_ASAP7_75t_SL U31024 ( .A(n24701), .B(n24675), .Y(n24702) );
  NAND2xp33_ASAP7_75t_SL U31025 ( .A(n27127), .B(n22378), .Y(n27126) );
  NAND2xp5_ASAP7_75t_SL U31026 ( .A(n30004), .B(n30003), .Y(n30005) );
  AOI22xp33_ASAP7_75t_SL U31027 ( .A1(uart1_r_THOLD__19__5_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__27__5_), .Y(n27701) );
  NAND2xp33_ASAP7_75t_SL U31028 ( .A(n26977), .B(n24667), .Y(n26978) );
  NAND2xp33_ASAP7_75t_SL U31029 ( .A(n23841), .B(n24678), .Y(n28558) );
  AOI21xp33_ASAP7_75t_SL U31030 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[45]), 
        .B(n24679), .Y(n30362) );
  INVxp67_ASAP7_75t_SL U31031 ( .A(n30958), .Y(n26737) );
  NAND2xp33_ASAP7_75t_SL U31032 ( .A(n26975), .B(n24667), .Y(n26976) );
  NAND2xp33_ASAP7_75t_SL U31033 ( .A(n25298), .B(n24672), .Y(n25297) );
  NAND2xp33_ASAP7_75t_SL U31034 ( .A(n25727), .B(n24670), .Y(n25728) );
  NAND2xp33_ASAP7_75t_SL U31035 ( .A(n25294), .B(n24673), .Y(n25293) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31036 ( .A1(n31565), .A2(n31586), .B(n31564), 
        .C(n24684), .Y(n31567) );
  AOI22xp33_ASAP7_75t_SL U31037 ( .A1(n28011), .A2(uart1_r_THOLD__22__0_), 
        .B1(uart1_r_THOLD__18__0_), .B2(n28010), .Y(n28012) );
  NAND2xp33_ASAP7_75t_SL U31038 ( .A(n30377), .B(n24664), .Y(n30378) );
  NAND2xp33_ASAP7_75t_SL U31039 ( .A(n29619), .B(n24661), .Y(n29620) );
  INVxp33_ASAP7_75t_SL U31040 ( .A(n30876), .Y(n32611) );
  NAND2xp33_ASAP7_75t_SL U31041 ( .A(n25749), .B(n24670), .Y(n25750) );
  NAND2xp33_ASAP7_75t_SL U31042 ( .A(n25719), .B(n24670), .Y(n25720) );
  OAI22xp33_ASAP7_75t_SL U31043 ( .A1(n29469), .A2(n30686), .B1(n29468), .B2(
        n29467), .Y(n25365) );
  NAND2xp33_ASAP7_75t_SL U31044 ( .A(n30828), .B(n24663), .Y(n30826) );
  AND2x2_ASAP7_75t_SL U31045 ( .A(n27037), .B(n22378), .Y(n27038) );
  NAND2xp33_ASAP7_75t_SL U31046 ( .A(n25813), .B(n24670), .Y(n25726) );
  AOI22xp33_ASAP7_75t_SL U31047 ( .A1(n28015), .A2(uart1_r_THOLD__6__0_), .B1(
        uart1_r_THOLD__14__0_), .B2(n28014), .Y(n28021) );
  INVxp33_ASAP7_75t_SL U31048 ( .A(n32455), .Y(n31806) );
  NAND2xp33_ASAP7_75t_SL U31049 ( .A(n25751), .B(n24670), .Y(n25752) );
  NAND2xp33_ASAP7_75t_SL U31050 ( .A(n27168), .B(n24669), .Y(n26189) );
  AOI21xp33_ASAP7_75t_SL U31051 ( .A1(n28017), .A2(uart1_r_THOLD__26__0_), .B(
        n28016), .Y(n28020) );
  NAND2xp33_ASAP7_75t_SL U31052 ( .A(n25230), .B(n24985), .Y(n30962) );
  NAND2xp5_ASAP7_75t_SL U31053 ( .A(n25853), .B(n25852), .Y(n25854) );
  NAND2xp33_ASAP7_75t_SL U31054 ( .A(n32063), .B(n24661), .Y(n32064) );
  NAND2xp33_ASAP7_75t_SL U31055 ( .A(n25362), .B(n24673), .Y(n25235) );
  NAND2xp5_ASAP7_75t_SL U31056 ( .A(n29347), .B(n30068), .Y(n29342) );
  NAND2xp33_ASAP7_75t_SL U31057 ( .A(n25543), .B(n24671), .Y(n25544) );
  AOI22xp33_ASAP7_75t_SL U31058 ( .A1(apbi[13]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[17]), .B2(n31494), .Y(n1766) );
  AND2x2_ASAP7_75t_SL U31059 ( .A(n29082), .B(n24678), .Y(n29083) );
  AOI22xp33_ASAP7_75t_SL U31060 ( .A1(apbi[16]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[20]), .B2(n31494), .Y(n1773) );
  NAND2xp33_ASAP7_75t_SL U31061 ( .A(n24374), .B(n24415), .Y(n24375) );
  INVxp67_ASAP7_75t_SL U31062 ( .A(n32860), .Y(n32874) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31063 ( .A1(n25685), .A2(n25684), .B(n25683), 
        .C(n25682), .Y(n25686) );
  NAND2xp33_ASAP7_75t_SL U31064 ( .A(n31678), .B(n24665), .Y(n31413) );
  INVxp67_ASAP7_75t_SL U31065 ( .A(DP_OP_1196_128_7433_n97), .Y(
        DP_OP_1196_128_7433_n95) );
  NAND2xp33_ASAP7_75t_SL U31066 ( .A(n26373), .B(n24669), .Y(n26374) );
  AOI22xp33_ASAP7_75t_SL U31067 ( .A1(apbi[28]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[32]), .B2(n31494), .Y(n1781) );
  AOI21xp33_ASAP7_75t_SL U31068 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__28_), .B(n25429), .Y(n26947) );
  INVxp33_ASAP7_75t_SL U31069 ( .A(add_x_735_A_29_), .Y(n26924) );
  NAND2xp33_ASAP7_75t_SL U31070 ( .A(n30230), .B(n24667), .Y(n30231) );
  OAI31xp33_ASAP7_75t_SRAM U31071 ( .A1(n26764), .A2(u0_0_dbgo_OPTYPE__1_), 
        .A3(n29180), .B(n26763), .Y(n26765) );
  NAND2xp33_ASAP7_75t_SL U31072 ( .A(n31348), .B(n24664), .Y(n31349) );
  AND2x2_ASAP7_75t_SL U31073 ( .A(n30607), .B(n24662), .Y(n30608) );
  INVx1_ASAP7_75t_SL U31074 ( .A(n26810), .Y(n31510) );
  NAND2xp33_ASAP7_75t_SL U31075 ( .A(n26842), .B(n24668), .Y(n26843) );
  AOI22xp33_ASAP7_75t_SL U31076 ( .A1(apbi[26]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[30]), .B2(n31494), .Y(n4615) );
  OAI21xp5_ASAP7_75t_SL U31077 ( .A1(n30239), .A2(n22376), .B(n26337), .Y(
        n26950) );
  NAND2xp33_ASAP7_75t_SL U31078 ( .A(n26852), .B(n24668), .Y(n26844) );
  NAND2xp33_ASAP7_75t_SL U31079 ( .A(n31514), .B(n24665), .Y(n31515) );
  NAND2xp5_ASAP7_75t_SL U31080 ( .A(n32885), .B(n32906), .Y(n32912) );
  NAND2xp33_ASAP7_75t_SL U31081 ( .A(n32115), .B(n24661), .Y(n32116) );
  NAND2xp33_ASAP7_75t_SL U31082 ( .A(n32117), .B(n24661), .Y(n32118) );
  INVxp67_ASAP7_75t_SL U31083 ( .A(n31849), .Y(n30979) );
  OAI21xp5_ASAP7_75t_SL U31084 ( .A1(n30450), .A2(n22376), .B(n25494), .Y(
        n30465) );
  AOI21xp33_ASAP7_75t_SL U31085 ( .A1(n31391), .A2(rf_do_a[0]), .B(n24680), 
        .Y(n31394) );
  NAND2xp33_ASAP7_75t_SL U31086 ( .A(n31812), .B(n30007), .Y(n29004) );
  AND2x2_ASAP7_75t_SL U31087 ( .A(n26912), .B(n24667), .Y(n26913) );
  NAND2xp33_ASAP7_75t_SL U31088 ( .A(n29086), .B(n24677), .Y(n29087) );
  NOR2xp33_ASAP7_75t_SL U31089 ( .A(n25942), .B(n27475), .Y(n26130) );
  NAND2xp33_ASAP7_75t_SL U31090 ( .A(n25537), .B(n24671), .Y(n25538) );
  NAND2xp33_ASAP7_75t_SL U31091 ( .A(n25539), .B(n24671), .Y(n25540) );
  NOR3xp33_ASAP7_75t_SRAM U31092 ( .A(n31450), .B(n31449), .C(n31448), .Y(
        n31454) );
  OAI21xp33_ASAP7_75t_SL U31093 ( .A1(n2927), .A2(n25332), .B(n25324), .Y(
        n25325) );
  NAND2xp33_ASAP7_75t_SL U31094 ( .A(n25541), .B(n24671), .Y(n25542) );
  INVxp67_ASAP7_75t_SL U31095 ( .A(n25028), .Y(n32457) );
  INVx1_ASAP7_75t_SL U31096 ( .A(n31461), .Y(n32243) );
  NAND2xp5_ASAP7_75t_SL U31097 ( .A(n31607), .B(n25331), .Y(n25330) );
  AOI21xp33_ASAP7_75t_SL U31098 ( .A1(n32489), .A2(n25333), .B(n25332), .Y(
        n25334) );
  NAND2xp5_ASAP7_75t_SL U31099 ( .A(n31933), .B(n32454), .Y(n32044) );
  AND2x2_ASAP7_75t_SL U31100 ( .A(n29023), .B(n24676), .Y(n29024) );
  NAND2xp33_ASAP7_75t_SL U31101 ( .A(n32292), .B(n32291), .Y(n32353) );
  OR4x1_ASAP7_75t_SL U31102 ( .A(n25165), .B(n25164), .C(n25163), .D(n25162), 
        .Y(n26338) );
  OAI21xp5_ASAP7_75t_SL U31103 ( .A1(n32838), .A2(n32860), .B(n32908), .Y(
        n32839) );
  OAI21xp5_ASAP7_75t_SL U31104 ( .A1(n30397), .A2(n22376), .B(n25167), .Y(
        n29899) );
  OAI21xp33_ASAP7_75t_SL U31105 ( .A1(n18844), .A2(n26804), .B(n26803), .Y(
        n26805) );
  NAND2xp33_ASAP7_75t_SL U31106 ( .A(n31984), .B(n24660), .Y(n31985) );
  NAND2xp33_ASAP7_75t_SL U31107 ( .A(n25359), .B(n24674), .Y(n24960) );
  NAND2xp33_ASAP7_75t_SL U31108 ( .A(n25172), .B(n24675), .Y(n24704) );
  NAND2xp33_ASAP7_75t_SL U31109 ( .A(n25675), .B(n24675), .Y(n24703) );
  NAND2xp33_ASAP7_75t_SL U31110 ( .A(n28451), .B(n24678), .Y(n28450) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31111 ( .A1(n29966), .A2(n33065), .B(n29965), 
        .C(n24694), .Y(n29968) );
  AOI21xp33_ASAP7_75t_SL U31112 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__30_), .B(n25643), .Y(n29613) );
  AND2x2_ASAP7_75t_SL U31113 ( .A(n29084), .B(n22378), .Y(n29085) );
  NAND2xp33_ASAP7_75t_SL U31114 ( .A(n26831), .B(n24668), .Y(n26832) );
  NAND2xp33_ASAP7_75t_SL U31115 ( .A(n31516), .B(n24665), .Y(n31517) );
  AND2x2_ASAP7_75t_SL U31116 ( .A(n25278), .B(n24673), .Y(n25277) );
  INVxp33_ASAP7_75t_SL U31117 ( .A(n29144), .Y(n26358) );
  AOI21xp33_ASAP7_75t_SL U31118 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[37]), 
        .B(n24679), .Y(n30419) );
  AOI21xp33_ASAP7_75t_SL U31119 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[38]), 
        .B(n24679), .Y(n30408) );
  NAND2xp33_ASAP7_75t_SL U31120 ( .A(n30413), .B(n24664), .Y(n30414) );
  AOI21xp33_ASAP7_75t_SL U31121 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[39]), 
        .B(n24679), .Y(n30398) );
  NAND2xp33_ASAP7_75t_SL U31122 ( .A(n30403), .B(n24664), .Y(n30404) );
  INVxp33_ASAP7_75t_SL U31123 ( .A(add_x_735_A_19_), .Y(n25828) );
  INVx1_ASAP7_75t_SL U31124 ( .A(n30180), .Y(n30186) );
  NAND2xp33_ASAP7_75t_SL U31125 ( .A(n30524), .B(n24666), .Y(n29823) );
  INVxp67_ASAP7_75t_SL U31126 ( .A(n30183), .Y(n30185) );
  NAND2xp33_ASAP7_75t_SL U31127 ( .A(n23848), .B(n24676), .Y(n28800) );
  INVxp33_ASAP7_75t_SL U31128 ( .A(DP_OP_1196_128_7433_n291), .Y(
        DP_OP_1196_128_7433_n289) );
  INVxp33_ASAP7_75t_SL U31129 ( .A(DP_OP_1196_128_7433_n290), .Y(
        DP_OP_1196_128_7433_n288) );
  NAND2xp33_ASAP7_75t_SL U31130 ( .A(n29049), .B(n24676), .Y(n29050) );
  NAND2xp33_ASAP7_75t_SL U31131 ( .A(n29825), .B(n24666), .Y(n29826) );
  NAND2xp33_ASAP7_75t_SL U31132 ( .A(n26247), .B(n24669), .Y(n26248) );
  NAND2xp33_ASAP7_75t_SL U31133 ( .A(n29827), .B(n24666), .Y(n29828) );
  NAND2xp33_ASAP7_75t_SL U31134 ( .A(n29829), .B(n24666), .Y(n29830) );
  NAND2xp33_ASAP7_75t_SL U31135 ( .A(n26245), .B(n24669), .Y(n26246) );
  NAND2xp33_ASAP7_75t_SL U31136 ( .A(n26243), .B(n24669), .Y(n26244) );
  NAND2xp33_ASAP7_75t_SL U31137 ( .A(n25296), .B(n24672), .Y(n25295) );
  NAND2xp33_ASAP7_75t_SL U31138 ( .A(n28653), .B(n24677), .Y(n28654) );
  NAND2xp33_ASAP7_75t_SL U31139 ( .A(n25290), .B(n24673), .Y(n25289) );
  NAND2xp33_ASAP7_75t_SL U31140 ( .A(n26241), .B(n24669), .Y(n26242) );
  AOI21xp33_ASAP7_75t_SL U31141 ( .A1(n24428), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__Y__2_), .B(n30455), .Y(n30456) );
  AOI22xp33_ASAP7_75t_SL U31142 ( .A1(apbi[27]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[31]), .B2(n31494), .Y(n4527) );
  NAND2xp33_ASAP7_75t_SL U31143 ( .A(n28594), .B(n24677), .Y(n28595) );
  NAND2xp5_ASAP7_75t_SL U31144 ( .A(n27981), .B(n27980), .Y(n27995) );
  BUFx6f_ASAP7_75t_SL U31145 ( .A(u0_0_leon3x0_p0_muli[18]), .Y(n24068) );
  NAND2xp33_ASAP7_75t_SL U31146 ( .A(n28596), .B(n24677), .Y(n28597) );
  NAND2xp33_ASAP7_75t_SL U31147 ( .A(n30459), .B(n24663), .Y(n30460) );
  AOI22xp33_ASAP7_75t_SL U31148 ( .A1(apbi[15]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[19]), .B2(n31494), .Y(n4636) );
  NAND2xp33_ASAP7_75t_SL U31149 ( .A(n23846), .B(n24677), .Y(n28609) );
  NAND2xp33_ASAP7_75t_SL U31150 ( .A(uart1_r_THOLD__25__0_), .B(n27998), .Y(
        n27983) );
  NAND2xp33_ASAP7_75t_SL U31151 ( .A(n25283), .B(n24673), .Y(n25282) );
  AOI22xp33_ASAP7_75t_SL U31152 ( .A1(n28011), .A2(uart1_r_THOLD__20__0_), 
        .B1(uart1_r_THOLD__24__0_), .B2(n28017), .Y(n27991) );
  NAND2xp33_ASAP7_75t_SL U31153 ( .A(n29079), .B(n24677), .Y(n29080) );
  AND2x2_ASAP7_75t_SL U31154 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__0_), .B(n24676), 
        .Y(n29015) );
  NAND2xp33_ASAP7_75t_SL U31155 ( .A(n31687), .B(n24666), .Y(n31685) );
  AND2x2_ASAP7_75t_SL U31156 ( .A(n26350), .B(n24669), .Y(n26349) );
  NAND2xp33_ASAP7_75t_SL U31157 ( .A(n30220), .B(n24665), .Y(n30221) );
  OAI21xp5_ASAP7_75t_SL U31158 ( .A1(n29180), .A2(n22376), .B(n25406), .Y(
        n31335) );
  NAND2xp33_ASAP7_75t_SL U31159 ( .A(n29088), .B(n24678), .Y(n29089) );
  NAND2xp33_ASAP7_75t_SL U31160 ( .A(n30441), .B(n24664), .Y(n30436) );
  AOI22xp33_ASAP7_75t_SL U31161 ( .A1(apbi[9]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[13]), .B2(n31494), .Y(n1804) );
  AOI21xp33_ASAP7_75t_SL U31162 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[36]), 
        .B(n24679), .Y(n30431) );
  NAND2xp33_ASAP7_75t_SL U31163 ( .A(n24957), .B(n24674), .Y(n24958) );
  NAND2xp33_ASAP7_75t_SL U31164 ( .A(n31943), .B(n24667), .Y(n31944) );
  NAND2xp33_ASAP7_75t_SL U31165 ( .A(n30454), .B(n24664), .Y(n30447) );
  AOI21xp33_ASAP7_75t_SL U31166 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[53]), 
        .B(n24680), .Y(n30278) );
  NAND2xp33_ASAP7_75t_SL U31167 ( .A(n30287), .B(n24664), .Y(n30283) );
  NAND2xp33_ASAP7_75t_SL U31168 ( .A(n32072), .B(n24661), .Y(n32073) );
  OAI21xp5_ASAP7_75t_SL U31169 ( .A1(n30392), .A2(n22376), .B(n25519), .Y(
        n30721) );
  OAI21xp5_ASAP7_75t_SL U31170 ( .A1(n30252), .A2(n22376), .B(n26393), .Y(
        n29778) );
  NAND2xp33_ASAP7_75t_SL U31171 ( .A(n31807), .B(n24666), .Y(n31808) );
  AOI21xp33_ASAP7_75t_SL U31172 ( .A1(n22376), .A2(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__23_), .B(n26415), .Y(n26523) );
  OAI21xp5_ASAP7_75t_SL U31173 ( .A1(n30267), .A2(n22376), .B(n26217), .Y(
        n29074) );
  AND2x2_ASAP7_75t_SL U31174 ( .A(n25273), .B(n24673), .Y(n25272) );
  INVxp33_ASAP7_75t_SL U31175 ( .A(n27066), .Y(n27148) );
  OAI21xp5_ASAP7_75t_SL U31176 ( .A1(n30285), .A2(n22376), .B(n26959), .Y(
        n27027) );
  NAND2xp33_ASAP7_75t_SL U31177 ( .A(n29102), .B(n24677), .Y(n29103) );
  OAI21xp5_ASAP7_75t_SL U31178 ( .A1(n30297), .A2(n22376), .B(n25753), .Y(
        n28529) );
  OAI21xp5_ASAP7_75t_SL U31179 ( .A1(n30306), .A2(n22376), .B(n25711), .Y(
        n28540) );
  NAND2xp33_ASAP7_75t_SL U31180 ( .A(n25292), .B(n24673), .Y(n25291) );
  NAND2xp33_ASAP7_75t_SL U31181 ( .A(n31511), .B(n24665), .Y(n31512) );
  NAND2xp33_ASAP7_75t_SL U31182 ( .A(n26840), .B(n24668), .Y(n26841) );
  OAI21xp5_ASAP7_75t_SL U31183 ( .A1(n30317), .A2(n22376), .B(n26702), .Y(
        n27275) );
  NAND2xp33_ASAP7_75t_SL U31184 ( .A(n32160), .B(n24665), .Y(n31513) );
  INVx2_ASAP7_75t_SL U31185 ( .A(u0_0_leon3x0_p0_muli[42]), .Y(n24693) );
  OAI21xp5_ASAP7_75t_SL U31186 ( .A1(n30328), .A2(n22376), .B(n26444), .Y(
        n28554) );
  NAND3xp33_ASAP7_75t_SRAM U31187 ( .A(n32092), .B(n32091), .C(n32090), .Y(
        n32093) );
  AOI22xp33_ASAP7_75t_SL U31188 ( .A1(apbi[25]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[29]), .B2(n31494), .Y(n4625) );
  NAND2xp33_ASAP7_75t_SL U31189 ( .A(n24952), .B(n24674), .Y(n24953) );
  NAND2xp33_ASAP7_75t_SL U31190 ( .A(n31254), .B(n24663), .Y(n31255) );
  NAND2xp5_ASAP7_75t_SL U31191 ( .A(n29660), .B(n29663), .Y(n29637) );
  NAND2xp33_ASAP7_75t_SL U31192 ( .A(n27045), .B(n22378), .Y(n27046) );
  AOI21xp33_ASAP7_75t_SL U31193 ( .A1(n31824), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__9_), .B(n24679), .Y(n27039) );
  AOI22xp33_ASAP7_75t_SL U31194 ( .A1(apbi[31]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[35]), .B2(n31494), .Y(n4771) );
  INVxp33_ASAP7_75t_SL U31195 ( .A(n32410), .Y(n32655) );
  NAND2xp33_ASAP7_75t_SL U31196 ( .A(n31786), .B(n24668), .Y(n26877) );
  INVxp33_ASAP7_75t_SL U31197 ( .A(n24717), .Y(n24716) );
  INVxp33_ASAP7_75t_SL U31198 ( .A(n32419), .Y(n32657) );
  NAND2xp33_ASAP7_75t_SL U31199 ( .A(n29231), .B(n24675), .Y(n29232) );
  AOI22xp33_ASAP7_75t_SL U31200 ( .A1(n31217), .A2(uart1_r_RHOLD__29__1_), 
        .B1(uart1_r_RHOLD__3__1_), .B2(n31216), .Y(n27442) );
  NAND2xp33_ASAP7_75t_SL U31201 ( .A(n31765), .B(n22378), .Y(n27043) );
  NAND2xp5_ASAP7_75t_SL U31202 ( .A(timer0_N65), .B(n24392), .Y(n24418) );
  NAND2xp33_ASAP7_75t_SL U31203 ( .A(n31518), .B(n24665), .Y(n31519) );
  NAND2xp33_ASAP7_75t_SL U31204 ( .A(n31537), .B(n24666), .Y(n31538) );
  AOI22xp33_ASAP7_75t_SL U31205 ( .A1(n31219), .A2(uart1_r_RHOLD__11__1_), 
        .B1(uart1_r_RHOLD__23__1_), .B2(n31218), .Y(n27441) );
  NAND2xp33_ASAP7_75t_SL U31206 ( .A(n25695), .B(n24675), .Y(n24917) );
  NAND2xp33_ASAP7_75t_SL U31207 ( .A(n27191), .B(n22378), .Y(n27178) );
  AOI22xp33_ASAP7_75t_SL U31208 ( .A1(apbi[8]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[12]), .B2(n31494), .Y(n4685) );
  NAND2xp5_ASAP7_75t_SL U31209 ( .A(n30955), .B(n24929), .Y(n24983) );
  INVx1_ASAP7_75t_SL U31210 ( .A(n31722), .Y(n31718) );
  NAND2xp33_ASAP7_75t_SL U31211 ( .A(n31864), .B(n24667), .Y(n31865) );
  AND2x2_ASAP7_75t_SL U31212 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__1_), .B(n24662), 
        .Y(n30649) );
  INVxp33_ASAP7_75t_SL U31213 ( .A(n28110), .Y(n28115) );
  INVx1_ASAP7_75t_SL U31214 ( .A(n24882), .Y(n24876) );
  NAND2xp5_ASAP7_75t_SL U31215 ( .A(n25497), .B(n30614), .Y(n26176) );
  NAND2xp33_ASAP7_75t_SL U31216 ( .A(n26214), .B(n24669), .Y(n26215) );
  NAND2xp33_ASAP7_75t_SL U31217 ( .A(n29037), .B(n24676), .Y(n29038) );
  NAND2xp33_ASAP7_75t_SL U31218 ( .A(n31866), .B(n24667), .Y(n31867) );
  NAND2xp5_ASAP7_75t_SL U31219 ( .A(n24882), .B(n25215), .Y(n24911) );
  NAND2xp33_ASAP7_75t_SL U31220 ( .A(n30292), .B(n24664), .Y(n30293) );
  NAND2xp33_ASAP7_75t_SL U31221 ( .A(n30585), .B(n24663), .Y(n30586) );
  NAND2xp33_ASAP7_75t_SL U31222 ( .A(n25356), .B(n24674), .Y(n24959) );
  NAND2xp33_ASAP7_75t_SL U31223 ( .A(n26212), .B(n24669), .Y(n26213) );
  NAND2xp33_ASAP7_75t_SL U31224 ( .A(n18799), .B(n24675), .Y(n24915) );
  INVxp33_ASAP7_75t_SL U31225 ( .A(n32371), .Y(n32635) );
  NAND2xp5_ASAP7_75t_SL U31226 ( .A(n28032), .B(n28033), .Y(n29952) );
  NAND2xp33_ASAP7_75t_SL U31227 ( .A(n27179), .B(n22378), .Y(n27180) );
  INVxp33_ASAP7_75t_SL U31228 ( .A(n32377), .Y(n32637) );
  NAND2xp33_ASAP7_75t_SL U31229 ( .A(n29765), .B(n24659), .Y(n29766) );
  INVxp33_ASAP7_75t_SL U31230 ( .A(n31262), .Y(n25398) );
  NAND2xp33_ASAP7_75t_SL U31231 ( .A(n25707), .B(n24670), .Y(n25708) );
  AOI21xp33_ASAP7_75t_SL U31232 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[49]), 
        .B(n24679), .Y(n30318) );
  NAND2xp33_ASAP7_75t_SL U31233 ( .A(n29774), .B(n24660), .Y(n29775) );
  NAND2xp33_ASAP7_75t_SL U31234 ( .A(n30323), .B(n24664), .Y(n30324) );
  NAND2xp33_ASAP7_75t_SL U31235 ( .A(n29776), .B(n24667), .Y(n29777) );
  AND2x2_ASAP7_75t_SL U31236 ( .A(n29098), .B(n24677), .Y(n29099) );
  AOI22xp33_ASAP7_75t_SL U31237 ( .A1(n28011), .A2(uart1_r_THOLD__22__6_), 
        .B1(uart1_r_THOLD__18__6_), .B2(n28010), .Y(n27640) );
  INVxp33_ASAP7_75t_SL U31238 ( .A(n32382), .Y(n32641) );
  AOI22xp33_ASAP7_75t_SL U31239 ( .A1(n28015), .A2(uart1_r_THOLD__6__6_), .B1(
        uart1_r_THOLD__14__6_), .B2(n28014), .Y(n27644) );
  AOI21xp33_ASAP7_75t_SL U31240 ( .A1(n28017), .A2(uart1_r_THOLD__26__6_), .B(
        n28016), .Y(n27643) );
  AOI21xp33_ASAP7_75t_SL U31241 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[50]), 
        .B(n24680), .Y(n30308) );
  INVxp33_ASAP7_75t_SL U31242 ( .A(n32384), .Y(n32643) );
  NAND2xp33_ASAP7_75t_SL U31243 ( .A(n30313), .B(n24664), .Y(n30314) );
  AOI22xp33_ASAP7_75t_SL U31244 ( .A1(apbi[14]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[18]), .B2(n31494), .Y(n2326) );
  NAND2xp5_ASAP7_75t_SL U31245 ( .A(n31027), .B(n29858), .Y(n28253) );
  NAND2xp5_ASAP7_75t_SL U31246 ( .A(n26507), .B(n26506), .Y(n26508) );
  NAND2xp33_ASAP7_75t_SL U31247 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__11_), 
        .B(n24581), .Y(n28685) );
  INVxp33_ASAP7_75t_SL U31248 ( .A(n31378), .Y(n32647) );
  NAND2xp5_ASAP7_75t_SL U31249 ( .A(n29434), .B(n29438), .Y(n29635) );
  NAND2xp33_ASAP7_75t_SL U31250 ( .A(n18891), .B(n29144), .Y(n27141) );
  INVxp33_ASAP7_75t_SL U31251 ( .A(n32399), .Y(n32649) );
  INVx1_ASAP7_75t_SL U31252 ( .A(n29450), .Y(n29634) );
  OAI21xp33_ASAP7_75t_SL U31253 ( .A1(n29438), .A2(n29437), .B(n29436), .Y(
        n29439) );
  NAND2xp33_ASAP7_75t_SL U31254 ( .A(n25313), .B(n24672), .Y(n25312) );
  NAND2xp33_ASAP7_75t_SL U31255 ( .A(n30517), .B(n24678), .Y(n28569) );
  NAND2xp33_ASAP7_75t_SL U31256 ( .A(n26829), .B(n24668), .Y(n26830) );
  NAND2xp33_ASAP7_75t_SL U31257 ( .A(n27051), .B(n22378), .Y(n27052) );
  INVxp33_ASAP7_75t_SL U31258 ( .A(n30904), .Y(n32651) );
  AOI22xp33_ASAP7_75t_SL U31259 ( .A1(n31215), .A2(uart1_r_RHOLD__28__1_), 
        .B1(uart1_r_RHOLD__1__1_), .B2(n31214), .Y(n27443) );
  NAND2xp33_ASAP7_75t_SL U31260 ( .A(n27049), .B(n22378), .Y(n27050) );
  AOI21xp33_ASAP7_75t_SL U31261 ( .A1(n31824), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__15_), .B(n24679), .Y(n26873) );
  AND2x2_ASAP7_75t_SL U31262 ( .A(n29092), .B(n24677), .Y(n29093) );
  INVxp33_ASAP7_75t_SL U31263 ( .A(n31509), .Y(n32653) );
  NAND2xp33_ASAP7_75t_SL U31264 ( .A(n27047), .B(n22378), .Y(n27048) );
  NAND2xp33_ASAP7_75t_SL U31265 ( .A(n28563), .B(n24678), .Y(n28564) );
  NAND2xp33_ASAP7_75t_SL U31266 ( .A(n30334), .B(n24664), .Y(n30335) );
  NAND2xp33_ASAP7_75t_SL U31267 ( .A(n25545), .B(n24671), .Y(n25546) );
  NAND2xp33_ASAP7_75t_SL U31268 ( .A(n25547), .B(n24671), .Y(n25548) );
  NAND2xp33_ASAP7_75t_SL U31269 ( .A(n32169), .B(n29206), .Y(n26806) );
  NAND2xp33_ASAP7_75t_SL U31270 ( .A(n27265), .B(n24679), .Y(n27266) );
  INVxp33_ASAP7_75t_SL U31271 ( .A(n25557), .Y(n25561) );
  INVxp33_ASAP7_75t_SL U31272 ( .A(n30671), .Y(n29168) );
  AOI31xp33_ASAP7_75t_SRAM U31273 ( .A1(n25705), .A2(n24991), .A3(n25080), .B(
        n24990), .Y(n24992) );
  NAND2xp33_ASAP7_75t_SL U31274 ( .A(n26723), .B(n24668), .Y(n26724) );
  AOI22xp33_ASAP7_75t_SL U31275 ( .A1(apbi[29]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[33]), .B2(n31494), .Y(n4665) );
  OAI21xp5_ASAP7_75t_SL U31276 ( .A1(u0_0_leon3x0_p0_c0mmu_a0_r_HLOCKEN_), 
        .A2(n25246), .B(n24896), .Y(n24974) );
  NAND2xp33_ASAP7_75t_SL U31277 ( .A(n26837), .B(n24668), .Y(n26838) );
  NAND2xp33_ASAP7_75t_SL U31278 ( .A(n29577), .B(n24661), .Y(n29578) );
  NAND2xp33_ASAP7_75t_SL U31279 ( .A(n28965), .B(n24674), .Y(n24996) );
  INVxp67_ASAP7_75t_SL U31280 ( .A(n25956), .Y(n25957) );
  NAND2xp5_ASAP7_75t_SL U31281 ( .A(n31949), .B(n30801), .Y(n4746) );
  AND2x2_ASAP7_75t_SL U31282 ( .A(n29096), .B(n22378), .Y(n29097) );
  NAND2xp33_ASAP7_75t_SL U31283 ( .A(n30923), .B(n24668), .Y(n26839) );
  NAND2xp33_ASAP7_75t_SL U31284 ( .A(n32650), .B(n24671), .Y(n25510) );
  AOI22xp33_ASAP7_75t_SL U31285 ( .A1(apbi[12]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[16]), .B2(n31494), .Y(n4754) );
  NAND2xp33_ASAP7_75t_SL U31286 ( .A(n32156), .B(n24666), .Y(n31521) );
  AOI22xp33_ASAP7_75t_SL U31287 ( .A1(apbi[30]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[34]), .B2(n31494), .Y(n4737) );
  NAND2xp33_ASAP7_75t_SL U31288 ( .A(n32652), .B(n24667), .Y(n26911) );
  INVxp33_ASAP7_75t_SL U31289 ( .A(n31824), .Y(n29888) );
  NAND2xp33_ASAP7_75t_SL U31290 ( .A(n24580), .B(n18909), .Y(n26362) );
  INVxp67_ASAP7_75t_SL U31291 ( .A(n25584), .Y(n25019) );
  NAND2xp33_ASAP7_75t_SL U31292 ( .A(n32656), .B(n24670), .Y(n25918) );
  AOI22xp33_ASAP7_75t_SL U31293 ( .A1(apbi[11]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[15]), .B2(n31494), .Y(n4521) );
  NAND2xp33_ASAP7_75t_SL U31294 ( .A(n32658), .B(n24662), .Y(n30596) );
  NAND2xp33_ASAP7_75t_SL U31295 ( .A(n31982), .B(n24659), .Y(n31983) );
  AOI21xp33_ASAP7_75t_SL U31296 ( .A1(n31824), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__TBA__17_), .B(n24679), .Y(n29025) );
  AOI22xp33_ASAP7_75t_SL U31297 ( .A1(apbi[17]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[21]), .B2(n31494), .Y(n4033) );
  OAI21xp33_ASAP7_75t_SL U31298 ( .A1(n30705), .A2(n29733), .B(n29732), .Y(
        n30709) );
  NAND2xp33_ASAP7_75t_SL U31299 ( .A(n31690), .B(n24676), .Y(n29029) );
  NAND2xp5_ASAP7_75t_SL U31300 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__15_), .B(n30207), .Y(n25046) );
  NAND2xp33_ASAP7_75t_SL U31301 ( .A(n29708), .B(n24662), .Y(n24700) );
  NAND2xp33_ASAP7_75t_SL U31302 ( .A(n25453), .B(n24671), .Y(n25454) );
  NAND2xp33_ASAP7_75t_SL U31303 ( .A(n26210), .B(n24669), .Y(n26211) );
  NAND2xp33_ASAP7_75t_SL U31304 ( .A(n30583), .B(n24663), .Y(n30584) );
  NAND2xp33_ASAP7_75t_SL U31305 ( .A(n31819), .B(n24666), .Y(n31820) );
  NAND2xp33_ASAP7_75t_SL U31306 ( .A(n25549), .B(n24671), .Y(n25550) );
  NAND2xp33_ASAP7_75t_SL U31307 ( .A(n31961), .B(n24674), .Y(n24955) );
  NAND2xp33_ASAP7_75t_SL U31308 ( .A(n26208), .B(n24669), .Y(n26209) );
  INVxp33_ASAP7_75t_SL U31309 ( .A(n32709), .Y(n31750) );
  AOI22xp33_ASAP7_75t_SL U31310 ( .A1(apbi[24]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[28]), .B2(n31494), .Y(n2273) );
  NAND2xp33_ASAP7_75t_SL U31311 ( .A(n28395), .B(n22378), .Y(n28396) );
  AOI22xp33_ASAP7_75t_SL U31312 ( .A1(n28015), .A2(uart1_r_THOLD__6__4_), .B1(
        uart1_r_THOLD__14__4_), .B2(n28014), .Y(n27777) );
  INVxp67_ASAP7_75t_SL U31313 ( .A(n25224), .Y(n25228) );
  AOI22xp33_ASAP7_75t_SL U31314 ( .A1(n28011), .A2(uart1_r_THOLD__22__4_), 
        .B1(uart1_r_THOLD__18__4_), .B2(n28010), .Y(n27779) );
  NAND2xp5_ASAP7_75t_SL U31315 ( .A(n27773), .B(n27772), .Y(n27782) );
  NAND2xp33_ASAP7_75t_SL U31316 ( .A(uart1_r_THOLD__19__4_), .B(n27999), .Y(
        n27769) );
  OAI21xp33_ASAP7_75t_SL U31317 ( .A1(n26761), .A2(n26789), .B(n29179), .Y(
        n26770) );
  AOI22xp33_ASAP7_75t_SL U31318 ( .A1(n28011), .A2(uart1_r_THOLD__20__4_), 
        .B1(uart1_r_THOLD__24__4_), .B2(n28017), .Y(n27763) );
  NAND2xp33_ASAP7_75t_SL U31319 ( .A(n28393), .B(n22378), .Y(n28394) );
  NAND2xp33_ASAP7_75t_SL U31320 ( .A(n25551), .B(n24671), .Y(n25552) );
  INVxp33_ASAP7_75t_SL U31321 ( .A(n24883), .Y(n24871) );
  NAND2xp33_ASAP7_75t_SL U31322 ( .A(n28391), .B(n22378), .Y(n28392) );
  NAND2xp5_ASAP7_75t_SL U31323 ( .A(n27758), .B(n27757), .Y(n27766) );
  NAND2xp33_ASAP7_75t_SL U31324 ( .A(uart1_r_THOLD__17__4_), .B(n27999), .Y(
        n27755) );
  NAND2xp33_ASAP7_75t_SL U31325 ( .A(n30719), .B(n24662), .Y(n30720) );
  NAND2xp33_ASAP7_75t_SL U31326 ( .A(n29094), .B(n24678), .Y(n29095) );
  NAND2xp33_ASAP7_75t_SL U31327 ( .A(n26833), .B(n24668), .Y(n26834) );
  NAND2xp33_ASAP7_75t_SL U31328 ( .A(n32137), .B(n24674), .Y(n24954) );
  AOI21xp33_ASAP7_75t_SL U31329 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[51]), 
        .B(n24679), .Y(n30298) );
  NAND2xp33_ASAP7_75t_SL U31330 ( .A(n28389), .B(n22378), .Y(n28390) );
  NAND2xp33_ASAP7_75t_SL U31331 ( .A(n32010), .B(n24660), .Y(n32011) );
  NAND2xp33_ASAP7_75t_SL U31332 ( .A(n30717), .B(n24662), .Y(n30718) );
  NAND2xp33_ASAP7_75t_SL U31333 ( .A(n26835), .B(n24668), .Y(n26836) );
  OAI21xp33_ASAP7_75t_SL U31334 ( .A1(n26794), .A2(n26793), .B(n26792), .Y(
        n26795) );
  INVxp67_ASAP7_75t_SL U31335 ( .A(DP_OP_1196_128_7433_n98), .Y(
        DP_OP_1196_128_7433_n96) );
  NAND2xp33_ASAP7_75t_SL U31336 ( .A(n30581), .B(n24663), .Y(n30582) );
  NAND2xp33_ASAP7_75t_SL U31337 ( .A(n32155), .B(n24666), .Y(n31520) );
  OAI21xp5_ASAP7_75t_SL U31338 ( .A1(n29733), .A2(n25948), .B(n25947), .Y(
        n29676) );
  NAND2xp33_ASAP7_75t_SL U31339 ( .A(n30715), .B(n24662), .Y(n30716) );
  NAND2xp33_ASAP7_75t_SL U31340 ( .A(n29173), .B(n24675), .Y(n29174) );
  NAND2xp33_ASAP7_75t_SL U31341 ( .A(n25887), .B(n24670), .Y(n25888) );
  NAND2xp33_ASAP7_75t_SL U31342 ( .A(n26721), .B(n24668), .Y(n26722) );
  NAND2xp33_ASAP7_75t_SL U31343 ( .A(n32012), .B(n24660), .Y(n32013) );
  NAND2xp33_ASAP7_75t_SL U31344 ( .A(n25080), .B(n24675), .Y(n24706) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U31345 ( .A1(n29715), .A2(n29714), .B(n29713), .C(
        n29712), .Y(n29725) );
  NAND2xp33_ASAP7_75t_SL U31346 ( .A(n25455), .B(n24671), .Y(n25456) );
  NAND2xp33_ASAP7_75t_SL U31347 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__23_), .B(
        n24669), .Y(n26442) );
  AOI22xp33_ASAP7_75t_SL U31348 ( .A1(uart1_r_THOLD__17__5_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__25__5_), .Y(n27693) );
  NAND2xp33_ASAP7_75t_SL U31349 ( .A(n30346), .B(n24664), .Y(n30347) );
  OAI21xp33_ASAP7_75t_SL U31350 ( .A1(n27986), .A2(n27704), .B(n27703), .Y(
        n27706) );
  NAND2xp33_ASAP7_75t_SL U31351 ( .A(n31389), .B(n24664), .Y(n31390) );
  AOI21xp33_ASAP7_75t_SL U31352 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[46]), 
        .B(n24679), .Y(n30352) );
  NAND2xp33_ASAP7_75t_SL U31353 ( .A(n25309), .B(n24672), .Y(n25308) );
  NAND2xp33_ASAP7_75t_SL U31354 ( .A(n26881), .B(n24668), .Y(n26882) );
  NAND2xp33_ASAP7_75t_SL U31355 ( .A(n23836), .B(n24678), .Y(n28467) );
  NAND2xp33_ASAP7_75t_SL U31356 ( .A(n30357), .B(n24664), .Y(n30358) );
  NAND2xp33_ASAP7_75t_SL U31357 ( .A(n32628), .B(n24669), .Y(n26584) );
  OR2x2_ASAP7_75t_SL U31358 ( .A(n25533), .B(n25988), .Y(n27328) );
  NAND2xp33_ASAP7_75t_SL U31359 ( .A(uart1_r_THOLD__25__6_), .B(n27998), .Y(
        n27625) );
  AOI22xp33_ASAP7_75t_SL U31360 ( .A1(n28011), .A2(uart1_r_THOLD__22__5_), 
        .B1(uart1_r_THOLD__18__5_), .B2(n28010), .Y(n27708) );
  AOI22xp33_ASAP7_75t_SL U31361 ( .A1(uart1_r_THOLD__19__2_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__27__2_), .Y(n27893) );
  AOI22xp33_ASAP7_75t_SL U31362 ( .A1(n28011), .A2(uart1_r_THOLD__20__1_), 
        .B1(uart1_r_THOLD__16__1_), .B2(n28010), .Y(n27414) );
  NAND2xp33_ASAP7_75t_SL U31363 ( .A(n25894), .B(n24675), .Y(n24923) );
  NAND2xp33_ASAP7_75t_SL U31364 ( .A(n28455), .B(n24678), .Y(n28456) );
  INVxp33_ASAP7_75t_SL U31365 ( .A(n32361), .Y(n32631) );
  AOI22xp33_ASAP7_75t_SL U31366 ( .A1(uart1_r_THOLD__19__3_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__27__3_), .Y(n27829) );
  NAND2xp33_ASAP7_75t_SL U31367 ( .A(n26879), .B(n24668), .Y(n26880) );
  NAND2xp33_ASAP7_75t_SL U31368 ( .A(n26883), .B(n24667), .Y(n26884) );
  NAND2xp5_ASAP7_75t_SL U31369 ( .A(n27623), .B(n27622), .Y(n27635) );
  AOI22xp33_ASAP7_75t_SL U31370 ( .A1(n28015), .A2(uart1_r_THOLD__4__1_), .B1(
        uart1_r_THOLD__12__1_), .B2(n28014), .Y(n27412) );
  AOI21xp33_ASAP7_75t_SL U31371 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[54]), 
        .B(n24679), .Y(n30268) );
  AOI22xp33_ASAP7_75t_SL U31372 ( .A1(n28011), .A2(uart1_r_THOLD__20__3_), 
        .B1(uart1_r_THOLD__16__3_), .B2(n28010), .Y(n27844) );
  AOI22xp33_ASAP7_75t_SL U31373 ( .A1(n28011), .A2(uart1_r_THOLD__22__1_), 
        .B1(uart1_r_THOLD__26__1_), .B2(n28017), .Y(n27419) );
  AOI21xp33_ASAP7_75t_SL U31374 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[47]), 
        .B(n24679), .Y(n30341) );
  NAND2xp33_ASAP7_75t_SL U31375 ( .A(n30273), .B(n24665), .Y(n30274) );
  INVxp33_ASAP7_75t_SL U31376 ( .A(n32354), .Y(n32629) );
  NAND2xp33_ASAP7_75t_SL U31377 ( .A(n28706), .B(n24676), .Y(n28707) );
  NAND2xp33_ASAP7_75t_SL U31378 ( .A(n25304), .B(n24672), .Y(n25303) );
  NAND2xp33_ASAP7_75t_SL U31379 ( .A(n31810), .B(n24674), .Y(n25001) );
  OAI21xp33_ASAP7_75t_SL U31380 ( .A1(n27986), .A2(n27840), .B(n27839), .Y(
        n27842) );
  NAND2xp33_ASAP7_75t_SL U31381 ( .A(n30258), .B(n24665), .Y(n30259) );
  NAND2xp33_ASAP7_75t_SL U31382 ( .A(n31812), .B(n24674), .Y(n25002) );
  INVxp33_ASAP7_75t_SL U31383 ( .A(n30155), .Y(n32615) );
  NAND2xp33_ASAP7_75t_SL U31384 ( .A(n29488), .B(n24660), .Y(n29489) );
  AOI21xp33_ASAP7_75t_SL U31385 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[48]), 
        .B(n24679), .Y(n30329) );
  NAND2xp33_ASAP7_75t_SL U31386 ( .A(n23839), .B(n22378), .Y(n27133) );
  AOI21xp5_ASAP7_75t_SL U31387 ( .A1(n25956), .A2(n25953), .B(n25954), .Y(
        n31251) );
  AOI22xp33_ASAP7_75t_SL U31388 ( .A1(n28015), .A2(uart1_r_THOLD__4__5_), .B1(
        uart1_r_THOLD__12__5_), .B2(n28014), .Y(n27694) );
  NAND2xp33_ASAP7_75t_SL U31389 ( .A(n30692), .B(n24660), .Y(n30693) );
  NAND2xp33_ASAP7_75t_SL U31390 ( .A(n28708), .B(n24676), .Y(n28709) );
  AOI22xp33_ASAP7_75t_SL U31391 ( .A1(n28011), .A2(uart1_r_THOLD__20__6_), 
        .B1(uart1_r_THOLD__24__6_), .B2(n28017), .Y(n27631) );
  INVxp33_ASAP7_75t_SL U31392 ( .A(n29670), .Y(n29672) );
  NAND2xp33_ASAP7_75t_SL U31393 ( .A(n24968), .B(n24674), .Y(n24969) );
  NAND2xp33_ASAP7_75t_SL U31394 ( .A(n28417), .B(n24678), .Y(n28418) );
  INVxp33_ASAP7_75t_SL U31395 ( .A(n32367), .Y(n32633) );
  NAND2xp33_ASAP7_75t_SL U31396 ( .A(n29486), .B(n24659), .Y(n29487) );
  AOI22xp33_ASAP7_75t_SL U31397 ( .A1(n28011), .A2(uart1_r_THOLD__20__5_), 
        .B1(uart1_r_THOLD__16__5_), .B2(n28010), .Y(n27696) );
  INVxp33_ASAP7_75t_SL U31398 ( .A(n30686), .Y(n30688) );
  AND2x2_ASAP7_75t_SL U31399 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__TT__1_), .B(
        n24661), .Y(n29671) );
  AOI22xp33_ASAP7_75t_SL U31400 ( .A1(n28011), .A2(uart1_r_THOLD__22__2_), 
        .B1(uart1_r_THOLD__26__2_), .B2(n28017), .Y(n27908) );
  AOI22xp33_ASAP7_75t_SL U31401 ( .A1(n28015), .A2(uart1_r_THOLD__6__3_), .B1(
        uart1_r_THOLD__14__3_), .B2(n28014), .Y(n27830) );
  NAND2xp33_ASAP7_75t_SL U31402 ( .A(n28754), .B(n24676), .Y(n28755) );
  NAND2xp33_ASAP7_75t_SL U31403 ( .A(n25420), .B(n25419), .Y(n25421) );
  AOI22xp33_ASAP7_75t_SL U31404 ( .A1(uart1_r_THOLD__19__1_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__27__1_), .Y(n27398) );
  AND2x2_ASAP7_75t_SL U31405 ( .A(n27025), .B(n24678), .Y(n27026) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31406 ( .A1(n31943), .A2(n25650), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_), .C(n24938), .Y(n24942) );
  NAND2xp33_ASAP7_75t_SL U31407 ( .A(n2929), .B(n31252), .Y(n27464) );
  NAND2xp33_ASAP7_75t_SL U31408 ( .A(n26981), .B(n24667), .Y(n26982) );
  NAND2xp33_ASAP7_75t_SL U31409 ( .A(n27183), .B(n22378), .Y(n27184) );
  NAND2xp33_ASAP7_75t_SL U31410 ( .A(n26368), .B(n24675), .Y(n25276) );
  NAND2xp33_ASAP7_75t_SL U31411 ( .A(n28698), .B(n24677), .Y(n28658) );
  AOI22xp33_ASAP7_75t_SL U31412 ( .A1(n28015), .A2(uart1_r_THOLD__6__1_), .B1(
        uart1_r_THOLD__14__1_), .B2(n28014), .Y(n27417) );
  INVxp33_ASAP7_75t_SL U31413 ( .A(n28785), .Y(n26268) );
  NAND2xp33_ASAP7_75t_SL U31414 ( .A(n26885), .B(n24667), .Y(n26886) );
  AOI22xp33_ASAP7_75t_SL U31415 ( .A1(n28011), .A2(uart1_r_THOLD__20__2_), 
        .B1(uart1_r_THOLD__24__2_), .B2(n28017), .Y(n27904) );
  BUFx6f_ASAP7_75t_SL U31416 ( .A(u0_0_leon3x0_p0_muli[27]), .Y(n24057) );
  NAND2xp33_ASAP7_75t_SL U31417 ( .A(n30797), .B(n24663), .Y(n30798) );
  INVxp33_ASAP7_75t_SL U31418 ( .A(n31032), .Y(n32627) );
  AOI22xp33_ASAP7_75t_SL U31419 ( .A1(n28015), .A2(uart1_r_THOLD__6__2_), .B1(
        uart1_r_THOLD__14__2_), .B2(n28014), .Y(n27906) );
  NAND2xp33_ASAP7_75t_SL U31420 ( .A(n28453), .B(n24678), .Y(n28454) );
  NAND2xp33_ASAP7_75t_SL U31421 ( .A(n24972), .B(n24674), .Y(n24973) );
  INVx1_ASAP7_75t_SL U31422 ( .A(n24430), .Y(n22420) );
  NAND2xp33_ASAP7_75t_SL U31423 ( .A(n23840), .B(n24677), .Y(n28579) );
  AOI22xp33_ASAP7_75t_SL U31424 ( .A1(apbi[10]), .A2(n31639), .B1(
        u0_0_leon3x0_p0_c0mmu_mcdi[14]), .B2(n31494), .Y(n4457) );
  AOI22xp33_ASAP7_75t_SL U31425 ( .A1(n28011), .A2(uart1_r_THOLD__22__3_), 
        .B1(uart1_r_THOLD__26__3_), .B2(n28017), .Y(n27832) );
  NAND2xp33_ASAP7_75t_SL U31426 ( .A(n25302), .B(n24672), .Y(n25301) );
  NAND2xp33_ASAP7_75t_SL U31427 ( .A(n25274), .B(n24673), .Y(n25275) );
  INVx1_ASAP7_75t_SL U31428 ( .A(n24681), .Y(n24676) );
  AOI22xp33_ASAP7_75t_SL U31429 ( .A1(uart1_r_THOLD__3__1_), .A2(n28003), .B1(
        n28002), .B2(uart1_r_THOLD__7__1_), .Y(n27396) );
  INVx1_ASAP7_75t_SL U31430 ( .A(n30774), .Y(n29958) );
  AOI22xp33_ASAP7_75t_SL U31431 ( .A1(uart1_r_THOLD__23__3_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__11__3_), .Y(n27827) );
  INVxp33_ASAP7_75t_SL U31432 ( .A(n31428), .Y(n31425) );
  AOI22xp33_ASAP7_75t_SL U31433 ( .A1(uart1_r_THOLD__3__3_), .A2(n28003), .B1(
        n28002), .B2(uart1_r_THOLD__7__3_), .Y(n27826) );
  AOI22xp33_ASAP7_75t_SL U31434 ( .A1(n28000), .A2(uart1_r_THOLD__11__1_), 
        .B1(uart1_r_THOLD__23__1_), .B2(n28001), .Y(n27397) );
  INVxp33_ASAP7_75t_SL U31435 ( .A(n28293), .Y(n28294) );
  NAND2xp33_ASAP7_75t_SL U31436 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__12_), .B(
        n29863), .Y(n28649) );
  AOI22xp33_ASAP7_75t_SL U31437 ( .A1(n27997), .A2(uart1_r_THOLD__13__6_), 
        .B1(uart1_r_THOLD__29__6_), .B2(n27996), .Y(n27622) );
  AOI22xp33_ASAP7_75t_SL U31438 ( .A1(n27997), .A2(uart1_r_THOLD__15__1_), 
        .B1(uart1_r_THOLD__31__1_), .B2(n27996), .Y(n27399) );
  NAND2xp33_ASAP7_75t_SL U31439 ( .A(n30161), .B(n30192), .Y(n24548) );
  NAND2xp33_ASAP7_75t_SL U31440 ( .A(n28180), .B(n30774), .Y(n28186) );
  NAND2xp5_ASAP7_75t_SL U31441 ( .A(n2992), .B(n25535), .Y(n25536) );
  OAI21xp33_ASAP7_75t_SL U31442 ( .A1(n25239), .A2(n25243), .B(n25242), .Y(
        n17285) );
  NAND2xp5_ASAP7_75t_SL U31443 ( .A(n24594), .B(n24603), .Y(n24596) );
  AOI22xp33_ASAP7_75t_SL U31444 ( .A1(n27997), .A2(uart1_r_THOLD__15__3_), 
        .B1(uart1_r_THOLD__31__3_), .B2(n27996), .Y(n27828) );
  INVxp67_ASAP7_75t_SL U31445 ( .A(n32054), .Y(n31382) );
  AOI22xp33_ASAP7_75t_SL U31446 ( .A1(uart1_r_THOLD__10__5_), .A2(n28009), 
        .B1(uart1_r_THOLD__2__5_), .B2(n28008), .Y(n27707) );
  AOI22xp33_ASAP7_75t_SL U31447 ( .A1(uart1_r_THOLD__10__3_), .A2(n28009), 
        .B1(uart1_r_THOLD__2__3_), .B2(n28008), .Y(n27831) );
  AOI22xp33_ASAP7_75t_SL U31448 ( .A1(uart1_r_THOLD__21__6_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__9__6_), .Y(n27624) );
  AOI22xp33_ASAP7_75t_SL U31449 ( .A1(n28009), .A2(uart1_r_THOLD__8__1_), .B1(
        uart1_r_THOLD__0__1_), .B2(n28008), .Y(n27413) );
  NAND4xp25_ASAP7_75t_SRAM U31450 ( .A(n31381), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), .C(n31380), .D(n31379), .Y(
        n31383) );
  AOI22xp33_ASAP7_75t_SL U31451 ( .A1(n28009), .A2(uart1_r_THOLD__10__1_), 
        .B1(uart1_r_THOLD__2__1_), .B2(n28008), .Y(n27418) );
  NAND2xp33_ASAP7_75t_SL U31452 ( .A(uart1_r_THOLD__6__5_), .B(n28015), .Y(
        n27703) );
  AOI22xp33_ASAP7_75t_SL U31453 ( .A1(uart1_r_THOLD__23__5_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__11__5_), .Y(n27699) );
  NAND2xp33_ASAP7_75t_SL U31454 ( .A(n26869), .B(n26868), .Y(n32090) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U31455 ( .A1(n32571), .A2(n32566), .B(n31551), .C(
        n31554), .Y(n31552) );
  AOI22xp33_ASAP7_75t_SL U31456 ( .A1(n27997), .A2(uart1_r_THOLD__13__0_), 
        .B1(uart1_r_THOLD__29__0_), .B2(n27996), .Y(n27980) );
  AOI22xp33_ASAP7_75t_SL U31457 ( .A1(uart1_r_THOLD__23__2_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__11__2_), .Y(n27892) );
  NAND2xp33_ASAP7_75t_SL U31458 ( .A(uart1_r_THOLD__30__0_), .B(n28018), .Y(
        n28019) );
  INVx1_ASAP7_75t_SL U31459 ( .A(n24681), .Y(n24663) );
  AOI22xp33_ASAP7_75t_SL U31460 ( .A1(n27997), .A2(uart1_r_THOLD__15__5_), 
        .B1(uart1_r_THOLD__31__5_), .B2(n27996), .Y(n27700) );
  AOI22xp33_ASAP7_75t_SL U31461 ( .A1(n27997), .A2(uart1_r_THOLD__15__2_), 
        .B1(uart1_r_THOLD__31__2_), .B2(n27996), .Y(n27891) );
  NAND2xp33_ASAP7_75t_SL U31462 ( .A(n27537), .B(n26089), .Y(n27534) );
  AOI22xp33_ASAP7_75t_SL U31463 ( .A1(uart1_r_THOLD__10__2_), .A2(n28009), 
        .B1(uart1_r_THOLD__2__2_), .B2(n28008), .Y(n27907) );
  AOI22xp33_ASAP7_75t_SL U31464 ( .A1(uart1_r_THOLD__8__5_), .A2(n28009), .B1(
        uart1_r_THOLD__0__5_), .B2(n28008), .Y(n27695) );
  AOI22xp33_ASAP7_75t_SL U31465 ( .A1(uart1_r_THOLD__3__2_), .A2(n28003), .B1(
        n28002), .B2(uart1_r_THOLD__7__2_), .Y(n27890) );
  INVx1_ASAP7_75t_SL U31466 ( .A(n29863), .Y(n30642) );
  AOI22xp33_ASAP7_75t_SL U31467 ( .A1(uart1_r_THOLD__10__0_), .A2(n28009), 
        .B1(uart1_r_THOLD__2__0_), .B2(n28008), .Y(n28013) );
  AOI22xp33_ASAP7_75t_SL U31468 ( .A1(uart1_r_THOLD__21__0_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__9__0_), .Y(n27982) );
  NAND2xp33_ASAP7_75t_SL U31469 ( .A(n25243), .B(n25242), .Y(n31939) );
  INVx1_ASAP7_75t_SL U31470 ( .A(n24681), .Y(n24648) );
  NAND2xp5_ASAP7_75t_SL U31471 ( .A(n25705), .B(n25075), .Y(n30958) );
  NAND2xp33_ASAP7_75t_SL U31472 ( .A(uart1_r_THOLD__4__3_), .B(n28015), .Y(
        n27839) );
  INVx1_ASAP7_75t_SL U31473 ( .A(n24681), .Y(n24662) );
  AOI22xp33_ASAP7_75t_SL U31474 ( .A1(n28008), .A2(uart1_r_THOLD__0__0_), .B1(
        uart1_r_THOLD__28__0_), .B2(n28018), .Y(n27989) );
  AOI22xp33_ASAP7_75t_SL U31475 ( .A1(uart1_r_THOLD__21__5_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__9__5_), .Y(n27691) );
  NAND2xp5_ASAP7_75t_SL U31476 ( .A(n31558), .B(n31554), .Y(n31556) );
  INVx1_ASAP7_75t_SL U31477 ( .A(n24681), .Y(n24661) );
  AOI22xp33_ASAP7_75t_SL U31478 ( .A1(uart1_r_THOLD__8__3_), .A2(n28009), .B1(
        uart1_r_THOLD__0__3_), .B2(n28008), .Y(n27843) );
  AOI22xp33_ASAP7_75t_SL U31479 ( .A1(uart1_r_THOLD__8__0_), .A2(n28009), .B1(
        uart1_r_THOLD__4__0_), .B2(n28015), .Y(n27990) );
  AOI22xp33_ASAP7_75t_SL U31480 ( .A1(uart1_r_THOLD__8__2_), .A2(n28009), .B1(
        uart1_r_THOLD__4__2_), .B2(n28015), .Y(n27903) );
  AOI22xp33_ASAP7_75t_SL U31481 ( .A1(n28008), .A2(uart1_r_THOLD__0__2_), .B1(
        uart1_r_THOLD__28__2_), .B2(n28018), .Y(n27902) );
  INVx1_ASAP7_75t_SL U31482 ( .A(n24681), .Y(n24659) );
  INVxp67_ASAP7_75t_SL U31483 ( .A(DP_OP_1196_128_7433_n266), .Y(
        DP_OP_1196_128_7433_n264) );
  OAI21xp5_ASAP7_75t_SL U31484 ( .A1(n2356), .A2(n31696), .B(n32717), .Y(
        n32709) );
  AND2x2_ASAP7_75t_SL U31485 ( .A(n24956), .B(n31574), .Y(n32270) );
  INVx1_ASAP7_75t_SL U31486 ( .A(timer0_N79), .Y(n24405) );
  NAND2xp5_ASAP7_75t_SL U31487 ( .A(sr1_r_SRHSEL_), .B(n32791), .Y(n31758) );
  NAND2xp5_ASAP7_75t_SL U31488 ( .A(n26464), .B(n26472), .Y(n28110) );
  OAI21xp5_ASAP7_75t_SL U31489 ( .A1(n24963), .A2(n25650), .B(n24962), .Y(
        n24985) );
  INVxp67_ASAP7_75t_SL U31490 ( .A(n25953), .Y(n25955) );
  INVxp33_ASAP7_75t_SL U31491 ( .A(n27065), .Y(n26675) );
  NAND2xp5_ASAP7_75t_SL U31492 ( .A(n24946), .B(n25671), .Y(n24949) );
  INVx1_ASAP7_75t_SL U31493 ( .A(n31400), .Y(n31342) );
  INVx1_ASAP7_75t_SL U31494 ( .A(n24682), .Y(n24680) );
  INVx1_ASAP7_75t_SL U31495 ( .A(n24681), .Y(n24647) );
  NAND3xp33_ASAP7_75t_SRAM U31496 ( .A(n29444), .B(n29443), .C(
        irqctrl0_r_ILEVEL__1_), .Y(n29451) );
  INVxp67_ASAP7_75t_SL U31497 ( .A(n25667), .Y(n25687) );
  INVxp67_ASAP7_75t_SL U31498 ( .A(DP_OP_1196_128_7433_n210), .Y(
        DP_OP_1196_128_7433_n208) );
  NAND2xp33_ASAP7_75t_SL U31499 ( .A(n25670), .B(n25231), .Y(n24947) );
  NAND2xp33_ASAP7_75t_SL U31500 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_), 
        .B(n25231), .Y(n24931) );
  INVx1_ASAP7_75t_SL U31501 ( .A(n27986), .Y(n28014) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31502 ( .A1(n25223), .A2(n32078), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), .C(n25222), .Y(n25224) );
  AOI22xp33_ASAP7_75t_SL U31503 ( .A1(uart1_r_THOLD__10__4_), .A2(n28009), 
        .B1(uart1_r_THOLD__2__4_), .B2(n28008), .Y(n27778) );
  INVxp33_ASAP7_75t_SL U31504 ( .A(n28018), .Y(n27774) );
  AOI22xp33_ASAP7_75t_SL U31505 ( .A1(uart1_r_THOLD__15__4_), .A2(n27997), 
        .B1(n27996), .B2(uart1_r_THOLD__31__4_), .Y(n27773) );
  AOI22xp33_ASAP7_75t_SL U31506 ( .A1(n28001), .A2(uart1_r_THOLD__23__4_), 
        .B1(uart1_r_THOLD__11__4_), .B2(n28000), .Y(n27768) );
  AOI22xp33_ASAP7_75t_SL U31507 ( .A1(n28008), .A2(uart1_r_THOLD__0__4_), .B1(
        uart1_r_THOLD__28__4_), .B2(n28018), .Y(n27761) );
  AOI22xp33_ASAP7_75t_SL U31508 ( .A1(uart1_r_THOLD__8__4_), .A2(n28009), .B1(
        uart1_r_THOLD__4__4_), .B2(n28015), .Y(n27762) );
  INVx1_ASAP7_75t_SL U31509 ( .A(n24681), .Y(n24668) );
  INVxp67_ASAP7_75t_SL U31510 ( .A(n28877), .Y(n25122) );
  AOI22xp33_ASAP7_75t_SL U31511 ( .A1(uart1_r_THOLD__13__4_), .A2(n27997), 
        .B1(n27996), .B2(uart1_r_THOLD__29__4_), .Y(n27758) );
  AOI22xp33_ASAP7_75t_SL U31512 ( .A1(n28001), .A2(uart1_r_THOLD__21__4_), 
        .B1(uart1_r_THOLD__9__4_), .B2(n28000), .Y(n27754) );
  INVxp67_ASAP7_75t_SL U31513 ( .A(n25176), .Y(n25497) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U31514 ( .A1(n32083), .A2(n32082), .B(n32081), .C(
        n32080), .Y(n32098) );
  INVxp33_ASAP7_75t_SL U31515 ( .A(n26087), .Y(n26088) );
  NAND2xp5_ASAP7_75t_SL U31516 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[0]), .B(n31697), 
        .Y(n25246) );
  INVx1_ASAP7_75t_SL U31517 ( .A(n24580), .Y(n27200) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31518 ( .A1(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_), .A2(n29711), .B(n29710), .C(
        n29709), .Y(n29712) );
  INVx1_ASAP7_75t_SL U31519 ( .A(n24681), .Y(n24665) );
  NAND2xp5_ASAP7_75t_SL U31520 ( .A(n28038), .B(n28037), .Y(n28039) );
  AOI22xp33_ASAP7_75t_SL U31521 ( .A1(uart1_r_THOLD__8__6_), .A2(n28009), .B1(
        uart1_r_THOLD__4__6_), .B2(n28015), .Y(n27630) );
  AOI22xp33_ASAP7_75t_SL U31522 ( .A1(n28008), .A2(uart1_r_THOLD__0__6_), .B1(
        uart1_r_THOLD__28__6_), .B2(n28018), .Y(n27629) );
  AOI22xp33_ASAP7_75t_SL U31523 ( .A1(n28000), .A2(uart1_r_THOLD__11__6_), 
        .B1(uart1_r_THOLD__23__6_), .B2(n28001), .Y(n27637) );
  AOI22xp33_ASAP7_75t_SL U31524 ( .A1(uart1_r_THOLD__10__6_), .A2(n28009), 
        .B1(uart1_r_THOLD__2__6_), .B2(n28008), .Y(n27641) );
  NAND2xp33_ASAP7_75t_SL U31525 ( .A(uart1_r_THOLD__30__6_), .B(n28018), .Y(
        n27642) );
  NAND2xp33_ASAP7_75t_SL U31526 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__4_), .B(
        n29863), .Y(n28861) );
  INVx1_ASAP7_75t_SL U31527 ( .A(n24681), .Y(n24664) );
  INVxp33_ASAP7_75t_SL U31528 ( .A(n25941), .Y(n27475) );
  AOI22xp33_ASAP7_75t_SL U31529 ( .A1(n31228), .A2(uart1_r_RHOLD__18__6_), 
        .B1(uart1_r_RHOLD__8__6_), .B2(n31227), .Y(n31232) );
  NOR2xp33_ASAP7_75t_SRAM U31530 ( .A(n27479), .B(n27460), .Y(n27461) );
  NAND2xp33_ASAP7_75t_SL U31531 ( .A(n25961), .B(n27459), .Y(n25956) );
  INVx1_ASAP7_75t_SL U31532 ( .A(n24681), .Y(n24667) );
  INVx1_ASAP7_75t_SL U31533 ( .A(n28934), .Y(n30612) );
  INVx1_ASAP7_75t_SL U31534 ( .A(n27771), .Y(n27998) );
  INVx1_ASAP7_75t_SL U31535 ( .A(n27985), .Y(n27999) );
  NAND2xp33_ASAP7_75t_SL U31536 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__13_), .B(
        n29863), .Y(n28603) );
  NAND2xp5_ASAP7_75t_SL U31537 ( .A(u0_0_leon3x0_p0_iu_r_E__CTRL__WICC_), .B(
        n27020), .Y(n29816) );
  NAND2xp33_ASAP7_75t_SL U31538 ( .A(n25586), .B(n31574), .Y(n25020) );
  INVxp33_ASAP7_75t_SL U31539 ( .A(n26574), .Y(n28737) );
  NAND2xp5_ASAP7_75t_SL U31540 ( .A(n29435), .B(n29436), .Y(n29633) );
  INVxp33_ASAP7_75t_SL U31541 ( .A(n29435), .Y(n29437) );
  INVxp33_ASAP7_75t_SL U31542 ( .A(n30806), .Y(n26502) );
  INVxp33_ASAP7_75t_SL U31543 ( .A(n29423), .Y(n29440) );
  AOI21xp33_ASAP7_75t_SL U31544 ( .A1(n29463), .A2(n29462), .B(n29461), .Y(
        n29464) );
  AOI21xp33_ASAP7_75t_SL U31545 ( .A1(n29459), .A2(n29458), .B(n29457), .Y(
        n29465) );
  INVx1_ASAP7_75t_SL U31546 ( .A(n24517), .Y(n22422) );
  NAND2xp5_ASAP7_75t_SL U31547 ( .A(u0_0_leon3x0_p0_div0_r_CNT__4_), .B(n24906), .Y(n31655) );
  NAND2xp5_ASAP7_75t_SL U31548 ( .A(n31664), .B(n28293), .Y(n31417) );
  AOI31xp33_ASAP7_75t_SRAM U31549 ( .A1(n25659), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), .A3(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__25_), .B(n25658), .Y(n25663) );
  INVxp33_ASAP7_75t_SL U31550 ( .A(n32289), .Y(n25409) );
  INVx3_ASAP7_75t_SL U31551 ( .A(n25491), .Y(n22423) );
  NAND2xp33_ASAP7_75t_SL U31552 ( .A(n32913), .B(n32909), .Y(n32910) );
  INVxp33_ASAP7_75t_SL U31553 ( .A(n24940), .Y(n24932) );
  NAND2xp33_ASAP7_75t_SL U31554 ( .A(n24926), .B(n24936), .Y(n24928) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31555 ( .A1(uart1_r_RIRQEN_), .A2(n1765), .B(
        n29361), .C(n31194), .Y(n29364) );
  AND2x4_ASAP7_75t_SL U31556 ( .A(n23531), .B(n23530), .Y(n23529) );
  INVx1_ASAP7_75t_SL U31557 ( .A(n30620), .Y(n25855) );
  NAND2xp33_ASAP7_75t_SL U31558 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__15_), 
        .B(n22376), .Y(n25166) );
  NAND2xp33_ASAP7_75t_SL U31559 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__7_), .B(
        n22376), .Y(n25167) );
  NOR2xp33_ASAP7_75t_SRAM U31560 ( .A(n31537), .B(n25681), .Y(n25683) );
  NAND2xp33_ASAP7_75t_SL U31561 ( .A(n32091), .B(n22379), .Y(n26826) );
  NAND2xp33_ASAP7_75t_SL U31562 ( .A(n31811), .B(n22379), .Y(n29670) );
  INVx1_ASAP7_75t_SL U31563 ( .A(n24681), .Y(n24674) );
  OAI21xp33_ASAP7_75t_SL U31564 ( .A1(n25665), .A2(n25655), .B(n25654), .Y(
        n25656) );
  INVxp67_ASAP7_75t_SL U31565 ( .A(n32048), .Y(n24845) );
  INVxp33_ASAP7_75t_SL U31566 ( .A(n25655), .Y(n25648) );
  NAND2xp5_ASAP7_75t_SL U31567 ( .A(n30804), .B(n30071), .Y(n29347) );
  INVx1_ASAP7_75t_SL U31568 ( .A(n31188), .Y(n30068) );
  NAND2xp33_ASAP7_75t_SL U31569 ( .A(n24858), .B(n32048), .Y(n25601) );
  AOI31xp33_ASAP7_75t_SRAM U31570 ( .A1(n25696), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__29_), .A3(n25695), .B(n25694), .Y(
        n25702) );
  AND4x1_ASAP7_75t_SL U31571 ( .A(n32717), .B(n32716), .C(n2356), .D(n2357), 
        .Y(n32718) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31572 ( .A1(n25666), .A2(n25698), .B(n25667), 
        .C(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), .Y(n25669) );
  NAND2xp33_ASAP7_75t_SL U31573 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__4_), .B(
        n29731), .Y(n29732) );
  INVxp67_ASAP7_75t_SL U31574 ( .A(DP_OP_1196_128_7433_n319), .Y(
        DP_OP_1196_128_7433_n317) );
  NAND2xp33_ASAP7_75t_SL U31575 ( .A(n26779), .B(n31862), .Y(n26803) );
  AOI22xp33_ASAP7_75t_SL U31576 ( .A1(n25583), .A2(n25582), .B1(n30197), .B2(
        n30192), .Y(n31579) );
  INVx1_ASAP7_75t_SL U31577 ( .A(n24681), .Y(n24675) );
  INVxp67_ASAP7_75t_SL U31578 ( .A(n29731), .Y(n29736) );
  AOI22xp33_ASAP7_75t_SL U31579 ( .A1(n31228), .A2(uart1_r_RHOLD__18__1_), 
        .B1(uart1_r_RHOLD__8__1_), .B2(n31227), .Y(n27453) );
  INVxp67_ASAP7_75t_SL U31580 ( .A(n32887), .Y(n32838) );
  NAND3xp33_ASAP7_75t_SRAM U31581 ( .A(n26791), .B(
        u0_0_leon3x0_p0_iu_r_X__RESULT__2_), .C(n29212), .Y(n26792) );
  NAND2xp33_ASAP7_75t_SL U31582 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__LD_), .B(
        n31868), .Y(n31869) );
  AOI21xp5_ASAP7_75t_SL U31583 ( .A1(n32887), .A2(n32913), .B(n32917), .Y(
        n32904) );
  NAND2xp33_ASAP7_75t_SL U31584 ( .A(n24937), .B(n24936), .Y(n24938) );
  NAND2xp33_ASAP7_75t_SL U31585 ( .A(n32496), .B(n32495), .Y(n32501) );
  NAND2xp33_ASAP7_75t_SL U31586 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__1_), .B(
        n29731), .Y(n25947) );
  NAND2xp33_ASAP7_75t_SL U31587 ( .A(n32482), .B(n32481), .Y(n32487) );
  INVxp33_ASAP7_75t_SL U31588 ( .A(n26190), .Y(n26194) );
  INVxp33_ASAP7_75t_SL U31589 ( .A(n26761), .Y(n26762) );
  INVxp67_ASAP7_75t_SL U31590 ( .A(n29964), .Y(n29965) );
  NAND2xp33_ASAP7_75t_SL U31591 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[1]), .B(n32474), .Y(n32479) );
  INVxp67_ASAP7_75t_SL U31592 ( .A(n31283), .Y(n30202) );
  NAND2xp33_ASAP7_75t_SL U31593 ( .A(n2927), .B(n32495), .Y(n32472) );
  NAND2xp5_ASAP7_75t_SL U31594 ( .A(n32489), .B(n32474), .Y(n32465) );
  OAI21xp5_ASAP7_75t_SL U31595 ( .A1(n26190), .A2(n26192), .B(
        u0_0_leon3x0_p0_iu_r_D__INULL_), .Y(n24883) );
  NAND2xp5_ASAP7_75t_SL U31596 ( .A(n3134), .B(n32289), .Y(n31461) );
  INVxp33_ASAP7_75t_SL U31597 ( .A(n31261), .Y(n31459) );
  NAND2xp5_ASAP7_75t_SL U31598 ( .A(n32138), .B(n32140), .Y(n31963) );
  NAND2xp33_ASAP7_75t_SL U31599 ( .A(n29702), .B(n30157), .Y(n30686) );
  NAND2xp33_ASAP7_75t_SL U31600 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__27_), 
        .B(n22376), .Y(n26337) );
  NAND2xp5_ASAP7_75t_SL U31601 ( .A(n25368), .B(n25367), .Y(n29472) );
  INVx1_ASAP7_75t_SL U31602 ( .A(n24681), .Y(n24672) );
  NAND2xp33_ASAP7_75t_SL U31603 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__2_), .B(
        n22376), .Y(n25494) );
  INVx1_ASAP7_75t_SL U31604 ( .A(n24681), .Y(n24669) );
  INVxp67_ASAP7_75t_SL U31605 ( .A(n32481), .Y(n25324) );
  AOI22xp33_ASAP7_75t_SL U31606 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__20_), 
        .A2(n29705), .B1(n29468), .B2(n25383), .Y(n29717) );
  INVx1_ASAP7_75t_SL U31607 ( .A(n24681), .Y(n24666) );
  NAND2xp33_ASAP7_75t_SL U31608 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__1_), .B(
        n22376), .Y(n25406) );
  INVx1_ASAP7_75t_SL U31609 ( .A(n24681), .Y(n24673) );
  INVxp33_ASAP7_75t_SL U31610 ( .A(n31323), .Y(n31324) );
  NAND2xp33_ASAP7_75t_SL U31611 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__24_), 
        .B(n22376), .Y(n26393) );
  NAND2xp33_ASAP7_75t_SL U31612 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__22_), 
        .B(n22376), .Y(n26217) );
  NAND2xp33_ASAP7_75t_SL U31613 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__20_), 
        .B(n22376), .Y(n26959) );
  NAND2xp33_ASAP7_75t_SL U31614 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__19_), 
        .B(n22376), .Y(n25753) );
  INVx2_ASAP7_75t_SL U31615 ( .A(n24051), .Y(n22425) );
  INVx2_ASAP7_75t_SL U31616 ( .A(n24049), .Y(n22426) );
  NAND2xp33_ASAP7_75t_SL U31617 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__17_), 
        .B(n22376), .Y(n26702) );
  NAND2xp33_ASAP7_75t_SL U31618 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__16_), 
        .B(n22376), .Y(n26444) );
  NAND2xp33_ASAP7_75t_SL U31619 ( .A(n3065), .B(n14803), .Y(n32565) );
  INVx1_ASAP7_75t_SL U31620 ( .A(n24681), .Y(n24671) );
  INVxp33_ASAP7_75t_SL U31621 ( .A(n25367), .Y(n25360) );
  INVxp67_ASAP7_75t_SL U31622 ( .A(n24718), .Y(n24715) );
  NAND2xp5_ASAP7_75t_SL U31623 ( .A(uart1_r_TRADDR__3_), .B(n27392), .Y(n27771) );
  INVx1_ASAP7_75t_SL U31624 ( .A(n27407), .Y(n28001) );
  NAND2xp5_ASAP7_75t_SL U31625 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__5_), 
        .B(n30179), .Y(n30181) );
  INVx1_ASAP7_75t_SL U31626 ( .A(n27409), .Y(n28003) );
  INVx1_ASAP7_75t_SL U31627 ( .A(n27410), .Y(n28002) );
  NAND2xp33_ASAP7_75t_SL U31628 ( .A(n4715), .B(n27426), .Y(n27437) );
  NAND2xp33_ASAP7_75t_SL U31629 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__22_), .B(
        n24428), .Y(n30269) );
  NAND2xp5_ASAP7_75t_SL U31630 ( .A(n27393), .B(n27392), .Y(n27985) );
  INVx1_ASAP7_75t_SL U31631 ( .A(n27405), .Y(n27996) );
  INVx1_ASAP7_75t_SL U31632 ( .A(n27408), .Y(n28000) );
  INVxp67_ASAP7_75t_SL U31633 ( .A(n25576), .Y(n25021) );
  INVx1_ASAP7_75t_SL U31634 ( .A(n26097), .Y(n26468) );
  NAND2xp33_ASAP7_75t_SL U31635 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_), 
        .B(n25680), .Y(n25655) );
  INVxp67_ASAP7_75t_SL U31636 ( .A(n29354), .Y(n29558) );
  AOI31xp33_ASAP7_75t_SRAM U31637 ( .A1(n25682), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_), .A3(n25881), .B(n25697), .Y(
        n25658) );
  NAND2xp33_ASAP7_75t_SL U31638 ( .A(n25670), .B(n25700), .Y(n24940) );
  NAND2xp5_ASAP7_75t_SL U31639 ( .A(n31980), .B(n25680), .Y(n25650) );
  INVxp67_ASAP7_75t_SL U31640 ( .A(n32753), .Y(n32752) );
  NAND2xp33_ASAP7_75t_SL U31641 ( .A(n31656), .B(n31420), .Y(n24886) );
  NOR2xp33_ASAP7_75t_SRAM U31642 ( .A(n32249), .B(n25399), .Y(n31261) );
  AOI22xp33_ASAP7_75t_SL U31643 ( .A1(u0_0_leon3x0_p0_divi[61]), .A2(n30430), 
        .B1(u0_0_leon3x0_p0_iu_r_W__S__Y__29_), .B2(n24428), .Y(n30228) );
  NAND2xp5_ASAP7_75t_SL U31644 ( .A(n24694), .B(n28180), .Y(n31188) );
  INVxp67_ASAP7_75t_SL U31645 ( .A(n29504), .Y(n28482) );
  INVx1_ASAP7_75t_SL U31646 ( .A(n30426), .Y(n31415) );
  NAND2xp33_ASAP7_75t_SL U31647 ( .A(n32157), .B(n26789), .Y(n26760) );
  NAND2xp5_ASAP7_75t_SL U31648 ( .A(n28824), .B(n26169), .Y(n28879) );
  AOI22xp33_ASAP7_75t_SL U31649 ( .A1(n30001), .A2(ahb0_r_HRDATAM__24_), .B1(
        ahb0_r_HRDATAS__24_), .B2(n30000), .Y(n26507) );
  NAND2xp33_ASAP7_75t_SL U31650 ( .A(n29696), .B(n25684), .Y(n29872) );
  INVxp33_ASAP7_75t_SL U31651 ( .A(n29698), .Y(n29224) );
  NAND2xp5_ASAP7_75t_SL U31652 ( .A(u0_0_leon3x0_p0_iu_r_W__S__ET_), .B(n33054), .Y(n26800) );
  NAND2xp33_ASAP7_75t_SL U31653 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__17_), .B(
        n24428), .Y(n30319) );
  INVxp33_ASAP7_75t_SL U31654 ( .A(n26789), .Y(n26794) );
  INVxp67_ASAP7_75t_SL U31655 ( .A(n25980), .Y(n25981) );
  NAND2xp33_ASAP7_75t_SL U31656 ( .A(n3704), .B(n24684), .Y(n31428) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U31657 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__3_), 
        .A2(n26137), .B(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__3_), .C(
        u0_0_leon3x0_p0_iu_r_X__MEXC_), .Y(n29889) );
  AOI22xp33_ASAP7_75t_SL U31658 ( .A1(n30001), .A2(ahb0_r_HRDATAM__12_), .B1(
        ahb0_r_HRDATAS__12_), .B2(n24574), .Y(n25420) );
  INVxp33_ASAP7_75t_SL U31659 ( .A(n27535), .Y(n27539) );
  NAND2xp5_ASAP7_75t_SL U31660 ( .A(n25451), .B(n25450), .Y(n26758) );
  INVxp33_ASAP7_75t_SL U31661 ( .A(n29966), .Y(n27531) );
  NOR3xp33_ASAP7_75t_SRAM U31662 ( .A(n31192), .B(uart1_v_RXDB__1_), .C(n29360), .Y(n29361) );
  INVxp33_ASAP7_75t_SL U31663 ( .A(DP_OP_1196_128_7433_n318), .Y(
        DP_OP_1196_128_7433_n316) );
  NAND4xp25_ASAP7_75t_SRAM U31664 ( .A(n29354), .B(n29353), .C(uart1_r_TIRQEN_), .D(n29352), .Y(n29355) );
  NAND2xp33_ASAP7_75t_SL U31665 ( .A(n25670), .B(n25230), .Y(n30957) );
  NAND2xp5_ASAP7_75t_SL U31666 ( .A(n30209), .B(n26137), .Y(n29733) );
  INVxp33_ASAP7_75t_SL U31667 ( .A(n25692), .Y(n25698) );
  OA21x2_ASAP7_75t_SRAM U31668 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__1_), 
        .A2(n33054), .B(n32153), .Y(rf_addr_w[1]) );
  AOI22xp33_ASAP7_75t_SL U31669 ( .A1(n30001), .A2(ahb0_r_HRDATAM__6_), .B1(
        ahb0_r_HRDATAS__6_), .B2(n30000), .Y(n25853) );
  NAND2xp5_ASAP7_75t_SL U31670 ( .A(n25731), .B(n33054), .Y(n25737) );
  INVxp33_ASAP7_75t_SL U31671 ( .A(n26778), .Y(n26779) );
  AOI22xp33_ASAP7_75t_SL U31672 ( .A1(n30001), .A2(ahb0_r_HRDATAM__5_), .B1(
        ahb0_r_HRDATAS__5_), .B2(n30000), .Y(n30004) );
  NAND2xp33_ASAP7_75t_SL U31673 ( .A(oen), .B(n32827), .Y(n32792) );
  INVxp67_ASAP7_75t_SL U31674 ( .A(n31192), .Y(n28235) );
  INVxp33_ASAP7_75t_SL U31675 ( .A(n31264), .Y(n32027) );
  NOR3xp33_ASAP7_75t_SRAM U31676 ( .A(n24961), .B(n24943), .C(n25670), .Y(
        n24926) );
  INVxp33_ASAP7_75t_SL U31677 ( .A(n32016), .Y(n32017) );
  INVxp33_ASAP7_75t_SL U31678 ( .A(n29951), .Y(n28028) );
  INVx1_ASAP7_75t_SL U31679 ( .A(n28680), .Y(n28771) );
  NOR2xp33_ASAP7_75t_SRAM U31680 ( .A(n32238), .B(n32237), .Y(n32240) );
  INVx1_ASAP7_75t_SL U31681 ( .A(n31325), .Y(n26071) );
  INVxp67_ASAP7_75t_SL U31682 ( .A(n24696), .Y(n24697) );
  NAND2xp33_ASAP7_75t_SL U31683 ( .A(n27428), .B(n27426), .Y(n27438) );
  NAND2xp33_ASAP7_75t_SL U31684 ( .A(uart1_v_RXDB__1_), .B(n29966), .Y(n27525)
         );
  NAND2xp5_ASAP7_75t_SL U31685 ( .A(uart1_r_TWADDR__4_), .B(n31325), .Y(n27321) );
  INVxp33_ASAP7_75t_SL U31686 ( .A(n31876), .Y(n25323) );
  OAI21xp33_ASAP7_75t_SRAM U31687 ( .A1(n32087), .A2(n31859), .B(n18815), .Y(
        n31860) );
  NOR2xp33_ASAP7_75t_SRAM U31688 ( .A(u0_0_leon3x0_p0_divo[31]), .B(n29109), 
        .Y(n29111) );
  AOI22xp33_ASAP7_75t_SL U31689 ( .A1(n25359), .A2(n30156), .B1(n25358), .B2(
        n25357), .Y(n25367) );
  INVxp33_ASAP7_75t_SL U31690 ( .A(n25357), .Y(n25361) );
  INVxp67_ASAP7_75t_SL U31691 ( .A(n26005), .Y(n26006) );
  INVxp33_ASAP7_75t_SL U31692 ( .A(n25230), .Y(n25668) );
  INVxp67_ASAP7_75t_SL U31693 ( .A(n1637), .Y(n25535) );
  NAND2xp5_ASAP7_75t_SL U31694 ( .A(n25984), .B(n26097), .Y(n25533) );
  NAND2xp5_ASAP7_75t_SL U31695 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__27_), 
        .B(n24708), .Y(n24709) );
  INVxp33_ASAP7_75t_SL U31696 ( .A(n27364), .Y(n27365) );
  INVxp33_ASAP7_75t_SL U31697 ( .A(n29421), .Y(n29405) );
  INVx1_ASAP7_75t_SL U31698 ( .A(n29865), .Y(n30644) );
  INVxp67_ASAP7_75t_SL U31699 ( .A(n26658), .Y(n31027) );
  INVxp33_ASAP7_75t_SL U31700 ( .A(n26195), .Y(n25174) );
  INVx1_ASAP7_75t_SL U31701 ( .A(n31396), .Y(n31336) );
  INVxp33_ASAP7_75t_SL U31702 ( .A(n27353), .Y(n27340) );
  INVxp33_ASAP7_75t_SL U31703 ( .A(n27333), .Y(n27334) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U31704 ( .A1(n32089), .A2(n32088), .B(n32087), 
        .C(n18815), .Y(n32092) );
  AOI211xp5_ASAP7_75t_SRAM U31705 ( .A1(n29705), .A2(n29703), .B(n29702), .C(
        n29706), .Y(n29713) );
  NAND2xp33_ASAP7_75t_SL U31706 ( .A(n32467), .B(n31876), .Y(n25333) );
  INVxp67_ASAP7_75t_SL U31707 ( .A(n27385), .Y(n27377) );
  NAND2xp5_ASAP7_75t_SL U31708 ( .A(n24694), .B(n27290), .Y(n29650) );
  INVxp67_ASAP7_75t_SL U31709 ( .A(n29391), .Y(n29654) );
  NOR2xp33_ASAP7_75t_SRAM U31710 ( .A(n32079), .B(n32078), .Y(n32080) );
  NOR2x1_ASAP7_75t_SL U31711 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__2_), .B(
        n25209), .Y(n31398) );
  INVxp33_ASAP7_75t_SL U31712 ( .A(n27369), .Y(n27361) );
  INVxp33_ASAP7_75t_SL U31713 ( .A(n27351), .Y(n27346) );
  INVxp33_ASAP7_75t_SL U31714 ( .A(n27338), .Y(n27330) );
  NAND2xp5_ASAP7_75t_SL U31715 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__0_), .B(
        n25079), .Y(n31400) );
  INVxp33_ASAP7_75t_SL U31716 ( .A(n30179), .Y(n30172) );
  INVx1_ASAP7_75t_SL U31717 ( .A(n24514), .Y(n22429) );
  INVx1_ASAP7_75t_SL U31718 ( .A(n27895), .Y(n27313) );
  INVxp33_ASAP7_75t_SL U31719 ( .A(n32826), .Y(n31710) );
  NAND2xp33_ASAP7_75t_SL U31720 ( .A(n30193), .B(n30195), .Y(n25578) );
  AOI21xp33_ASAP7_75t_SL U31721 ( .A1(n25576), .A2(u0_0_leon3x0_p0_dci[41]), 
        .B(u0_0_leon3x0_p0_dci[38]), .Y(n25577) );
  NOR2xp33_ASAP7_75t_SRAM U31722 ( .A(n31754), .B(n31753), .Y(n31711) );
  NAND2xp5_ASAP7_75t_SL U31723 ( .A(n22919), .B(n25919), .Y(n31664) );
  INVx1_ASAP7_75t_SL U31724 ( .A(n31721), .Y(n31720) );
  NAND2xp33_ASAP7_75t_SL U31725 ( .A(n25379), .B(n29701), .Y(n25387) );
  NAND2xp5_ASAP7_75t_SL U31726 ( .A(n32827), .B(n32826), .Y(n32828) );
  NAND2xp33_ASAP7_75t_SL U31727 ( .A(n25379), .B(n29706), .Y(n29468) );
  NOR2x1_ASAP7_75t_SL U31728 ( .A(n24979), .B(n32249), .Y(n31574) );
  INVxp33_ASAP7_75t_SL U31729 ( .A(n29452), .Y(n29454) );
  INVxp33_ASAP7_75t_SL U31730 ( .A(n29460), .Y(n29463) );
  INVxp33_ASAP7_75t_SL U31731 ( .A(n32097), .Y(n24999) );
  INVxp33_ASAP7_75t_SL U31732 ( .A(n25653), .Y(n25703) );
  NAND2xp5_ASAP7_75t_SL U31733 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ENABLE_), .B(
        n32564), .Y(n14803) );
  INVx1_ASAP7_75t_SL U31734 ( .A(n31740), .Y(n31760) );
  INVxp67_ASAP7_75t_SL U31735 ( .A(n32102), .Y(n31381) );
  INVx1_ASAP7_75t_SL U31736 ( .A(timer0_N91), .Y(n22430) );
  NAND2xp33_ASAP7_75t_SL U31737 ( .A(irqctrl0_r_ILEVEL__5_), .B(n29422), .Y(
        n29445) );
  INVxp33_ASAP7_75t_SL U31738 ( .A(n32886), .Y(n32836) );
  AOI21xp5_ASAP7_75t_SL U31739 ( .A1(n32087), .A2(n26815), .B(n32084), .Y(
        n25215) );
  NAND2xp33_ASAP7_75t_SL U31740 ( .A(n24613), .B(n24626), .Y(n24614) );
  NAND2xp33_ASAP7_75t_SL U31741 ( .A(n4388), .B(n24694), .Y(n32041) );
  NAND2xp33_ASAP7_75t_SL U31742 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(
        u0_0_leon3x0_p0_iu_v_A__CWP__1_), .Y(n26778) );
  NAND2xp33_ASAP7_75t_SL U31743 ( .A(n2926), .B(n25239), .Y(n17284) );
  OR2x2_ASAP7_75t_SL U31744 ( .A(n25985), .B(n12995), .Y(n31639) );
  NAND2xp33_ASAP7_75t_SL U31745 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__19_), 
        .B(n26753), .Y(n25605) );
  INVxp33_ASAP7_75t_SL U31746 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .Y(n29186) );
  INVxp33_ASAP7_75t_SL U31747 ( .A(n25558), .Y(n25564) );
  OAI21xp5_ASAP7_75t_SL U31748 ( .A1(irqctrl0_r_IFORCE__0__11_), .A2(
        irqctrl0_r_IPEND__11_), .B(n29412), .Y(n29433) );
  INVxp67_ASAP7_75t_SL U31749 ( .A(n26367), .Y(n26366) );
  INVxp67_ASAP7_75t_SL U31750 ( .A(n24944), .Y(n25649) );
  NAND2xp33_ASAP7_75t_SL U31751 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__0_), 
        .B(n25705), .Y(n24993) );
  INVxp67_ASAP7_75t_SL U31752 ( .A(n32772), .Y(n32767) );
  INVxp67_ASAP7_75t_SL U31753 ( .A(n29431), .Y(n29408) );
  INVxp33_ASAP7_75t_SL U31754 ( .A(n29429), .Y(n29410) );
  INVxp33_ASAP7_75t_SL U31755 ( .A(DP_OP_1196_128_7433_n129), .Y(
        DP_OP_1196_128_7433_n131) );
  OAI21xp33_ASAP7_75t_SL U31756 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[30]), .A2(
        n32656), .B(n32661), .Y(n31265) );
  INVxp33_ASAP7_75t_SL U31757 ( .A(DP_OP_1196_128_7433_n308), .Y(
        DP_OP_1196_128_7433_n310) );
  AOI21xp5_ASAP7_75t_SL U31758 ( .A1(n31668), .A2(n2811), .B(
        u0_0_leon3x0_p0_div0_r_ZERO2_), .Y(n29110) );
  NAND2xp5_ASAP7_75t_SL U31759 ( .A(n26790), .B(n26787), .Y(n26769) );
  NAND2xp5_ASAP7_75t_SL U31760 ( .A(n25412), .B(n24982), .Y(n25238) );
  NAND2xp5_ASAP7_75t_SL U31761 ( .A(n18842), .B(n30909), .Y(n30908) );
  INVxp33_ASAP7_75t_SL U31762 ( .A(n29746), .Y(n29748) );
  INVxp67_ASAP7_75t_SL U31763 ( .A(n31379), .Y(n26816) );
  NAND2xp5_ASAP7_75t_SL U31764 ( .A(n31754), .B(n4391), .Y(n24698) );
  NAND2xp5_ASAP7_75t_SL U31765 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), 
        .B(n25670), .Y(n24963) );
  NAND2xp5_ASAP7_75t_SL U31766 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), 
        .B(n31537), .Y(n25692) );
  NAND2xp5_ASAP7_75t_SL U31767 ( .A(n3132), .B(n32250), .Y(n25399) );
  NAND2xp5_ASAP7_75t_SL U31768 ( .A(u0_0_leon3x0_p0_iu_v_X__DCI__LOCK_), .B(
        n25604), .Y(n31264) );
  INVxp33_ASAP7_75t_SL U31769 ( .A(DP_OP_1196_128_7433_n122), .Y(
        DP_OP_1196_128_7433_n120) );
  INVxp67_ASAP7_75t_SL U31770 ( .A(DP_OP_1196_128_7433_n301), .Y(
        DP_OP_1196_128_7433_n299) );
  NAND2xp5_ASAP7_75t_SL U31771 ( .A(n31656), .B(n29112), .Y(n28292) );
  NAND3xp33_ASAP7_75t_SRAM U31772 ( .A(n31537), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_), .C(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__30_), .Y(n24922) );
  INVxp67_ASAP7_75t_SL U31773 ( .A(n27540), .Y(n26129) );
  NAND2xp5_ASAP7_75t_SL U31774 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_), 
        .B(n31962), .Y(n26195) );
  INVxp33_ASAP7_75t_SL U31775 ( .A(n25705), .Y(n25651) );
  NOR2xp33_ASAP7_75t_SRAM U31776 ( .A(n31962), .B(n31961), .Y(n32139) );
  NAND2xp5_ASAP7_75t_SL U31777 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .B(
        n25894), .Y(n26169) );
  NAND2xp33_ASAP7_75t_SL U31778 ( .A(uart1_r_RXTICK_), .B(n30804), .Y(n29335)
         );
  NAND3xp33_ASAP7_75t_SRAM U31779 ( .A(n30873), .B(uart1_uarto_TXEN_), .C(
        uart1_r_TFIFOIRQEN_), .Y(n29363) );
  NAND2xp33_ASAP7_75t_SL U31780 ( .A(uart1_r_TRADDR__2_), .B(n27395), .Y(
        n27410) );
  NAND2xp5_ASAP7_75t_SL U31781 ( .A(n30873), .B(n28045), .Y(n29354) );
  NAND2xp5_ASAP7_75t_SL U31782 ( .A(u0_0_leon3x0_p0_iu_de_icc_2_), .B(n24712), 
        .Y(n24713) );
  NAND2xp5_ASAP7_75t_SL U31783 ( .A(n22919), .B(u0_0_leon3x0_p0_div0_r_NEG_), 
        .Y(n31667) );
  INVx1_ASAP7_75t_SL U31784 ( .A(n25665), .Y(n29696) );
  NAND2xp33_ASAP7_75t_SRAM U31785 ( .A(n18842), .B(n32079), .Y(n23898) );
  NAND2xp5_ASAP7_75t_SL U31786 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__31_), 
        .B(n30909), .Y(n32097) );
  INVx1_ASAP7_75t_SL U31787 ( .A(n28824), .Y(n25403) );
  NOR2x1_ASAP7_75t_SL U31788 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__2_), .B(
        n28931), .Y(n25901) );
  NAND2xp5_ASAP7_75t_SL U31789 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), 
        .B(n24878), .Y(n32082) );
  NAND2xp5_ASAP7_75t_SL U31790 ( .A(n25159), .B(n25158), .Y(n25163) );
  INVxp33_ASAP7_75t_SL U31791 ( .A(n29112), .Y(n31653) );
  NAND2xp5_ASAP7_75t_SL U31792 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__1_), .B(
        n26872), .Y(n26732) );
  NAND2xp5_ASAP7_75t_SL U31793 ( .A(n25161), .B(n25160), .Y(n25162) );
  NAND2xp33_ASAP7_75t_SL U31794 ( .A(u0_0_leon3x0_p0_iu_r_A__DIVSTART_), .B(
        n31811), .Y(n28285) );
  INVxp67_ASAP7_75t_SL U31795 ( .A(n24852), .Y(n24853) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U31796 ( .A1(u0_0_leon3x0_p0_ici[60]), .A2(n32504), 
        .B(n31902), .C(n32677), .Y(n31903) );
  NAND2xp5_ASAP7_75t_SL U31797 ( .A(n27394), .B(n27395), .Y(n27409) );
  INVxp33_ASAP7_75t_SL U31798 ( .A(n29972), .Y(n27529) );
  NAND2xp5_ASAP7_75t_SL U31799 ( .A(n30905), .B(n24844), .Y(n32102) );
  NAND2xp5_ASAP7_75t_SL U31800 ( .A(n25554), .B(n29178), .Y(n25555) );
  INVxp67_ASAP7_75t_SL U31801 ( .A(n29419), .Y(n29407) );
  NOR2xp33_ASAP7_75t_SRAM U31802 ( .A(n4325), .B(n28372), .Y(n28373) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U31803 ( .A1(u0_0_leon3x0_p0_ici[60]), .A2(n32475), 
        .B(n31899), .C(n32677), .Y(n31900) );
  NAND2xp33_ASAP7_75t_SL U31804 ( .A(u0_0_leon3x0_p0_divi[31]), .B(n32012), 
        .Y(n23103) );
  OAI22xp33_ASAP7_75t_SL U31805 ( .A1(uart1_r_RXF__3_), .A2(n29944), .B1(
        uart1_r_TICK_), .B2(uart1_r_RXF__4_), .Y(n4677) );
  NAND3xp33_ASAP7_75t_SRAM U31806 ( .A(n29359), .B(uart1_r_IRQPEND_), .C(
        n30804), .Y(n29370) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U31807 ( .A1(u0_0_leon3x0_p0_ici[60]), .A2(n32463), 
        .B(n31898), .C(u0_0_leon3x0_p0_ici[61]), .Y(n31901) );
  OAI22xp33_ASAP7_75t_SL U31808 ( .A1(uart1_r_RXF__2_), .A2(n29944), .B1(
        uart1_r_TICK_), .B2(uart1_r_RXF__3_), .Y(n4679) );
  INVxp33_ASAP7_75t_SL U31809 ( .A(n29469), .Y(n29470) );
  NAND2xp33_ASAP7_75t_SL U31810 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_), 
        .B(n29817), .Y(n24726) );
  OAI22xp33_ASAP7_75t_SL U31811 ( .A1(uart1_r_RXF__1_), .A2(n29944), .B1(
        uart1_r_TICK_), .B2(uart1_r_RXF__2_), .Y(n4681) );
  INVx1_ASAP7_75t_SL U31812 ( .A(n26013), .Y(n26016) );
  NOR2xp33_ASAP7_75t_SRAM U31813 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), 
        .B(n32084), .Y(n32089) );
  INVxp33_ASAP7_75t_SL U31814 ( .A(n31964), .Y(n24707) );
  INVx1_ASAP7_75t_SL U31815 ( .A(n24541), .Y(n22432) );
  NAND2xp5_ASAP7_75t_SL U31816 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), 
        .B(n25675), .Y(n30956) );
  INVx1_ASAP7_75t_SL U31817 ( .A(n24873), .Y(n24727) );
  NOR2xp33_ASAP7_75t_SRAM U31818 ( .A(n32713), .B(n29708), .Y(n29703) );
  NAND2xp5_ASAP7_75t_SL U31819 ( .A(n24591), .B(n24606), .Y(n24593) );
  INVxp67_ASAP7_75t_SL U31820 ( .A(DP_OP_1196_128_7433_n327), .Y(
        DP_OP_1196_128_7433_n325) );
  INVx1_ASAP7_75t_SL U31821 ( .A(n31404), .Y(n30430) );
  NAND2xp5_ASAP7_75t_SL U31822 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__30_), 
        .B(n32051), .Y(n32091) );
  NAND2xp5_ASAP7_75t_SL U31823 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__1_), 
        .B(n24920), .Y(n24989) );
  INVx1_ASAP7_75t_SL U31824 ( .A(n30955), .Y(n24961) );
  NAND2xp5_ASAP7_75t_SL U31825 ( .A(timer0_vtimers_1__ENABLE_), .B(n24683), 
        .Y(n26463) );
  NAND2xp33_ASAP7_75t_SL U31826 ( .A(n30200), .B(n3055), .Y(n30201) );
  NAND2xp5_ASAP7_75t_SL U31827 ( .A(sr1_r_BSTATE__0_), .B(n31715), .Y(n31740)
         );
  NOR2x1_ASAP7_75t_SL U31828 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__0_), .B(
        n25208), .Y(n31391) );
  NAND2xp5_ASAP7_75t_SL U31829 ( .A(sr1_r_BSTATE__1_), .B(n31732), .Y(n31753)
         );
  NAND2x1_ASAP7_75t_SL U31830 ( .A(n25129), .B(n28824), .Y(n28830) );
  NAND2xp5_ASAP7_75t_SL U31831 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__1_), .B(
        n25074), .Y(n25209) );
  NAND2xp5_ASAP7_75t_SL U31832 ( .A(n4724), .B(n31724), .Y(n31714) );
  INVxp67_ASAP7_75t_SL U31833 ( .A(n25129), .Y(n25130) );
  NAND2xp5_ASAP7_75t_SL U31834 ( .A(n27355), .B(n27320), .Y(n27338) );
  INVx1_ASAP7_75t_SL U31835 ( .A(n25937), .Y(n26869) );
  NAND2xp33_ASAP7_75t_SL U31836 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), 
        .B(n32083), .Y(n25225) );
  INVx1_ASAP7_75t_SL U31837 ( .A(n29147), .Y(n24632) );
  INVx1_ASAP7_75t_SL U31838 ( .A(n28931), .Y(n29148) );
  NAND2xp5_ASAP7_75t_SL U31839 ( .A(uart1_r_TWADDR__2_), .B(n27320), .Y(n27333) );
  AND3x1_ASAP7_75t_SRAM U31840 ( .A(n25670), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_), .C(
        u0_0_leon3x0_p0_iu_v_E__ET_), .Y(n25666) );
  NAND2xp33_ASAP7_75t_SL U31841 ( .A(n24688), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__31_), .Y(n25124) );
  NAND2xp5_ASAP7_75t_SL U31842 ( .A(n2929), .B(n26501), .Y(n27477) );
  NAND2xp33_ASAP7_75t_SL U31843 ( .A(n24694), .B(n29960), .Y(n28187) );
  NAND2xp33_ASAP7_75t_SL U31844 ( .A(n3135), .B(n30204), .Y(n31578) );
  NAND2xp33_ASAP7_75t_SL U31845 ( .A(n31982), .B(n25356), .Y(n25358) );
  NAND2xp33_ASAP7_75t_SL U31846 ( .A(n32069), .B(n31441), .Y(n24705) );
  NAND2xp5_ASAP7_75t_SL U31847 ( .A(n2867), .B(n27536), .Y(n28189) );
  INVx2_ASAP7_75t_SL U31848 ( .A(n24527), .Y(n22433) );
  AOI22xp33_ASAP7_75t_SL U31849 ( .A1(n4752), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__PIL__1_), .B1(n4763), .B2(n30697), .Y(
        n25371) );
  NAND2xp5_ASAP7_75t_SL U31850 ( .A(n30980), .B(n26075), .Y(n25971) );
  INVxp33_ASAP7_75t_SL U31851 ( .A(DP_OP_1196_128_7433_n278), .Y(
        DP_OP_1196_128_7433_n280) );
  INVxp67_ASAP7_75t_SL U31852 ( .A(DP_OP_1196_128_7433_n271), .Y(
        DP_OP_1196_128_7433_n269) );
  NOR3xp33_ASAP7_75t_SRAM U31853 ( .A(n31848), .B(n2931), .C(n2929), .Y(n27474) );
  NAND2xp5_ASAP7_75t_SL U31854 ( .A(n3134), .B(n31594), .Y(n32249) );
  NAND2xp5_ASAP7_75t_SL U31855 ( .A(n31258), .B(n25586), .Y(n25587) );
  INVxp33_ASAP7_75t_SL U31856 ( .A(n26757), .Y(n26759) );
  NAND2xp33_ASAP7_75t_SL U31857 ( .A(u0_0_leon3x0_p0_iu_de_icc_0_), .B(n30952), 
        .Y(n30954) );
  NAND2xp33_ASAP7_75t_SL U31858 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__29_), 
        .B(n24685), .Y(n24546) );
  AOI22xp33_ASAP7_75t_SL U31859 ( .A1(uart1_uarto_SCALER__0_), .A2(n24608), 
        .B1(uart1_uarto_SCALER__1_), .B2(n24609), .Y(uart1_scaler_1_) );
  NAND2xp33_ASAP7_75t_SL U31860 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__6_), .B(n32583), .Y(n32591) );
  NAND2xp33_ASAP7_75t_SL U31861 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_), .B(
        n28965), .Y(n25120) );
  NOR3xp33_ASAP7_75t_SRAM U31862 ( .A(n25677), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__10_), .C(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__11_), .Y(n25678) );
  NAND2xp33_ASAP7_75t_SL U31863 ( .A(
        u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_), .B(n31883), .Y(n32562) );
  NAND2xp33_ASAP7_75t_SL U31864 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__18_), 
        .B(n29576), .Y(n25169) );
  OAI21xp33_ASAP7_75t_SL U31865 ( .A1(u0_0_leon3x0_p0_iu_r_E__ALUOP__2_), .A2(
        n26482), .B(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .Y(n28680) );
  NAND2xp33_ASAP7_75t_SL U31866 ( .A(read), .B(n32832), .Y(n32826) );
  NAND2xp33_ASAP7_75t_SL U31867 ( .A(n4517), .B(n29947), .Y(n29945) );
  NAND2xp5_ASAP7_75t_SL U31868 ( .A(n24617), .B(n24625), .Y(n24620) );
  NAND2xp33_ASAP7_75t_SL U31869 ( .A(n25177), .B(n29147), .Y(n28734) );
  INVx1_ASAP7_75t_SL U31870 ( .A(n25208), .Y(n25079) );
  NOR2x1_ASAP7_75t_SL U31871 ( .A(n28965), .B(n25123), .Y(n28894) );
  OAI21xp33_ASAP7_75t_SL U31872 ( .A1(n3068), .A2(n32033), .B(n31703), .Y(
        n32732) );
  NAND2xp5_ASAP7_75t_SL U31873 ( .A(n2933), .B(n32482), .Y(n32503) );
  NAND2xp5_ASAP7_75t_SL U31874 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__0_), 
        .B(n32583), .Y(n32566) );
  NAND2xp33_ASAP7_75t_SL U31875 ( .A(n32467), .B(n32482), .Y(n32510) );
  NOR2x1_ASAP7_75t_SL U31876 ( .A(n31848), .B(n27479), .Y(n31325) );
  INVxp33_ASAP7_75t_SL U31877 ( .A(n32771), .Y(n32779) );
  NAND2xp5_ASAP7_75t_SL U31878 ( .A(n3068), .B(n32244), .Y(n31303) );
  NAND2xp5_ASAP7_75t_SL U31879 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[1]), .B(n32496), 
        .Y(n32511) );
  OR2x2_ASAP7_75t_SL U31880 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUSEL__1_), .B(
        n25123), .Y(n30637) );
  INVxp33_ASAP7_75t_SL U31881 ( .A(DP_OP_1196_128_7433_n222), .Y(
        DP_OP_1196_128_7433_n224) );
  INVxp33_ASAP7_75t_SL U31882 ( .A(DP_OP_1196_128_7433_n245), .Y(
        DP_OP_1196_128_7433_n243) );
  INVxp67_ASAP7_75t_SL U31883 ( .A(n32238), .Y(n25006) );
  AOI22xp33_ASAP7_75t_SL U31884 ( .A1(timer0_r_SCALER__0_), .A2(n24627), .B1(
        timer0_r_SCALER__1_), .B2(n24628), .Y(timer0_scaler_1_) );
  NAND2xp5_ASAP7_75t_SL U31885 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__WY_), .B(
        n31389), .Y(n30446) );
  NAND2xp33_ASAP7_75t_SL U31886 ( .A(u0_0_leon3x0_p0_dci[41]), .B(n25583), .Y(
        n25581) );
  NAND2xp5_ASAP7_75t_SL U31887 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__31_), 
        .B(n25170), .Y(n25366) );
  INVxp33_ASAP7_75t_SL U31888 ( .A(DP_OP_1196_128_7433_n196), .Y(
        DP_OP_1196_128_7433_n198) );
  NAND2xp5_ASAP7_75t_SL U31889 ( .A(n32461), .B(n32482), .Y(n32490) );
  OR2x2_ASAP7_75t_SL U31890 ( .A(n2867), .B(n27536), .Y(n28180) );
  INVxp67_ASAP7_75t_SL U31891 ( .A(n30156), .Y(n30158) );
  INVxp67_ASAP7_75t_SL U31892 ( .A(DP_OP_1196_128_7433_n189), .Y(
        DP_OP_1196_128_7433_n187) );
  NOR2xp33_ASAP7_75t_SL U31893 ( .A(u0_0_leon3x0_p0_dci[37]), .B(n25583), .Y(
        n25574) );
  INVx1_ASAP7_75t_SL U31894 ( .A(n25961), .Y(n25635) );
  NAND2xp5_ASAP7_75t_SL U31895 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__WY_), .B(
        n26365), .Y(n30426) );
  NAND2xp5_ASAP7_75t_SL U31896 ( .A(n4715), .B(n27427), .Y(n27439) );
  NOR2xp33_ASAP7_75t_SL U31897 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_), 
        .B(n29708), .Y(n25379) );
  INVxp33_ASAP7_75t_SL U31898 ( .A(DP_OP_1196_128_7433_n252), .Y(
        DP_OP_1196_128_7433_n254) );
  NAND2xp5_ASAP7_75t_SL U31899 ( .A(n2931), .B(n31529), .Y(n26658) );
  INVx1_ASAP7_75t_SL U31900 ( .A(n29706), .Y(n25384) );
  NAND2xp5_ASAP7_75t_SL U31901 ( .A(n30204), .B(n30161), .Y(n30193) );
  INVxp67_ASAP7_75t_SL U31902 ( .A(DP_OP_1196_128_7433_n215), .Y(
        DP_OP_1196_128_7433_n213) );
  NAND2xp5_ASAP7_75t_SL U31903 ( .A(n3067), .B(n32570), .Y(n29995) );
  NAND2xp5_ASAP7_75t_SL U31904 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[1]), .B(n32467), 
        .Y(n31318) );
  NAND2xp33_ASAP7_75t_SL U31905 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__19_), 
        .B(n25362), .Y(n25363) );
  INVx1_ASAP7_75t_SL U31906 ( .A(n25382), .Y(n25364) );
  AND3x1_ASAP7_75t_SL U31907 ( .A(n25961), .B(n2925), .C(n26501), .Y(n25962)
         );
  INVxp67_ASAP7_75t_SL U31908 ( .A(n32482), .Y(n32459) );
  NAND2xp33_ASAP7_75t_SL U31909 ( .A(n27428), .B(n27427), .Y(n27450) );
  INVxp67_ASAP7_75t_SL U31910 ( .A(n31604), .Y(n24976) );
  INVx1_ASAP7_75t_SL U31911 ( .A(u0_0_leon3x0_p0_divo[22]), .Y(n28507) );
  INVxp33_ASAP7_75t_SL U31912 ( .A(n4371), .Y(n25951) );
  INVxp67_ASAP7_75t_SL U31913 ( .A(apbi[31]), .Y(n26474) );
  INVxp67_ASAP7_75t_SL U31914 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__24_), .Y(
        n29774) );
  INVx1_ASAP7_75t_SL U31915 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__22_), .Y(
        n26224) );
  INVx1_ASAP7_75t_SL U31916 ( .A(u0_0_leon3x0_p0_ici[85]), .Y(n31786) );
  XNOR2xp5_ASAP7_75t_SRAM U31917 ( .A(it_q[10]), .B(u0_0_leon3x0_p0_ici[72]), 
        .Y(n31918) );
  INVx1_ASAP7_75t_SL U31918 ( .A(u0_0_leon3x0_p0_mulo[6]), .Y(n26285) );
  INVx1_ASAP7_75t_SL U31919 ( .A(u0_0_leon3x0_p0_iu_r_E__SHLEFT_), .Y(n26140)
         );
  INVx1_ASAP7_75t_SL U31920 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[28]), .Y(n32654)
         );
  XNOR2xp5_ASAP7_75t_SRAM U31921 ( .A(it_q[9]), .B(u0_0_leon3x0_p0_ici[71]), 
        .Y(n31919) );
  NOR2xp33_ASAP7_75t_SRAM U31922 ( .A(uart1_r_RSHIFT__3_), .B(
        uart1_r_RSHIFT__1_), .Y(n28228) );
  INVxp67_ASAP7_75t_SL U31923 ( .A(uart1_r_RIRQEN_), .Y(n29346) );
  INVx1_ASAP7_75t_SL U31924 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__26_), .Y(n29801)
         );
  XNOR2xp5_ASAP7_75t_SRAM U31925 ( .A(it_q[13]), .B(u0_0_leon3x0_p0_ici[75]), 
        .Y(n31917) );
  INVx1_ASAP7_75t_SL U31926 ( .A(u0_0_leon3x0_p0_div0_v_ZERO2_), .Y(n31668) );
  INVx1_ASAP7_75t_SL U31927 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__0_), .Y(
        n31423) );
  INVxp67_ASAP7_75t_SL U31928 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__17_), .Y(
        n27271) );
  INVxp67_ASAP7_75t_SL U31929 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__14_), .Y(
        n27181) );
  INVxp67_ASAP7_75t_SL U31930 ( .A(timer0_r_RELOAD__5_), .Y(n25867) );
  NAND2xp5_ASAP7_75t_SL U31931 ( .A(u0_0_dbgo_OPTYPE__2_), .B(
        u0_0_dbgo_OPTYPE__5_), .Y(n25449) );
  XNOR2xp5_ASAP7_75t_SRAM U31932 ( .A(it_q[14]), .B(u0_0_leon3x0_p0_ici[76]), 
        .Y(n31910) );
  NOR2xp33_ASAP7_75t_SRAM U31933 ( .A(uart1_r_RSHIFT__0_), .B(
        uart1_r_RSHIFT__6_), .Y(n28227) );
  INVx1_ASAP7_75t_SL U31934 ( .A(u0_0_leon3x0_p0_iu_r_W__S__ICC__1_), .Y(
        n30669) );
  INVxp67_ASAP7_75t_SL U31935 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__6_), .Y(
        n31518) );
  INVx1_ASAP7_75t_SL U31936 ( .A(u0_0_leon3x0_p0_ici[76]), .Y(n31834) );
  INVx1_ASAP7_75t_SL U31937 ( .A(timer0_vtimers_1__RELOAD__24_), .Y(n26520) );
  INVx1_ASAP7_75t_SL U31938 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__5_), .Y(
        n29684) );
  INVx1_ASAP7_75t_SL U31939 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__31_), .Y(
        n31680) );
  INVx1_ASAP7_75t_SL U31940 ( .A(u0_0_leon3x0_p0_div0_r_X__27_), .Y(n28282) );
  INVx1_ASAP7_75t_SL U31941 ( .A(irqctrl0_r_IMASK__0__8_), .Y(n29409) );
  INVx1_ASAP7_75t_SL U31942 ( .A(u0_0_dbgo_OPTYPE__3_), .Y(n31984) );
  XNOR2xp5_ASAP7_75t_SRAM U31943 ( .A(it_q[21]), .B(u0_0_leon3x0_p0_ici[83]), 
        .Y(n31920) );
  NOR2xp33_ASAP7_75t_SRAM U31944 ( .A(uart1_r_RSHIFT__7_), .B(
        uart1_r_RSHIFT__4_), .Y(n28230) );
  INVxp33_ASAP7_75t_SL U31945 ( .A(u0_0_leon3x0_p0_iu_r_M__IRQEN2_), .Y(n30692) );
  INVx1_ASAP7_75t_SL U31946 ( .A(ahb0_r_CFGA11_), .Y(n30975) );
  INVxp67_ASAP7_75t_SL U31947 ( .A(u0_0_leon3x0_p0_ici[11]), .Y(n27183) );
  INVxp67_ASAP7_75t_SL U31948 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__16_), .Y(
        n27231) );
  NAND2xp5_ASAP7_75t_SL U31949 ( .A(n2929), .B(n2931), .Y(n27479) );
  INVx1_ASAP7_75t_SL U31950 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__22_), .Y(n28513)
         );
  INVx1_ASAP7_75t_SL U31951 ( .A(u0_0_leon3x0_p0_mulo[33]), .Y(n25273) );
  INVx1_ASAP7_75t_SL U31952 ( .A(u0_0_leon3x0_p0_iu_r_E__SHCNT__3_), .Y(n30817) );
  INVxp67_ASAP7_75t_SL U31953 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__26_), .Y(
        n28393) );
  INVx1_ASAP7_75t_SL U31954 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__2_), 
        .Y(n32668) );
  INVx1_ASAP7_75t_SL U31955 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[29]), .Y(n32656)
         );
  INVx1_ASAP7_75t_SL U31956 ( .A(u0_0_leon3x0_p0_mulo[43]), .Y(n25290) );
  INVx1_ASAP7_75t_SL U31957 ( .A(u0_0_leon3x0_p0_div0_r_X__13_), .Y(n28330) );
  INVxp67_ASAP7_75t_SL U31958 ( .A(uart1_r_IRQPEND_), .Y(n29345) );
  INVxp67_ASAP7_75t_SL U31959 ( .A(irqctrl0_r_IMASK__0__15_), .Y(n29386) );
  XNOR2xp5_ASAP7_75t_SRAM U31960 ( .A(it_q[15]), .B(u0_0_leon3x0_p0_ici[77]), 
        .Y(n31911) );
  INVxp67_ASAP7_75t_SL U31961 ( .A(u0_0_leon3x0_p0_divi[51]), .Y(n30292) );
  INVxp67_ASAP7_75t_SL U31962 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__24_), .Y(
        n29765) );
  INVx1_ASAP7_75t_SL U31963 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__7_), .Y(
        n30397) );
  INVx1_ASAP7_75t_SL U31964 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__23_), .Y(n28472)
         );
  INVx1_ASAP7_75t_SL U31965 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[44]), .Y(n30973)
         );
  INVx1_ASAP7_75t_SL U31966 ( .A(u0_0_leon3x0_p0_divo[31]), .Y(n31673) );
  INVx1_ASAP7_75t_SL U31967 ( .A(u0_0_leon3x0_p0_div0_r_X__3_), .Y(n29691) );
  INVxp67_ASAP7_75t_SL U31968 ( .A(timer0_r_RELOAD__4_), .Y(n25878) );
  INVx1_ASAP7_75t_SL U31969 ( .A(u0_0_leon3x0_p0_divo[23]), .Y(n28316) );
  INVx1_ASAP7_75t_SL U31970 ( .A(u0_0_leon3x0_p0_div0_r_X__12_), .Y(n27222) );
  INVxp67_ASAP7_75t_SL U31971 ( .A(irqctrl0_r_IMASK__0__1_), .Y(n27298) );
  INVx1_ASAP7_75t_SL U31972 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[30]), .Y(n32658)
         );
  INVxp67_ASAP7_75t_SL U31973 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[46]), .Y(n30527)
         );
  INVxp67_ASAP7_75t_SL U31974 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__14_), .Y(
        n27179) );
  INVx1_ASAP7_75t_SL U31975 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[35]), .Y(n32976)
         );
  INVx1_ASAP7_75t_SL U31976 ( .A(timer0_vtimers_1__RELOAD__12_), .Y(n26610) );
  INVxp33_ASAP7_75t_SL U31977 ( .A(uart1_r_BREAKIRQEN_), .Y(n29360) );
  INVx1_ASAP7_75t_SL U31978 ( .A(u0_0_leon3x0_p0_mulo[46]), .Y(n25296) );
  XNOR2xp5_ASAP7_75t_SRAM U31979 ( .A(it_q[8]), .B(u0_0_leon3x0_p0_ici[70]), 
        .Y(n31912) );
  INVx1_ASAP7_75t_SL U31980 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__3_), .Y(
        n32681) );
  INVx1_ASAP7_75t_SL U31981 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .Y(n25177) );
  INVxp67_ASAP7_75t_SL U31982 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__8_), .Y(n28754) );
  XNOR2xp5_ASAP7_75t_SRAM U31983 ( .A(it_q[27]), .B(u0_0_leon3x0_p0_ici[89]), 
        .Y(n31909) );
  NOR2xp33_ASAP7_75t_SRAM U31984 ( .A(uart1_r_RSHIFT__5_), .B(
        uart1_r_RSHIFT__2_), .Y(n28229) );
  INVxp33_ASAP7_75t_SL U31985 ( .A(uart1_r_TCNT__4_), .Y(n29352) );
  INVxp33_ASAP7_75t_SL U31986 ( .A(u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__0_), .Y(
        n24968) );
  XNOR2xp5_ASAP7_75t_SRAM U31987 ( .A(it_q[17]), .B(u0_0_leon3x0_p0_ici[79]), 
        .Y(n31913) );
  INVxp67_ASAP7_75t_SL U31988 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__13_), .Y(
        n28594) );
  XNOR2xp5_ASAP7_75t_SRAM U31989 ( .A(it_q[23]), .B(u0_0_leon3x0_p0_ici[85]), 
        .Y(n31908) );
  INVx1_ASAP7_75t_SL U31990 ( .A(u0_0_leon3x0_p0_divi[37]), .Y(n30413) );
  INVx1_ASAP7_75t_SL U31991 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[31]), .Y(n32661)
         );
  INVx1_ASAP7_75t_SL U31992 ( .A(u0_0_leon3x0_p0_ici[74]), .Y(n30533) );
  INVxp33_ASAP7_75t_SL U31993 ( .A(n4635), .Y(n31030) );
  INVx1_ASAP7_75t_SL U31994 ( .A(timer0_vtimers_1__RELOAD__7_), .Y(n30874) );
  INVx1_ASAP7_75t_SL U31995 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__18_), .Y(
        n28538) );
  XNOR2xp5_ASAP7_75t_SRAM U31996 ( .A(it_q[25]), .B(u0_0_leon3x0_p0_ici[87]), 
        .Y(n31907) );
  INVxp67_ASAP7_75t_SL U31997 ( .A(sr1_r_MCFG2__RMW_), .Y(n32741) );
  INVx1_ASAP7_75t_SL U31998 ( .A(timer0_vtimers_1__RELOAD__4_), .Y(n26639) );
  NAND2xp33_ASAP7_75t_SL U31999 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), .B(
        u0_0_leon3x0_p0_iu_r_X__ICC__1_), .Y(n30668) );
  INVx1_ASAP7_75t_SL U32000 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[5]), .Y(n32843) );
  INVx1_ASAP7_75t_SL U32001 ( .A(u0_0_leon3x0_p0_mulo[51]), .Y(n25306) );
  NAND2xp5_ASAP7_75t_SL U32002 ( .A(n4388), .B(apb0_r_STATE__0_), .Y(n12995)
         );
  INVxp33_ASAP7_75t_SL U32003 ( .A(n1634), .Y(n29859) );
  INVxp67_ASAP7_75t_SL U32004 ( .A(u0_0_leon3x0_p0_ici[23]), .Y(n28395) );
  INVx1_ASAP7_75t_SL U32005 ( .A(timer0_vtimers_1__RELOAD__10_), .Y(n26619) );
  XNOR2xp5_ASAP7_75t_SRAM U32006 ( .A(it_q[11]), .B(u0_0_leon3x0_p0_ici[73]), 
        .Y(n31914) );
  INVx1_ASAP7_75t_SL U32007 ( .A(u0_0_leon3x0_p0_mulo[20]), .Y(n27025) );
  INVx1_ASAP7_75t_SL U32008 ( .A(u0_0_leon3x0_p0_mulo[14]), .Y(n29096) );
  INVx1_ASAP7_75t_SL U32009 ( .A(u0_0_leon3x0_p0_divo[27]), .Y(n28304) );
  INVx1_ASAP7_75t_SL U32010 ( .A(timer0_vtimers_1__RELOAD__31_), .Y(n26477) );
  INVx1_ASAP7_75t_SL U32011 ( .A(sr1_r_MCFG2__RAMBANKSZ__1_), .Y(n32774) );
  INVxp67_ASAP7_75t_SL U32012 ( .A(dataout[19]), .Y(n32895) );
  INVxp67_ASAP7_75t_SL U32013 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__17_), .Y(
        n27284) );
  NAND2xp33_ASAP7_75t_SL U32014 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), .B(
        u0_0_leon3x0_p0_iu_r_X__ICC__2_), .Y(n29165) );
  INVxp67_ASAP7_75t_SL U32015 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__26_), .Y(
        n28389) );
  INVxp33_ASAP7_75t_SL U32016 ( .A(u0_0_leon3x0_p0_iu_r_E__YMSB_), .Y(n31406)
         );
  INVx1_ASAP7_75t_SL U32017 ( .A(apbi[41]), .Y(n25526) );
  INVxp67_ASAP7_75t_SL U32018 ( .A(u0_0_leon3x0_p0_divo[12]), .Y(n28648) );
  INVxp33_ASAP7_75t_SL U32019 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__19_), .Y(
        n27033) );
  INVx1_ASAP7_75t_SL U32020 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__5_), .Y(
        n29728) );
  INVx1_ASAP7_75t_SL U32021 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__13_), .Y(
        n30361) );
  INVx1_ASAP7_75t_SL U32022 ( .A(apbi[40]), .Y(n25525) );
  INVxp67_ASAP7_75t_SL U32023 ( .A(u0_0_leon3x0_p0_ici[25]), .Y(n28266) );
  INVxp67_ASAP7_75t_SL U32024 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__12_), .Y(
        n29619) );
  INVxp33_ASAP7_75t_SL U32025 ( .A(u0_0_leon3x0_p0_iu_r_X__MEXC_), .Y(n30209)
         );
  INVxp67_ASAP7_75t_SL U32026 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[17]), .Y(n26601)
         );
  INVxp67_ASAP7_75t_SL U32027 ( .A(dataout[18]), .Y(n32893) );
  INVx1_ASAP7_75t_SL U32028 ( .A(u0_0_leon3x0_p0_ici[73]), .Y(n30517) );
  INVxp33_ASAP7_75t_SL U32029 ( .A(n1771), .Y(n26662) );
  INVx1_ASAP7_75t_SL U32030 ( .A(u0_0_leon3x0_p0_div0_r_X__18_), .Y(n28320) );
  INVxp67_ASAP7_75t_SL U32031 ( .A(uart1_r_TSHIFT__2_), .Y(n28027) );
  INVxp67_ASAP7_75t_SL U32032 ( .A(dataout[17]), .Y(n32891) );
  INVxp33_ASAP7_75t_SL U32033 ( .A(u0_0_leon3x0_p0_iu_r_A__WOVF_), .Y(n29697)
         );
  INVxp67_ASAP7_75t_SL U32034 ( .A(irqctrl0_r_IMASK__0__10_), .Y(n29259) );
  INVx1_ASAP7_75t_SL U32035 ( .A(u0_0_leon3x0_p0_mulo[29]), .Y(n29023) );
  INVxp67_ASAP7_75t_SL U32036 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__16_), .Y(
        n27229) );
  INVxp67_ASAP7_75t_SL U32037 ( .A(apbi[16]), .Y(n26655) );
  INVx1_ASAP7_75t_SL U32038 ( .A(u0_0_leon3x0_p0_iu_r_A__JMPL_), .Y(n31810) );
  INVxp33_ASAP7_75t_SL U32039 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__LD_), .Y(
        n31866) );
  INVx1_ASAP7_75t_SL U32040 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__5_), .Y(
        n30418) );
  INVx1_ASAP7_75t_SL U32041 ( .A(u0_0_leon3x0_p0_divo[15]), .Y(n28333) );
  INVx1_ASAP7_75t_SL U32042 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__24_), .Y(
        n29782) );
  INVx1_ASAP7_75t_SL U32043 ( .A(timer0_vtimers_1__RELOAD__16_), .Y(n26659) );
  INVx1_ASAP7_75t_SL U32044 ( .A(u0_0_leon3x0_p0_div0_r_X__29_), .Y(n28298) );
  INVxp67_ASAP7_75t_SL U32045 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__20_), .Y(
        n30286) );
  INVx1_ASAP7_75t_SL U32046 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__2_), .Y(n25210) );
  INVx1_ASAP7_75t_SL U32047 ( .A(u0_0_leon3x0_p0_divo[29]), .Y(n28302) );
  INVx1_ASAP7_75t_SL U32048 ( .A(u0_0_leon3x0_p0_mulo[41]), .Y(n25286) );
  INVxp67_ASAP7_75t_SL U32049 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[49]), .Y(n30534)
         );
  INVxp67_ASAP7_75t_SL U32050 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[20]), .Y(n26448)
         );
  INVxp67_ASAP7_75t_SL U32051 ( .A(u0_0_leon3x0_p0_iu_r_W__S__PIL__1_), .Y(
        n27136) );
  INVx1_ASAP7_75t_SL U32052 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__6_), .Y(
        n30407) );
  INVx1_ASAP7_75t_SL U32053 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__27_), .Y(
        n26910) );
  INVxp33_ASAP7_75t_SL U32054 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__9_), .Y(n30124) );
  INVx1_ASAP7_75t_SL U32055 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__17_), .Y(
        n27279) );
  INVx1_ASAP7_75t_SL U32056 ( .A(u0_0_leon3x0_p0_divo[11]), .Y(n28697) );
  INVx1_ASAP7_75t_SL U32057 ( .A(u0_0_leon3x0_p0_div0_r_X__2_), .Y(n28357) );
  INVx1_ASAP7_75t_SL U32058 ( .A(u0_0_leon3x0_p0_mulo[2]), .Y(n29106) );
  INVxp67_ASAP7_75t_SL U32059 ( .A(u0_0_leon3x0_p0_iu_r_W__S__WIM__2_), .Y(
        n29196) );
  INVxp67_ASAP7_75t_SL U32060 ( .A(ahbso_0__HRDATA__9_), .Y(n32859) );
  INVxp67_ASAP7_75t_SL U32061 ( .A(dataout[16]), .Y(n32889) );
  INVxp67_ASAP7_75t_SL U32062 ( .A(apbi[28]), .Y(n31496) );
  INVx1_ASAP7_75t_SL U32063 ( .A(u0_0_leon3x0_p0_mulo[0]), .Y(n29107) );
  INVxp67_ASAP7_75t_SL U32064 ( .A(ahbso_0__HRDATA__15_), .Y(n32873) );
  INVx1_ASAP7_75t_SL U32065 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__20_), .Y(
        n27009) );
  INVx1_ASAP7_75t_SL U32066 ( .A(uart1_r_RSEMPTY_), .Y(n26075) );
  INVxp33_ASAP7_75t_SL U32067 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[63]), .Y(n31688)
         );
  INVx1_ASAP7_75t_SL U32068 ( .A(u0_0_leon3x0_p0_mulo[15]), .Y(n28563) );
  INVxp67_ASAP7_75t_SL U32069 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__31_), .Y(
        n31407) );
  INVxp67_ASAP7_75t_SL U32070 ( .A(ahbso_0__HRDATA__14_), .Y(n32870) );
  INVxp67_ASAP7_75t_SL U32071 ( .A(n4928), .Y(n26823) );
  INVx1_ASAP7_75t_SL U32072 ( .A(u0_0_leon3x0_p0_muli[10]), .Y(n31661) );
  INVx1_ASAP7_75t_SL U32073 ( .A(u0_0_leon3x0_p0_ici[71]), .Y(n30526) );
  INVxp67_ASAP7_75t_SL U32074 ( .A(irqctrl0_r_IFORCE__0__12_), .Y(n29244) );
  INVx1_ASAP7_75t_SL U32075 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__29_), .Y(
        n30224) );
  INVxp67_ASAP7_75t_SL U32076 ( .A(ahbso_0__HRDATA__11_), .Y(n32864) );
  INVx1_ASAP7_75t_SL U32077 ( .A(uart1_v_RXF__1_), .Y(n4783) );
  INVxp33_ASAP7_75t_SL U32078 ( .A(ahbso_0__HRDATA__13_), .Y(n32868) );
  INVx1_ASAP7_75t_SL U32079 ( .A(u0_0_leon3x0_p0_ici[70]), .Y(n30524) );
  INVx1_ASAP7_75t_SL U32080 ( .A(u0_0_leon3x0_p0_ici[68]), .Y(n32586) );
  INVx1_ASAP7_75t_SL U32081 ( .A(uart1_r_RXCLK__1_), .Y(n28181) );
  INVx1_ASAP7_75t_SL U32082 ( .A(sr1_r_BUSW__1_), .Y(n32833) );
  INVxp67_ASAP7_75t_SL U32083 ( .A(sr1_r_MCFG2__RAMWIDTH__1_), .Y(n32721) );
  INVx1_ASAP7_75t_SL U32084 ( .A(u0_0_leon3x0_p0_ici[61]), .Y(n32677) );
  NAND2xp5_ASAP7_75t_SL U32085 ( .A(uart1_r_RXCLK__0_), .B(uart1_r_TICK_), .Y(
        n28182) );
  INVxp33_ASAP7_75t_SL U32086 ( .A(ahbso_0__HRDATA__12_), .Y(n32866) );
  INVx1_ASAP7_75t_SL U32087 ( .A(u0_0_leon3x0_p0_iu_r_W__S__ICC__0_), .Y(
        n27018) );
  NOR2xp33_ASAP7_75t_SRAM U32088 ( .A(apbi[35]), .B(apbi[34]), .Y(n27476) );
  XNOR2xp5_ASAP7_75t_SRAM U32089 ( .A(it_q[12]), .B(u0_0_leon3x0_p0_ici[74]), 
        .Y(n31924) );
  INVxp67_ASAP7_75t_SL U32090 ( .A(dataout[23]), .Y(n32905) );
  XNOR2xp5_ASAP7_75t_SRAM U32091 ( .A(it_q[22]), .B(u0_0_leon3x0_p0_ici[84]), 
        .Y(n31923) );
  INVxp33_ASAP7_75t_SL U32092 ( .A(n4456), .Y(n30987) );
  INVxp67_ASAP7_75t_SL U32093 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__26_), .Y(
        n28391) );
  INVxp33_ASAP7_75t_SL U32094 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__1_), .Y(
        n32138) );
  INVxp33_ASAP7_75t_SL U32095 ( .A(n2271), .Y(n26505) );
  INVxp67_ASAP7_75t_SL U32096 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[48]), .Y(n30518)
         );
  INVx1_ASAP7_75t_SL U32097 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__21_), .Y(n28523)
         );
  XNOR2xp5_ASAP7_75t_SRAM U32098 ( .A(it_q[26]), .B(u0_0_leon3x0_p0_ici[88]), 
        .Y(n31922) );
  INVx1_ASAP7_75t_SL U32099 ( .A(u0_0_leon3x0_p0_mulo[40]), .Y(n25285) );
  INVx1_ASAP7_75t_SL U32100 ( .A(uart1_r_PARSEL_), .Y(n29950) );
  NAND2xp5_ASAP7_75t_SL U32101 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__30_), 
        .B(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__31_), .Y(n25151) );
  INVx2_ASAP7_75t_SL U32102 ( .A(uart1_r_RSHIFT__0_), .Y(n29956) );
  INVx1_ASAP7_75t_SL U32103 ( .A(u0_0_leon3x0_p0_mulo[47]), .Y(n25298) );
  INVx1_ASAP7_75t_SL U32104 ( .A(u0_0_leon3x0_p0_ici[75]), .Y(n30540) );
  INVxp67_ASAP7_75t_SL U32105 ( .A(u0_0_leon3x0_p0_ici[9]), .Y(n29829) );
  XNOR2xp5_ASAP7_75t_SRAM U32106 ( .A(it_q[16]), .B(u0_0_leon3x0_p0_ici[78]), 
        .Y(n31921) );
  INVx1_ASAP7_75t_SL U32107 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__21_), .Y(n31539)
         );
  XNOR2xp5_ASAP7_75t_SRAM U32108 ( .A(it_q[19]), .B(u0_0_leon3x0_p0_ici[81]), 
        .Y(n31927) );
  INVxp67_ASAP7_75t_SL U32109 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__28_), .Y(
        n28262) );
  INVx1_ASAP7_75t_SL U32110 ( .A(u0_0_leon3x0_p0_mulo[4]), .Y(n29104) );
  NAND2xp33_ASAP7_75t_SL U32111 ( .A(u0_0_leon3x0_p0_iu_r_W__S__CWP__0_), .B(
        u0_0_leon3x0_p0_iu_r_W__S__CWP__1_), .Y(n26790) );
  INVxp67_ASAP7_75t_SL U32112 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__12_), .Y(
        n28653) );
  INVx1_ASAP7_75t_SL U32113 ( .A(u0_0_leon3x0_p0_iu_r_X__NPC__2_), .Y(n25731)
         );
  INVxp33_ASAP7_75t_SL U32114 ( .A(n4517), .Y(n29946) );
  NAND2xp33_ASAP7_75t_SL U32115 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_), 
        .B(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_), .Y(n32015) );
  INVx1_ASAP7_75t_SL U32116 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__20_), .Y(n27013)
         );
  INVx1_ASAP7_75t_SL U32117 ( .A(u0_0_leon3x0_p0_iu_r_M__WCWP_), .Y(n26783) );
  INVx1_ASAP7_75t_SL U32118 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__0_), .Y(
        n32152) );
  INVxp67_ASAP7_75t_SL U32119 ( .A(u0_0_leon3x0_p0_ici[14]), .Y(n27273) );
  INVxp67_ASAP7_75t_SL U32120 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__7_), .Y(n25058) );
  INVx1_ASAP7_75t_SL U32121 ( .A(uart1_r_IRQCNT__3_), .Y(n29340) );
  INVx1_ASAP7_75t_SL U32122 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__2_), .Y(
        n29640) );
  INVxp67_ASAP7_75t_SL U32123 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_UNDERRUN_), 
        .Y(n25567) );
  INVx1_ASAP7_75t_SL U32124 ( .A(uart1_r_TPAR_), .Y(n29953) );
  INVxp33_ASAP7_75t_SL U32125 ( .A(n4518), .Y(n29947) );
  INVx1_ASAP7_75t_SL U32126 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__2_), .Y(
        n32155) );
  INVxp33_ASAP7_75t_SL U32127 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__11_), .Y(n30881) );
  NOR2xp33_ASAP7_75t_SRAM U32128 ( .A(uart1_r_RSHIFT__0_), .B(uart1_r_PAREN_), 
        .Y(n29972) );
  INVx1_ASAP7_75t_SL U32129 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__3_), .Y(
        n32156) );
  INVxp67_ASAP7_75t_SL U32130 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__1_), .Y(
        n26831) );
  INVxp33_ASAP7_75t_SL U32131 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__1_), 
        .Y(n32571) );
  INVx1_ASAP7_75t_SL U32132 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__6_), .Y(
        n32570) );
  NAND2xp33_ASAP7_75t_SL U32133 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), .B(
        u0_0_leon3x0_p0_iu_r_X__ICC__3_), .Y(n29811) );
  INVx1_ASAP7_75t_SL U32134 ( .A(u0_0_leon3x0_p0_iu_r_W__S__CWP__0_), .Y(
        n32157) );
  INVx1_ASAP7_75t_SL U32135 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__24_), .Y(n30251)
         );
  INVxp67_ASAP7_75t_SL U32136 ( .A(irqctrl0_r_IMASK__0__3_), .Y(n28246) );
  INVx1_ASAP7_75t_SL U32137 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__20_), .Y(n27088)
         );
  INVxp67_ASAP7_75t_SL U32138 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[15]), .Y(n28135)
         );
  INVxp33_ASAP7_75t_SL U32139 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__24_), .Y(
        n30255) );
  INVx1_ASAP7_75t_SL U32140 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__14_), .Y(
        n30351) );
  INVx1_ASAP7_75t_SL U32141 ( .A(u0_0_leon3x0_p0_iu_r_W__S__CWP__1_), .Y(
        n32158) );
  INVx1_ASAP7_75t_SL U32142 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[31]), .Y(n32942)
         );
  AND2x2_ASAP7_75t_SRAM U32143 ( .A(n4325), .B(n3725), .Y(n24899) );
  INVxp67_ASAP7_75t_SL U32144 ( .A(dataout[22]), .Y(n32901) );
  INVx1_ASAP7_75t_SL U32145 ( .A(n2925), .Y(n31848) );
  INVxp67_ASAP7_75t_SL U32146 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__1_), .Y(
        n31516) );
  INVxp33_ASAP7_75t_SL U32147 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__30_), 
        .Y(n24957) );
  INVx1_ASAP7_75t_SL U32148 ( .A(u0_0_leon3x0_p0_iu_r_W__S__CWP__2_), .Y(
        n32159) );
  INVx1_ASAP7_75t_SL U32149 ( .A(timer0_vtimers_1__RELOAD__17_), .Y(n26550) );
  INVxp67_ASAP7_75t_SL U32150 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__30_), .Y(
        n30583) );
  INVx1_ASAP7_75t_SL U32151 ( .A(u0_0_leon3x0_p0_ici[72]), .Y(n30506) );
  INVx1_ASAP7_75t_SL U32152 ( .A(u0_0_leon3x0_p0_divo[24]), .Y(n28310) );
  INVx1_ASAP7_75t_SL U32153 ( .A(u0_0_leon3x0_p0_divo[14]), .Y(n28334) );
  INVxp67_ASAP7_75t_SL U32154 ( .A(uart1_r_BRATE__0_), .Y(n28176) );
  INVxp67_ASAP7_75t_SL U32155 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__28_), .Y(
        n28264) );
  INVxp67_ASAP7_75t_SL U32156 ( .A(apbi[17]), .Y(n26547) );
  INVx1_ASAP7_75t_SL U32157 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__9_), .Y(
        n27129) );
  INVx1_ASAP7_75t_SL U32158 ( .A(u0_0_leon3x0_p0_mulo[27]), .Y(n26912) );
  INVxp67_ASAP7_75t_SL U32159 ( .A(dataout[21]), .Y(n32899) );
  INVx1_ASAP7_75t_SL U32160 ( .A(uart1_r_IRQCNT__0_), .Y(n29334) );
  INVxp67_ASAP7_75t_SL U32161 ( .A(n4701), .Y(n28031) );
  INVxp33_ASAP7_75t_SL U32162 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__2_), 
        .Y(n31551) );
  INVx1_ASAP7_75t_SL U32163 ( .A(timer0_vtimers_1__RELOAD__11_), .Y(n28121) );
  INVx1_ASAP7_75t_SL U32164 ( .A(timer0_vtimers_1__RESTART_), .Y(n26465) );
  INVxp67_ASAP7_75t_SL U32165 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[21]), .Y(n27287)
         );
  INVxp67_ASAP7_75t_SL U32166 ( .A(u0_0_leon3x0_p0_iu_r_W__S__ET_), .Y(n33055)
         );
  INVx1_ASAP7_75t_SL U32167 ( .A(u0_0_leon3x0_p0_iu_r_W__S__ICC__3_), .Y(
        n29812) );
  INVxp67_ASAP7_75t_SL U32168 ( .A(timer0_vtimers_1__LOAD_), .Y(n26464) );
  INVxp67_ASAP7_75t_SL U32169 ( .A(dataout[20]), .Y(n32897) );
  INVxp67_ASAP7_75t_SL U32170 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__29_), 
        .Y(n25543) );
  INVxp67_ASAP7_75t_SL U32171 ( .A(u0_0_leon3x0_p0_ici[27]), .Y(n30585) );
  INVx1_ASAP7_75t_SL U32172 ( .A(u0_0_leon3x0_p0_div0_r_X__26_), .Y(n28276) );
  NAND2xp33_ASAP7_75t_SL U32173 ( .A(n18819), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .Y(n32085) );
  INVx1_ASAP7_75t_SL U32174 ( .A(u0_0_leon3x0_p0_mulo[3]), .Y(n29105) );
  INVxp67_ASAP7_75t_SL U32175 ( .A(u0_0_leon3x0_p0_divo[0]), .Y(n29011) );
  INVx1_ASAP7_75t_SL U32176 ( .A(u0_0_leon3x0_p0_ici[60]), .Y(n32669) );
  INVx1_ASAP7_75t_SL U32177 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__4_), .Y(
        n30429) );
  INVx1_ASAP7_75t_SL U32178 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__20_), .Y(n32535) );
  INVx1_ASAP7_75t_SL U32179 ( .A(u0_0_leon3x0_p0_divi[35]), .Y(n30441) );
  INVxp67_ASAP7_75t_SL U32180 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__3_), .Y(
        n30440) );
  INVx1_ASAP7_75t_SL U32181 ( .A(n1765), .Y(n30804) );
  INVx1_ASAP7_75t_SL U32182 ( .A(n2924), .Y(n32761) );
  INVxp67_ASAP7_75t_SL U32183 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__12_), .Y(
        n28623) );
  INVxp67_ASAP7_75t_SL U32184 ( .A(n1769), .Y(n25388) );
  INVx1_ASAP7_75t_SL U32185 ( .A(n4838), .Y(n27194) );
  INVxp67_ASAP7_75t_SL U32186 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__TRAP_), .Y(
        n31444) );
  INVx1_ASAP7_75t_SL U32187 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__19_), .Y(n30296)
         );
  INVxp33_ASAP7_75t_SL U32188 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__14_), .Y(
        n27218) );
  INVx1_ASAP7_75t_SL U32189 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__22_), .Y(n32538) );
  INVx1_ASAP7_75t_SL U32190 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__ANNUL_), .Y(
        n25604) );
  INVx1_ASAP7_75t_SL U32191 ( .A(timer0_vtimers_1__RELOAD__2_), .Y(n26646) );
  INVxp67_ASAP7_75t_SL U32192 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__25_), 
        .Y(n25539) );
  INVxp67_ASAP7_75t_SL U32193 ( .A(irqctrl0_r_ILEVEL__5_), .Y(n29287) );
  INVxp67_ASAP7_75t_SL U32194 ( .A(address[18]), .Y(n33021) );
  INVx1_ASAP7_75t_SL U32195 ( .A(irqctrl0_r_IFORCE__0__6_), .Y(n29312) );
  INVx1_ASAP7_75t_SL U32196 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_), .Y(
        n31980) );
  INVx1_ASAP7_75t_SL U32197 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__29_), .Y(
        n32063) );
  INVx1_ASAP7_75t_SL U32198 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_), .Y(
        n25670) );
  INVx1_ASAP7_75t_SL U32199 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__21_), .Y(
        n25362) );
  INVxp33_ASAP7_75t_SL U32200 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__25_), 
        .Y(n25541) );
  INVxp67_ASAP7_75t_SL U32201 ( .A(address[17]), .Y(n33018) );
  INVx1_ASAP7_75t_SL U32202 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__4_), 
        .Y(n30174) );
  INVxp67_ASAP7_75t_SL U32203 ( .A(irqctrl0_r_IMASK__0__13_), .Y(n30805) );
  INVx1_ASAP7_75t_SL U32204 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__30_), .Y(
        n25170) );
  INVxp67_ASAP7_75t_SL U32205 ( .A(address[16]), .Y(n33015) );
  INVxp67_ASAP7_75t_SL U32206 ( .A(address[15]), .Y(n33012) );
  INVx1_ASAP7_75t_SL U32207 ( .A(u0_0_leon3x0_p0_muli[8]), .Y(n25172) );
  INVxp67_ASAP7_75t_SL U32208 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__21_), .Y(
        n27047) );
  INVxp67_ASAP7_75t_SL U32209 ( .A(n3046), .Y(n31451) );
  INVxp67_ASAP7_75t_SL U32210 ( .A(address[14]), .Y(n33009) );
  NAND2xp5_ASAP7_75t_SL U32211 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), 
        .B(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_), .Y(n25697) );
  INVx1_ASAP7_75t_SL U32212 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__23_), .Y(n32541) );
  INVxp67_ASAP7_75t_SL U32213 ( .A(address[12]), .Y(n33005) );
  INVx1_ASAP7_75t_SL U32214 ( .A(n4520), .Y(n33068) );
  INVx1_ASAP7_75t_SL U32215 ( .A(n3055), .Y(n33067) );
  INVx1_ASAP7_75t_SL U32216 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__16_), .Y(n30327)
         );
  INVx1_ASAP7_75t_SL U32217 ( .A(u0_0_leon3x0_p0_divo[20]), .Y(n28321) );
  INVxp67_ASAP7_75t_SL U32218 ( .A(address[4]), .Y(n32987) );
  INVx1_ASAP7_75t_SL U32219 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), .Y(
        n25695) );
  INVxp67_ASAP7_75t_SL U32220 ( .A(n3132), .Y(n25512) );
  NOR2xp33_ASAP7_75t_SL U32221 ( .A(n4316), .B(u0_0_leon3x0_p0_dci[1]), .Y(
        n32290) );
  INVxp67_ASAP7_75t_SL U32222 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__21_), .Y(
        n27045) );
  INVx1_ASAP7_75t_SL U32223 ( .A(u0_0_leon3x0_p0_mulo[45]), .Y(n25294) );
  NAND2xp33_ASAP7_75t_SL U32224 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_), 
        .B(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .Y(n24944) );
  INVx1_ASAP7_75t_SL U32225 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__15_), .Y(n30338)
         );
  INVxp67_ASAP7_75t_SL U32226 ( .A(u0_0_leon3x0_p0_ici[83]), .Y(n29036) );
  INVx1_ASAP7_75t_SL U32227 ( .A(n3134), .Y(n31586) );
  INVxp67_ASAP7_75t_SL U32228 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__16_), .Y(
        n26680) );
  INVxp67_ASAP7_75t_SL U32229 ( .A(irqctrl0_r_IMASK__0__6_), .Y(n29304) );
  INVx1_ASAP7_75t_SL U32230 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__2_), .Y(
        n28952) );
  INVx1_ASAP7_75t_SL U32231 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__14_), .Y(n30350)
         );
  INVx1_ASAP7_75t_SL U32232 ( .A(u0_0_leon3x0_p0_div0_r_X__16_), .Y(n27264) );
  INVxp33_ASAP7_75t_SL U32233 ( .A(n4385), .Y(n31855) );
  INVx1_ASAP7_75t_SL U32234 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__8_), .Y(
        n30730) );
  NAND2xp5_ASAP7_75t_SL U32235 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUSEL__1_), .Y(n29000) );
  INVx1_ASAP7_75t_SL U32236 ( .A(u0_0_leon3x0_p0_divo[18]), .Y(n28324) );
  INVxp67_ASAP7_75t_SL U32237 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__12_), .Y(
        n29825) );
  INVx1_ASAP7_75t_SL U32238 ( .A(u0_0_leon3x0_p0_dci[3]), .Y(n32236) );
  INVx1_ASAP7_75t_SL U32239 ( .A(apbi[15]), .Y(n29389) );
  NAND2xp33_ASAP7_75t_SL U32240 ( .A(ahb0_r_HTRANS__1_), .B(ahb0_r_DEFSLV_), 
        .Y(n31802) );
  INVx1_ASAP7_75t_SL U32241 ( .A(timer0_vtimers_1__RELOAD__8_), .Y(n26626) );
  INVxp67_ASAP7_75t_SL U32242 ( .A(uart1_r_TCNT__1_), .Y(n31851) );
  INVxp67_ASAP7_75t_SL U32243 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__21_), .Y(
        n27049) );
  NAND2xp5_ASAP7_75t_SL U32244 ( .A(ahb0_r_HTRANS__1_), .B(n4832), .Y(n32038)
         );
  INVx1_ASAP7_75t_SL U32245 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__14_), .Y(
        n29575) );
  INVx1_ASAP7_75t_SL U32246 ( .A(apbi[13]), .Y(n29236) );
  INVx1_ASAP7_75t_SL U32247 ( .A(timer0_vtimers_1__RELOAD__21_), .Y(n31852) );
  INVx1_ASAP7_75t_SL U32248 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__18_), .Y(
        n25815) );
  INVxp67_ASAP7_75t_SL U32249 ( .A(u0_0_leon3x0_p0_ici[82]), .Y(n29773) );
  INVx1_ASAP7_75t_SL U32250 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[2]), .Y(n32733) );
  INVxp67_ASAP7_75t_SL U32251 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__12_), .Y(
        n29049) );
  INVx1_ASAP7_75t_SL U32252 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__17_), .Y(
        n29576) );
  INVx1_ASAP7_75t_SL U32253 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__13_), .Y(
        n25881) );
  INVx1_ASAP7_75t_SL U32254 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[0]), .Y(n32713)
         );
  NAND2xp5_ASAP7_75t_SL U32255 ( .A(irqo[1]), .B(n3325), .Y(n29316) );
  INVxp67_ASAP7_75t_SL U32256 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__17_), .Y(
        n23551) );
  INVx1_ASAP7_75t_SL U32257 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__17_), .Y(n27257)
         );
  INVx1_ASAP7_75t_SL U32258 ( .A(u0_0_leon3x0_p0_muli[2]), .Y(n30458) );
  INVx1_ASAP7_75t_SL U32259 ( .A(u0_0_leon3x0_p0_div0_r_X__1_), .Y(n30463) );
  INVx1_ASAP7_75t_SL U32260 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[1]), .Y(n32734)
         );
  INVx1_ASAP7_75t_SL U32261 ( .A(irqo[0]), .Y(n28833) );
  INVx1_ASAP7_75t_SL U32262 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[11]), .Y(n32857)
         );
  INVxp67_ASAP7_75t_SL U32263 ( .A(irqctrl0_r_IFORCE__0__11_), .Y(n25965) );
  INVx1_ASAP7_75t_SL U32264 ( .A(apbi[21]), .Y(n31842) );
  INVxp67_ASAP7_75t_SL U32265 ( .A(u0_0_leon3x0_p0_ici[13]), .Y(n27235) );
  INVxp67_ASAP7_75t_SL U32266 ( .A(irqctrl0_r_ILEVEL__8_), .Y(n29270) );
  INVx1_ASAP7_75t_SL U32267 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[2]), .Y(n32602)
         );
  INVxp67_ASAP7_75t_SL U32268 ( .A(timer0_r_RELOAD__3_), .Y(n29511) );
  INVx1_ASAP7_75t_SL U32269 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__25_), .Y(n30247)
         );
  INVxp33_ASAP7_75t_SL U32270 ( .A(n4497), .Y(n31535) );
  INVx1_ASAP7_75t_SL U32271 ( .A(u0_0_leon3x0_p0_dci[5]), .Y(n31694) );
  INVx1_ASAP7_75t_SL U32272 ( .A(uart1_r_TRADDR__3_), .Y(n27393) );
  INVx1_ASAP7_75t_SL U32273 ( .A(n2933), .Y(n32467) );
  INVx1_ASAP7_75t_SL U32274 ( .A(timer0_vtimers_1__RELOAD__20_), .Y(n31532) );
  INVxp33_ASAP7_75t_SL U32275 ( .A(uart1_r_PAREN_), .Y(n28034) );
  INVx1_ASAP7_75t_SL U32276 ( .A(n2927), .Y(n32496) );
  INVx1_ASAP7_75t_SL U32277 ( .A(uart1_r_TRADDR__2_), .Y(n27394) );
  INVxp33_ASAP7_75t_SL U32278 ( .A(n1775), .Y(n31507) );
  INVx1_ASAP7_75t_SL U32279 ( .A(timer0_vtimers_1__RELOAD__0_), .Y(n26654) );
  INVxp67_ASAP7_75t_SL U32280 ( .A(u0_0_leon3x0_p0_iu_r_M__DIVZ_), .Y(n29467)
         );
  INVxp67_ASAP7_75t_SL U32281 ( .A(address[27]), .Y(n33050) );
  INVxp67_ASAP7_75t_SL U32282 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[19]), .Y(n26589)
         );
  INVx1_ASAP7_75t_SL U32283 ( .A(uart1_r_TRADDR__1_), .Y(n28016) );
  INVx1_ASAP7_75t_SL U32284 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__1_), 
        .Y(n32461) );
  INVxp67_ASAP7_75t_SL U32285 ( .A(address[26]), .Y(n33047) );
  INVxp67_ASAP7_75t_SL U32286 ( .A(address[25]), .Y(n33044) );
  INVxp67_ASAP7_75t_SL U32287 ( .A(n2963), .Y(n25013) );
  INVxp67_ASAP7_75t_SL U32288 ( .A(address[24]), .Y(n33041) );
  INVx1_ASAP7_75t_SL U32289 ( .A(u0_0_leon3x0_p0_mulo[16]), .Y(n27224) );
  INVx1_ASAP7_75t_SL U32290 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_), .Y(
        n31982) );
  INVxp33_ASAP7_75t_SL U32291 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), 
        .Y(n25356) );
  INVx1_ASAP7_75t_SL U32292 ( .A(u0_0_leon3x0_p0_divo[19]), .Y(n28323) );
  INVx1_ASAP7_75t_SL U32293 ( .A(u0_0_leon3x0_p0_iu_r_D__PV_), .Y(n30681) );
  INVx1_ASAP7_75t_SL U32294 ( .A(apbi[0]), .Y(n28108) );
  INVx1_ASAP7_75t_SL U32295 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DFRZ_), 
        .Y(n30012) );
  INVx1_ASAP7_75t_SL U32296 ( .A(timer0_vtimers_1__RELOAD__28_), .Y(n31504) );
  INVxp67_ASAP7_75t_SL U32297 ( .A(irqi_0__IRL__0_), .Y(n25370) );
  NAND2xp5_ASAP7_75t_SL U32298 ( .A(uart1_r_TRADDR__2_), .B(uart1_r_TRADDR__3_), .Y(n27390) );
  INVx1_ASAP7_75t_SL U32299 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__27_), .Y(n30238)
         );
  INVxp33_ASAP7_75t_SL U32300 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__20_), .Y(
        n26967) );
  INVx1_ASAP7_75t_SL U32301 ( .A(n4763), .Y(n29645) );
  INVxp67_ASAP7_75t_SL U32302 ( .A(uart1_r_RWADDR__1_), .Y(n26009) );
  INVx1_ASAP7_75t_SL U32303 ( .A(u0_0_leon3x0_p0_iu_v_X__DCI__SIGNED_), .Y(
        n25050) );
  INVx1_ASAP7_75t_SL U32304 ( .A(n3327), .Y(n30694) );
  INVx1_ASAP7_75t_SL U32305 ( .A(u0_0_leon3x0_p0_divi[34]), .Y(n30454) );
  INVx1_ASAP7_75t_SL U32306 ( .A(u0_0_leon3x0_p0_iu_r_W__S__PIL__0_), .Y(
        n30700) );
  OAI21xp33_ASAP7_75t_SL U32307 ( .A1(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .A2(
        u0_0_leon3x0_p0_iu_r_E__ALUOP__2_), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .Y(n25129) );
  INVx1_ASAP7_75t_SL U32308 ( .A(u0_0_leon3x0_p0_mulo[32]), .Y(n26350) );
  INVx1_ASAP7_75t_SL U32309 ( .A(u0_0_leon3x0_p0_muli[4]), .Y(n30428) );
  INVx1_ASAP7_75t_SL U32310 ( .A(n3328), .Y(n30697) );
  INVx1_ASAP7_75t_SL U32311 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__14_), .Y(
        n25115) );
  NAND2xp5_ASAP7_75t_SL U32312 ( .A(u0_0_leon3x0_p0_iu_v_M__IRQEN2_), .B(
        u0_0_leon3x0_p0_iu_r_M__IRQEN2_), .Y(n25377) );
  INVx1_ASAP7_75t_SL U32313 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__28_), .Y(n30234)
         );
  INVx1_ASAP7_75t_SL U32314 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__23_), .Y(n30262)
         );
  INVx1_ASAP7_75t_SL U32315 ( .A(n4774), .Y(n29882) );
  INVxp33_ASAP7_75t_SL U32316 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__16_), .Y(
        n26692) );
  INVx1_ASAP7_75t_SL U32317 ( .A(timer0_vtimers_1__RELOAD__1_), .Y(n26650) );
  INVx1_ASAP7_75t_SL U32318 ( .A(apbi[20]), .Y(n31526) );
  INVxp67_ASAP7_75t_SL U32319 ( .A(address[23]), .Y(n33037) );
  INVxp67_ASAP7_75t_SL U32320 ( .A(address[22]), .Y(n33034) );
  INVxp67_ASAP7_75t_SL U32321 ( .A(address[21]), .Y(n33030) );
  INVx1_ASAP7_75t_SL U32322 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[1]), .Y(n32489) );
  INVxp67_ASAP7_75t_SL U32323 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[24]), .Y(n31522)
         );
  INVx1_ASAP7_75t_SL U32324 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__20_), .Y(
        n29708) );
  INVxp33_ASAP7_75t_SL U32325 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__13_), .Y(
        n26160) );
  INVx1_ASAP7_75t_SL U32326 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__19_), .Y(
        n29705) );
  INVx1_ASAP7_75t_SL U32327 ( .A(u0_0_leon3x0_p0_mulo[12]), .Y(n29098) );
  NAND2xp5_ASAP7_75t_SL U32328 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__30_), 
        .B(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__31_), .Y(n25396) );
  INVxp67_ASAP7_75t_SL U32329 ( .A(u0_0_leon3x0_p0_dci[0]), .Y(n30797) );
  INVx1_ASAP7_75t_SL U32330 ( .A(sr1_r_MCFG2__RAMBANKSZ__0_), .Y(n32784) );
  INVx1_ASAP7_75t_SL U32331 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[39]), .Y(n31017)
         );
  INVx1_ASAP7_75t_SL U32332 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__16_), .Y(
        n28552) );
  INVxp67_ASAP7_75t_SL U32333 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__17_), .Y(
        n27255) );
  INVx1_ASAP7_75t_SL U32334 ( .A(timer0_vtimers_1__RELOAD__13_), .Y(n30803) );
  INVxp33_ASAP7_75t_SL U32335 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__4_), .Y(
        n30433) );
  INVxp67_ASAP7_75t_SL U32336 ( .A(address[20]), .Y(n33027) );
  INVx1_ASAP7_75t_SL U32337 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__4_), .Y(
        n31260) );
  INVx1_ASAP7_75t_SL U32338 ( .A(u0_0_leon3x0_p0_divi[45]), .Y(n30357) );
  INVx1_ASAP7_75t_SL U32339 ( .A(u0_0_leon3x0_p0_dci[2]), .Y(n31573) );
  INVxp67_ASAP7_75t_SL U32340 ( .A(address[19]), .Y(n33024) );
  INVxp33_ASAP7_75t_SL U32341 ( .A(n2846), .Y(n28089) );
  INVx1_ASAP7_75t_SL U32342 ( .A(uart1_r_TCNT__0_), .Y(n31531) );
  INVxp33_ASAP7_75t_SL U32343 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__21_), .Y(
        n26335) );
  INVxp67_ASAP7_75t_SL U32344 ( .A(u0_0_leon3x0_p0_ici[78]), .Y(n29043) );
  INVxp67_ASAP7_75t_SL U32345 ( .A(u0_0_leon3x0_p0_divi[38]), .Y(n30403) );
  INVx1_ASAP7_75t_SL U32346 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PV_), .Y(n30684) );
  INVx1_ASAP7_75t_SL U32347 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[14]), .Y(n32626)
         );
  INVxp67_ASAP7_75t_SL U32348 ( .A(apbi[29]), .Y(n26492) );
  INVx1_ASAP7_75t_SL U32349 ( .A(u0_0_leon3x0_p0_dci[38]), .Y(n25583) );
  INVx1_ASAP7_75t_SL U32350 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__15_), .Y(
        n28572) );
  INVxp67_ASAP7_75t_SL U32351 ( .A(u0_0_dbgo_SU_), .Y(n30118) );
  INVx1_ASAP7_75t_SL U32352 ( .A(n2386), .Y(n27445) );
  INVx1_ASAP7_75t_SL U32353 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[15]), .Y(n32628)
         );
  INVxp67_ASAP7_75t_SL U32354 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__17_), .Y(
        n27260) );
  INVx1_ASAP7_75t_SL U32355 ( .A(irqctrl0_r_IMASK__0__5_), .Y(n29404) );
  INVx1_ASAP7_75t_SL U32356 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[16]), .Y(n32630)
         );
  INVxp67_ASAP7_75t_SL U32357 ( .A(ramoen[2]), .Y(n32804) );
  INVxp67_ASAP7_75t_SL U32358 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__0_), 
        .Y(n32258) );
  INVx1_ASAP7_75t_SL U32359 ( .A(irqctrl0_r_IMASK__0__4_), .Y(n29402) );
  INVx1_ASAP7_75t_SL U32360 ( .A(u0_0_leon3x0_p0_dci[41]), .Y(n30204) );
  INVx1_ASAP7_75t_SL U32361 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__28_), .Y(
        n26916) );
  INVxp33_ASAP7_75t_SL U32362 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__5_), .Y(n26318) );
  INVx1_ASAP7_75t_SL U32363 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[17]), .Y(n32632)
         );
  INVxp67_ASAP7_75t_SL U32364 ( .A(irqctrl0_r_IFORCE__0__10_), .Y(n29266) );
  INVx1_ASAP7_75t_SL U32365 ( .A(u0_0_leon3x0_p0_div0_r_X__15_), .Y(n27223) );
  NAND2xp5_ASAP7_75t_SL U32366 ( .A(n2388), .B(n2387), .Y(n27469) );
  INVx1_ASAP7_75t_SL U32367 ( .A(u0_0_leon3x0_p0_ici[79]), .Y(n31765) );
  INVxp67_ASAP7_75t_SL U32368 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__16_), .Y(
        n27233) );
  INVx1_ASAP7_75t_SL U32369 ( .A(u0_0_dbgo_OPTYPE__0_), .Y(n26755) );
  INVx1_ASAP7_75t_SL U32370 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[6]), .Y(n32845) );
  INVxp33_ASAP7_75t_SL U32371 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__16_), .Y(
        n30331) );
  INVx1_ASAP7_75t_SL U32372 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[18]), .Y(n32634)
         );
  OAI21xp33_ASAP7_75t_SL U32373 ( .A1(irqctrl0_r_IPEND__6_), .A2(
        irqctrl0_r_IFORCE__0__6_), .B(irqctrl0_r_IMASK__0__6_), .Y(n29419) );
  INVxp67_ASAP7_75t_SL U32374 ( .A(irqctrl0_r_IPEND__2_), .Y(n29377) );
  INVx1_ASAP7_75t_SL U32375 ( .A(u0_0_leon3x0_p0_mulo[59]), .Y(n25319) );
  INVx1_ASAP7_75t_SL U32376 ( .A(irqctrl0_r_ILEVEL__6_), .Y(n29420) );
  INVxp67_ASAP7_75t_SL U32377 ( .A(u0_0_leon3x0_p0_ici[26]), .Y(n29577) );
  INVxp67_ASAP7_75t_SL U32378 ( .A(irqctrl0_r_IFORCE__0__2_), .Y(n29378) );
  INVx1_ASAP7_75t_SL U32379 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[19]), .Y(n32636)
         );
  INVxp33_ASAP7_75t_SL U32380 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__29_), .Y(
        n25417) );
  INVx1_ASAP7_75t_SL U32381 ( .A(n3133), .Y(n32445) );
  NOR2xp33_ASAP7_75t_SRAM U32382 ( .A(uart1_r_TCNT__3_), .B(uart1_r_TCNT__5_), 
        .Y(n29353) );
  INVxp67_ASAP7_75t_SL U32383 ( .A(u0_0_leon3x0_p0_ici[84]), .Y(n29034) );
  NAND2xp5_ASAP7_75t_SL U32384 ( .A(u0_0_leon3x0_p0_dci[40]), .B(
        u0_0_leon3x0_p0_dci[39]), .Y(n25575) );
  INVx1_ASAP7_75t_SL U32385 ( .A(u0_0_leon3x0_p0_mulo[36]), .Y(n25280) );
  INVx1_ASAP7_75t_SL U32386 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[20]), .Y(n32638)
         );
  INVx1_ASAP7_75t_SL U32387 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__17_), .Y(n30320)
         );
  NAND2xp33_ASAP7_75t_SL U32388 ( .A(irqctrl0_r_IMASK__0__12_), .B(
        irqctrl0_r_ILEVEL__12_), .Y(n29425) );
  NAND2xp5_ASAP7_75t_SL U32389 ( .A(uart1_r_RWADDR__0_), .B(uart1_r_RWADDR__1_), .Y(n26001) );
  INVx1_ASAP7_75t_SL U32390 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__IFRZ_), 
        .Y(n31467) );
  INVx1_ASAP7_75t_SL U32391 ( .A(u0_0_leon3x0_p0_mulo[9]), .Y(n27127) );
  INVxp67_ASAP7_75t_SL U32392 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__30_), .Y(
        n25887) );
  INVxp67_ASAP7_75t_SL U32393 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__27_), .Y(
        n26889) );
  INVx1_ASAP7_75t_SL U32394 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[21]), .Y(n32640)
         );
  INVx1_ASAP7_75t_SL U32395 ( .A(u0_0_leon3x0_p0_mulo[21]), .Y(n27037) );
  INVxp67_ASAP7_75t_SL U32396 ( .A(uart1_r_TSEMPTY_), .Y(n29366) );
  INVx1_ASAP7_75t_SL U32397 ( .A(n3067), .Y(n32437) );
  INVx1_ASAP7_75t_SL U32398 ( .A(u0_0_leon3x0_p0_iu_r_E__SHCNT__0_), .Y(n30487) );
  INVx1_ASAP7_75t_SL U32399 ( .A(irqctrl0_r_ILEVEL__3_), .Y(n29416) );
  INVx1_ASAP7_75t_SL U32400 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[22]), .Y(n32642)
         );
  INVxp67_ASAP7_75t_SL U32401 ( .A(u0_0_leon3x0_p0_divi[48]), .Y(n30323) );
  INVx1_ASAP7_75t_SL U32402 ( .A(u0_0_leon3x0_p0_divo[17]), .Y(n28327) );
  INVx1_ASAP7_75t_SL U32403 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[23]), .Y(n32644)
         );
  INVxp67_ASAP7_75t_SL U32404 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__30_), .Y(
        n30581) );
  NAND2xp5_ASAP7_75t_SL U32405 ( .A(uart1_r_TXCLK__0_), .B(uart1_r_TICK_), .Y(
        n26084) );
  INVxp67_ASAP7_75t_SL U32406 ( .A(ramoen[3]), .Y(n32812) );
  INVx1_ASAP7_75t_SL U32407 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[24]), .Y(n32646)
         );
  INVxp33_ASAP7_75t_SL U32408 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__2_), .Y(n28946) );
  INVx1_ASAP7_75t_SL U32409 ( .A(u0_0_leon3x0_p0_div0_r_X__0_), .Y(n28353) );
  INVxp67_ASAP7_75t_SL U32410 ( .A(u0_0_leon3x0_p0_divi[49]), .Y(n30313) );
  INVx1_ASAP7_75t_SL U32411 ( .A(u0_0_dbgo_OPTYPE__1_), .Y(n29212) );
  INVx1_ASAP7_75t_SL U32412 ( .A(u0_0_leon3x0_p0_ici[77]), .Y(n30828) );
  INVx1_ASAP7_75t_SL U32413 ( .A(apbi[10]), .Y(n30978) );
  INVx1_ASAP7_75t_SL U32414 ( .A(u0_0_leon3x0_p0_dci[4]), .Y(n32730) );
  INVxp33_ASAP7_75t_SL U32415 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__19_), 
        .Y(n24701) );
  INVx1_ASAP7_75t_SL U32416 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__0_), 
        .Y(n32150) );
  INVxp33_ASAP7_75t_SL U32417 ( .A(ramsn[3]), .Y(n32814) );
  INVx1_ASAP7_75t_SL U32418 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[25]), .Y(n32648)
         );
  INVx1_ASAP7_75t_SL U32419 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_NOMDS_), .Y(
        n25586) );
  INVxp67_ASAP7_75t_SL U32420 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__26_), .Y(
        n26236) );
  INVx1_ASAP7_75t_SL U32421 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__0_), .Y(
        n32148) );
  INVxp67_ASAP7_75t_SL U32422 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__12_), .Y(
        n29827) );
  INVxp67_ASAP7_75t_SL U32423 ( .A(u0_0_leon3x0_p0_ici[21]), .Y(n29776) );
  INVx1_ASAP7_75t_SL U32424 ( .A(u0_0_leon3x0_p0_mulo[37]), .Y(n25281) );
  INVx1_ASAP7_75t_SL U32425 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[26]), .Y(n32650)
         );
  INVx1_ASAP7_75t_SL U32426 ( .A(u0_0_leon3x0_p0_mulo[10]), .Y(n27168) );
  INVxp33_ASAP7_75t_SL U32427 ( .A(irqctrl0_r_IPEND__15_), .Y(n31024) );
  INVx1_ASAP7_75t_SL U32428 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__1_), .Y(
        n32145) );
  INVx1_ASAP7_75t_SL U32429 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[27]), .Y(n32652)
         );
  INVx1_ASAP7_75t_SL U32430 ( .A(irqctrl0_r_IMASK__0__12_), .Y(n29399) );
  INVx1_ASAP7_75t_SL U32431 ( .A(u0_0_leon3x0_p0_mulo[44]), .Y(n25292) );
  INVx1_ASAP7_75t_SL U32432 ( .A(u0_0_leon3x0_p0_mulo[56]), .Y(n25314) );
  INVx1_ASAP7_75t_SL U32433 ( .A(n4948), .Y(n33057) );
  INVxp67_ASAP7_75t_SL U32434 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), 
        .Y(n32010) );
  INVxp33_ASAP7_75t_SL U32435 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__WY_), .Y(
        n25274) );
  INVxp33_ASAP7_75t_SL U32436 ( .A(uart1_r_THOLD__12__2_), .Y(n27900) );
  INVx1_ASAP7_75t_SL U32437 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[3]), .Y(n32604)
         );
  INVxp67_ASAP7_75t_SL U32438 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__6_), .Y(
        n26241) );
  INVxp67_ASAP7_75t_SL U32439 ( .A(u0_0_leon3x0_p0_ici[18]), .Y(n27051) );
  INVxp67_ASAP7_75t_SL U32440 ( .A(u0_0_leon3x0_p0_ici[80]), .Y(n29040) );
  INVxp67_ASAP7_75t_SL U32441 ( .A(timer0_r_RELOAD__6_), .Y(n25864) );
  INVx1_ASAP7_75t_SL U32442 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__28_), .Y(
        n28271) );
  INVxp67_ASAP7_75t_SL U32443 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__6_), .Y(
        n26243) );
  INVx1_ASAP7_75t_SL U32444 ( .A(u0_0_leon3x0_p0_muli[5]), .Y(n30417) );
  INVxp67_ASAP7_75t_SL U32445 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__6_), .Y(
        n26245) );
  INVx1_ASAP7_75t_SL U32446 ( .A(u0_0_leon3x0_p0_div0_r_X__11_), .Y(n28335) );
  INVx1_ASAP7_75t_SL U32447 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[33]), .Y(n32958)
         );
  INVxp67_ASAP7_75t_SL U32448 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__23_), .Y(
        n29037) );
  INVxp67_ASAP7_75t_SL U32449 ( .A(ramoen[0]), .Y(n32793) );
  INVx1_ASAP7_75t_SL U32450 ( .A(u0_0_leon3x0_p0_dco_HIT_), .Y(n32244) );
  INVxp67_ASAP7_75t_SL U32451 ( .A(u0_0_leon3x0_p0_ici[3]), .Y(n26247) );
  INVx1_ASAP7_75t_SL U32452 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[4]), .Y(n32606)
         );
  NAND2xp5_ASAP7_75t_SL U32453 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__0_), 
        .B(u0_0_leon3x0_p0_c0mmu_dcache0_r_SIZE__1_), .Y(n32245) );
  INVx1_ASAP7_75t_SL U32454 ( .A(u0_0_leon3x0_p0_div0_r_X__17_), .Y(n28322) );
  INVxp67_ASAP7_75t_SL U32455 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__19_), .Y(
        n25768) );
  INVx1_ASAP7_75t_SL U32456 ( .A(u0_0_leon3x0_p0_mulo[28]), .Y(n28277) );
  INVx1_ASAP7_75t_SL U32457 ( .A(u0_0_leon3x0_p0_mulo[1]), .Y(n26752) );
  INVx1_ASAP7_75t_SL U32458 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[5]), .Y(n32608)
         );
  INVxp67_ASAP7_75t_SL U32459 ( .A(irqctrl0_r_IFORCE__0__8_), .Y(n29274) );
  INVx1_ASAP7_75t_SL U32460 ( .A(u0_0_leon3x0_p0_div0_r_X__5_), .Y(n29906) );
  INVx1_ASAP7_75t_SL U32461 ( .A(u0_0_leon3x0_p0_divo[28]), .Y(n28303) );
  INVxp67_ASAP7_75t_SL U32462 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__12_), .Y(
        n30371) );
  INVx1_ASAP7_75t_SL U32463 ( .A(u0_0_leon3x0_p0_mulo[13]), .Y(n27191) );
  INVx1_ASAP7_75t_SL U32464 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[6]), .Y(n32610)
         );
  INVx1_ASAP7_75t_SL U32465 ( .A(u0_0_leon3x0_p0_divo[13]), .Y(n28336) );
  INVxp67_ASAP7_75t_SL U32466 ( .A(u0_0_leon3x0_p0_ici[81]), .Y(n29066) );
  INVxp67_ASAP7_75t_SL U32467 ( .A(u0_0_leon3x0_p0_divi[43]), .Y(n30377) );
  INVx1_ASAP7_75t_SL U32468 ( .A(irqctrl0_r_ILEVEL__10_), .Y(n30984) );
  INVx1_ASAP7_75t_SL U32469 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[7]), .Y(n32612)
         );
  INVxp67_ASAP7_75t_SL U32470 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__9_), .Y(n27175) );
  INVx1_ASAP7_75t_SL U32471 ( .A(u0_0_leon3x0_p0_div0_r_X__6_), .Y(n29924) );
  INVx1_ASAP7_75t_SL U32472 ( .A(u0_0_leon3x0_p0_mulo[5]), .Y(n29102) );
  INVx1_ASAP7_75t_SL U32473 ( .A(timer0_vtimers_1__RELOAD__29_), .Y(n29988) );
  INVxp67_ASAP7_75t_SL U32474 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__30_), .Y(
        n30215) );
  INVx1_ASAP7_75t_SL U32475 ( .A(u0_0_leon3x0_p0_divo[16]), .Y(n28329) );
  INVx1_ASAP7_75t_SL U32476 ( .A(timer0_vtimers_1__RELOAD__5_), .Y(n30106) );
  INVx1_ASAP7_75t_SL U32477 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[8]), .Y(n32614)
         );
  INVxp67_ASAP7_75t_SL U32478 ( .A(u0_0_leon3x0_p0_dci[37]), .Y(n30119) );
  INVx1_ASAP7_75t_SL U32479 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__30_), .Y(n30594)
         );
  OAI21xp5_ASAP7_75t_SL U32480 ( .A1(irqctrl0_r_IPEND__9_), .A2(
        irqctrl0_r_IFORCE__0__9_), .B(irqctrl0_r_IMASK__0__9_), .Y(n29429) );
  INVx1_ASAP7_75t_SL U32481 ( .A(irqctrl0_r_ILEVEL__9_), .Y(n29430) );
  INVx1_ASAP7_75t_SL U32482 ( .A(u0_0_leon3x0_p0_div0_r_X__4_), .Y(n29692) );
  INVx1_ASAP7_75t_SL U32483 ( .A(u0_0_leon3x0_p0_mulo[52]), .Y(n25307) );
  INVxp67_ASAP7_75t_SL U32484 ( .A(uart1_r_RWADDR__0_), .Y(n28193) );
  INVx1_ASAP7_75t_SL U32485 ( .A(u0_0_leon3x0_p0_divi[44]), .Y(n30372) );
  INVx1_ASAP7_75t_SL U32486 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[9]), .Y(n32616)
         );
  INVxp33_ASAP7_75t_SL U32487 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__13_), .Y(
        n26181) );
  INVxp67_ASAP7_75t_SL U32488 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__17_), .Y(
        n27258) );
  INVx1_ASAP7_75t_SL U32489 ( .A(u0_0_leon3x0_p0_iu_v_E__SU_), .Y(n29219) );
  INVx1_ASAP7_75t_SL U32490 ( .A(u0_0_leon3x0_p0_divo[21]), .Y(n28319) );
  INVxp33_ASAP7_75t_SL U32491 ( .A(uart1_r_PARERR_), .Y(n30065) );
  INVxp33_ASAP7_75t_SL U32492 ( .A(u0_0_leon3x0_p0_iu_r_W__S__Y__14_), .Y(
        n30354) );
  INVxp67_ASAP7_75t_SL U32493 ( .A(u0_0_leon3x0_p0_dci[39]), .Y(n25585) );
  INVx1_ASAP7_75t_SL U32494 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__30_), .Y(
        n30574) );
  INVx1_ASAP7_75t_SL U32495 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[10]), .Y(n32618)
         );
  OAI21xp5_ASAP7_75t_SL U32496 ( .A1(irqctrl0_r_IPEND__14_), .A2(
        irqctrl0_r_IFORCE__0__14_), .B(irqctrl0_r_IMASK__0__14_), .Y(n29631)
         );
  INVx1_ASAP7_75t_SL U32497 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[11]), .Y(n32620)
         );
  INVx1_ASAP7_75t_SL U32498 ( .A(irqctrl0_r_ILEVEL__14_), .Y(n30552) );
  INVx1_ASAP7_75t_SL U32499 ( .A(n4715), .Y(n27428) );
  INVx1_ASAP7_75t_SL U32500 ( .A(apbi[11]), .Y(n28116) );
  INVx1_ASAP7_75t_SL U32501 ( .A(u0_0_leon3x0_p0_mulo[7]), .Y(n29101) );
  OAI21xp5_ASAP7_75t_SL U32502 ( .A1(irqctrl0_r_IPEND__15_), .A2(
        irqctrl0_r_IFORCE__0__15_), .B(irqctrl0_r_IMASK__0__15_), .Y(n29632)
         );
  INVx1_ASAP7_75t_SL U32503 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__7_), .Y(
        n29898) );
  INVxp67_ASAP7_75t_SL U32504 ( .A(ramoen[1]), .Y(n32797) );
  INVx1_ASAP7_75t_SL U32505 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[12]), .Y(n32622)
         );
  INVxp67_ASAP7_75t_SL U32506 ( .A(u0_0_leon3x0_p0_ici[10]), .Y(n28596) );
  INVx1_ASAP7_75t_SL U32507 ( .A(irqctrl0_r_ILEVEL__15_), .Y(n29428) );
  INVx1_ASAP7_75t_SL U32508 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__13_), .Y(
        n28593) );
  INVx1_ASAP7_75t_SL U32509 ( .A(timer0_vtimers_1__RELOAD__15_), .Y(n31021) );
  INVxp67_ASAP7_75t_SL U32510 ( .A(timer0_r_RELOAD__2_), .Y(n29518) );
  OAI21xp5_ASAP7_75t_SL U32511 ( .A1(irqctrl0_r_IPEND__13_), .A2(
        irqctrl0_r_IFORCE__0__13_), .B(irqctrl0_r_IMASK__0__13_), .Y(n29629)
         );
  INVxp33_ASAP7_75t_SL U32512 ( .A(ramsn[1]), .Y(n32798) );
  INVx1_ASAP7_75t_SL U32513 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[13]), .Y(n32624)
         );
  INVx1_ASAP7_75t_SL U32514 ( .A(irqctrl0_r_ILEVEL__13_), .Y(n29426) );
  INVx1_ASAP7_75t_SL U32515 ( .A(u0_0_leon3x0_p0_iu_r_E__JMPL_), .Y(n31812) );
  INVxp67_ASAP7_75t_SL U32516 ( .A(u0_0_leon3x0_p0_divi[46]), .Y(n30346) );
  INVx1_ASAP7_75t_SL U32517 ( .A(u0_0_leon3x0_p0_muli[0]), .Y(n30610) );
  INVx1_ASAP7_75t_SL U32518 ( .A(u0_0_leon3x0_p0_iu_r_E__CTRL__WICC_), .Y(
        n30952) );
  INVx1_ASAP7_75t_SL U32519 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__25_), .Y(
        n30248) );
  INVx1_ASAP7_75t_SL U32520 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__22_), .Y(
        n28509) );
  INVxp33_ASAP7_75t_SL U32521 ( .A(n4363), .Y(n32007) );
  INVx1_ASAP7_75t_SL U32522 ( .A(oen), .Y(n31752) );
  INVxp67_ASAP7_75t_SL U32523 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__19_), .Y(
        n25745) );
  INVxp67_ASAP7_75t_SL U32524 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[12]), .Y(n30521)
         );
  INVx1_ASAP7_75t_SL U32525 ( .A(u0_0_leon3x0_p0_mulo[34]), .Y(n25278) );
  INVx1_ASAP7_75t_SL U32526 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[40]), .Y(n30800)
         );
  INVxp67_ASAP7_75t_SL U32527 ( .A(irqctrl0_r_IFORCE__0__4_), .Y(n29321) );
  INVxp67_ASAP7_75t_SL U32528 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[13]), .Y(n30131)
         );
  INVxp67_ASAP7_75t_SL U32529 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__3_), .Y(
        n26837) );
  INVx1_ASAP7_75t_SL U32530 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[3]), .Y(n31703) );
  INVx1_ASAP7_75t_SL U32531 ( .A(timer0_r_DISHLT_), .Y(n30147) );
  INVxp67_ASAP7_75t_SL U32532 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[23]), .Y(n26539)
         );
  INVxp67_ASAP7_75t_SL U32533 ( .A(apbi[25]), .Y(n31368) );
  INVx1_ASAP7_75t_SL U32534 ( .A(uart1_r_RCNT__5_), .Y(n30980) );
  INVx1_ASAP7_75t_SL U32535 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__4_), .Y(
        n30920) );
  INVxp67_ASAP7_75t_SL U32536 ( .A(u0_0_leon3x0_p0_divo[25]), .Y(n28452) );
  NAND2xp5_ASAP7_75t_SL U32537 ( .A(uart1_r_TWADDR__0_), .B(uart1_r_TWADDR__1_), .Y(n27373) );
  INVx1_ASAP7_75t_SL U32538 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[27]), .Y(n31997)
         );
  INVxp67_ASAP7_75t_SL U32539 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[55]), .Y(n31774)
         );
  NAND2xp33_ASAP7_75t_SL U32540 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__0_), .Y(n24740) );
  INVxp67_ASAP7_75t_SL U32541 ( .A(uart1_r_THOLD__4__3_), .Y(n27792) );
  INVxp67_ASAP7_75t_SL U32542 ( .A(sr1_r_MCFG1__ROMWWS__2_), .Y(n31195) );
  INVxp33_ASAP7_75t_SL U32543 ( .A(n4614), .Y(n31331) );
  INVx1_ASAP7_75t_SL U32544 ( .A(n2926), .Y(n25243) );
  INVxp67_ASAP7_75t_SL U32545 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__WY_), .Y(
        n31385) );
  INVx1_ASAP7_75t_SL U32546 ( .A(u0_0_leon3x0_p0_div0_r_X__20_), .Y(n28306) );
  INVxp67_ASAP7_75t_SL U32547 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[51]), .Y(n31835)
         );
  INVxp67_ASAP7_75t_SL U32548 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__18_), .Y(
        n25719) );
  INVx1_ASAP7_75t_SL U32549 ( .A(n2972), .Y(n31999) );
  INVxp67_ASAP7_75t_SL U32550 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__19_), .Y(
        n25747) );
  INVx1_ASAP7_75t_SL U32551 ( .A(ahb0_r_HADDR__9_), .Y(n25412) );
  INVx1_ASAP7_75t_SL U32552 ( .A(apbi[22]), .Y(n31641) );
  INVxp67_ASAP7_75t_SL U32553 ( .A(uart1_r_THOLD__7__7_), .Y(n27571) );
  INVxp33_ASAP7_75t_SL U32554 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__WREG_), .Y(
        n30925) );
  INVx1_ASAP7_75t_SL U32555 ( .A(u0_0_leon3x0_p0_mulo[35]), .Y(n25279) );
  INVx1_ASAP7_75t_SL U32556 ( .A(ahb0_r_HADDR__6_), .Y(n25240) );
  INVxp67_ASAP7_75t_SL U32557 ( .A(sr1_r_MCFG1__ROMWWS__3_), .Y(n30868) );
  INVxp67_ASAP7_75t_SL U32558 ( .A(uart1_r_THOLD__7__6_), .Y(n27612) );
  INVx1_ASAP7_75t_SL U32559 ( .A(ahb0_r_HADDR__7_), .Y(n25241) );
  INVxp67_ASAP7_75t_SL U32560 ( .A(uart1_r_THOLD__5__3_), .Y(n27796) );
  INVx1_ASAP7_75t_SL U32561 ( .A(uart1_r_TWADDR__2_), .Y(n27355) );
  INVx1_ASAP7_75t_SL U32562 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__3_), .Y(
        n30923) );
  INVx1_ASAP7_75t_SL U32563 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__0_), .Y(
        n26819) );
  INVx1_ASAP7_75t_SL U32564 ( .A(ahb0_r_HADDR__5_), .Y(n31949) );
  INVxp33_ASAP7_75t_SL U32565 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[62]), .Y(n31691)
         );
  INVxp67_ASAP7_75t_SL U32566 ( .A(uart1_r_THOLD__7__5_), .Y(n27680) );
  INVxp67_ASAP7_75t_SL U32567 ( .A(uart1_r_THOLD__6__7_), .Y(n27567) );
  INVx1_ASAP7_75t_SL U32568 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__5_), .Y(n28815)
         );
  INVxp67_ASAP7_75t_SL U32569 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__19_), .Y(
        n25749) );
  INVx1_ASAP7_75t_SL U32570 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__2_), .Y(n32169)
         );
  INVx1_ASAP7_75t_SL U32571 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__11_), .Y(
        n28699) );
  NAND2xp5_ASAP7_75t_SL U32572 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .Y(n26815) );
  INVxp67_ASAP7_75t_SL U32573 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__0_), .Y(
        n29231) );
  INVxp67_ASAP7_75t_SL U32574 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_), 
        .Y(n30907) );
  INVx1_ASAP7_75t_SL U32575 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__0_), .Y(
        n30927) );
  INVx1_ASAP7_75t_SL U32576 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[0]), .Y(n32033) );
  INVxp67_ASAP7_75t_SL U32577 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[47]), .Y(n30511)
         );
  INVxp67_ASAP7_75t_SL U32578 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__14_), 
        .Y(n24789) );
  INVx1_ASAP7_75t_SL U32579 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__18_), .Y(
        n25813) );
  INVxp67_ASAP7_75t_SL U32580 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RD__5_), .Y(
        n31514) );
  INVxp67_ASAP7_75t_SL U32581 ( .A(uart1_r_THOLD__7__4_), .Y(n27744) );
  INVxp67_ASAP7_75t_SL U32582 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__31_), .Y(
        n26721) );
  INVxp67_ASAP7_75t_SL U32583 ( .A(uart1_r_THOLD__6__3_), .Y(n27812) );
  INVxp67_ASAP7_75t_SL U32584 ( .A(u0_0_leon3x0_p0_ici[5]), .Y(n30719) );
  INVxp67_ASAP7_75t_SL U32585 ( .A(uart1_r_THOLD__5__7_), .Y(n27541) );
  INVx1_ASAP7_75t_SL U32586 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__23_), .Y(
        n29071) );
  INVxp67_ASAP7_75t_SL U32587 ( .A(uart1_r_THOLD__7__3_), .Y(n27816) );
  NAND2xp33_ASAP7_75t_SL U32588 ( .A(uart1_v_RXDB__1_), .B(uart1_r_RXTICK_), 
        .Y(n29337) );
  INVx1_ASAP7_75t_SL U32589 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__28_), .Y(
        n25234) );
  INVx1_ASAP7_75t_SL U32590 ( .A(u0_0_leon3x0_p0_mulo[22]), .Y(n29079) );
  INVx1_ASAP7_75t_SL U32591 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__23_), .Y(
        n31981) );
  INVxp67_ASAP7_75t_SL U32592 ( .A(uart1_r_TWADDR__4_), .Y(n27327) );
  INVxp33_ASAP7_75t_SL U32593 ( .A(sr1_r_BSTATE__1_), .Y(n31715) );
  INVx1_ASAP7_75t_SL U32594 ( .A(uart1_r_RCNT__0_), .Y(n31327) );
  INVxp67_ASAP7_75t_SL U32595 ( .A(sr1_r_MCFG1__ROMRWS__0_), .Y(n28057) );
  INVxp67_ASAP7_75t_SL U32596 ( .A(u0_0_leon3x0_p0_ici[16]), .Y(n25751) );
  INVx1_ASAP7_75t_SL U32597 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__6_), .Y(
        n30935) );
  INVx1_ASAP7_75t_SL U32598 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[30]), .Y(n32934)
         );
  INVx1_ASAP7_75t_SL U32599 ( .A(u0_0_leon3x0_p0_divo[2]), .Y(n28364) );
  INVx1_ASAP7_75t_SL U32600 ( .A(u0_0_leon3x0_p0_mulo[38]), .Y(n25283) );
  INVx1_ASAP7_75t_SL U32601 ( .A(u0_0_leon3x0_p0_divi[52]), .Y(n30287) );
  INVxp33_ASAP7_75t_SL U32602 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__2_), 
        .Y(n30170) );
  INVxp67_ASAP7_75t_SL U32603 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[16]), .Y(n29848)
         );
  INVxp67_ASAP7_75t_SL U32604 ( .A(uart1_r_THOLD__4__7_), .Y(n27557) );
  INVx1_ASAP7_75t_SL U32605 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_), .Y(
        n30906) );
  INVxp67_ASAP7_75t_SL U32606 ( .A(u0_0_leon3x0_p0_iu_r_E__CWP__1_), .Y(n31348) );
  INVxp67_ASAP7_75t_SL U32607 ( .A(uart1_r_THOLD__7__2_), .Y(n27880) );
  INVxp67_ASAP7_75t_SL U32608 ( .A(sr1_r_BSTATE__0_), .Y(n31732) );
  INVxp67_ASAP7_75t_SL U32609 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__25_), .Y(
        n28417) );
  INVxp67_ASAP7_75t_SL U32610 ( .A(uart1_r_THOLD__3__7_), .Y(n27575) );
  INVxp67_ASAP7_75t_SL U32611 ( .A(uart1_r_THOLD__7__1_), .Y(n27371) );
  INVxp67_ASAP7_75t_SL U32612 ( .A(u0_0_leon3x0_p0_ici[17]), .Y(n26981) );
  INVx1_ASAP7_75t_SL U32613 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[43]), .Y(n31056)
         );
  INVx1_ASAP7_75t_SL U32614 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__1_), .Y(n26777)
         );
  INVx1_ASAP7_75t_SL U32615 ( .A(apbi[12]), .Y(n29851) );
  INVx1_ASAP7_75t_SL U32616 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__12_), .Y(
        n25938) );
  INVxp67_ASAP7_75t_SL U32617 ( .A(uart1_r_THOLD__2__7_), .Y(n27565) );
  INVxp67_ASAP7_75t_SL U32618 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[10]), .Y(n30530)
         );
  INVxp67_ASAP7_75t_SL U32619 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[27]), .Y(n26526)
         );
  XNOR2xp5_ASAP7_75t_SRAM U32620 ( .A(dt_q[9]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[13]), .Y(n31274) );
  INVxp67_ASAP7_75t_SL U32621 ( .A(uart1_r_THOLD__0__5_), .Y(n27654) );
  INVx1_ASAP7_75t_SL U32622 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[4]), .Y(n32841) );
  INVx1_ASAP7_75t_SL U32623 ( .A(u0_0_leon3x0_p0_mulo[17]), .Y(n27265) );
  INVx1_ASAP7_75t_SL U32624 ( .A(sr1_sdi_HSIZE__0_), .Y(n32834) );
  INVxp67_ASAP7_75t_SL U32625 ( .A(u0_0_leon3x0_p0_ici[28]), .Y(n26723) );
  INVxp67_ASAP7_75t_SL U32626 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[12]), .Y(n25522)
         );
  NAND2xp33_ASAP7_75t_SL U32627 ( .A(n2292), .B(n2356), .Y(n31716) );
  INVx1_ASAP7_75t_SL U32628 ( .A(u0_0_leon3x0_p0_ici[89]), .Y(n31687) );
  XNOR2xp5_ASAP7_75t_SRAM U32629 ( .A(dt_q[18]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[22]), .Y(n31267) );
  INVx1_ASAP7_75t_SL U32630 ( .A(u0_0_leon3x0_p0_mulo[24]), .Y(n29088) );
  INVxp33_ASAP7_75t_SL U32631 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__28_), 
        .Y(n25455) );
  INVx1_ASAP7_75t_SL U32632 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__5_), .Y(
        n26842) );
  INVxp33_ASAP7_75t_SL U32633 ( .A(n2867), .Y(n25970) );
  XNOR2xp5_ASAP7_75t_SRAM U32634 ( .A(dt_q[25]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[29]), .Y(n31268) );
  INVx1_ASAP7_75t_SL U32635 ( .A(u0_0_leon3x0_p0_mulo[8]), .Y(n29100) );
  INVx1_ASAP7_75t_SL U32636 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[28]), .Y(n32916)
         );
  INVx1_ASAP7_75t_SL U32637 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[45]), .Y(n31790)
         );
  INVxp67_ASAP7_75t_SL U32638 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__9_), .Y(
        n26208) );
  INVx1_ASAP7_75t_SL U32639 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__0_), .Y(
        n26829) );
  INVxp67_ASAP7_75t_SL U32640 ( .A(u0_0_leon3x0_p0_ici[22]), .Y(n28455) );
  INVx1_ASAP7_75t_SL U32641 ( .A(sr1_sdi_HSIZE__1_), .Y(n32835) );
  INVxp67_ASAP7_75t_SL U32642 ( .A(u0_0_leon3x0_p0_ici[7]), .Y(n28708) );
  NAND2xp33_ASAP7_75t_SL U32643 ( .A(sr1_r_BSTATE__1_), .B(sr1_r_BSTATE__0_), 
        .Y(n32710) );
  XNOR2xp5_ASAP7_75t_SRAM U32644 ( .A(dt_q[27]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[31]), .Y(n31269) );
  INVx1_ASAP7_75t_SL U32645 ( .A(timer0_vtimers_1__RELOAD__25_), .Y(n31373) );
  INVx1_ASAP7_75t_SL U32646 ( .A(u0_0_leon3x0_p0_divo[5]), .Y(n28356) );
  INVxp67_ASAP7_75t_SL U32647 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__28_), 
        .Y(n25545) );
  INVx1_ASAP7_75t_SL U32648 ( .A(u0_0_leon3x0_p0_div0_r_X__28_), .Y(n29022) );
  INVxp33_ASAP7_75t_SL U32649 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__BURST_), 
        .Y(n26664) );
  INVx1_ASAP7_75t_SL U32650 ( .A(u0_0_leon3x0_p0_div0_r_X__23_), .Y(n29792) );
  INVxp67_ASAP7_75t_SL U32651 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[15]), .Y(n31792)
         );
  NAND2xp5_ASAP7_75t_SL U32652 ( .A(u0_0_leon3x0_p0_iu_v_M__MUL_), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__LD_), .Y(n24814) );
  INVxp67_ASAP7_75t_SL U32653 ( .A(uart1_r_THOLD__6__6_), .Y(n27608) );
  INVx1_ASAP7_75t_SL U32654 ( .A(apbi[19]), .Y(n26544) );
  INVx1_ASAP7_75t_SL U32655 ( .A(uart1_r_RCNT__2_), .Y(n31503) );
  INVx1_ASAP7_75t_SL U32656 ( .A(u0_0_leon3x0_p0_mulo[53]), .Y(n25309) );
  INVxp67_ASAP7_75t_SL U32657 ( .A(uart1_r_THOLD__5__6_), .Y(n27582) );
  INVx1_ASAP7_75t_SL U32658 ( .A(uart1_r_RXTICK_), .Y(n29960) );
  INVxp67_ASAP7_75t_SL U32659 ( .A(n2307), .Y(n28286) );
  INVxp67_ASAP7_75t_SL U32660 ( .A(sr1_r_AREA__0_), .Y(n31744) );
  INVx1_ASAP7_75t_SL U32661 ( .A(timer0_vtimers_1__RELOAD__22_), .Y(n31646) );
  INVxp67_ASAP7_75t_SL U32662 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__28_), 
        .Y(n25547) );
  INVxp67_ASAP7_75t_SL U32663 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__6_), 
        .Y(n31254) );
  INVxp67_ASAP7_75t_SL U32664 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__25_), .Y(
        n28453) );
  INVxp67_ASAP7_75t_SL U32665 ( .A(uart1_r_THOLD__4__6_), .Y(n27598) );
  INVx1_ASAP7_75t_SL U32666 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__8_), .Y(
        n28720) );
  INVxp67_ASAP7_75t_SL U32667 ( .A(uart1_r_THOLD__3__6_), .Y(n27616) );
  INVx1_ASAP7_75t_SL U32668 ( .A(u0_0_leon3x0_p0_mulo[31]), .Y(n30607) );
  INVx1_ASAP7_75t_SL U32669 ( .A(u0_0_leon3x0_p0_div0_r_X__22_), .Y(n28309) );
  INVx1_ASAP7_75t_SL U32670 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__1_), .Y(
        n29180) );
  INVxp33_ASAP7_75t_SL U32671 ( .A(uart1_r_THOLD__12__6_), .Y(n27627) );
  INVxp67_ASAP7_75t_SL U32672 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[11]), .Y(n30514)
         );
  INVxp67_ASAP7_75t_SL U32673 ( .A(uart1_r_THOLD__2__6_), .Y(n27606) );
  INVx1_ASAP7_75t_SL U32674 ( .A(u0_0_leon3x0_p0_iu_r_D__INULL_), .Y(n30502)
         );
  INVxp67_ASAP7_75t_SL U32675 ( .A(n3878), .Y(n30791) );
  INVx1_ASAP7_75t_SL U32676 ( .A(apbi[24]), .Y(n29277) );
  INVx1_ASAP7_75t_SL U32677 ( .A(uart1_r_RCNT__1_), .Y(n30898) );
  INVxp67_ASAP7_75t_SL U32678 ( .A(sr1_r_MCFG1__ROMWIDTH__1_), .Y(n30137) );
  INVxp67_ASAP7_75t_SL U32679 ( .A(uart1_r_THOLD__1__6_), .Y(n27586) );
  INVx1_ASAP7_75t_SL U32680 ( .A(u0_0_leon3x0_p0_mulo[50]), .Y(n25304) );
  INVxp67_ASAP7_75t_SL U32681 ( .A(n4930), .Y(n28255) );
  INVx1_ASAP7_75t_SL U32682 ( .A(u0_0_leon3x0_p0_mulo[23]), .Y(n29090) );
  INVxp67_ASAP7_75t_SL U32683 ( .A(uart1_r_THOLD__0__3_), .Y(n27790) );
  INVx1_ASAP7_75t_SL U32684 ( .A(u0_0_leon3x0_p0_mulo[49]), .Y(n25302) );
  INVxp33_ASAP7_75t_SL U32685 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[58]), .Y(n31784)
         );
  INVx1_ASAP7_75t_SL U32686 ( .A(timer0_vtimers_1__RELOAD__19_), .Y(n32005) );
  INVx1_ASAP7_75t_SL U32687 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__9_), .Y(
        n30388) );
  INVxp67_ASAP7_75t_SL U32688 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[13]), .Y(n30537)
         );
  INVx1_ASAP7_75t_SL U32689 ( .A(u0_0_leon3x0_p0_c0mmu_a0_r_NBA_), .Y(n24896)
         );
  INVxp67_ASAP7_75t_SL U32690 ( .A(uart1_r_THOLD__1__3_), .Y(n27800) );
  INVxp67_ASAP7_75t_SL U32691 ( .A(sr1_r_SRHSEL_), .Y(n31738) );
  INVxp33_ASAP7_75t_SL U32692 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__7_), .Y(
        n28767) );
  INVx1_ASAP7_75t_SL U32693 ( .A(u0_0_leon3x0_p0_divo[4]), .Y(n28860) );
  INVxp67_ASAP7_75t_SL U32694 ( .A(uart1_r_THOLD__0__6_), .Y(n27596) );
  INVxp67_ASAP7_75t_SL U32695 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__20_), 
        .Y(n26753) );
  INVx1_ASAP7_75t_SL U32696 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__5_), .Y(
        n30120) );
  INVx1_ASAP7_75t_SL U32697 ( .A(u0_0_leon3x0_p0_mulo[63]), .Y(n29082) );
  INVx1_ASAP7_75t_SL U32698 ( .A(apbi[9]), .Y(n30139) );
  INVx1_ASAP7_75t_SL U32699 ( .A(u0_0_leon3x0_p0_mulo[58]), .Y(n25317) );
  INVxp67_ASAP7_75t_SL U32700 ( .A(uart1_r_THOLD__2__3_), .Y(n27810) );
  NAND2xp5_ASAP7_75t_SL U32701 ( .A(u0_0_leon3x0_p0_c0mmu_a0_r_NBA_), .B(
        u0_0_leon3x0_p0_c0mmu_a0_r_NBO__0_), .Y(n24897) );
  INVxp33_ASAP7_75t_SL U32702 ( .A(n2838), .Y(n30105) );
  INVx1_ASAP7_75t_SL U32703 ( .A(read), .Y(n31751) );
  INVxp67_ASAP7_75t_SL U32704 ( .A(uart1_r_THOLD__3__3_), .Y(n27820) );
  INVx1_ASAP7_75t_SL U32705 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__19_), .Y(
        n28527) );
  INVx1_ASAP7_75t_SL U32706 ( .A(uart1_r_RCNT__4_), .Y(n31940) );
  INVx1_ASAP7_75t_SL U32707 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), .Y(
        n32083) );
  INVxp67_ASAP7_75t_SL U32708 ( .A(u0_0_leon3x0_p0_iu_r_A__CTRL__TT__0_), .Y(
        n31807) );
  INVxp67_ASAP7_75t_SL U32709 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WY_), .Y(
        n26368) );
  INVxp67_ASAP7_75t_SL U32710 ( .A(uart1_r_THOLD__3__2_), .Y(n27884) );
  INVxp67_ASAP7_75t_SL U32711 ( .A(uart1_r_THOLD__1__0_), .Y(n27923) );
  INVx1_ASAP7_75t_SL U32712 ( .A(n2935), .Y(n32673) );
  INVxp33_ASAP7_75t_SL U32713 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__23_), .Y(
        n26521) );
  INVxp33_ASAP7_75t_SL U32714 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_OVERRUN_), 
        .Y(n31895) );
  INVx1_ASAP7_75t_SL U32715 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[34]), .Y(n32966)
         );
  INVx1_ASAP7_75t_SL U32716 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__11_), .Y(n30382)
         );
  INVx1_ASAP7_75t_SL U32717 ( .A(u0_0_leon3x0_p0_divi[32]), .Y(n26746) );
  NAND2xp5_ASAP7_75t_SL U32718 ( .A(u0_0_leon3x0_p0_iu_r_E__MULSTEP_), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__WY_), .Y(n31404) );
  OAI21xp33_ASAP7_75t_SL U32719 ( .A1(u0_0_leon3x0_p0_iu_r_E__BP_), .A2(
        u0_0_leon3x0_p0_iu_r_A__BP_), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), .Y(n24859) );
  INVxp67_ASAP7_75t_SL U32720 ( .A(uart1_r_THOLD__4__2_), .Y(n27866) );
  INVxp67_ASAP7_75t_SL U32721 ( .A(uart1_r_THOLD__2__0_), .Y(n27953) );
  INVxp67_ASAP7_75t_SL U32722 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__23_), .Y(
        n30263) );
  INVx1_ASAP7_75t_SL U32723 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[7]), .Y(n32847) );
  INVx1_ASAP7_75t_SL U32724 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__10_), .Y(
        n28713) );
  INVxp67_ASAP7_75t_SL U32725 ( .A(uart1_r_THOLD__6__1_), .Y(n27366) );
  INVx1_ASAP7_75t_SL U32726 ( .A(u0_0_leon3x0_p0_ici[69]), .Y(n30974) );
  INVxp67_ASAP7_75t_SL U32727 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[26]), .Y(n31634)
         );
  INVx1_ASAP7_75t_SL U32728 ( .A(u0_0_leon3x0_p0_iu_r_X__INTACK_), .Y(n29741)
         );
  INVxp67_ASAP7_75t_SL U32729 ( .A(u0_0_leon3x0_p0_ici[15]), .Y(n25729) );
  INVxp67_ASAP7_75t_SL U32730 ( .A(u0_0_leon3x0_p0_c0mmu_a0_r_BG_), .Y(n24977)
         );
  INVxp67_ASAP7_75t_SL U32731 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[25]), .Y(n29291)
         );
  INVx1_ASAP7_75t_SL U32732 ( .A(u0_0_leon3x0_p0_mulo[18]), .Y(n29094) );
  INVx1_ASAP7_75t_SL U32733 ( .A(n2736), .Y(n29307) );
  INVxp67_ASAP7_75t_SL U32734 ( .A(uart1_r_THOLD__5__1_), .Y(n27341) );
  NAND2xp5_ASAP7_75t_SL U32735 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__4_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__TT__0_), .Y(n25946) );
  INVxp67_ASAP7_75t_SL U32736 ( .A(uart1_r_THOLD__5__2_), .Y(n27850) );
  INVx1_ASAP7_75t_SL U32737 ( .A(u0_0_leon3x0_p0_mulo[57]), .Y(n25315) );
  INVx1_ASAP7_75t_SL U32738 ( .A(u0_0_leon3x0_p0_mulo[55]), .Y(n25313) );
  INVxp67_ASAP7_75t_SL U32739 ( .A(irqo[1]), .Y(n29646) );
  INVx1_ASAP7_75t_SL U32740 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__0_), .Y(
        n24920) );
  INVxp67_ASAP7_75t_SL U32741 ( .A(uart1_r_THOLD__4__1_), .Y(n27335) );
  INVxp67_ASAP7_75t_SL U32742 ( .A(uart1_r_THOLD__6__2_), .Y(n27876) );
  INVx1_ASAP7_75t_SL U32743 ( .A(apbi[14]), .Y(n30547) );
  INVxp67_ASAP7_75t_SL U32744 ( .A(uart1_r_THOLD__3__1_), .Y(n27378) );
  INVx1_ASAP7_75t_SL U32745 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__30_), .Y(
        n30590) );
  INVx1_ASAP7_75t_SL U32746 ( .A(apbi[18]), .Y(n29570) );
  INVx1_ASAP7_75t_SL U32747 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_), .Y(
        n31962) );
  INVxp67_ASAP7_75t_SL U32748 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[36]), .Y(n32714)
         );
  INVx1_ASAP7_75t_SL U32749 ( .A(u0_0_leon3x0_p0_divo[26]), .Y(n28305) );
  INVx1_ASAP7_75t_SL U32750 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__25_), .Y(
        n25537) );
  INVx1_ASAP7_75t_SL U32751 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__23_), .Y(
        n32219) );
  NAND2xp5_ASAP7_75t_SL U32752 ( .A(u0_0_leon3x0_p0_muli[8]), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__23_), .Y(n31964) );
  INVxp67_ASAP7_75t_SL U32753 ( .A(irqctrl0_r_IMASK__0__14_), .Y(n25640) );
  INVxp67_ASAP7_75t_SL U32754 ( .A(uart1_r_THOLD__3__0_), .Y(n27969) );
  NAND2xp33_ASAP7_75t_SL U32755 ( .A(u0_0_leon3x0_p0_iu_de_icc_1_), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_), .Y(n24724) );
  INVxp67_ASAP7_75t_SL U32756 ( .A(uart1_r_THOLD__2__1_), .Y(n27362) );
  INVx1_ASAP7_75t_SL U32757 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__TRAP_), .Y(
        n31441) );
  INVx1_ASAP7_75t_SL U32758 ( .A(timer0_vtimers_1__RELOAD__14_), .Y(n30549) );
  INVx1_ASAP7_75t_SL U32759 ( .A(irqctrl0_r_IFORCE__0__14_), .Y(n29655) );
  INVx1_ASAP7_75t_SL U32760 ( .A(u0_0_leon3x0_p0_muli[1]), .Y(n26369) );
  INVx1_ASAP7_75t_SL U32761 ( .A(timer0_vtimers_1__RELOAD__18_), .Y(n29573) );
  INVxp67_ASAP7_75t_SL U32762 ( .A(u0_0_leon3x0_p0_iu_de_icc_3_), .Y(n29817)
         );
  INVxp67_ASAP7_75t_SL U32763 ( .A(uart1_r_THOLD__1__1_), .Y(n27347) );
  INVxp33_ASAP7_75t_SL U32764 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__1_), .Y(
        n26729) );
  INVxp67_ASAP7_75t_SL U32765 ( .A(uart1_r_THOLD__0__1_), .Y(n27331) );
  INVx1_ASAP7_75t_SL U32766 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__22_), .Y(
        n32216) );
  INVx1_ASAP7_75t_SL U32767 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__25_), .Y(
        n25689) );
  INVx1_ASAP7_75t_SL U32768 ( .A(u0_0_leon3x0_p0_mulo[42]), .Y(n25288) );
  INVxp67_ASAP7_75t_SL U32769 ( .A(uart1_r_THOLD__4__0_), .Y(n27943) );
  INVx1_ASAP7_75t_SL U32770 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__26_), .Y(
        n24714) );
  INVx1_ASAP7_75t_SL U32771 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__20_), .Y(
        n32213) );
  INVxp67_ASAP7_75t_SL U32772 ( .A(u0_0_leon3x0_p0_divi[41]), .Y(n30390) );
  NAND2xp5_ASAP7_75t_SL U32773 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__1_), 
        .B(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__2_), .Y(n31559) );
  INVx1_ASAP7_75t_SL U32774 ( .A(u0_0_leon3x0_p0_iu_de_icc_1_), .Y(n30677) );
  INVxp67_ASAP7_75t_SL U32775 ( .A(apbi[26]), .Y(n26498) );
  INVxp67_ASAP7_75t_SL U32776 ( .A(uart1_r_THOLD__5__0_), .Y(n27916) );
  INVx1_ASAP7_75t_SL U32777 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__0_), .Y(n26872) );
  INVxp67_ASAP7_75t_SL U32778 ( .A(uart1_r_THOLD__6__0_), .Y(n27956) );
  INVx1_ASAP7_75t_SL U32779 ( .A(u0_0_leon3x0_p0_iu_r_E__BP_), .Y(n25453) );
  OAI21xp5_ASAP7_75t_SL U32780 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__0_), 
        .A2(u0_0_leon3x0_p0_iu_r_M__MUL_), .B(
        u0_0_leon3x0_p0_iu_r_M__CTRL__WICC_), .Y(n24850) );
  INVx1_ASAP7_75t_SL U32781 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__14_), .Y(
        n28585) );
  INVxp67_ASAP7_75t_SL U32782 ( .A(u0_0_leon3x0_p0_iu_r_A__BP_), .Y(n24720) );
  INVx1_ASAP7_75t_SL U32783 ( .A(u0_0_leon3x0_p0_mulo[26]), .Y(n29086) );
  INVx1_ASAP7_75t_SL U32784 ( .A(u0_0_leon3x0_p0_mulo[30]), .Y(n29084) );
  INVx1_ASAP7_75t_SL U32785 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__8_), .Y(
        n30392) );
  INVxp67_ASAP7_75t_SL U32786 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__3_), 
        .Y(n30168) );
  INVxp67_ASAP7_75t_SL U32787 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__TT__2_), .Y(
        n25707) );
  INVxp67_ASAP7_75t_SL U32788 ( .A(uart1_r_THOLD__7__0_), .Y(n27963) );
  INVxp67_ASAP7_75t_SL U32789 ( .A(uart1_r_THOLD__1__7_), .Y(n27545) );
  INVxp67_ASAP7_75t_SL U32790 ( .A(sr1_r_MCFG1__ROMRWS__1_), .Y(n26131) );
  INVx1_ASAP7_75t_SL U32791 ( .A(irqctrl0_r_IMASK__0__2_), .Y(n29400) );
  INVxp33_ASAP7_75t_SL U32792 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__1_), .Y(
        n31819) );
  INVx1_ASAP7_75t_SL U32793 ( .A(sr1_r_WS__0_), .Y(n31724) );
  INVx1_ASAP7_75t_SL U32794 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__21_), .Y(
        n28520) );
  INVx1_ASAP7_75t_SL U32795 ( .A(u0_0_leon3x0_p0_divo[30]), .Y(n28301) );
  INVx1_ASAP7_75t_SL U32796 ( .A(apbi[8]), .Y(n29744) );
  INVxp67_ASAP7_75t_SL U32797 ( .A(uart1_r_THOLD__0__7_), .Y(n27555) );
  INVx1_ASAP7_75t_SL U32798 ( .A(u0_0_leon3x0_p0_divo[33]), .Y(n31675) );
  INVxp67_ASAP7_75t_SL U32799 ( .A(timer0_r_RELOAD__1_), .Y(n26133) );
  INVx1_ASAP7_75t_SL U32800 ( .A(timer0_vtimers_1__RELOAD__3_), .Y(n28254) );
  INVx1_ASAP7_75t_SL U32801 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__3_), .Y(n28904)
         );
  INVxp67_ASAP7_75t_SL U32802 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__18_), .Y(
        n25727) );
  INVxp67_ASAP7_75t_SL U32803 ( .A(n2267), .Y(n27322) );
  INVx1_ASAP7_75t_SL U32804 ( .A(u0_0_leon3x0_p0_divo[1]), .Y(n28370) );
  INVx1_ASAP7_75t_SL U32805 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .Y(
        n31537) );
  INVxp67_ASAP7_75t_SL U32806 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__1_), 
        .Y(n30165) );
  INVx1_ASAP7_75t_SL U32807 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[29]), .Y(n32926)
         );
  INVx1_ASAP7_75t_SL U32808 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_), .Y(
        n25675) );
  INVx1_ASAP7_75t_SL U32809 ( .A(timer0_vtimers_1__RELOAD__26_), .Y(n31328) );
  INVx1_ASAP7_75t_SL U32810 ( .A(uart1_r_DPAR_), .Y(n30066) );
  INVx1_ASAP7_75t_SL U32811 ( .A(u0_0_leon3x0_p0_divi[33]), .Y(n30459) );
  INVx1_ASAP7_75t_SL U32812 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_), .Y(
        n31958) );
  INVxp67_ASAP7_75t_SL U32813 ( .A(u0_0_leon3x0_p0_divi[31]), .Y(n26738) );
  INVx1_ASAP7_75t_SL U32814 ( .A(timer0_vtimers_1__RELOAD__9_), .Y(n30151) );
  INVxp67_ASAP7_75t_SL U32815 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__2_), .Y(
        n25104) );
  AOI21xp33_ASAP7_75t_SL U32816 ( .A1(u0_0_leon3x0_p0_iu_r_A__CTRL__WICC_), 
        .A2(u0_0_leon3x0_p0_iu_r_A__MULSTART_), .B(
        u0_0_leon3x0_p0_iu_r_A__NOBP_), .Y(n24851) );
  INVxp67_ASAP7_75t_SL U32817 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__8_), .Y(
        n30717) );
  INVxp67_ASAP7_75t_SL U32818 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__WY_), .Y(
        n31389) );
  INVx1_ASAP7_75t_SL U32819 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[38]), .Y(n31948)
         );
  INVx1_ASAP7_75t_SL U32820 ( .A(u0_0_leon3x0_p0_div0_r_X__14_), .Y(n28328) );
  INVxp67_ASAP7_75t_SL U32821 ( .A(u0_0_leon3x0_p0_iu_r_E__MULSTEP_), .Y(
        n26365) );
  INVxp67_ASAP7_75t_SL U32822 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WREG_), .Y(
        n24952) );
  INVx1_ASAP7_75t_SL U32823 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__22_), .Y(n30270)
         );
  INVxp67_ASAP7_75t_SL U32824 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[57]), .Y(n31776)
         );
  INVx1_ASAP7_75t_SL U32825 ( .A(n4076), .Y(n32023) );
  INVx1_ASAP7_75t_SL U32826 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__2_), .Y(n28956)
         );
  INVx1_ASAP7_75t_SL U32827 ( .A(timer0_vtimers_1__RELOAD__6_), .Y(n31244) );
  INVxp33_ASAP7_75t_SL U32828 ( .A(u0_0_leon3x0_p0_c0mmu_a0_r_HLOCKEN_), .Y(
        n25244) );
  INVx1_ASAP7_75t_SL U32829 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), .Y(
        n31858) );
  INVxp67_ASAP7_75t_SL U32830 ( .A(n3325), .Y(n27294) );
  INVx1_ASAP7_75t_SL U32831 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[9]), .Y(n32851) );
  INVxp67_ASAP7_75t_SL U32832 ( .A(uart1_r_THOLD__0__2_), .Y(n27864) );
  INVxp67_ASAP7_75t_SL U32833 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[18]), .Y(n25631)
         );
  INVx1_ASAP7_75t_SL U32834 ( .A(u0_0_leon3x0_p0_mulo[48]), .Y(n25300) );
  INVxp67_ASAP7_75t_SL U32835 ( .A(u0_0_leon3x0_p0_divi[61]), .Y(n30220) );
  INVx1_ASAP7_75t_SL U32836 ( .A(u0_0_leon3x0_p0_divi[62]), .Y(n31678) );
  INVxp67_ASAP7_75t_SL U32837 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__20_), .Y(
        n26979) );
  INVxp67_ASAP7_75t_SL U32838 ( .A(uart1_r_TWADDR__1_), .Y(n27343) );
  INVxp67_ASAP7_75t_SL U32839 ( .A(uart1_r_THOLD__1__2_), .Y(n27854) );
  INVx1_ASAP7_75t_SL U32840 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__27_), .Y(
        n30905) );
  INVxp67_ASAP7_75t_SL U32841 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[22]), .Y(n25843)
         );
  INVx1_ASAP7_75t_SL U32842 ( .A(timer0_vtimers_1__RELOAD__27_), .Y(n30899) );
  INVxp67_ASAP7_75t_SL U32843 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__TRAP_), .Y(
        n31804) );
  INVx1_ASAP7_75t_SL U32844 ( .A(sr1_r_HBURST__0_), .Y(n31698) );
  INVxp33_ASAP7_75t_SL U32845 ( .A(n4531), .Y(n30902) );
  INVxp33_ASAP7_75t_SL U32846 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__14_), .Y(n25613) );
  INVxp67_ASAP7_75t_SL U32847 ( .A(sr1_r_MCFG1__ROMRWS__3_), .Y(n28236) );
  INVxp67_ASAP7_75t_SL U32848 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__0_), .Y(
        n25095) );
  INVxp67_ASAP7_75t_SL U32849 ( .A(apbi[30]), .Y(n26479) );
  INVx1_ASAP7_75t_SL U32850 ( .A(u0_0_leon3x0_p0_mulo[61]), .Y(n25322) );
  INVxp67_ASAP7_75t_SL U32851 ( .A(irqctrl0_r_IFORCE__0__3_), .Y(n28242) );
  INVxp67_ASAP7_75t_SL U32852 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__20_), .Y(
        n26977) );
  INVx1_ASAP7_75t_SL U32853 ( .A(u0_0_leon3x0_p0_div0_r_X__31_), .Y(n28295) );
  INVxp67_ASAP7_75t_SL U32854 ( .A(uart1_r_THOLD__2__2_), .Y(n27874) );
  NAND2xp5_ASAP7_75t_SL U32855 ( .A(n18819), .B(n18842), .Y(n24878) );
  INVxp33_ASAP7_75t_SL U32856 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__1_), .Y(
        n30941) );
  INVxp67_ASAP7_75t_SL U32857 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[28]), .Y(n25251)
         );
  INVx1_ASAP7_75t_SL U32858 ( .A(u0_0_leon3x0_p0_mulo[54]), .Y(n25311) );
  INVx1_ASAP7_75t_SL U32859 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[42]), .Y(n31971)
         );
  INVx1_ASAP7_75t_SL U32860 ( .A(timer0_vtimers_1__RELOAD__30_), .Y(n31941) );
  INVxp67_ASAP7_75t_SL U32861 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__20_), .Y(
        n26975) );
  INVx1_ASAP7_75t_SL U32862 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[41]), .Y(n30737)
         );
  INVxp67_ASAP7_75t_SL U32863 ( .A(uart1_r_THOLD__0__0_), .Y(n27940) );
  INVxp67_ASAP7_75t_SL U32864 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__8_), .Y(
        n30715) );
  INVxp67_ASAP7_75t_SL U32865 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[50]), .Y(n30541)
         );
  INVxp67_ASAP7_75t_SL U32866 ( .A(uart1_r_THOLD__2__4_), .Y(n27738) );
  INVx1_ASAP7_75t_SL U32867 ( .A(u0_0_leon3x0_p0_div0_r_X__24_), .Y(n29793) );
  INVx1_ASAP7_75t_SL U32868 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__3_), .Y(
        n30439) );
  INVx1_ASAP7_75t_SL U32869 ( .A(u0_0_leon3x0_p0_divo[8]), .Y(n28749) );
  INVxp67_ASAP7_75t_SL U32870 ( .A(u0_0_leon3x0_p0_ici[86]), .Y(n29032) );
  XNOR2xp5_ASAP7_75t_SRAM U32871 ( .A(dt_q[19]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[23]), .Y(n31287) );
  INVxp67_ASAP7_75t_SL U32872 ( .A(irqctrl0_r_IFORCE__0__5_), .Y(n29299) );
  INVx1_ASAP7_75t_SL U32873 ( .A(u0_0_leon3x0_p0_mulo[39]), .Y(n25284) );
  INVxp67_ASAP7_75t_SL U32874 ( .A(uart1_r_THOLD__1__4_), .Y(n27718) );
  INVxp67_ASAP7_75t_SL U32875 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__3_), .Y(
        n29486) );
  INVxp67_ASAP7_75t_SL U32876 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__7_), .Y(
        n31511) );
  INVx1_ASAP7_75t_SL U32877 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__11_), .Y(
        n30696) );
  INVx1_ASAP7_75t_SL U32878 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[20]), .Y(n31761)
         );
  XNOR2xp5_ASAP7_75t_SRAM U32879 ( .A(dt_q[16]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[20]), .Y(n31288) );
  INVxp67_ASAP7_75t_SL U32880 ( .A(uart1_r_THOLD__0__4_), .Y(n27728) );
  INVx1_ASAP7_75t_SL U32881 ( .A(u0_0_leon3x0_p0_mulo[25]), .Y(n28451) );
  INVx1_ASAP7_75t_SL U32882 ( .A(n2962), .Y(n31607) );
  INVxp33_ASAP7_75t_SL U32883 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__8_), .Y(n29760) );
  INVxp67_ASAP7_75t_SL U32884 ( .A(u0_0_leon3x0_p0_ici[0]), .Y(n29488) );
  INVxp67_ASAP7_75t_SL U32885 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[54]), .Y(n31766)
         );
  INVxp67_ASAP7_75t_SL U32886 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__7_), .Y(
        n26840) );
  INVxp67_ASAP7_75t_SL U32887 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__27_), 
        .Y(n25551) );
  INVxp33_ASAP7_75t_SL U32888 ( .A(uart1_r_THOLD__12__4_), .Y(n27759) );
  INVx1_ASAP7_75t_SL U32889 ( .A(u0_0_leon3x0_p0_div0_r_X__8_), .Y(n27176) );
  INVxp67_ASAP7_75t_SL U32890 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FLUSH2_), 
        .Y(n30200) );
  INVxp67_ASAP7_75t_SL U32891 ( .A(u0_0_leon3x0_p0_ici[24]), .Y(n26885) );
  INVxp67_ASAP7_75t_SL U32892 ( .A(u0_0_leon3x0_p0_ici[6]), .Y(n26214) );
  INVxp67_ASAP7_75t_SL U32893 ( .A(uart1_r_BRATE__3_), .Y(n28160) );
  INVxp33_ASAP7_75t_SL U32894 ( .A(n4414), .Y(n31978) );
  INVxp67_ASAP7_75t_SL U32895 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[37]), .Y(n32737)
         );
  INVx1_ASAP7_75t_SL U32896 ( .A(sr1_r_BUSW__0_), .Y(n32884) );
  INVxp67_ASAP7_75t_SL U32897 ( .A(uart1_r_THOLD__6__5_), .Y(n27676) );
  INVx1_ASAP7_75t_SL U32898 ( .A(n3880), .Y(n31883) );
  INVxp67_ASAP7_75t_SL U32899 ( .A(u0_0_leon3x0_p0_iu_v_E__CWP__0_), .Y(n32115) );
  INVx1_ASAP7_75t_SL U32900 ( .A(u0_0_leon3x0_p0_div0_r_X__9_), .Y(n27177) );
  INVxp67_ASAP7_75t_SL U32901 ( .A(uart1_r_THOLD__5__5_), .Y(n27660) );
  XNOR2xp5_ASAP7_75t_SRAM U32902 ( .A(n31278), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[21]), .Y(n31279) );
  INVx1_ASAP7_75t_SL U32903 ( .A(u0_0_leon3x0_p0_mulo[19]), .Y(n29092) );
  INVx1_ASAP7_75t_SL U32904 ( .A(n2861), .Y(n28184) );
  INVx1_ASAP7_75t_SL U32905 ( .A(u0_0_leon3x0_p0_divo[10]), .Y(n28344) );
  INVx1_ASAP7_75t_SL U32906 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[17]), .Y(n31768)
         );
  INVxp67_ASAP7_75t_SL U32907 ( .A(sr1_r_MCFG1__IOWIDTH__1_), .Y(n31499) );
  INVxp67_ASAP7_75t_SL U32908 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__31_), 
        .Y(n31959) );
  INVx1_ASAP7_75t_SL U32909 ( .A(u0_0_leon3x0_p0_mulo[11]), .Y(n28698) );
  INVx1_ASAP7_75t_SL U32910 ( .A(u0_0_leon3x0_p0_ici[63]), .Y(n32567) );
  INVxp67_ASAP7_75t_SL U32911 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__31_), .Y(
        n26373) );
  INVxp67_ASAP7_75t_SL U32912 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__28_), .Y(
        n30235) );
  INVx1_ASAP7_75t_SL U32913 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[23]), .Y(n31778)
         );
  INVxp67_ASAP7_75t_SL U32914 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[52]), .Y(n30829)
         );
  INVx1_ASAP7_75t_SL U32915 ( .A(n4519), .Y(n28032) );
  INVx1_ASAP7_75t_SL U32916 ( .A(u0_0_leon3x0_p0_ici[66]), .Y(n32577) );
  XNOR2xp5_ASAP7_75t_SRAM U32917 ( .A(dt_q[11]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[15]), .Y(n31289) );
  INVxp33_ASAP7_75t_SL U32918 ( .A(uart1_r_THOLD__12__0_), .Y(n27987) );
  INVx1_ASAP7_75t_SL U32919 ( .A(u0_0_leon3x0_p0_ici[67]), .Y(n32580) );
  INVx1_ASAP7_75t_SL U32920 ( .A(uart1_r_TICK_), .Y(n29944) );
  INVx1_ASAP7_75t_SL U32921 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__12_), .Y(
        n30370) );
  INVx1_ASAP7_75t_SL U32922 ( .A(u0_0_leon3x0_p0_iu_r_X__Y__26_), .Y(n30243)
         );
  INVx1_ASAP7_75t_SL U32923 ( .A(u0_0_leon3x0_p0_ici[65]), .Y(n32574) );
  INVx1_ASAP7_75t_SL U32924 ( .A(u0_0_leon3x0_p0_mulo[60]), .Y(n25321) );
  INVx1_ASAP7_75t_SL U32925 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[32]), .Y(n32950)
         );
  INVx1_ASAP7_75t_SL U32926 ( .A(u0_0_leon3x0_p0_ici[64]), .Y(n31018) );
  INVxp67_ASAP7_75t_SL U32927 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[24]), .Y(n25257)
         );
  INVxp67_ASAP7_75t_SL U32928 ( .A(uart1_r_THOLD__6__4_), .Y(n27740) );
  INVxp67_ASAP7_75t_SL U32929 ( .A(uart1_r_THOLD__5__4_), .Y(n27714) );
  INVx1_ASAP7_75t_SL U32930 ( .A(n1723), .Y(address[1]) );
  INVx1_ASAP7_75t_SL U32931 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__5_), .Y(
        n26852) );
  INVx1_ASAP7_75t_SL U32932 ( .A(n1724), .Y(address[0]) );
  INVx1_ASAP7_75t_SL U32933 ( .A(u0_0_leon3x0_p0_divo[9]), .Y(n28347) );
  INVxp67_ASAP7_75t_SL U32934 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__18_), .Y(
        n25841) );
  INVx1_ASAP7_75t_SL U32935 ( .A(u0_0_leon3x0_p0_div0_r_X__25_), .Y(n29794) );
  INVxp67_ASAP7_75t_SL U32936 ( .A(u0_0_leon3x0_p0_ici[88]), .Y(n25890) );
  INVxp67_ASAP7_75t_SL U32937 ( .A(uart1_r_THOLD__4__4_), .Y(n27730) );
  INVxp67_ASAP7_75t_SL U32938 ( .A(uart1_r_THOLD__3__4_), .Y(n27748) );
  INVx1_ASAP7_75t_SL U32939 ( .A(u0_0_leon3x0_p0_iu_r_W__S__ICC__2_), .Y(
        n29166) );
  INVx1_ASAP7_75t_SL U32940 ( .A(u0_0_leon3x0_p0_ici[87]), .Y(n31690) );
  XNOR2xp5_ASAP7_75t_SRAM U32941 ( .A(dt_q[14]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[18]), .Y(n31285) );
  INVxp67_ASAP7_75t_SL U32942 ( .A(u0_0_leon3x0_p0_iu_r_X__ICC__2_), .Y(n29132) );
  INVxp33_ASAP7_75t_SL U32943 ( .A(uart1_r_THOLD__30__4_), .Y(n27775) );
  INVx1_ASAP7_75t_SL U32944 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[22]), .Y(n31782)
         );
  XNOR2xp5_ASAP7_75t_SRAM U32945 ( .A(dt_q[13]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[17]), .Y(n31286) );
  INVxp33_ASAP7_75t_SL U32946 ( .A(uart1_r_TCNT__3_), .Y(n31974) );
  INVxp33_ASAP7_75t_SL U32947 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__1_), .Y(
        n30606) );
  XNOR2xp5_ASAP7_75t_SRAM U32948 ( .A(dt_q[15]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[19]), .Y(n31271) );
  INVxp67_ASAP7_75t_SL U32949 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__10_), .Y(
        n23549) );
  INVx1_ASAP7_75t_SL U32950 ( .A(u0_0_leon3x0_p0_mulo[62]), .Y(n26371) );
  INVxp33_ASAP7_75t_SL U32951 ( .A(n4573), .Y(n31649) );
  INVx1_ASAP7_75t_SL U32952 ( .A(n3065), .Y(n32583) );
  INVx1_ASAP7_75t_SL U32953 ( .A(u0_0_leon3x0_p0_div0_r_X__7_), .Y(n29926) );
  INVxp67_ASAP7_75t_SL U32954 ( .A(irqctrl0_r_IMASK__0__9_), .Y(n29249) );
  INVxp67_ASAP7_75t_SL U32955 ( .A(u0_0_leon3x0_p0_iu_r_E__CWP__0_), .Y(n32117) );
  INVx1_ASAP7_75t_SL U32956 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__26_), .Y(
        n28400) );
  XNOR2xp5_ASAP7_75t_SRAM U32957 ( .A(dt_q[10]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[14]), .Y(n31272) );
  INVx1_ASAP7_75t_SL U32958 ( .A(timer0_vtimers_1__RELOAD__23_), .Y(n31975) );
  INVx1_ASAP7_75t_SL U32959 ( .A(n2883), .Y(uart1_uarto_SCALER__11_) );
  INVx1_ASAP7_75t_SL U32960 ( .A(n3725), .Y(n31658) );
  INVxp67_ASAP7_75t_SL U32961 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[16]), .Y(n30832)
         );
  INVx1_ASAP7_75t_SL U32962 ( .A(u0_0_leon3x0_p0_iu_r_W__RESULT__1_), .Y(
        n30643) );
  NAND2xp5_ASAP7_75t_SL U32963 ( .A(u0_0_leon3x0_p0_div0_r_CNT__0_), .B(
        u0_0_leon3x0_p0_div0_r_CNT__1_), .Y(n24900) );
  INVxp33_ASAP7_75t_SL U32964 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_), .Y(
        n29135) );
  INVx1_ASAP7_75t_SL U32965 ( .A(u0_0_leon3x0_p0_div0_r_X__21_), .Y(n28312) );
  INVxp67_ASAP7_75t_SL U32966 ( .A(uart1_r_THOLD__2__5_), .Y(n27674) );
  INVx1_ASAP7_75t_SL U32967 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[8]), .Y(n32849) );
  INVxp67_ASAP7_75t_SL U32968 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__27_), .Y(
        n26881) );
  INVxp67_ASAP7_75t_SL U32969 ( .A(uart1_r_BRATE__4_), .Y(n28156) );
  INVxp67_ASAP7_75t_SL U32970 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__9_), .Y(
        n26212) );
  INVxp33_ASAP7_75t_SL U32971 ( .A(n4624), .Y(n31376) );
  INVxp33_ASAP7_75t_SL U32972 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__10_), .Y(n31000) );
  INVx1_ASAP7_75t_SL U32973 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__4_), .Y(
        n25005) );
  INVx1_ASAP7_75t_SL U32974 ( .A(u0_0_leon3x0_p0_div0_r_X__30_), .Y(n28283) );
  INVx1_ASAP7_75t_SL U32975 ( .A(u0_0_leon3x0_p0_divo[7]), .Y(n28794) );
  INVx1_ASAP7_75t_SL U32976 ( .A(uart1_r_TCNT__5_), .Y(n31372) );
  INVx1_ASAP7_75t_SL U32977 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__10_), .Y(n28715)
         );
  NAND2xp33_ASAP7_75t_SL U32978 ( .A(apbi[45]), .B(apbi[43]), .Y(n17251) );
  INVxp67_ASAP7_75t_SL U32979 ( .A(uart1_r_THOLD__3__5_), .Y(n27684) );
  INVx1_ASAP7_75t_SL U32980 ( .A(u0_0_leon3x0_p0_div0_r_X__10_), .Y(n28337) );
  INVxp67_ASAP7_75t_SL U32981 ( .A(uart1_r_THOLD__4__5_), .Y(n27656) );
  INVxp67_ASAP7_75t_SL U32982 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__9_), .Y(
        n26210) );
  INVx1_ASAP7_75t_SL U32983 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__10_), .Y(
        n30699) );
  INVxp67_ASAP7_75t_SL U32984 ( .A(u0_0_leon3x0_p0_div0_r_CNT__3_), .Y(n24885)
         );
  INVx1_ASAP7_75t_SL U32985 ( .A(u0_0_leon3x0_p0_iu_r_X__RESULT__2_), .Y(
        n30450) );
  INVxp67_ASAP7_75t_SL U32986 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__PC__27_), .Y(
        n26879) );
  INVx1_ASAP7_75t_SL U32987 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__11_), .Y(
        n32592) );
  INVx1_ASAP7_75t_SL U32988 ( .A(u0_0_leon3x0_p0_c0mmu_mcdi[10]), .Y(n32853)
         );
  INVxp67_ASAP7_75t_SL U32989 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__27_), .Y(
        n26883) );
  INVxp67_ASAP7_75t_SL U32990 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__2_), .Y(
        n26835) );
  INVxp67_ASAP7_75t_SL U32991 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__2_), .Y(
        n26833) );
  INVxp67_ASAP7_75t_SL U32992 ( .A(uart1_r_THOLD__1__5_), .Y(n27664) );
  INVxp67_ASAP7_75t_SL U32993 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__PC__10_), .Y(
        n28706) );
  INVx1_ASAP7_75t_SL U32994 ( .A(uart1_r_TCNT__2_), .Y(n31645) );
  INVx1_ASAP7_75t_SL U32995 ( .A(apbi[23]), .Y(n26530) );
  INVxp67_ASAP7_75t_SL U32996 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[14]), .Y(n30544)
         );
  INVxp33_ASAP7_75t_SL U32997 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_NOFLUSH_), 
        .Y(n30184) );
  INVx1_ASAP7_75t_SL U32998 ( .A(u0_0_leon3x0_p0_div0_r_X__19_), .Y(n27036) );
  INVx1_ASAP7_75t_SL U32999 ( .A(it_q[2]), .Y(n32475) );
  INVx1_ASAP7_75t_SL U33000 ( .A(dt_q[7]), .Y(n31266) );
  INVx1_ASAP7_75t_SL U33001 ( .A(it_q[6]), .Y(n32504) );
  INVx1_ASAP7_75t_SL U33002 ( .A(it_q[3]), .Y(n32483) );
  INVx1_ASAP7_75t_SL U33003 ( .A(it_q[7]), .Y(n32514) );
  INVx1_ASAP7_75t_SL U33004 ( .A(dt_q[26]), .Y(n31277) );
  INVx1_ASAP7_75t_SL U33005 ( .A(it_q[0]), .Y(n32463) );
  INVx1_ASAP7_75t_SL U33006 ( .A(dc_q[9]), .Y(n30127) );
  INVx1_ASAP7_75t_SL U33007 ( .A(ic_q[9]), .Y(n30125) );
  INVx1_ASAP7_75t_SL U33008 ( .A(it_q[5]), .Y(n32497) );
  INVx1_ASAP7_75t_SL U33009 ( .A(ic_q[1]), .Y(n31353) );
  INVx1_ASAP7_75t_SL U33010 ( .A(it_q[4]), .Y(n32491) );
  INVx1_ASAP7_75t_SL U33011 ( .A(it_q[1]), .Y(n32468) );
  XNOR2xp5_ASAP7_75t_SL U33012 ( .A(mult_x_1196_n2173), .B(mult_x_1196_n2544), 
        .Y(n22435) );
  HB1xp67_ASAP7_75t_SL U33013 ( .A(u0_0_leon3x0_p0_muli[47]), .Y(n22436) );
  XNOR2xp5_ASAP7_75t_SL U33014 ( .A(mult_x_1196_n1640), .B(n22437), .Y(
        mult_x_1196_n1599) );
  XOR2xp5_ASAP7_75t_SL U33015 ( .A(mult_x_1196_n1638), .B(mult_x_1196_n1642), 
        .Y(n22437) );
  INVx8_ASAP7_75t_SL U33016 ( .A(n23645), .Y(n24012) );
  NAND2x1_ASAP7_75t_SL U33017 ( .A(mult_x_1196_n1391), .B(mult_x_1196_n1358), 
        .Y(mult_x_1196_n565) );
  XOR2xp5_ASAP7_75t_SL U33018 ( .A(n22438), .B(n23027), .Y(n22483) );
  INVx1_ASAP7_75t_SL U33019 ( .A(mult_x_1196_n1900), .Y(n22438) );
  NOR2x1p5_ASAP7_75t_SL U33020 ( .A(mult_x_1196_n3145), .B(n23992), .Y(n23430)
         );
  NAND2xp5_ASAP7_75t_SL U33021 ( .A(n22884), .B(n22883), .Y(n22879) );
  XOR2xp5_ASAP7_75t_SL U33022 ( .A(n22440), .B(n22836), .Y(n22883) );
  INVx1_ASAP7_75t_SL U33023 ( .A(mult_x_1196_n1308), .Y(n22440) );
  INVx1_ASAP7_75t_SL U33024 ( .A(n22500), .Y(n22502) );
  XNOR2xp5_ASAP7_75t_SL U33025 ( .A(n24292), .B(n23029), .Y(n22500) );
  INVx3_ASAP7_75t_SL U33026 ( .A(n23972), .Y(n23973) );
  HB1xp67_ASAP7_75t_SL U33027 ( .A(mult_x_1196_n646), .Y(n22441) );
  NOR2x1_ASAP7_75t_SL U33028 ( .A(n22258), .B(mult_x_1196_n323), .Y(n22443) );
  XOR2xp5_ASAP7_75t_SL U33029 ( .A(n22336), .B(n23583), .Y(n23250) );
  XNOR2x2_ASAP7_75t_SL U33030 ( .A(n23251), .B(n22666), .Y(n23583) );
  INVxp67_ASAP7_75t_SL U33031 ( .A(n25089), .Y(n23568) );
  INVx1_ASAP7_75t_SL U33032 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__15_), .Y(
        n26562) );
  XOR2x2_ASAP7_75t_SL U33033 ( .A(n24064), .B(n23397), .Y(mult_x_1196_n3165)
         );
  AND2x4_ASAP7_75t_SL U33034 ( .A(n22919), .B(u0_0_leon3x0_p0_muli[36]), .Y(
        u0_0_leon3x0_p0_muli[37]) );
  XOR2x2_ASAP7_75t_SL U33035 ( .A(n23383), .B(n23382), .Y(mult_x_1196_n1572)
         );
  BUFx2_ASAP7_75t_SL U33036 ( .A(n23465), .Y(n22450) );
  NAND2x1p5_ASAP7_75t_SL U33037 ( .A(n22444), .B(n23696), .Y(mult_x_1196_n2295) );
  NAND2x1p5_ASAP7_75t_SL U33038 ( .A(n22446), .B(n22445), .Y(n22444) );
  INVx1_ASAP7_75t_SL U33039 ( .A(mult_x_1196_n2861), .Y(n22445) );
  INVx1_ASAP7_75t_SL U33040 ( .A(mult_x_1196_n2385), .Y(n22447) );
  INVx3_ASAP7_75t_SL U33041 ( .A(add_x_735_A_32_), .Y(n23974) );
  INVx5_ASAP7_75t_SL U33042 ( .A(n23622), .Y(add_x_735_A_26_) );
  XNOR2x2_ASAP7_75t_SL U33043 ( .A(u0_0_leon3x0_p0_muli[48]), .B(n23482), .Y(
        n24037) );
  NAND2xp5_ASAP7_75t_SL U33044 ( .A(n25101), .B(n25102), .Y(n23482) );
  OAI22x1_ASAP7_75t_SL U33045 ( .A1(n24007), .A2(mult_x_1196_n3068), .B1(
        n24005), .B2(mult_x_1196_n3067), .Y(mult_x_1196_n2496) );
  MAJIxp5_ASAP7_75t_SL U33046 ( .A(mult_x_1196_n2426), .B(n22452), .C(
        mult_x_1196_n2550), .Y(mult_x_1196_n1735) );
  OAI21xp5_ASAP7_75t_SL U33047 ( .A1(mult_x_1196_n3158), .A2(n23994), .B(
        n22453), .Y(n22452) );
  NAND2xp5_ASAP7_75t_SL U33048 ( .A(n22388), .B(n22454), .Y(n22453) );
  OAI21xp5_ASAP7_75t_SL U33049 ( .A1(n22456), .A2(n22805), .B(n22455), .Y(
        mult_x_1196_n1972) );
  NAND2xp5_ASAP7_75t_SL U33050 ( .A(mult_x_1196_n2010), .B(mult_x_1196_n2012), 
        .Y(n22455) );
  XNOR2xp5_ASAP7_75t_SL U33051 ( .A(n22249), .B(n22858), .Y(n22805) );
  OAI22x1_ASAP7_75t_SL U33052 ( .A1(mult_x_1196_n2986), .A2(n23311), .B1(
        mult_x_1196_n2985), .B2(n24012), .Y(n23874) );
  AO21x1_ASAP7_75t_SL U33053 ( .A1(n24171), .A2(n23262), .B(n22748), .Y(
        mult_x_1196_n2657) );
  XNOR2xp5_ASAP7_75t_SL U33054 ( .A(mult_x_1196_n1965), .B(n22729), .Y(n22457)
         );
  MAJIxp5_ASAP7_75t_SL U33055 ( .A(mult_x_1196_n1574), .B(mult_x_1196_n1566), 
        .C(mult_x_1196_n1568), .Y(n22994) );
  XOR2xp5_ASAP7_75t_SL U33056 ( .A(n22458), .B(n22873), .Y(mult_x_1196_n1574)
         );
  INVx1_ASAP7_75t_SL U33057 ( .A(mult_x_1196_n2325), .Y(n22458) );
  MAJIxp5_ASAP7_75t_SL U33058 ( .A(n23710), .B(mult_x_1196_n2540), .C(
        mult_x_1196_n2480), .Y(n23306) );
  NAND2xp5_ASAP7_75t_SL U33059 ( .A(mult_x_1196_n2133), .B(mult_x_1196_n1866), 
        .Y(n24131) );
  NAND2x1_ASAP7_75t_SL U33060 ( .A(n22460), .B(n22459), .Y(n23435) );
  MAJIxp5_ASAP7_75t_SL U33061 ( .A(mult_x_1196_n1948), .B(mult_x_1196_n2135), 
        .C(mult_x_1196_n2467), .Y(n22608) );
  XNOR2xp5_ASAP7_75t_SL U33062 ( .A(n22461), .B(mult_x_1196_n2527), .Y(
        mult_x_1196_n1948) );
  INVx1_ASAP7_75t_SL U33063 ( .A(mult_x_1196_n2687), .Y(n22461) );
  XNOR2x1_ASAP7_75t_SL U33064 ( .A(n22462), .B(n22570), .Y(mult_x_1196_n1363)
         );
  XNOR2x1_ASAP7_75t_SL U33065 ( .A(mult_x_1196_n1361), .B(n22463), .Y(n22462)
         );
  BUFx6f_ASAP7_75t_SL U33066 ( .A(n23116), .Y(n22464) );
  OAI22xp5_ASAP7_75t_SL U33067 ( .A1(n24287), .A2(n18414), .B1(
        mult_x_1196_n3178), .B2(n23992), .Y(mult_x_1196_n2140) );
  MAJIxp5_ASAP7_75t_SL U33068 ( .A(mult_x_1196_n2580), .B(mult_x_1196_n2548), 
        .C(n23867), .Y(mult_x_1196_n1671) );
  OAI21xp5_ASAP7_75t_SL U33069 ( .A1(mult_x_1196_n3156), .A2(n23081), .B(
        n22465), .Y(mult_x_1196_n2580) );
  NAND2xp5_ASAP7_75t_SL U33070 ( .A(n22388), .B(n22466), .Y(n22465) );
  INVx1_ASAP7_75t_SL U33071 ( .A(mult_x_1196_n3155), .Y(n22466) );
  BUFx6f_ASAP7_75t_SL U33072 ( .A(n18919), .Y(n23100) );
  BUFx2_ASAP7_75t_SL U33073 ( .A(n24076), .Y(n22578) );
  INVx1_ASAP7_75t_SL U33074 ( .A(n23639), .Y(n23643) );
  MAJIxp5_ASAP7_75t_SL U33075 ( .A(n22469), .B(mult_x_1196_n2129), .C(
        mult_x_1196_n2359), .Y(mult_x_1196_n1636) );
  XOR2xp5_ASAP7_75t_SL U33076 ( .A(n22471), .B(n22470), .Y(mult_x_1196_n1637)
         );
  INVx1_ASAP7_75t_SL U33077 ( .A(mult_x_1196_n2359), .Y(n22470) );
  HB1xp67_ASAP7_75t_SL U33078 ( .A(n18380), .Y(n22472) );
  MAJIxp5_ASAP7_75t_SL U33079 ( .A(n23750), .B(n22292), .C(n22473), .Y(
        mult_x_1196_n1751) );
  MAJIxp5_ASAP7_75t_SL U33080 ( .A(mult_x_1196_n2333), .B(n24182), .C(
        mult_x_1196_n2649), .Y(n23750) );
  XOR2xp5_ASAP7_75t_SL U33081 ( .A(mult_x_1196_n2637), .B(mult_x_1196_n2231), 
        .Y(n23420) );
  AO21x1_ASAP7_75t_SL U33082 ( .A1(n23984), .A2(n24082), .B(mult_x_1196_n3213), 
        .Y(mult_x_1196_n2637) );
  INVx4_ASAP7_75t_SL U33083 ( .A(n22285), .Y(n23972) );
  XNOR2x1_ASAP7_75t_SL U33084 ( .A(n22474), .B(n22529), .Y(mult_x_1196_n1198)
         );
  INVx1_ASAP7_75t_SL U33085 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__11_), .Y(
        n25138) );
  NAND2x1p5_ASAP7_75t_SL U33086 ( .A(n23489), .B(n23516), .Y(n23998) );
  MAJIxp5_ASAP7_75t_SL U33087 ( .A(n24297), .B(n23924), .C(n22943), .Y(
        mult_x_1196_n1200) );
  MAJIxp5_ASAP7_75t_SL U33088 ( .A(mult_x_1196_n1235), .B(mult_x_1196_n1253), 
        .C(mult_x_1196_n1249), .Y(n23924) );
  HB1xp67_ASAP7_75t_SL U33089 ( .A(mult_x_1196_n1809), .Y(n22475) );
  BUFx2_ASAP7_75t_SL U33090 ( .A(n24038), .Y(n22509) );
  XNOR2x1_ASAP7_75t_SL U33091 ( .A(n22476), .B(n22477), .Y(mult_x_1196_n1597)
         );
  XOR2x1_ASAP7_75t_SL U33092 ( .A(mult_x_1196_n1610), .B(mult_x_1196_n1604), 
        .Y(n22476) );
  XNOR2x1_ASAP7_75t_SL U33093 ( .A(mult_x_1196_n2006), .B(n22478), .Y(
        mult_x_1196_n2004) );
  BUFx3_ASAP7_75t_SL U33094 ( .A(n23985), .Y(n22953) );
  XOR2xp5_ASAP7_75t_SL U33095 ( .A(mult_x_1196_n1553), .B(mult_x_1196_n1510), 
        .Y(n23503) );
  XOR2xp5_ASAP7_75t_SL U33096 ( .A(mult_x_1196_n1563), .B(n23372), .Y(
        mult_x_1196_n1510) );
  XNOR2xp5_ASAP7_75t_SL U33097 ( .A(mult_x_1196_n1187), .B(n23174), .Y(n23173)
         );
  OAI21xp5_ASAP7_75t_SL U33098 ( .A1(mult_x_1196_n2256), .A2(n22479), .B(
        n23652), .Y(mult_x_1196_n1187) );
  NAND2xp5_ASAP7_75t_SL U33099 ( .A(mult_x_1196_n2410), .B(mult_x_1196_n2506), 
        .Y(n22480) );
  NAND2x1_ASAP7_75t_SL U33100 ( .A(mult_x_1196_n1427), .B(mult_x_1196_n1426), 
        .Y(mult_x_1196_n579) );
  XNOR2x1_ASAP7_75t_SL U33101 ( .A(add_x_735_A_25_), .B(n24692), .Y(n24028) );
  HB1xp67_ASAP7_75t_SL U33102 ( .A(mult_x_1196_n1863), .Y(n22484) );
  INVx1_ASAP7_75t_SL U33103 ( .A(mult_x_1196_n2551), .Y(n23340) );
  OAI22xp5_ASAP7_75t_SL U33104 ( .A1(n23997), .A2(mult_x_1196_n3126), .B1(
        mult_x_1196_n3127), .B2(n24000), .Y(mult_x_1196_n2551) );
  XOR2xp5_ASAP7_75t_SL U33105 ( .A(n22253), .B(mult_x_1196_n1766), .Y(n22485)
         );
  XOR2xp5_ASAP7_75t_SL U33106 ( .A(mult_x_1196_n2622), .B(mult_x_1196_n2402), 
        .Y(n23762) );
  OAI22xp5_ASAP7_75t_SL U33107 ( .A1(n23522), .A2(mult_x_1196_n3198), .B1(
        mult_x_1196_n3197), .B2(n23987), .Y(mult_x_1196_n2622) );
  NOR2x1p5_ASAP7_75t_SL U33108 ( .A(mult_x_1196_n1191), .B(n24311), .Y(
        mult_x_1196_n519) );
  HB1xp67_ASAP7_75t_SL U33109 ( .A(mult_x_1196_n1448), .Y(n22486) );
  HB1xp67_ASAP7_75t_SL U33110 ( .A(n24022), .Y(n22487) );
  XOR2x2_ASAP7_75t_SL U33111 ( .A(n24070), .B(n23076), .Y(mult_x_1196_n2797)
         );
  OAI21x1_ASAP7_75t_SL U33112 ( .A1(n22322), .A2(n18410), .B(n24275), .Y(
        mult_x_1196_n1459) );
  MAJIxp5_ASAP7_75t_SL U33113 ( .A(mult_x_1196_n2383), .B(mult_x_1196_n2539), 
        .C(n22794), .Y(mult_x_1196_n1348) );
  OAI21xp5_ASAP7_75t_SL U33114 ( .A1(mult_x_1196_n2987), .A2(n24014), .B(
        n22301), .Y(n22794) );
  INVx2_ASAP7_75t_SL U33115 ( .A(mult_x_1196_n1094), .Y(n24097) );
  XNOR2xp5_ASAP7_75t_SL U33116 ( .A(mult_x_1196_n2000), .B(n23438), .Y(n23039)
         );
  XNOR2xp5_ASAP7_75t_SL U33117 ( .A(n22489), .B(n22488), .Y(mult_x_1196_n1274)
         );
  XOR2xp5_ASAP7_75t_SL U33118 ( .A(n22348), .B(mult_x_1196_n1284), .Y(n22488)
         );
  INVx1_ASAP7_75t_SL U33119 ( .A(n22799), .Y(n22489) );
  XNOR2x1_ASAP7_75t_SL U33120 ( .A(mult_x_1196_n2334), .B(n22732), .Y(n22731)
         );
  NOR2x1p5_ASAP7_75t_SL U33121 ( .A(n22492), .B(n22491), .Y(mult_x_1196_n464)
         );
  XNOR2xp5_ASAP7_75t_SL U33122 ( .A(n24057), .B(n23955), .Y(mult_x_1196_n3226)
         );
  INVx1_ASAP7_75t_SL U33123 ( .A(u0_0_leon3x0_p0_muli[47]), .Y(n23707) );
  INVx4_ASAP7_75t_SL U33124 ( .A(n23962), .Y(n23396) );
  NAND2xp33_ASAP7_75t_SL U33125 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__27_), 
        .B(n18911), .Y(n25140) );
  BUFx6f_ASAP7_75t_SL U33126 ( .A(n23983), .Y(n23358) );
  XNOR2xp5_ASAP7_75t_SL U33127 ( .A(mult_x_1196_n2606), .B(n24211), .Y(n22703)
         );
  OAI22x1_ASAP7_75t_SL U33128 ( .A1(mult_x_1196_n3181), .A2(n23987), .B1(
        mult_x_1196_n3182), .B2(n23989), .Y(mult_x_1196_n2606) );
  NAND2x1p5_ASAP7_75t_SL U33129 ( .A(n22298), .B(n23273), .Y(mult_x_1196_n1927) );
  XNOR2xp5_ASAP7_75t_SL U33130 ( .A(mult_x_1196_n2135), .B(n22790), .Y(n22494)
         );
  OAI22xp5_ASAP7_75t_SL U33131 ( .A1(mult_x_1196_n3102), .A2(n23100), .B1(
        n24002), .B2(mult_x_1196_n3101), .Y(mult_x_1196_n2526) );
  MAJIxp5_ASAP7_75t_SL U33132 ( .A(n22981), .B(mult_x_1196_n2390), .C(
        mult_x_1196_n2300), .Y(mult_x_1196_n1603) );
  OAI21x1_ASAP7_75t_SL U33133 ( .A1(add_x_735_n256), .A2(add_x_735_n254), .B(
        add_x_735_n255), .Y(add_x_735_n253) );
  XOR2x2_ASAP7_75t_SL U33134 ( .A(n22993), .B(mult_x_1196_n1527), .Y(
        mult_x_1196_n1517) );
  XNOR2xp5_ASAP7_75t_SL U33135 ( .A(mult_x_1196_n1264), .B(mult_x_1196_n1274), 
        .Y(n23196) );
  INVx1_ASAP7_75t_SL U33136 ( .A(n22497), .Y(n22495) );
  XOR2xp5_ASAP7_75t_SL U33137 ( .A(n22496), .B(mult_x_1196_n926), .Y(
        mult_x_1196_n924) );
  XOR2xp5_ASAP7_75t_SL U33138 ( .A(n22497), .B(mult_x_1196_n944), .Y(n22496)
         );
  MAJx2_ASAP7_75t_SL U33139 ( .A(mult_x_1196_n2277), .B(n23275), .C(
        mult_x_1196_n2152), .Y(n22497) );
  XNOR2xp5_ASAP7_75t_SL U33140 ( .A(n22498), .B(mult_x_1196_n1643), .Y(n22785)
         );
  XNOR2xp5_ASAP7_75t_SL U33141 ( .A(n24123), .B(n24124), .Y(mult_x_1196_n1643)
         );
  INVx1_ASAP7_75t_SL U33142 ( .A(mult_x_1196_n1639), .Y(n22498) );
  MAJIxp5_ASAP7_75t_SL U33143 ( .A(mult_x_1196_n1039), .B(n22257), .C(
        mult_x_1196_n1020), .Y(mult_x_1196_n1016) );
  NAND2xp5_ASAP7_75t_SL U33144 ( .A(mult_x_1196_n1036), .B(mult_x_1196_n1017), 
        .Y(mult_x_1196_n451) );
  INVx1_ASAP7_75t_SL U33145 ( .A(mult_x_1196_n1023), .Y(n22499) );
  MAJIxp5_ASAP7_75t_SL U33146 ( .A(n22500), .B(mult_x_1196_n1209), .C(
        mult_x_1196_n1178), .Y(mult_x_1196_n1169) );
  XNOR2xp5_ASAP7_75t_SL U33147 ( .A(mult_x_1196_n1209), .B(n22502), .Y(n22501)
         );
  NAND2xp5_ASAP7_75t_SL U33148 ( .A(n23265), .B(n23653), .Y(n23652) );
  HB1xp67_ASAP7_75t_SL U33149 ( .A(mult_x_1196_n594), .Y(n22503) );
  HB1xp67_ASAP7_75t_SL U33150 ( .A(n24198), .Y(n22504) );
  XOR2xp5_ASAP7_75t_SL U33151 ( .A(n23932), .B(mult_x_1196_n2521), .Y(
        mult_x_1196_n1819) );
  NOR2x1_ASAP7_75t_SL U33152 ( .A(mult_x_1196_n564), .B(mult_x_1196_n557), .Y(
        mult_x_1196_n555) );
  XNOR2x2_ASAP7_75t_SL U33153 ( .A(mult_x_1196_n1336), .B(n22505), .Y(n22884)
         );
  XNOR2xp5_ASAP7_75t_SL U33154 ( .A(mult_x_1196_n1344), .B(n22311), .Y(n22505)
         );
  AOI21xp5_ASAP7_75t_SL U33155 ( .A1(n23106), .A2(mult_x_1196_n1790), .B(
        mult_x_1196_n1794), .Y(n23096) );
  MAJIxp5_ASAP7_75t_SL U33156 ( .A(mult_x_1196_n1818), .B(mult_x_1196_n2520), 
        .C(n23659), .Y(mult_x_1196_n1794) );
  XNOR2x1_ASAP7_75t_SL U33157 ( .A(n22863), .B(n22506), .Y(mult_x_1196_n2070)
         );
  INVx1_ASAP7_75t_SL U33158 ( .A(n22862), .Y(n22506) );
  XOR2xp5_ASAP7_75t_SL U33159 ( .A(mult_x_1196_n2140), .B(n23563), .Y(n22862)
         );
  BUFx3_ASAP7_75t_SL U33160 ( .A(n23993), .Y(n23994) );
  INVx1_ASAP7_75t_SL U33161 ( .A(mult_x_1196_n1322), .Y(n23856) );
  MAJIxp5_ASAP7_75t_SL U33162 ( .A(n23156), .B(mult_x_1196_n2493), .C(
        mult_x_1196_n2585), .Y(mult_x_1196_n1814) );
  OAI21xp5_ASAP7_75t_SL U33163 ( .A1(mult_x_1196_n3161), .A2(n23994), .B(
        n22507), .Y(mult_x_1196_n2585) );
  NAND2xp5_ASAP7_75t_SL U33164 ( .A(n22388), .B(n22508), .Y(n22507) );
  XNOR2xp5_ASAP7_75t_SL U33165 ( .A(n18936), .B(mult_x_1196_n1833), .Y(n23133)
         );
  NOR2x1p5_ASAP7_75t_SL U33166 ( .A(n23935), .B(n22227), .Y(n22580) );
  XNOR2x2_ASAP7_75t_SL U33167 ( .A(n23217), .B(n23518), .Y(mult_x_1196_n1712)
         );
  AOI21x1_ASAP7_75t_SL U33168 ( .A1(mult_x_1196_n2130), .A2(mult_x_1196_n1712), 
        .B(n23728), .Y(n23727) );
  HB1xp67_ASAP7_75t_SL U33169 ( .A(mult_x_1196_n655), .Y(n22510) );
  INVx3_ASAP7_75t_SL U33170 ( .A(n23983), .Y(n24120) );
  BUFx6f_ASAP7_75t_SL U33171 ( .A(u0_0_leon3x0_p0_muli[17]), .Y(n24070) );
  XNOR2xp5_ASAP7_75t_SL U33172 ( .A(mult_x_1196_n1069), .B(n22512), .Y(
        mult_x_1196_n1064) );
  XOR2xp5_ASAP7_75t_SL U33173 ( .A(mult_x_1196_n1090), .B(mult_x_1196_n1072), 
        .Y(n22512) );
  NAND2xp5_ASAP7_75t_SL U33174 ( .A(mult_x_1196_n465), .B(n23674), .Y(n23675)
         );
  BUFx2_ASAP7_75t_SL U33175 ( .A(mult_x_1196_n1500), .Y(n22514) );
  XOR2x2_ASAP7_75t_SL U33176 ( .A(n24693), .B(n23424), .Y(n23571) );
  XOR2xp5_ASAP7_75t_SL U33177 ( .A(n23183), .B(n22515), .Y(n23377) );
  XNOR2xp5_ASAP7_75t_SL U33178 ( .A(n24243), .B(mult_x_1196_n2629), .Y(n22515)
         );
  XNOR2xp5_ASAP7_75t_SL U33179 ( .A(n18315), .B(n22516), .Y(mult_x_1196_n1479)
         );
  XOR2xp5_ASAP7_75t_SL U33180 ( .A(mult_x_1196_n1524), .B(mult_x_1196_n1488), 
        .Y(n22516) );
  INVx2_ASAP7_75t_SL U33181 ( .A(n22928), .Y(n23197) );
  OR2x2_ASAP7_75t_SL U33182 ( .A(mult_x_1196_n948), .B(mult_x_1196_n963), .Y(
        mult_x_1196_n785) );
  XOR2xp5_ASAP7_75t_SL U33183 ( .A(mult_x_1196_n1348), .B(n22594), .Y(
        mult_x_1196_n1310) );
  XNOR2xp5_ASAP7_75t_SL U33184 ( .A(mult_x_1196_n2375), .B(n22518), .Y(
        mult_x_1196_n1100) );
  XOR2xp5_ASAP7_75t_SL U33185 ( .A(mult_x_1196_n2439), .B(mult_x_1196_n2407), 
        .Y(n22518) );
  MAJx2_ASAP7_75t_SL U33186 ( .A(mult_x_1196_n2374), .B(n23255), .C(
        mult_x_1196_n2342), .Y(mult_x_1196_n1049) );
  MAJIxp5_ASAP7_75t_SL U33187 ( .A(mult_x_1196_n2149), .B(mult_x_1196_n2242), 
        .C(n22520), .Y(mult_x_1196_n898) );
  XNOR2xp5_ASAP7_75t_SL U33188 ( .A(mult_x_1196_n2149), .B(n22519), .Y(
        mult_x_1196_n899) );
  XOR2xp5_ASAP7_75t_SL U33189 ( .A(n22520), .B(mult_x_1196_n2242), .Y(n22519)
         );
  OAI22xp5_ASAP7_75t_SL U33190 ( .A1(n24031), .A2(mult_x_1196_n2840), .B1(
        n24030), .B2(mult_x_1196_n2839), .Y(n22520) );
  MAJIxp5_ASAP7_75t_SL U33191 ( .A(n23537), .B(n23538), .C(mult_x_1196_n1006), 
        .Y(n23928) );
  INVx2_ASAP7_75t_SL U33192 ( .A(mult_x_1196_n360), .Y(mult_x_1196_n358) );
  BUFx6f_ASAP7_75t_SL U33193 ( .A(n23972), .Y(n23479) );
  MAJIxp5_ASAP7_75t_SL U33194 ( .A(n23928), .B(n22365), .C(mult_x_1196_n982), 
        .Y(mult_x_1196_n978) );
  XOR2xp5_ASAP7_75t_SL U33195 ( .A(n22522), .B(mult_x_1196_n982), .Y(
        mult_x_1196_n979) );
  XNOR2xp5_ASAP7_75t_SL U33196 ( .A(n22365), .B(n23928), .Y(n22522) );
  MAJIxp5_ASAP7_75t_SL U33197 ( .A(mult_x_1196_n928), .B(mult_x_1196_n940), 
        .C(mult_x_1196_n937), .Y(mult_x_1196_n921) );
  XNOR2xp5_ASAP7_75t_SL U33198 ( .A(mult_x_1196_n924), .B(n22362), .Y(n22524)
         );
  XNOR2xp5_ASAP7_75t_SL U33199 ( .A(mult_x_1196_n937), .B(n22526), .Y(n22525)
         );
  XOR2xp5_ASAP7_75t_SL U33200 ( .A(mult_x_1196_n940), .B(n22527), .Y(n22526)
         );
  NOR2x1_ASAP7_75t_SL U33201 ( .A(mult_x_1196_n1103), .B(n24251), .Y(n22656)
         );
  NOR2x1_ASAP7_75t_SL U33202 ( .A(mult_x_1196_n2886), .B(n24026), .Y(n24126)
         );
  BUFx2_ASAP7_75t_SL U33203 ( .A(mult_x_1196_n794), .Y(n22663) );
  XOR2xp5_ASAP7_75t_SL U33204 ( .A(mult_x_1196_n874), .B(n22530), .Y(n23245)
         );
  OAI22xp5_ASAP7_75t_SL U33205 ( .A1(mult_x_1196_n2879), .A2(n24026), .B1(
        mult_x_1196_n2878), .B2(n24025), .Y(n22531) );
  INVx1_ASAP7_75t_SL U33206 ( .A(mult_x_1196_n2371), .Y(n22532) );
  NOR2x1_ASAP7_75t_SL U33207 ( .A(n22534), .B(n23277), .Y(n23792) );
  NOR2x1_ASAP7_75t_SL U33208 ( .A(mult_x_1196_n3168), .B(n24230), .Y(n22534)
         );
  INVx1_ASAP7_75t_SL U33209 ( .A(n22537), .Y(n22535) );
  XNOR2xp5_ASAP7_75t_SL U33210 ( .A(n22537), .B(mult_x_1196_n1763), .Y(n22536)
         );
  INVx3_ASAP7_75t_SL U33211 ( .A(add_x_735_A_16_), .Y(n23963) );
  OAI21xp5_ASAP7_75t_SL U33212 ( .A1(mult_x_1196_n557), .A2(mult_x_1196_n565), 
        .B(mult_x_1196_n558), .Y(mult_x_1196_n556) );
  XNOR2x1_ASAP7_75t_SL U33213 ( .A(n22539), .B(n23939), .Y(n24286) );
  HB1xp67_ASAP7_75t_SL U33214 ( .A(mult_x_1196_n575), .Y(n22541) );
  XNOR2xp5_ASAP7_75t_SL U33215 ( .A(n23403), .B(n22542), .Y(n23241) );
  XNOR2xp5_ASAP7_75t_SL U33216 ( .A(n22250), .B(n23912), .Y(n22542) );
  XOR2xp5_ASAP7_75t_SL U33217 ( .A(mult_x_1196_n2607), .B(mult_x_1196_n2127), 
        .Y(n22646) );
  OAI21x1_ASAP7_75t_SL U33218 ( .A1(mult_x_1196_n3133), .A2(n18397), .B(n22601), .Y(n23519) );
  XNOR2xp5_ASAP7_75t_SL U33219 ( .A(n24062), .B(n23955), .Y(mult_x_1196_n3231)
         );
  AOI21x1_ASAP7_75t_SL U33220 ( .A1(n24254), .A2(mult_x_1196_n771), .B(n23246), 
        .Y(mult_x_1196_n766) );
  MAJIxp5_ASAP7_75t_SL U33221 ( .A(n23606), .B(n23192), .C(n23108), .Y(n23691)
         );
  INVx4_ASAP7_75t_SL U33222 ( .A(add_x_735_A_12_), .Y(n23961) );
  NOR2x1_ASAP7_75t_SL U33223 ( .A(n24121), .B(mult_x_1196_n3232), .Y(n23189)
         );
  XNOR2xp5_ASAP7_75t_SL U33224 ( .A(n24063), .B(n23955), .Y(mult_x_1196_n3232)
         );
  XNOR2xp5_ASAP7_75t_SL U33225 ( .A(mult_x_1196_n2294), .B(mult_x_1196_n2230), 
        .Y(n22544) );
  INVx1_ASAP7_75t_SL U33226 ( .A(n23865), .Y(n22545) );
  MAJIxp5_ASAP7_75t_SL U33227 ( .A(mult_x_1196_n1658), .B(n22547), .C(
        mult_x_1196_n1691), .Y(mult_x_1196_n1653) );
  MAJIxp5_ASAP7_75t_SL U33228 ( .A(n23238), .B(mult_x_1196_n1699), .C(
        mult_x_1196_n1697), .Y(n22547) );
  NOR2x1_ASAP7_75t_SL U33229 ( .A(n22549), .B(n22548), .Y(n24431) );
  INVx1_ASAP7_75t_SL U33230 ( .A(n24687), .Y(n22548) );
  INVx1_ASAP7_75t_SL U33231 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__0_), .Y(n22549)
         );
  OAI22x1_ASAP7_75t_SL U33232 ( .A1(mult_x_1196_n2892), .A2(n24026), .B1(
        mult_x_1196_n2891), .B2(n22983), .Y(n23742) );
  NAND2xp5_ASAP7_75t_SL U33233 ( .A(n22551), .B(n23388), .Y(n23392) );
  AOI31xp67_ASAP7_75t_SL U33234 ( .A1(n23926), .A2(n23385), .A3(n23391), .B(
        n23390), .Y(n22551) );
  NAND2x1p5_ASAP7_75t_SL U33235 ( .A(n24016), .B(n23143), .Y(n24018) );
  BUFx2_ASAP7_75t_SL U33236 ( .A(n24029), .Y(n22743) );
  INVx6_ASAP7_75t_SL U33237 ( .A(n22962), .Y(n24030) );
  NAND2xp5_ASAP7_75t_SL U33238 ( .A(mult_x_1196_n1455), .B(n22552), .Y(n22771)
         );
  NAND2xp5_ASAP7_75t_SL U33239 ( .A(mult_x_1196_n1487), .B(n23318), .Y(n22552)
         );
  XOR2x2_ASAP7_75t_SL U33240 ( .A(mult_x_1196_n1373), .B(mult_x_1196_n1345), 
        .Y(n23057) );
  XNOR2x1_ASAP7_75t_SL U33241 ( .A(n22739), .B(n23057), .Y(n22905) );
  OAI22xp5_ASAP7_75t_SL U33242 ( .A1(n22961), .A2(n23637), .B1(n24005), .B2(
        mult_x_1196_n3076), .Y(mult_x_1196_n2137) );
  HB1xp67_ASAP7_75t_SL U33243 ( .A(n18985), .Y(n22553) );
  MAJx2_ASAP7_75t_SL U33244 ( .A(mult_x_1196_n1156), .B(mult_x_1196_n1158), 
        .C(mult_x_1196_n1154), .Y(mult_x_1196_n1092) );
  MAJx2_ASAP7_75t_SL U33245 ( .A(mult_x_1196_n1605), .B(mult_x_1196_n1609), 
        .C(mult_x_1196_n1603), .Y(n22589) );
  XOR2xp5_ASAP7_75t_SL U33246 ( .A(n22554), .B(n22753), .Y(mult_x_1196_n1037)
         );
  INVx1_ASAP7_75t_SL U33247 ( .A(n23495), .Y(n22554) );
  XNOR2xp5_ASAP7_75t_SL U33248 ( .A(mult_x_1196_n1966), .B(mult_x_1196_n1962), 
        .Y(n22555) );
  INVx1_ASAP7_75t_SL U33249 ( .A(mult_x_1196_n1474), .Y(n24095) );
  MAJIxp5_ASAP7_75t_SL U33250 ( .A(n22728), .B(mult_x_1196_n1516), .C(n23268), 
        .Y(mult_x_1196_n1474) );
  XNOR2xp5_ASAP7_75t_SL U33251 ( .A(n22559), .B(mult_x_1196_n943), .Y(n22558)
         );
  NAND2xp5_ASAP7_75t_SL U33252 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__25_), .B(
        n18910), .Y(n24553) );
  AND2x4_ASAP7_75t_SL U33253 ( .A(n23623), .B(n24553), .Y(n23622) );
  MAJIxp5_ASAP7_75t_SL U33254 ( .A(mult_x_1196_n1148), .B(mult_x_1196_n1175), 
        .C(n22560), .Y(mult_x_1196_n1141) );
  INVx1_ASAP7_75t_SL U33255 ( .A(n22562), .Y(n22560) );
  XNOR2xp5_ASAP7_75t_SL U33256 ( .A(n22562), .B(mult_x_1196_n1175), .Y(n22561)
         );
  XOR2xp5_ASAP7_75t_SL U33257 ( .A(n23175), .B(n23173), .Y(n22562) );
  INVx2_ASAP7_75t_SL U33258 ( .A(mult_x_1196_n488), .Y(mult_x_1196_n793) );
  INVx2_ASAP7_75t_SL U33259 ( .A(mult_x_1196_n1440), .Y(n22967) );
  XOR2xp5_ASAP7_75t_SL U33260 ( .A(mult_x_1196_n2490), .B(n22564), .Y(
        mult_x_1196_n1738) );
  NAND2x1p5_ASAP7_75t_SL U33261 ( .A(n23638), .B(mult_x_1196_n60), .Y(n24006)
         );
  XOR2xp5_ASAP7_75t_SL U33262 ( .A(mult_x_1196_n2302), .B(n23332), .Y(n23331)
         );
  OAI22xp5_ASAP7_75t_SL U33263 ( .A1(mult_x_1196_n2868), .A2(n23449), .B1(
        n22743), .B2(mult_x_1196_n2867), .Y(mult_x_1196_n2302) );
  MAJIxp5_ASAP7_75t_SL U33264 ( .A(n23647), .B(mult_x_1196_n1536), .C(
        mult_x_1196_n1534), .Y(n23337) );
  MAJx2_ASAP7_75t_SL U33265 ( .A(mult_x_1196_n1707), .B(mult_x_1196_n1666), 
        .C(mult_x_1196_n1709), .Y(mult_x_1196_n1629) );
  OAI21x1_ASAP7_75t_SL U33266 ( .A1(add_x_735_n216), .A2(n18894), .B(
        add_x_735_n217), .Y(add_x_735_n215) );
  INVx1_ASAP7_75t_SL U33267 ( .A(mult_x_1196_n3233), .Y(n24171) );
  XNOR2xp5_ASAP7_75t_SL U33268 ( .A(n23030), .B(mult_x_1196_n1188), .Y(n23029)
         );
  XNOR2x1_ASAP7_75t_SL U33269 ( .A(n23124), .B(n22648), .Y(mult_x_1196_n1440)
         );
  BUFx2_ASAP7_75t_SL U33270 ( .A(n24037), .Y(n22936) );
  XNOR2x2_ASAP7_75t_SL U33271 ( .A(n22899), .B(n22898), .Y(mult_x_1196_n1376)
         );
  XOR2xp5_ASAP7_75t_SL U33272 ( .A(mult_x_1196_n1435), .B(n22602), .Y(n24089)
         );
  XNOR2xp5_ASAP7_75t_SL U33273 ( .A(add_x_735_A_25_), .B(add_x_735_A_26_), .Y(
        n24113) );
  NOR2x1p5_ASAP7_75t_SL U33274 ( .A(n23313), .B(n23312), .Y(n23428) );
  INVx1_ASAP7_75t_SL U33275 ( .A(n22757), .Y(n22566) );
  NAND2xp5_ASAP7_75t_SL U33276 ( .A(n22567), .B(n22388), .Y(n24267) );
  INVx8_ASAP7_75t_SL U33277 ( .A(n23935), .Y(n23967) );
  MAJIxp5_ASAP7_75t_SL U33278 ( .A(mult_x_1196_n1128), .B(mult_x_1196_n1126), 
        .C(mult_x_1196_n1130), .Y(mult_x_1196_n1095) );
  XNOR2xp5_ASAP7_75t_SL U33279 ( .A(mult_x_1196_n1130), .B(n22568), .Y(
        mult_x_1196_n1096) );
  XNOR2xp5_ASAP7_75t_SL U33280 ( .A(n22569), .B(mult_x_1196_n1128), .Y(n22568)
         );
  INVx1_ASAP7_75t_SL U33281 ( .A(mult_x_1196_n1126), .Y(n22569) );
  XNOR2x1_ASAP7_75t_SL U33282 ( .A(n22773), .B(mult_x_1196_n1198), .Y(
        mult_x_1196_n1191) );
  XNOR2xp5_ASAP7_75t_SL U33283 ( .A(n22751), .B(n22643), .Y(n24309) );
  BUFx2_ASAP7_75t_SL U33284 ( .A(n23860), .Y(n22772) );
  XNOR2xp5_ASAP7_75t_SL U33285 ( .A(mult_x_1196_n2275), .B(n22572), .Y(
        mult_x_1196_n913) );
  MAJIxp5_ASAP7_75t_SL U33286 ( .A(mult_x_1196_n2275), .B(mult_x_1196_n2150), 
        .C(n22573), .Y(mult_x_1196_n912) );
  OAI22xp5_ASAP7_75t_SL U33287 ( .A1(mult_x_1196_n2777), .A2(n22509), .B1(
        mult_x_1196_n2776), .B2(n22481), .Y(n22573) );
  BUFx6f_ASAP7_75t_SL U33288 ( .A(n24006), .Y(n24007) );
  XNOR2x1_ASAP7_75t_SL U33289 ( .A(n22574), .B(n23470), .Y(mult_x_1196_n1509)
         );
  XNOR2x1_ASAP7_75t_SL U33290 ( .A(mult_x_1196_n1548), .B(mult_x_1196_n1517), 
        .Y(n22574) );
  MAJIxp5_ASAP7_75t_SL U33291 ( .A(n22576), .B(mult_x_1196_n1214), .C(n22577), 
        .Y(mult_x_1196_n1172) );
  XOR2xp5_ASAP7_75t_SL U33292 ( .A(mult_x_1196_n1214), .B(n22576), .Y(n22575)
         );
  XNOR2xp5_ASAP7_75t_SL U33293 ( .A(n23202), .B(mult_x_1196_n1218), .Y(n22576)
         );
  MAJIxp5_ASAP7_75t_SL U33294 ( .A(n22310), .B(mult_x_1196_n1219), .C(
        mult_x_1196_n1223), .Y(n22577) );
  OAI21x1_ASAP7_75t_SL U33295 ( .A1(mult_x_1196_n2863), .A2(n24031), .B(n23773), .Y(n24227) );
  NOR2x1p5_ASAP7_75t_SL U33296 ( .A(n22269), .B(n23850), .Y(n25644) );
  INVx1_ASAP7_75t_SL U33297 ( .A(n22580), .Y(n22579) );
  OAI22x1_ASAP7_75t_SL U33298 ( .A1(mult_x_1196_n2922), .A2(n24021), .B1(
        n24020), .B2(mult_x_1196_n2921), .Y(mult_x_1196_n2350) );
  INVx2_ASAP7_75t_SL U33299 ( .A(mult_x_1196_n3098), .Y(n22583) );
  OAI21x1_ASAP7_75t_SL U33300 ( .A1(mult_x_1196_n2925), .A2(n24022), .B(n22352), .Y(mult_x_1196_n2353) );
  MAJIxp5_ASAP7_75t_SL U33301 ( .A(mult_x_1196_n1100), .B(mult_x_1196_n1104), 
        .C(mult_x_1196_n1092), .Y(mult_x_1196_n1093) );
  OAI22x1_ASAP7_75t_SL U33302 ( .A1(n24287), .A2(mult_x_1196_n3150), .B1(
        n23992), .B2(mult_x_1196_n3149), .Y(mult_x_1196_n2574) );
  MAJIxp5_ASAP7_75t_SL U33303 ( .A(mult_x_1196_n1265), .B(mult_x_1196_n1267), 
        .C(mult_x_1196_n1234), .Y(mult_x_1196_n1229) );
  XNOR2xp5_ASAP7_75t_SL U33304 ( .A(mult_x_1196_n1234), .B(n22585), .Y(
        mult_x_1196_n1230) );
  XNOR2xp5_ASAP7_75t_SL U33305 ( .A(n22586), .B(mult_x_1196_n1265), .Y(n22585)
         );
  INVx1_ASAP7_75t_SL U33306 ( .A(mult_x_1196_n1267), .Y(n22586) );
  NAND2x1p5_ASAP7_75t_SL U33307 ( .A(mult_x_1196_n3320), .B(mult_x_1196_n96), 
        .Y(mult_x_1196_n99) );
  XNOR2x1_ASAP7_75t_SL U33308 ( .A(n22587), .B(n22722), .Y(mult_x_1196_n1750)
         );
  XOR2x2_ASAP7_75t_SL U33309 ( .A(mult_x_1196_n1755), .B(mult_x_1196_n1781), 
        .Y(n22587) );
  BUFx10_ASAP7_75t_SL U33310 ( .A(add_x_735_A_24_), .Y(n23089) );
  MAJx2_ASAP7_75t_SL U33311 ( .A(n23319), .B(n22370), .C(n23317), .Y(
        mult_x_1196_n1361) );
  MAJIxp5_ASAP7_75t_SL U33312 ( .A(mult_x_1196_n2295), .B(mult_x_1196_n2385), 
        .C(mult_x_1196_n2605), .Y(mult_x_1196_n1418) );
  XNOR2xp5_ASAP7_75t_SL U33313 ( .A(mult_x_1196_n2605), .B(n22588), .Y(
        mult_x_1196_n1419) );
  MAJIxp5_ASAP7_75t_SL U33314 ( .A(mult_x_1196_n966), .B(mult_x_1196_n962), 
        .C(mult_x_1196_n981), .Y(mult_x_1196_n963) );
  XNOR2xp5_ASAP7_75t_SL U33315 ( .A(mult_x_1196_n962), .B(mult_x_1196_n981), 
        .Y(n22590) );
  HB1xp67_ASAP7_75t_SL U33316 ( .A(mult_x_1196_n695), .Y(n22592) );
  OAI21x1_ASAP7_75t_SL U33317 ( .A1(mult_x_1196_n2836), .A2(n24034), .B(n22715), .Y(n23332) );
  XNOR2xp5_ASAP7_75t_SL U33318 ( .A(mult_x_1196_n2473), .B(mult_x_1196_n2409), 
        .Y(n22593) );
  BUFx2_ASAP7_75t_SL U33319 ( .A(n23989), .Y(n22802) );
  OR2x2_ASAP7_75t_SL U33320 ( .A(n23996), .B(mult_x_1196_n3132), .Y(n22601) );
  INVx1_ASAP7_75t_SL U33321 ( .A(mult_x_1196_n1512), .Y(n23466) );
  XNOR2xp5_ASAP7_75t_SL U33322 ( .A(n23503), .B(n22775), .Y(mult_x_1196_n1512)
         );
  OAI22xp5_ASAP7_75t_SL U33323 ( .A1(n22599), .A2(n22598), .B1(n26224), .B2(
        n24686), .Y(u0_0_leon3x0_p0_muli[47]) );
  INVx1_ASAP7_75t_SL U33324 ( .A(n18862), .Y(n22598) );
  HB1xp67_ASAP7_75t_SL U33325 ( .A(mult_x_1196_n1476), .Y(n22600) );
  MAJx2_ASAP7_75t_SL U33326 ( .A(n23243), .B(n18590), .C(mult_x_1196_n1473), 
        .Y(mult_x_1196_n1427) );
  NAND2x1p5_ASAP7_75t_SL U33327 ( .A(n23126), .B(n22582), .Y(n22917) );
  XNOR2xp5_ASAP7_75t_SL U33328 ( .A(n24213), .B(mult_x_1196_n2298), .Y(
        mult_x_1196_n1531) );
  XNOR2xp5_ASAP7_75t_SL U33329 ( .A(mult_x_1196_n1448), .B(mult_x_1196_n1446), 
        .Y(n22602) );
  XOR2xp5_ASAP7_75t_SL U33330 ( .A(n22603), .B(n23804), .Y(mult_x_1196_n1178)
         );
  INVx1_ASAP7_75t_SL U33331 ( .A(mult_x_1196_n1186), .Y(n22603) );
  XOR2xp5_ASAP7_75t_SL U33332 ( .A(mult_x_1196_n1568), .B(mult_x_1196_n1566), 
        .Y(n24115) );
  XNOR2xp5_ASAP7_75t_SL U33333 ( .A(n22605), .B(n22604), .Y(mult_x_1196_n1568)
         );
  XNOR2xp5_ASAP7_75t_SL U33334 ( .A(mult_x_1196_n2389), .B(mult_x_1196_n2235), 
        .Y(n22604) );
  INVx1_ASAP7_75t_SL U33335 ( .A(mult_x_1196_n2545), .Y(n22605) );
  NAND2xp5_ASAP7_75t_SL U33336 ( .A(mult_x_1196_n2564), .B(mult_x_1196_n2596), 
        .Y(n22607) );
  OAI21xp5_ASAP7_75t_SL U33337 ( .A1(mult_x_1196_n3140), .A2(n23999), .B(
        n22288), .Y(mult_x_1196_n2564) );
  XNOR2x1_ASAP7_75t_SL U33338 ( .A(n22959), .B(n24283), .Y(n22822) );
  XOR2x2_ASAP7_75t_SL U33339 ( .A(n22822), .B(n22823), .Y(mult_x_1196_n1979)
         );
  MAJIxp5_ASAP7_75t_SL U33340 ( .A(n22609), .B(mult_x_1196_n1928), .C(n22608), 
        .Y(mult_x_1196_n1916) );
  NAND2xp5_ASAP7_75t_SL U33341 ( .A(n23605), .B(n23592), .Y(n22609) );
  NAND2x1_ASAP7_75t_SL U33342 ( .A(n24303), .B(n24286), .Y(mult_x_1196_n547)
         );
  XNOR2x1_ASAP7_75t_SL U33343 ( .A(n18927), .B(n24047), .Y(mult_x_1196_n3250)
         );
  XOR2xp5_ASAP7_75t_SL U33344 ( .A(n22613), .B(n22612), .Y(n22611) );
  INVx1_ASAP7_75t_SL U33345 ( .A(mult_x_1196_n2437), .Y(n22613) );
  XNOR2xp5_ASAP7_75t_SL U33346 ( .A(n22614), .B(mult_x_1196_n1050), .Y(n22809)
         );
  MAJIxp5_ASAP7_75t_SL U33347 ( .A(mult_x_1196_n1049), .B(mult_x_1196_n2219), 
        .C(mult_x_1196_n2437), .Y(mult_x_1196_n1050) );
  INVx1_ASAP7_75t_SL U33348 ( .A(mult_x_1196_n1029), .Y(n22614) );
  INVx1_ASAP7_75t_SL U33349 ( .A(mult_x_1196_n871), .Y(mult_x_1196_n858) );
  XNOR2x2_ASAP7_75t_SL U33350 ( .A(n22704), .B(n22668), .Y(n23920) );
  XOR2xp5_ASAP7_75t_SL U33351 ( .A(mult_x_1196_n1411), .B(n22615), .Y(
        mult_x_1196_n1372) );
  XNOR2xp5_ASAP7_75t_SL U33352 ( .A(n22308), .B(mult_x_1196_n1378), .Y(n22615)
         );
  BUFx3_ASAP7_75t_SL U33353 ( .A(n23985), .Y(n22647) );
  MAJIxp5_ASAP7_75t_SL U33354 ( .A(n22617), .B(mult_x_1196_n1839), .C(
        mult_x_1196_n1817), .Y(mult_x_1196_n1806) );
  XNOR2xp5_ASAP7_75t_SL U33355 ( .A(mult_x_1196_n1817), .B(n22616), .Y(
        mult_x_1196_n1807) );
  XOR2xp5_ASAP7_75t_SL U33356 ( .A(mult_x_1196_n1839), .B(n22617), .Y(n22616)
         );
  XNOR2xp5_ASAP7_75t_SL U33357 ( .A(mult_x_1196_n2585), .B(n22777), .Y(n22617)
         );
  NAND2xp33_ASAP7_75t_SRAM U33358 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__16_), 
        .B(n24685), .Y(n25094) );
  NOR2x1_ASAP7_75t_SL U33359 ( .A(n22792), .B(mult_x_1196_n3054), .Y(n24223)
         );
  AO21x2_ASAP7_75t_SL U33360 ( .A1(n24165), .A2(n24151), .B(n24166), .Y(n24280) );
  XOR2xp5_ASAP7_75t_SL U33361 ( .A(mult_x_1196_n1887), .B(mult_x_1196_n1883), 
        .Y(n22618) );
  XNOR2xp5_ASAP7_75t_SL U33362 ( .A(n22619), .B(n22623), .Y(mult_x_1196_n1847)
         );
  XOR2xp5_ASAP7_75t_SL U33363 ( .A(n22620), .B(mult_x_1196_n1876), .Y(n22619)
         );
  INVx1_ASAP7_75t_SL U33364 ( .A(n22622), .Y(n22621) );
  NAND2xp5_ASAP7_75t_SL U33365 ( .A(mult_x_1196_n1883), .B(mult_x_1196_n1887), 
        .Y(n22622) );
  XNOR2x2_ASAP7_75t_SL U33366 ( .A(n23419), .B(n23420), .Y(mult_x_1196_n1415)
         );
  XOR2xp5_ASAP7_75t_SL U33367 ( .A(mult_x_1196_n2449), .B(mult_x_1196_n2353), 
        .Y(n22829) );
  XNOR2xp5_ASAP7_75t_SL U33368 ( .A(n22626), .B(n22768), .Y(n22767) );
  INVx1_ASAP7_75t_SL U33369 ( .A(mult_x_1196_n1096), .Y(n22626) );
  XNOR2xp5_ASAP7_75t_SL U33370 ( .A(n22628), .B(n22627), .Y(mult_x_1196_n955)
         );
  XOR2xp5_ASAP7_75t_SL U33371 ( .A(mult_x_1196_n2185), .B(mult_x_1196_n975), 
        .Y(n22627) );
  INVx1_ASAP7_75t_SL U33372 ( .A(n22629), .Y(n22628) );
  MAJIxp5_ASAP7_75t_SL U33373 ( .A(mult_x_1196_n975), .B(n22629), .C(
        mult_x_1196_n953), .Y(mult_x_1196_n954) );
  MAJIxp5_ASAP7_75t_SL U33374 ( .A(mult_x_1196_n2279), .B(n24169), .C(
        mult_x_1196_n2154), .Y(n22629) );
  INVx8_ASAP7_75t_SL U33375 ( .A(n24019), .Y(n24020) );
  OR2x2_ASAP7_75t_SL U33376 ( .A(mult_x_1196_n2323), .B(n24084), .Y(n24215) );
  OAI22xp5_ASAP7_75t_SL U33377 ( .A1(mult_x_1196_n3087), .A2(n18920), .B1(
        mult_x_1196_n3086), .B2(n24002), .Y(n24084) );
  MAJIxp5_ASAP7_75t_SL U33378 ( .A(mult_x_1196_n2292), .B(mult_x_1196_n2199), 
        .C(mult_x_1196_n2228), .Y(mult_x_1196_n1316) );
  XNOR2xp5_ASAP7_75t_SL U33379 ( .A(n22631), .B(n22630), .Y(mult_x_1196_n1317)
         );
  XNOR2xp5_ASAP7_75t_SL U33380 ( .A(mult_x_1196_n2199), .B(mult_x_1196_n2292), 
        .Y(n22630) );
  INVx1_ASAP7_75t_SL U33381 ( .A(mult_x_1196_n2228), .Y(n22631) );
  BUFx2_ASAP7_75t_SL U33382 ( .A(add_x_735_A_26_), .Y(n22897) );
  OAI21x1_ASAP7_75t_SL U33383 ( .A1(mult_x_1196_n3180), .A2(n23522), .B(n22317), .Y(mult_x_1196_n2604) );
  MAJIxp5_ASAP7_75t_SL U33384 ( .A(mult_x_1196_n949), .B(n22340), .C(n22632), 
        .Y(mult_x_1196_n932) );
  INVx1_ASAP7_75t_SL U33385 ( .A(n22633), .Y(n22632) );
  XNOR2xp5_ASAP7_75t_SL U33386 ( .A(n22360), .B(n22634), .Y(n22633) );
  XNOR2xp5_ASAP7_75t_SL U33387 ( .A(mult_x_1196_n954), .B(mult_x_1196_n951), 
        .Y(n22634) );
  NOR2x2_ASAP7_75t_SL U33388 ( .A(mult_x_1196_n3109), .B(n18654), .Y(n23598)
         );
  MAJx2_ASAP7_75t_SL U33389 ( .A(mult_x_1196_n2622), .B(n24148), .C(
        mult_x_1196_n2402), .Y(n23502) );
  NOR2x1_ASAP7_75t_SL U33390 ( .A(mult_x_1196_n645), .B(mult_x_1196_n640), .Y(
        mult_x_1196_n638) );
  MAJIxp5_ASAP7_75t_SL U33391 ( .A(mult_x_1196_n2086), .B(mult_x_1196_n2698), 
        .C(n23078), .Y(mult_x_1196_n2080) );
  OAI22xp5_ASAP7_75t_SL U33392 ( .A1(mult_x_1196_n3274), .A2(n23982), .B1(
        n23980), .B2(mult_x_1196_n3273), .Y(mult_x_1196_n2698) );
  NAND2xp5_ASAP7_75t_SL U33393 ( .A(n22636), .B(n22791), .Y(n24170) );
  XNOR2x1_ASAP7_75t_SL U33394 ( .A(n22844), .B(n22843), .Y(n24312) );
  NAND2x1p5_ASAP7_75t_SL U33395 ( .A(mult_x_1196_n39), .B(
        u0_0_leon3x0_p0_muli[44]), .Y(n24109) );
  NAND2xp5_ASAP7_75t_SL U33396 ( .A(n23158), .B(n23159), .Y(n23157) );
  XNOR2x1_ASAP7_75t_SL U33397 ( .A(n23660), .B(n22871), .Y(n22870) );
  XNOR2xp5_ASAP7_75t_SL U33398 ( .A(n22637), .B(n23544), .Y(n23543) );
  INVx1_ASAP7_75t_SL U33399 ( .A(mult_x_1196_n2690), .Y(n22637) );
  OAI22xp5_ASAP7_75t_SL U33400 ( .A1(mult_x_1196_n3266), .A2(n18319), .B1(
        n22389), .B2(mult_x_1196_n3265), .Y(mult_x_1196_n2690) );
  MAJx2_ASAP7_75t_SL U33401 ( .A(n23304), .B(mult_x_1196_n1480), .C(
        mult_x_1196_n1526), .Y(mult_x_1196_n1435) );
  XNOR2xp5_ASAP7_75t_SL U33402 ( .A(mult_x_1196_n2363), .B(n23379), .Y(n23378)
         );
  XNOR2x2_ASAP7_75t_SL U33403 ( .A(n23380), .B(n23378), .Y(mult_x_1196_n1762)
         );
  NAND2x1p5_ASAP7_75t_SL U33404 ( .A(n24024), .B(n23705), .Y(n24027) );
  INVx1_ASAP7_75t_SL U33405 ( .A(n18539), .Y(mult_x_1196_n623) );
  OR2x2_ASAP7_75t_SL U33406 ( .A(n24270), .B(n18918), .Y(mult_x_1196_n810) );
  NAND2x1_ASAP7_75t_SL U33407 ( .A(n24217), .B(n24219), .Y(n23273) );
  NAND2x1_ASAP7_75t_SL U33408 ( .A(mult_x_1196_n2687), .B(mult_x_1196_n2527), 
        .Y(n24217) );
  XNOR2xp5_ASAP7_75t_SL U33409 ( .A(mult_x_1196_n1408), .B(mult_x_1196_n1405), 
        .Y(n22668) );
  XNOR2x1_ASAP7_75t_SL U33410 ( .A(n24101), .B(n23095), .Y(n24302) );
  XNOR2x2_ASAP7_75t_SL U33411 ( .A(n23457), .B(n23456), .Y(mult_x_1196_n1488)
         );
  INVxp33_ASAP7_75t_SRAM U33412 ( .A(n18918), .Y(n24150) );
  AND2x2_ASAP7_75t_SL U33413 ( .A(n24270), .B(n18918), .Y(mult_x_1196_n626) );
  NOR2x1_ASAP7_75t_SL U33414 ( .A(mult_x_1196_n1796), .B(mult_x_1196_n1772), 
        .Y(mult_x_1196_n645) );
  XNOR2xp5_ASAP7_75t_SL U33415 ( .A(n22820), .B(n22639), .Y(mult_x_1196_n2022)
         );
  XNOR2xp5_ASAP7_75t_SL U33416 ( .A(mult_x_1196_n2029), .B(n22821), .Y(n22639)
         );
  XNOR2xp5_ASAP7_75t_SL U33417 ( .A(n22641), .B(mult_x_1196_n1858), .Y(n22690)
         );
  XOR2xp5_ASAP7_75t_SL U33418 ( .A(n22640), .B(n23602), .Y(mult_x_1196_n1858)
         );
  INVx1_ASAP7_75t_SL U33419 ( .A(mult_x_1196_n1884), .Y(n22640) );
  INVx1_ASAP7_75t_SL U33420 ( .A(mult_x_1196_n1862), .Y(n22641) );
  BUFx5_ASAP7_75t_SL U33421 ( .A(n23979), .Y(n22642) );
  XOR2xp5_ASAP7_75t_SL U33422 ( .A(mult_x_1196_n1836), .B(n24306), .Y(n22643)
         );
  XOR2xp5_ASAP7_75t_SL U33423 ( .A(n22645), .B(n23460), .Y(mult_x_1196_n1708)
         );
  INVx1_ASAP7_75t_SL U33424 ( .A(mult_x_1196_n2581), .Y(n22645) );
  XNOR2x1_ASAP7_75t_SL U33425 ( .A(n23062), .B(n23063), .Y(mult_x_1196_n1610)
         );
  OAI22x1_ASAP7_75t_SL U33426 ( .A1(n24007), .A2(mult_x_1196_n3050), .B1(
        n24005), .B2(mult_x_1196_n3049), .Y(mult_x_1196_n2478) );
  XNOR2x1_ASAP7_75t_SL U33427 ( .A(n23874), .B(mult_x_1196_n2478), .Y(n23873)
         );
  NOR2x1_ASAP7_75t_SL U33428 ( .A(n24025), .B(mult_x_1196_n2902), .Y(n24202)
         );
  XNOR2xp5_ASAP7_75t_SL U33429 ( .A(n23565), .B(n22646), .Y(mult_x_1196_n1501)
         );
  INVx4_ASAP7_75t_SL U33430 ( .A(n23995), .Y(n23996) );
  INVx1_ASAP7_75t_SL U33431 ( .A(n22890), .Y(n22893) );
  NAND2xp5_ASAP7_75t_SL U33432 ( .A(n22650), .B(n22649), .Y(n22890) );
  NAND2xp5_ASAP7_75t_SL U33433 ( .A(n23262), .B(n24172), .Y(n22649) );
  XNOR2xp5_ASAP7_75t_SL U33434 ( .A(n22338), .B(mult_x_1196_n1139), .Y(n23866)
         );
  XOR2xp5_ASAP7_75t_SL U33435 ( .A(mult_x_1196_n1349), .B(n22896), .Y(n24155)
         );
  XNOR2xp5_ASAP7_75t_SL U33436 ( .A(n22794), .B(n22793), .Y(mult_x_1196_n1349)
         );
  XNOR2x1_ASAP7_75t_SL U33437 ( .A(n22831), .B(n22210), .Y(mult_x_1196_n1772)
         );
  INVx6_ASAP7_75t_SL U33438 ( .A(n24688), .Y(n24689) );
  BUFx3_ASAP7_75t_SL U33439 ( .A(n23849), .Y(n23829) );
  XNOR2x1_ASAP7_75t_SL U33440 ( .A(n22934), .B(mult_x_1196_n1471), .Y(
        mult_x_1196_n1473) );
  INVx1_ASAP7_75t_SL U33441 ( .A(mult_x_1196_n2538), .Y(n22923) );
  OAI22xp5_ASAP7_75t_SL U33442 ( .A1(mult_x_1196_n3114), .A2(n23999), .B1(
        n23997), .B2(mult_x_1196_n3113), .Y(mult_x_1196_n2538) );
  AOI21xp5_ASAP7_75t_SL U33443 ( .A1(mult_x_1196_n1103), .A2(n24251), .B(
        mult_x_1196_n1101), .Y(n22657) );
  NAND2x1_ASAP7_75t_SL U33444 ( .A(n22659), .B(n22658), .Y(n24307) );
  INVx1_ASAP7_75t_SL U33445 ( .A(mult_x_1196_n2030), .Y(n22658) );
  INVx1_ASAP7_75t_SL U33446 ( .A(mult_x_1196_n2043), .Y(n22659) );
  INVx2_ASAP7_75t_SL U33447 ( .A(n24079), .Y(n24078) );
  XNOR2x1_ASAP7_75t_SL U33448 ( .A(n22991), .B(n23132), .Y(n22901) );
  OAI22x1_ASAP7_75t_SL U33449 ( .A1(n23522), .A2(mult_x_1196_n3191), .B1(
        mult_x_1196_n3190), .B2(n23987), .Y(mult_x_1196_n2615) );
  OAI22x1_ASAP7_75t_SL U33450 ( .A1(mult_x_1196_n2924), .A2(n24022), .B1(
        mult_x_1196_n2923), .B2(n24020), .Y(mult_x_1196_n2352) );
  XNOR2x1_ASAP7_75t_SL U33451 ( .A(mult_x_1196_n1979), .B(n22960), .Y(n23567)
         );
  MAJIxp5_ASAP7_75t_SL U33452 ( .A(n22660), .B(mult_x_1196_n1005), .C(
        mult_x_1196_n987), .Y(mult_x_1196_n981) );
  MAJx2_ASAP7_75t_SL U33453 ( .A(n22789), .B(mult_x_1196_n1009), .C(
        mult_x_1196_n1002), .Y(n22660) );
  NAND2xp33_ASAP7_75t_SRAM U33454 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__20_), 
        .B(n24685), .Y(n25089) );
  XNOR2xp5_ASAP7_75t_SL U33455 ( .A(mult_x_1196_n2128), .B(n22661), .Y(
        mult_x_1196_n1566) );
  XOR2xp5_ASAP7_75t_SL U33456 ( .A(mult_x_1196_n2357), .B(mult_x_1196_n2453), 
        .Y(n22661) );
  NOR2x1_ASAP7_75t_SL U33457 ( .A(n23257), .B(n23256), .Y(mult_x_1196_n2059)
         );
  OAI21x1_ASAP7_75t_SL U33458 ( .A1(mult_x_1196_n3049), .A2(n18561), .B(n22276), .Y(n23680) );
  MAJIxp5_ASAP7_75t_SL U33459 ( .A(n22662), .B(mult_x_1196_n1811), .C(n18936), 
        .Y(n23860) );
  INVx1_ASAP7_75t_SL U33460 ( .A(mult_x_1196_n1833), .Y(n22662) );
  MAJIxp5_ASAP7_75t_SL U33461 ( .A(n23591), .B(mult_x_1196_n1832), .C(n22484), 
        .Y(mult_x_1196_n1833) );
  NOR2x1p5_ASAP7_75t_SL U33462 ( .A(n23152), .B(n23151), .Y(mult_x_1196_n1255)
         );
  INVx8_ASAP7_75t_SL U33463 ( .A(n24004), .Y(n24005) );
  BUFx2_ASAP7_75t_SL U33464 ( .A(n24027), .Y(n23708) );
  OAI22x1_ASAP7_75t_SL U33465 ( .A1(n18837), .A2(n25815), .B1(n23559), .B2(
        n23844), .Y(u0_0_leon3x0_p0_muli[26]) );
  INVx1_ASAP7_75t_SL U33466 ( .A(mult_x_1196_n2238), .Y(n22665) );
  XNOR2xp5_ASAP7_75t_SL U33467 ( .A(mult_x_1196_n1630), .B(mult_x_1196_n1599), 
        .Y(n22666) );
  MAJIxp5_ASAP7_75t_SL U33468 ( .A(mult_x_1196_n1011), .B(mult_x_1196_n1032), 
        .C(mult_x_1196_n1013), .Y(mult_x_1196_n1005) );
  XNOR2xp5_ASAP7_75t_SL U33469 ( .A(mult_x_1196_n1011), .B(n22667), .Y(
        mult_x_1196_n1006) );
  XOR2xp5_ASAP7_75t_SL U33470 ( .A(mult_x_1196_n1032), .B(mult_x_1196_n1013), 
        .Y(n22667) );
  XNOR2x1_ASAP7_75t_SL U33471 ( .A(mult_x_1196_n1460), .B(mult_x_1196_n1455), 
        .Y(n23783) );
  MAJIxp5_ASAP7_75t_SL U33472 ( .A(n22669), .B(mult_x_1196_n1633), .C(
        mult_x_1196_n1659), .Y(mult_x_1196_n1624) );
  XNOR2xp5_ASAP7_75t_SL U33473 ( .A(mult_x_1196_n1659), .B(n22670), .Y(
        mult_x_1196_n1625) );
  XNOR2xp5_ASAP7_75t_SL U33474 ( .A(n22671), .B(mult_x_1196_n1633), .Y(n22670)
         );
  INVx8_ASAP7_75t_SL U33475 ( .A(n23639), .Y(n24076) );
  XNOR2xp5_ASAP7_75t_SL U33476 ( .A(n23373), .B(n23104), .Y(mult_x_1196_n1866)
         );
  MAJIxp5_ASAP7_75t_SL U33477 ( .A(mult_x_1196_n994), .B(mult_x_1196_n990), 
        .C(n22672), .Y(mult_x_1196_n984) );
  INVx1_ASAP7_75t_SL U33478 ( .A(n22674), .Y(n22672) );
  XOR2xp5_ASAP7_75t_SL U33479 ( .A(n22674), .B(mult_x_1196_n990), .Y(n22673)
         );
  MAJIxp5_ASAP7_75t_SL U33480 ( .A(n22988), .B(n24253), .C(mult_x_1196_n1028), 
        .Y(n22674) );
  INVx1_ASAP7_75t_SL U33481 ( .A(mult_x_1196_n994), .Y(n22675) );
  MAJx2_ASAP7_75t_SL U33482 ( .A(mult_x_1196_n882), .B(mult_x_1196_n878), .C(
        mult_x_1196_n893), .Y(mult_x_1196_n867) );
  MAJIxp5_ASAP7_75t_SL U33483 ( .A(mult_x_1196_n1975), .B(mult_x_1196_n1954), 
        .C(mult_x_1196_n1961), .Y(mult_x_1196_n1955) );
  INVx1_ASAP7_75t_SL U33484 ( .A(mult_x_1196_n1954), .Y(n22677) );
  HB1xp67_ASAP7_75t_SL U33485 ( .A(n23123), .Y(n22678) );
  INVx8_ASAP7_75t_SL U33486 ( .A(n23959), .Y(n23960) );
  INVx1_ASAP7_75t_SL U33487 ( .A(mult_x_1196_n2013), .Y(n22680) );
  NAND2xp5_ASAP7_75t_SL U33488 ( .A(n23125), .B(n23288), .Y(n24235) );
  XOR2xp5_ASAP7_75t_SL U33489 ( .A(n22681), .B(mult_x_1196_n2182), .Y(
        mult_x_1196_n915) );
  XNOR2xp5_ASAP7_75t_SL U33490 ( .A(n22682), .B(mult_x_1196_n929), .Y(n22681)
         );
  OAI22xp5_ASAP7_75t_SL U33491 ( .A1(mult_x_1196_n2809), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2808), .Y(n22682) );
  MAJIxp5_ASAP7_75t_SL U33492 ( .A(mult_x_1196_n2229), .B(mult_x_1196_n2447), 
        .C(mult_x_1196_n2351), .Y(mult_x_1196_n1346) );
  XOR2xp5_ASAP7_75t_SL U33493 ( .A(n22684), .B(mult_x_1196_n1353), .Y(n22683)
         );
  XNOR2xp5_ASAP7_75t_SL U33494 ( .A(mult_x_1196_n2351), .B(n22685), .Y(n22684)
         );
  XOR2xp5_ASAP7_75t_SL U33495 ( .A(mult_x_1196_n2229), .B(mult_x_1196_n2447), 
        .Y(n22685) );
  MAJIxp5_ASAP7_75t_SL U33496 ( .A(n22687), .B(mult_x_1196_n1552), .C(
        mult_x_1196_n1593), .Y(mult_x_1196_n1553) );
  XOR2xp5_ASAP7_75t_SL U33497 ( .A(mult_x_1196_n1593), .B(n22686), .Y(
        mult_x_1196_n1554) );
  XNOR2xp5_ASAP7_75t_SL U33498 ( .A(mult_x_1196_n1552), .B(n22687), .Y(n22686)
         );
  XNOR2xp5_ASAP7_75t_SL U33499 ( .A(n23349), .B(n23348), .Y(n22687) );
  XOR2xp5_ASAP7_75t_SL U33500 ( .A(mult_x_1196_n1606), .B(mult_x_1196_n1602), 
        .Y(n22689) );
  BUFx6f_ASAP7_75t_SL U33501 ( .A(n24018), .Y(n23142) );
  OAI22x1_ASAP7_75t_SL U33502 ( .A1(n23522), .A2(mult_x_1196_n3183), .B1(
        mult_x_1196_n3182), .B2(n24106), .Y(mult_x_1196_n2607) );
  OR2x2_ASAP7_75t_SL U33503 ( .A(mult_x_1196_n393), .B(n23475), .Y(
        mult_x_1196_n387) );
  INVx1_ASAP7_75t_SL U33504 ( .A(mult_x_1196_n489), .Y(mult_x_1196_n491) );
  INVx8_ASAP7_75t_SL U33505 ( .A(n24151), .Y(n23992) );
  INVx4_ASAP7_75t_SL U33506 ( .A(n23704), .Y(n23116) );
  MAJx2_ASAP7_75t_SL U33507 ( .A(n23912), .B(n23814), .C(mult_x_1196_n2232), 
        .Y(n23419) );
  XNOR2x1_ASAP7_75t_SL U33508 ( .A(n23753), .B(n18396), .Y(n23752) );
  XOR2xp5_ASAP7_75t_SL U33509 ( .A(mult_x_1196_n1251), .B(mult_x_1196_n1247), 
        .Y(n24103) );
  MAJIxp5_ASAP7_75t_SL U33510 ( .A(n24288), .B(mult_x_1196_n1559), .C(
        mult_x_1196_n1557), .Y(mult_x_1196_n1548) );
  INVx1_ASAP7_75t_SL U33511 ( .A(mult_x_1196_n2069), .Y(n22691) );
  XNOR2xp5_ASAP7_75t_SL U33512 ( .A(n22692), .B(mult_x_1196_n2257), .Y(
        mult_x_1196_n1223) );
  XNOR2xp5_ASAP7_75t_SL U33513 ( .A(mult_x_1196_n2196), .B(mult_x_1196_n1255), 
        .Y(n22692) );
  BUFx2_ASAP7_75t_SL U33514 ( .A(n24089), .Y(n22693) );
  INVx1_ASAP7_75t_SL U33515 ( .A(mult_x_1196_n2138), .Y(n22860) );
  OAI21x1_ASAP7_75t_SL U33516 ( .A1(n18435), .A2(mult_x_1196_n3110), .B(n22695), .Y(mult_x_1196_n2138) );
  INVx1_ASAP7_75t_SL U33517 ( .A(n22696), .Y(n22695) );
  XNOR2x1_ASAP7_75t_SL U33518 ( .A(n22828), .B(n22208), .Y(mult_x_1196_n1648)
         );
  MAJIxp5_ASAP7_75t_SL U33519 ( .A(n24296), .B(mult_x_1196_n2055), .C(
        mult_x_1196_n2051), .Y(mult_x_1196_n2043) );
  NAND2xp5_ASAP7_75t_SL U33520 ( .A(mult_x_1196_n2044), .B(mult_x_1196_n2052), 
        .Y(mult_x_1196_n728) );
  XOR2xp5_ASAP7_75t_SL U33521 ( .A(mult_x_1196_n2051), .B(mult_x_1196_n2055), 
        .Y(n22699) );
  XNOR2xp5_ASAP7_75t_SL U33522 ( .A(n22700), .B(n18538), .Y(mult_x_1196_n1811)
         );
  XOR2xp5_ASAP7_75t_SL U33523 ( .A(mult_x_1196_n2132), .B(mult_x_1196_n2365), 
        .Y(n22700) );
  MAJIxp5_ASAP7_75t_SL U33524 ( .A(mult_x_1196_n1819), .B(mult_x_1196_n2365), 
        .C(mult_x_1196_n2132), .Y(mult_x_1196_n1810) );
  BUFx2_ASAP7_75t_SL U33525 ( .A(n23449), .Y(n22780) );
  MAJIxp5_ASAP7_75t_SL U33526 ( .A(mult_x_1196_n896), .B(mult_x_1196_n898), 
        .C(mult_x_1196_n886), .Y(mult_x_1196_n881) );
  XOR2xp5_ASAP7_75t_SL U33527 ( .A(n22702), .B(n22701), .Y(mult_x_1196_n882)
         );
  INVx1_ASAP7_75t_SL U33528 ( .A(mult_x_1196_n896), .Y(n22702) );
  INVx1_ASAP7_75t_SL U33529 ( .A(n22974), .Y(n22704) );
  BUFx3_ASAP7_75t_SL U33530 ( .A(n24024), .Y(n22983) );
  OAI22x1_ASAP7_75t_SL U33531 ( .A1(mult_x_1196_n3095), .A2(n23100), .B1(
        n24002), .B2(mult_x_1196_n3094), .Y(mult_x_1196_n2519) );
  NOR2x1p5_ASAP7_75t_SL U33532 ( .A(n22226), .B(n23587), .Y(n23588) );
  OAI22xp5_ASAP7_75t_SL U33533 ( .A1(mult_x_1196_n2952), .A2(n24017), .B1(
        mult_x_1196_n2953), .B2(n23141), .Y(mult_x_1196_n2381) );
  OAI22xp5_ASAP7_75t_SL U33534 ( .A1(mult_x_1196_n2959), .A2(n24017), .B1(
        mult_x_1196_n2960), .B2(n23141), .Y(mult_x_1196_n2388) );
  MAJIxp5_ASAP7_75t_SL U33535 ( .A(mult_x_1196_n2663), .B(n23402), .C(
        mult_x_1196_n2599), .Y(mult_x_1196_n2057) );
  XNOR2xp5_ASAP7_75t_SL U33536 ( .A(n23298), .B(n22707), .Y(n23035) );
  XOR2xp5_ASAP7_75t_SL U33537 ( .A(mult_x_1196_n1442), .B(mult_x_1196_n1439), 
        .Y(n22707) );
  MAJIxp5_ASAP7_75t_SL U33538 ( .A(mult_x_1196_n2422), .B(n22708), .C(
        mult_x_1196_n2578), .Y(mult_x_1196_n1605) );
  OAI22xp5_ASAP7_75t_SL U33539 ( .A1(n23637), .A2(mult_x_1196_n3058), .B1(
        n24005), .B2(mult_x_1196_n3057), .Y(n22708) );
  OAI22x1_ASAP7_75t_SL U33540 ( .A1(mult_x_1196_n3205), .A2(n23072), .B1(
        mult_x_1196_n3204), .B2(n23987), .Y(mult_x_1196_n2629) );
  OAI22x1_ASAP7_75t_SL U33541 ( .A1(mult_x_1196_n3091), .A2(n24002), .B1(
        n23100), .B2(mult_x_1196_n3092), .Y(mult_x_1196_n2516) );
  MAJx2_ASAP7_75t_SL U33542 ( .A(mult_x_1196_n1336), .B(mult_x_1196_n1344), 
        .C(n22311), .Y(mult_x_1196_n1264) );
  MAJIxp5_ASAP7_75t_SL U33543 ( .A(mult_x_1196_n2608), .B(mult_x_1196_n2544), 
        .C(mult_x_1196_n2173), .Y(mult_x_1196_n1534) );
  XNOR2xp5_ASAP7_75t_SL U33544 ( .A(n23305), .B(n22719), .Y(n23304) );
  INVx1_ASAP7_75t_SL U33545 ( .A(mult_x_1196_n1748), .Y(n23343) );
  INVx1_ASAP7_75t_SL U33546 ( .A(n23917), .Y(n22710) );
  OAI22xp5_ASAP7_75t_SL U33547 ( .A1(mult_x_1196_n2756), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2755), .Y(n23286) );
  XOR2xp5_ASAP7_75t_SL U33548 ( .A(n22711), .B(mult_x_1196_n2354), .Y(n22851)
         );
  INVx1_ASAP7_75t_SL U33549 ( .A(mult_x_1196_n2171), .Y(n22711) );
  NAND2x2_ASAP7_75t_SL U33550 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__24_), .B(
        n22986), .Y(n23741) );
  XNOR2xp5_ASAP7_75t_SL U33551 ( .A(n22713), .B(n22712), .Y(mult_x_1196_n1557)
         );
  XNOR2xp5_ASAP7_75t_SL U33552 ( .A(mult_x_1196_n1572), .B(mult_x_1196_n1570), 
        .Y(n22712) );
  INVx1_ASAP7_75t_SL U33553 ( .A(n24284), .Y(n22713) );
  INVx2_ASAP7_75t_SL U33554 ( .A(mult_x_1196_n2172), .Y(n22714) );
  XOR2xp5_ASAP7_75t_SL U33555 ( .A(mult_x_1196_n2576), .B(n24212), .Y(n24213)
         );
  XOR2x2_ASAP7_75t_SL U33556 ( .A(mult_x_1196_n1619), .B(mult_x_1196_n1579), 
        .Y(n23092) );
  XOR2x2_ASAP7_75t_SL U33557 ( .A(mult_x_1196_n1624), .B(n22857), .Y(
        mult_x_1196_n1579) );
  MAJIxp5_ASAP7_75t_SL U33558 ( .A(n23525), .B(n22343), .C(mult_x_1196_n1625), 
        .Y(mult_x_1196_n1619) );
  NOR2x1_ASAP7_75t_SL U33559 ( .A(mult_x_1196_n1931), .B(mult_x_1196_n1911), 
        .Y(mult_x_1196_n683) );
  NAND2xp5_ASAP7_75t_SL U33560 ( .A(n24032), .B(n22716), .Y(n22715) );
  XOR2xp5_ASAP7_75t_SL U33561 ( .A(n23726), .B(n22846), .Y(mult_x_1196_n1660)
         );
  NAND2x1p5_ASAP7_75t_SL U33562 ( .A(mult_x_1196_n2513), .B(mult_x_1196_n2673), 
        .Y(n23071) );
  INVx2_ASAP7_75t_SL U33563 ( .A(n23071), .Y(n23069) );
  MAJx2_ASAP7_75t_SL U33564 ( .A(mult_x_1196_n1496), .B(n23411), .C(n22514), 
        .Y(mult_x_1196_n1406) );
  BUFx6f_ASAP7_75t_SL U33565 ( .A(n24687), .Y(n22986) );
  MAJIxp5_ASAP7_75t_SL U33566 ( .A(n22271), .B(mult_x_1196_n2537), .C(n23680), 
        .Y(mult_x_1196_n1283) );
  OAI21xp5_ASAP7_75t_SL U33567 ( .A1(n23999), .A2(mult_x_1196_n3113), .B(
        n22717), .Y(mult_x_1196_n2537) );
  NAND2xp5_ASAP7_75t_SL U33568 ( .A(n23995), .B(n22718), .Y(n22717) );
  AOI21x1_ASAP7_75t_SL U33569 ( .A1(mult_x_1196_n391), .A2(mult_x_1196_n425), 
        .B(mult_x_1196_n392), .Y(mult_x_1196_n390) );
  OAI22x1_ASAP7_75t_SL U33570 ( .A1(mult_x_1196_n3251), .A2(n23981), .B1(
        n22389), .B2(mult_x_1196_n3250), .Y(mult_x_1196_n2675) );
  INVx1_ASAP7_75t_SL U33571 ( .A(mult_x_1196_n1609), .Y(n24105) );
  XNOR2xp5_ASAP7_75t_SL U33572 ( .A(n24255), .B(mult_x_1196_n1528), .Y(n22719)
         );
  XNOR2xp5_ASAP7_75t_SL U33573 ( .A(mult_x_1196_n1454), .B(n23748), .Y(n23272)
         );
  XNOR2x1_ASAP7_75t_SL U33574 ( .A(n23434), .B(mult_x_1196_n2392), .Y(n23433)
         );
  XNOR2x1_ASAP7_75t_SL U33575 ( .A(n23433), .B(n23432), .Y(mult_x_1196_n1670)
         );
  BUFx10_ASAP7_75t_SL U33576 ( .A(u0_0_leon3x0_p0_muli[32]), .Y(n24052) );
  MAJIxp5_ASAP7_75t_SL U33577 ( .A(n24179), .B(mult_x_1196_n2163), .C(
        mult_x_1196_n2378), .Y(n23174) );
  OAI22xp5_ASAP7_75t_SL U33578 ( .A1(mult_x_1196_n2950), .A2(n23141), .B1(
        n22694), .B2(mult_x_1196_n2949), .Y(mult_x_1196_n2378) );
  XNOR2xp5_ASAP7_75t_SL U33579 ( .A(n24278), .B(mult_x_1196_n1750), .Y(n23398)
         );
  INVx1_ASAP7_75t_SL U33580 ( .A(n23326), .Y(n22722) );
  XNOR2xp5_ASAP7_75t_SL U33581 ( .A(n23127), .B(n23321), .Y(n23720) );
  OAI21x1_ASAP7_75t_SL U33582 ( .A1(n28623), .A2(n23830), .B(n28622), .Y(
        u0_0_leon3x0_p0_muli[22]) );
  OAI21x1_ASAP7_75t_SL U33583 ( .A1(mult_x_1196_n2831), .A2(n24034), .B(n22309), .Y(n24180) );
  NAND2xp5_ASAP7_75t_SL U33584 ( .A(mult_x_1196_n1472), .B(mult_x_1196_n1434), 
        .Y(n22724) );
  NOR2xp33_ASAP7_75t_SL U33585 ( .A(mult_x_1196_n1434), .B(mult_x_1196_n1472), 
        .Y(n22726) );
  NAND2x1_ASAP7_75t_SL U33586 ( .A(mult_x_1196_n3323), .B(n23444), .Y(
        mult_x_1196_n72) );
  BUFx5_ASAP7_75t_SL U33587 ( .A(add_x_735_A_12_), .Y(n23091) );
  OAI22x1_ASAP7_75t_SL U33588 ( .A1(mult_x_1196_n3151), .A2(n23992), .B1(
        n24230), .B2(mult_x_1196_n3152), .Y(mult_x_1196_n2576) );
  XOR2xp5_ASAP7_75t_SL U33589 ( .A(n23000), .B(n22571), .Y(mult_x_1196_n1542)
         );
  XNOR2xp5_ASAP7_75t_SL U33590 ( .A(n22727), .B(mult_x_1196_n1730), .Y(n22803)
         );
  INVx1_ASAP7_75t_SL U33591 ( .A(mult_x_1196_n1732), .Y(n22727) );
  OAI21x1_ASAP7_75t_SL U33592 ( .A1(mult_x_1196_n613), .A2(mult_x_1196_n617), 
        .B(mult_x_1196_n614), .Y(mult_x_1196_n612) );
  MAJIxp5_ASAP7_75t_SL U33593 ( .A(mult_x_1196_n2607), .B(mult_x_1196_n2127), 
        .C(n23565), .Y(mult_x_1196_n1500) );
  MAJx2_ASAP7_75t_SL U33594 ( .A(mult_x_1196_n1904), .B(n23501), .C(
        mult_x_1196_n1906), .Y(mult_x_1196_n1872) );
  INVx1_ASAP7_75t_SL U33595 ( .A(n23482), .Y(n23483) );
  INVx1_ASAP7_75t_SL U33596 ( .A(mult_x_1196_n904), .Y(mult_x_1196_n888) );
  MAJIxp5_ASAP7_75t_SL U33597 ( .A(n22729), .B(mult_x_1196_n1965), .C(
        mult_x_1196_n1963), .Y(mult_x_1196_n1957) );
  MAJIxp5_ASAP7_75t_SL U33598 ( .A(n24283), .B(mult_x_1196_n1985), .C(n18304), 
        .Y(n22729) );
  XNOR2xp5_ASAP7_75t_SL U33599 ( .A(n23866), .B(mult_x_1196_n1112), .Y(
        mult_x_1196_n1105) );
  OAI22x1_ASAP7_75t_SL U33600 ( .A1(n24080), .A2(mult_x_1196_n3215), .B1(
        mult_x_1196_n3214), .B2(n23984), .Y(n23565) );
  MAJIxp5_ASAP7_75t_SL U33601 ( .A(mult_x_1196_n2650), .B(mult_x_1196_n2334), 
        .C(n22730), .Y(mult_x_1196_n1839) );
  INVx1_ASAP7_75t_SL U33602 ( .A(n22732), .Y(n22730) );
  HB1xp67_ASAP7_75t_SL U33603 ( .A(n23816), .Y(n22735) );
  AND2x2_ASAP7_75t_SL U33604 ( .A(add_x_735_A_12_), .B(n23747), .Y(n22965) );
  OAI22xp5_ASAP7_75t_SL U33605 ( .A1(mult_x_1196_n2956), .A2(n24017), .B1(
        mult_x_1196_n2957), .B2(n23142), .Y(mult_x_1196_n2385) );
  XNOR2xp5_ASAP7_75t_SL U33606 ( .A(mult_x_1196_n1312), .B(n22798), .Y(n22736)
         );
  XNOR2x1_ASAP7_75t_SL U33607 ( .A(n22980), .B(n22982), .Y(mult_x_1196_n1604)
         );
  NOR2x2_ASAP7_75t_SL U33608 ( .A(mult_x_1196_n2999), .B(n23311), .Y(n23879)
         );
  INVx8_ASAP7_75t_SL U33609 ( .A(n24076), .Y(n23658) );
  BUFx5_ASAP7_75t_SL U33610 ( .A(mult_x_1196_n39), .Y(add_x_735_A_10_) );
  XNOR2xp5_ASAP7_75t_SL U33611 ( .A(n22895), .B(n22737), .Y(mult_x_1196_n1650)
         );
  XNOR2xp5_ASAP7_75t_SL U33612 ( .A(n22738), .B(mult_x_1196_n1660), .Y(n22737)
         );
  INVx1_ASAP7_75t_SL U33613 ( .A(mult_x_1196_n1694), .Y(n22738) );
  BUFx2_ASAP7_75t_SL U33614 ( .A(n23142), .Y(n22779) );
  INVx2_ASAP7_75t_SL U33615 ( .A(add_x_735_A_20_), .Y(n23936) );
  INVx1_ASAP7_75t_SL U33616 ( .A(n23956), .Y(n23958) );
  OAI22x1_ASAP7_75t_SL U33617 ( .A1(mult_x_1196_n3186), .A2(n23072), .B1(
        mult_x_1196_n3185), .B2(n23987), .Y(n23330) );
  MAJIxp5_ASAP7_75t_SL U33618 ( .A(mult_x_1196_n967), .B(mult_x_1196_n955), 
        .C(mult_x_1196_n969), .Y(mult_x_1196_n949) );
  MAJIxp5_ASAP7_75t_SL U33619 ( .A(n22741), .B(mult_x_1196_n946), .C(
        mult_x_1196_n965), .Y(mult_x_1196_n947) );
  XNOR2xp5_ASAP7_75t_SL U33620 ( .A(mult_x_1196_n965), .B(n22740), .Y(
        mult_x_1196_n948) );
  XOR2xp5_ASAP7_75t_SL U33621 ( .A(mult_x_1196_n946), .B(n22741), .Y(n22740)
         );
  XNOR2xp5_ASAP7_75t_SL U33622 ( .A(mult_x_1196_n967), .B(n22742), .Y(n22741)
         );
  XOR2xp5_ASAP7_75t_SL U33623 ( .A(mult_x_1196_n969), .B(mult_x_1196_n955), 
        .Y(n22742) );
  MAJIxp5_ASAP7_75t_SL U33624 ( .A(mult_x_1196_n2619), .B(mult_x_1196_n2495), 
        .C(mult_x_1196_n2651), .Y(mult_x_1196_n1863) );
  OAI21xp5_ASAP7_75t_SL U33625 ( .A1(mult_x_1196_n3004), .A2(n24014), .B(
        n22305), .Y(n23760) );
  MAJIxp5_ASAP7_75t_SL U33626 ( .A(n22208), .B(n22745), .C(n22744), .Y(
        mult_x_1196_n1614) );
  INVx1_ASAP7_75t_SL U33627 ( .A(n18354), .Y(n22745) );
  XNOR2x1_ASAP7_75t_SL U33628 ( .A(n24216), .B(n22746), .Y(mult_x_1196_n1460)
         );
  INVx2_ASAP7_75t_SL U33629 ( .A(n24215), .Y(n22746) );
  XOR2x2_ASAP7_75t_SL U33630 ( .A(n22851), .B(mult_x_1196_n2386), .Y(
        mult_x_1196_n1455) );
  XNOR2xp5_ASAP7_75t_SL U33631 ( .A(n22747), .B(n23822), .Y(n23820) );
  OAI22xp5_ASAP7_75t_SL U33632 ( .A1(mult_x_1196_n2996), .A2(n24012), .B1(
        mult_x_1196_n2997), .B2(n23311), .Y(n23822) );
  INVx1_ASAP7_75t_SL U33633 ( .A(mult_x_1196_n2393), .Y(n22747) );
  INVx2_ASAP7_75t_SL U33634 ( .A(mult_x_1196_n3329), .Y(n24232) );
  MAJx2_ASAP7_75t_SL U33635 ( .A(mult_x_1196_n1837), .B(mult_x_1196_n1835), 
        .C(n23049), .Y(mult_x_1196_n1780) );
  NOR2x1_ASAP7_75t_SL U33636 ( .A(n23984), .B(mult_x_1196_n3232), .Y(n22748)
         );
  XNOR2x2_ASAP7_75t_SL U33637 ( .A(mult_x_1196_n2361), .B(n23679), .Y(n23678)
         );
  XOR2xp5_ASAP7_75t_SL U33638 ( .A(mult_x_1196_n1787), .B(n22869), .Y(n24077)
         );
  INVx1_ASAP7_75t_SL U33639 ( .A(mult_x_1196_n3150), .Y(n24165) );
  XNOR2xp5_ASAP7_75t_SL U33640 ( .A(n22750), .B(n22749), .Y(mult_x_1196_n1719)
         );
  XOR2xp5_ASAP7_75t_SL U33641 ( .A(mult_x_1196_n1749), .B(n22213), .Y(n22749)
         );
  BUFx2_ASAP7_75t_SL U33642 ( .A(n24268), .Y(n22751) );
  HB1xp67_ASAP7_75t_SL U33643 ( .A(mult_x_1196_n549), .Y(n22752) );
  XOR2xp5_ASAP7_75t_SL U33644 ( .A(n22372), .B(mult_x_1196_n1061), .Y(n22753)
         );
  OAI21x1_ASAP7_75t_SL U33645 ( .A1(mult_x_1196_n696), .A2(mult_x_1196_n708), 
        .B(mult_x_1196_n697), .Y(mult_x_1196_n695) );
  AOI21x1_ASAP7_75t_SL U33646 ( .A1(mult_x_1196_n695), .A2(mult_x_1196_n687), 
        .B(mult_x_1196_n688), .Y(n23454) );
  BUFx2_ASAP7_75t_SL U33647 ( .A(mult_x_1196_n1721), .Y(n22827) );
  INVx1_ASAP7_75t_SL U33648 ( .A(n22755), .Y(n22754) );
  MAJIxp5_ASAP7_75t_SL U33649 ( .A(n22755), .B(mult_x_1196_n1565), .C(
        mult_x_1196_n1567), .Y(mult_x_1196_n1526) );
  MAJIxp5_ASAP7_75t_SL U33650 ( .A(n22872), .B(mult_x_1196_n2325), .C(
        mult_x_1196_n2206), .Y(n22755) );
  INVx2_ASAP7_75t_SL U33651 ( .A(n22897), .Y(n24691) );
  INVx1_ASAP7_75t_SL U33652 ( .A(mult_x_1196_n2584), .Y(n22757) );
  NOR2x1_ASAP7_75t_SL U33653 ( .A(mult_x_1196_n546), .B(mult_x_1196_n539), .Y(
        mult_x_1196_n533) );
  XNOR2xp5_ASAP7_75t_SL U33654 ( .A(n22759), .B(n23526), .Y(n23541) );
  MAJx2_ASAP7_75t_SL U33655 ( .A(n23691), .B(mult_x_1196_n1737), .C(
        mult_x_1196_n1733), .Y(mult_x_1196_n1661) );
  BUFx3_ASAP7_75t_SL U33656 ( .A(n24028), .Y(n22962) );
  XNOR2x1_ASAP7_75t_SL U33657 ( .A(n23525), .B(n22343), .Y(n23524) );
  XNOR2x1_ASAP7_75t_SL U33658 ( .A(n23524), .B(n23528), .Y(mult_x_1196_n1620)
         );
  NOR2x1_ASAP7_75t_SL U33659 ( .A(n23040), .B(n24285), .Y(mult_x_1196_n539) );
  INVx1_ASAP7_75t_SL U33660 ( .A(mult_x_1196_n1260), .Y(n23040) );
  MAJIxp5_ASAP7_75t_SL U33661 ( .A(mult_x_1196_n2246), .B(n22763), .C(
        mult_x_1196_n2336), .Y(mult_x_1196_n958) );
  XOR2xp5_ASAP7_75t_SL U33662 ( .A(n22763), .B(mult_x_1196_n2336), .Y(n22762)
         );
  OAI22xp5_ASAP7_75t_SL U33663 ( .A1(mult_x_1196_n2780), .A2(n22412), .B1(
        mult_x_1196_n2779), .B2(n22391), .Y(n22763) );
  NAND2xp5_ASAP7_75t_SL U33664 ( .A(mult_x_1196_n1922), .B(n22765), .Y(n22764)
         );
  INVx1_ASAP7_75t_SL U33665 ( .A(mult_x_1196_n1937), .Y(n22765) );
  OAI21xp5_ASAP7_75t_SL U33666 ( .A1(n23831), .A2(n28523), .B(n27056), .Y(
        u0_0_leon3x0_p0_muli[29]) );
  XNOR2xp5_ASAP7_75t_SL U33667 ( .A(n24692), .B(n23707), .Y(n23706) );
  OAI22x1_ASAP7_75t_SL U33668 ( .A1(mult_x_1196_n2898), .A2(n22983), .B1(
        mult_x_1196_n2899), .B2(n23116), .Y(mult_x_1196_n2327) );
  XOR2xp5_ASAP7_75t_SL U33669 ( .A(mult_x_1196_n1125), .B(mult_x_1196_n1131), 
        .Y(n22766) );
  MAJIxp5_ASAP7_75t_SL U33670 ( .A(n22768), .B(mult_x_1196_n1119), .C(
        mult_x_1196_n1096), .Y(mult_x_1196_n1088) );
  XNOR2xp5_ASAP7_75t_SL U33671 ( .A(mult_x_1196_n1119), .B(n22767), .Y(
        mult_x_1196_n1089) );
  MAJIxp5_ASAP7_75t_SL U33672 ( .A(n22314), .B(mult_x_1196_n1125), .C(
        mult_x_1196_n1131), .Y(n22768) );
  OR2x2_ASAP7_75t_SL U33673 ( .A(n24232), .B(n23983), .Y(n24082) );
  MAJIxp5_ASAP7_75t_SL U33674 ( .A(mult_x_1196_n1383), .B(n23523), .C(
        mult_x_1196_n1381), .Y(mult_x_1196_n1344) );
  XNOR2xp5_ASAP7_75t_SL U33675 ( .A(n22770), .B(mult_x_1196_n1381), .Y(n22769)
         );
  INVx1_ASAP7_75t_SL U33676 ( .A(n23523), .Y(n22770) );
  OAI21xp5_ASAP7_75t_SL U33677 ( .A1(n23318), .A2(mult_x_1196_n1487), .B(
        n22771), .Y(n23320) );
  NOR2x1p5_ASAP7_75t_SL U33678 ( .A(n23871), .B(n23872), .Y(n23870) );
  MAJIxp5_ASAP7_75t_SL U33679 ( .A(mult_x_1196_n1198), .B(n22346), .C(n18989), 
        .Y(mult_x_1196_n1194) );
  XOR2xp5_ASAP7_75t_SL U33680 ( .A(n23323), .B(n23325), .Y(mult_x_1196_n2018)
         );
  OAI21xp5_ASAP7_75t_SL U33681 ( .A1(n22377), .A2(n22776), .B(n25310), .Y(
        n4199) );
  XOR2xp5_ASAP7_75t_SL U33682 ( .A(n22223), .B(n23763), .Y(n22776) );
  XOR2xp5_ASAP7_75t_SL U33683 ( .A(mult_x_1196_n2493), .B(n23156), .Y(n22777)
         );
  MAJIxp5_ASAP7_75t_SL U33684 ( .A(mult_x_1196_n2646), .B(mult_x_1196_n2272), 
        .C(mult_x_1196_n2330), .Y(mult_x_1196_n1739) );
  XNOR2xp5_ASAP7_75t_SL U33685 ( .A(mult_x_1196_n2330), .B(mult_x_1196_n2272), 
        .Y(n22778) );
  MAJIxp5_ASAP7_75t_SL U33686 ( .A(mult_x_1196_n1639), .B(mult_x_1196_n1643), 
        .C(mult_x_1196_n1629), .Y(mult_x_1196_n1630) );
  INVx1_ASAP7_75t_SL U33687 ( .A(n22784), .Y(n22782) );
  XNOR2xp5_ASAP7_75t_SL U33688 ( .A(mult_x_1196_n1662), .B(n22784), .Y(n22783)
         );
  XOR2xp5_ASAP7_75t_SL U33689 ( .A(mult_x_1196_n1629), .B(n22785), .Y(n22784)
         );
  XNOR2xp5_ASAP7_75t_SL U33690 ( .A(mult_x_1196_n1245), .B(mult_x_1196_n1273), 
        .Y(n22786) );
  INVx1_ASAP7_75t_SL U33691 ( .A(mult_x_1196_n1242), .Y(n22787) );
  OAI22x1_ASAP7_75t_SL U33692 ( .A1(mult_x_1196_n2891), .A2(n24026), .B1(
        mult_x_1196_n2890), .B2(n22983), .Y(mult_x_1196_n2319) );
  MAJx2_ASAP7_75t_SL U33693 ( .A(n23039), .B(mult_x_1196_n1994), .C(
        mult_x_1196_n2005), .Y(mult_x_1196_n1969) );
  XNOR2xp5_ASAP7_75t_SL U33694 ( .A(mult_x_1196_n1009), .B(n22788), .Y(
        mult_x_1196_n1004) );
  XNOR2xp5_ASAP7_75t_SL U33695 ( .A(mult_x_1196_n1015), .B(n22789), .Y(n22788)
         );
  MAJIxp5_ASAP7_75t_SL U33696 ( .A(n23284), .B(mult_x_1196_n1054), .C(
        mult_x_1196_n1052), .Y(n22789) );
  INVx1_ASAP7_75t_SL U33697 ( .A(mult_x_1196_n2467), .Y(n22790) );
  INVx3_ASAP7_75t_SL U33698 ( .A(mult_x_1196_n96), .Y(n24019) );
  OAI21xp5_ASAP7_75t_SL U33699 ( .A1(n24196), .A2(mult_x_1196_n748), .B(n24198), .Y(mult_x_1196_n735) );
  INVx2_ASAP7_75t_SL U33700 ( .A(mult_x_1196_n1670), .Y(n23527) );
  XNOR2x1_ASAP7_75t_SL U33701 ( .A(mult_x_1196_n2418), .B(mult_x_1196_n2574), 
        .Y(n24216) );
  OR3x1_ASAP7_75t_SL U33702 ( .A(n23496), .B(mult_x_1196_n393), .C(n22404), 
        .Y(n23575) );
  INVx1_ASAP7_75t_SL U33703 ( .A(n24189), .Y(n24245) );
  BUFx3_ASAP7_75t_SL U33704 ( .A(n23993), .Y(n24230) );
  XOR2xp5_ASAP7_75t_SL U33705 ( .A(mult_x_1196_n2383), .B(mult_x_1196_n2539), 
        .Y(n22793) );
  MAJIxp5_ASAP7_75t_SL U33706 ( .A(mult_x_1196_n2151), .B(mult_x_1196_n2183), 
        .C(n22795), .Y(mult_x_1196_n925) );
  XOR2xp5_ASAP7_75t_SL U33707 ( .A(n22797), .B(n22796), .Y(mult_x_1196_n926)
         );
  XNOR2xp5_ASAP7_75t_SL U33708 ( .A(mult_x_1196_n929), .B(mult_x_1196_n2183), 
        .Y(n22797) );
  OAI22xp5_ASAP7_75t_SL U33709 ( .A1(mult_x_1196_n2778), .A2(n24038), .B1(
        n22391), .B2(mult_x_1196_n2777), .Y(mult_x_1196_n929) );
  MAJIxp5_ASAP7_75t_SL U33710 ( .A(mult_x_1196_n1284), .B(n22348), .C(
        mult_x_1196_n1282), .Y(mult_x_1196_n1273) );
  MAJIxp5_ASAP7_75t_SL U33711 ( .A(mult_x_1196_n1269), .B(mult_x_1196_n1280), 
        .C(mult_x_1196_n1312), .Y(mult_x_1196_n1270) );
  INVx1_ASAP7_75t_SL U33712 ( .A(mult_x_1196_n1280), .Y(n22798) );
  INVx1_ASAP7_75t_SL U33713 ( .A(mult_x_1196_n1282), .Y(n22799) );
  INVx1_ASAP7_75t_SL U33714 ( .A(mult_x_1196_n701), .Y(mult_x_1196_n699) );
  OAI21xp5_ASAP7_75t_SL U33715 ( .A1(mult_x_1196_n3175), .A2(n23994), .B(
        n22800), .Y(mult_x_1196_n2599) );
  NAND2xp5_ASAP7_75t_SL U33716 ( .A(n22388), .B(n22801), .Y(n22800) );
  MAJIxp5_ASAP7_75t_SL U33717 ( .A(n24308), .B(mult_x_1196_n1732), .C(
        mult_x_1196_n1730), .Y(mult_x_1196_n1721) );
  XNOR2xp5_ASAP7_75t_SL U33718 ( .A(n22805), .B(n22804), .Y(mult_x_1196_n1994)
         );
  XOR2xp5_ASAP7_75t_SL U33719 ( .A(n22808), .B(mult_x_1196_n1249), .Y(n22807)
         );
  INVx1_ASAP7_75t_SL U33720 ( .A(mult_x_1196_n1253), .Y(n22808) );
  XOR2xp5_ASAP7_75t_SL U33721 ( .A(n24142), .B(mult_x_1196_n1025), .Y(n24143)
         );
  XNOR2xp5_ASAP7_75t_SL U33722 ( .A(n22364), .B(n22809), .Y(mult_x_1196_n1025)
         );
  NAND2xp33_ASAP7_75t_SRAM U33723 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__26_), 
        .B(n24685), .Y(n25109) );
  NAND2xp5_ASAP7_75t_SL U33724 ( .A(n22653), .B(n24302), .Y(n22811) );
  NOR2x1_ASAP7_75t_SL U33725 ( .A(n22653), .B(n24302), .Y(n22812) );
  XNOR2xp5_ASAP7_75t_SL U33726 ( .A(n23680), .B(n22271), .Y(n24187) );
  MAJIxp5_ASAP7_75t_SL U33727 ( .A(mult_x_1196_n2655), .B(mult_x_1196_n2623), 
        .C(n23646), .Y(mult_x_1196_n1945) );
  OAI22xp5_ASAP7_75t_SL U33728 ( .A1(n23984), .A2(mult_x_1196_n3230), .B1(
        n24121), .B2(mult_x_1196_n3231), .Y(mult_x_1196_n2655) );
  NOR2x1_ASAP7_75t_SL U33729 ( .A(mult_x_1196_n2729), .B(n24043), .Y(
        mult_x_1196_n2167) );
  XNOR2xp5_ASAP7_75t_SL U33730 ( .A(n23797), .B(n22813), .Y(mult_x_1196_n1949)
         );
  INVx1_ASAP7_75t_SL U33731 ( .A(mult_x_1196_n1956), .Y(n22813) );
  OAI22x1_ASAP7_75t_SL U33732 ( .A1(mult_x_1196_n2762), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2761), .Y(mult_x_1196_n2199) );
  OAI22xp5_ASAP7_75t_SL U33733 ( .A1(mult_x_1196_n3197), .A2(n23989), .B1(
        n24106), .B2(mult_x_1196_n3196), .Y(n22814) );
  BUFx6f_ASAP7_75t_SL U33734 ( .A(n24009), .Y(n22815) );
  INVx1_ASAP7_75t_SL U33735 ( .A(mult_x_1196_n752), .Y(mult_x_1196_n750) );
  BUFx3_ASAP7_75t_SL U33736 ( .A(n23993), .Y(n23081) );
  MAJIxp5_ASAP7_75t_SL U33737 ( .A(n23940), .B(mult_x_1196_n2289), .C(
        mult_x_1196_n2315), .Y(mult_x_1196_n1218) );
  XNOR2xp5_ASAP7_75t_SL U33738 ( .A(mult_x_1196_n1219), .B(n22816), .Y(n24199)
         );
  INVx1_ASAP7_75t_SL U33739 ( .A(mult_x_1196_n1223), .Y(n22816) );
  XNOR2xp5_ASAP7_75t_SL U33740 ( .A(n23940), .B(n22817), .Y(mult_x_1196_n1219)
         );
  XOR2xp5_ASAP7_75t_SL U33741 ( .A(mult_x_1196_n2315), .B(mult_x_1196_n2289), 
        .Y(n22817) );
  OAI21x1_ASAP7_75t_SL U33742 ( .A1(mult_x_1196_n579), .A2(mult_x_1196_n575), 
        .B(n24201), .Y(mult_x_1196_n570) );
  AOI21x1_ASAP7_75t_SL U33743 ( .A1(mult_x_1196_n555), .A2(mult_x_1196_n570), 
        .B(mult_x_1196_n556), .Y(mult_x_1196_n550) );
  MAJIxp5_ASAP7_75t_SL U33744 ( .A(mult_x_1196_n2024), .B(mult_x_1196_n2013), 
        .C(n22818), .Y(mult_x_1196_n2005) );
  INVx1_ASAP7_75t_SL U33745 ( .A(n22819), .Y(n22818) );
  INVx1_ASAP7_75t_SL U33746 ( .A(mult_x_1196_n2027), .Y(n22820) );
  MAJIxp5_ASAP7_75t_SL U33747 ( .A(n22861), .B(mult_x_1196_n2138), .C(
        mult_x_1196_n2565), .Y(n22821) );
  INVx1_ASAP7_75t_SL U33748 ( .A(mult_x_1196_n2078), .Y(mult_x_1196_n2067) );
  AND2x4_ASAP7_75t_SL U33749 ( .A(mult_x_1196_n2067), .B(mult_x_1196_n2070), 
        .Y(mult_x_1196_n744) );
  INVx1_ASAP7_75t_SL U33750 ( .A(mult_x_1196_n1985), .Y(n22823) );
  XOR2xp5_ASAP7_75t_SL U33751 ( .A(n22826), .B(n22825), .Y(mult_x_1196_n1961)
         );
  XNOR2xp5_ASAP7_75t_SL U33752 ( .A(n23052), .B(n23051), .Y(n22825) );
  INVx1_ASAP7_75t_SL U33753 ( .A(mult_x_1196_n1982), .Y(n22826) );
  BUFx6f_ASAP7_75t_SL U33754 ( .A(n24107), .Y(n23072) );
  NAND2xp33_ASAP7_75t_SRAM U33755 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__28_), 
        .B(n24685), .Y(n25102) );
  NOR2x1_ASAP7_75t_SL U33756 ( .A(mult_x_1196_n2733), .B(n24043), .Y(
        mult_x_1196_n2171) );
  XOR2xp5_ASAP7_75t_SL U33757 ( .A(mult_x_1196_n1685), .B(mult_x_1196_n1650), 
        .Y(n22828) );
  XNOR2xp5_ASAP7_75t_SL U33758 ( .A(mult_x_1196_n1974), .B(n23784), .Y(
        mult_x_1196_n1968) );
  XOR2xp5_ASAP7_75t_SL U33759 ( .A(n22209), .B(n24300), .Y(mult_x_1196_n1438)
         );
  NOR2x1p5_ASAP7_75t_SL U33760 ( .A(n23880), .B(n23879), .Y(n23878) );
  MAJIxp5_ASAP7_75t_SL U33761 ( .A(n24211), .B(n23749), .C(n24224), .Y(n23748)
         );
  MAJIxp5_ASAP7_75t_SL U33762 ( .A(mult_x_1196_n2353), .B(mult_x_1196_n2417), 
        .C(mult_x_1196_n2449), .Y(mult_x_1196_n1416) );
  XNOR2xp5_ASAP7_75t_SL U33763 ( .A(mult_x_1196_n1417), .B(mult_x_1196_n1406), 
        .Y(n24174) );
  NAND2x1_ASAP7_75t_SL U33764 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__21_), .B(
        n18910), .Y(n22830) );
  MAJIxp5_ASAP7_75t_SL U33765 ( .A(n23377), .B(mult_x_1196_n2050), .C(
        mult_x_1196_n2048), .Y(mult_x_1196_n2034) );
  MAJIxp5_ASAP7_75t_SL U33766 ( .A(mult_x_1196_n1775), .B(mult_x_1196_n1777), 
        .C(n22210), .Y(mult_x_1196_n1771) );
  XOR2xp5_ASAP7_75t_SL U33767 ( .A(mult_x_1196_n1777), .B(mult_x_1196_n1775), 
        .Y(n22831) );
  XOR2xp5_ASAP7_75t_SL U33768 ( .A(mult_x_1196_n1281), .B(n22832), .Y(
        mult_x_1196_n1242) );
  XNOR2xp5_ASAP7_75t_SL U33769 ( .A(mult_x_1196_n2153), .B(mult_x_1196_n2278), 
        .Y(n23347) );
  INVx1_ASAP7_75t_SL U33770 ( .A(mult_x_1196_n1709), .Y(n22833) );
  XNOR2xp5_ASAP7_75t_SL U33771 ( .A(mult_x_1196_n2583), .B(mult_x_1196_n2615), 
        .Y(n23341) );
  BUFx6f_ASAP7_75t_SL U33772 ( .A(n22255), .Y(n23981) );
  BUFx6f_ASAP7_75t_SL U33773 ( .A(mult_x_1196_n9), .Y(n23982) );
  XOR2xp5_ASAP7_75t_SL U33774 ( .A(mult_x_1196_n2048), .B(n23377), .Y(n23376)
         );
  MAJIxp5_ASAP7_75t_SL U33775 ( .A(mult_x_1196_n1034), .B(mult_x_1196_n2249), 
        .C(n22839), .Y(mult_x_1196_n1014) );
  XOR2xp5_ASAP7_75t_SL U33776 ( .A(mult_x_1196_n2249), .B(n22839), .Y(n22838)
         );
  OAI22xp5_ASAP7_75t_SL U33777 ( .A1(n24040), .A2(mult_x_1196_n2750), .B1(
        n24041), .B2(mult_x_1196_n2751), .Y(n22839) );
  INVx1_ASAP7_75t_SL U33778 ( .A(mult_x_1196_n1612), .Y(n22841) );
  NOR2x1_ASAP7_75t_SL U33779 ( .A(n22251), .B(mult_x_1196_n2836), .Y(n23493)
         );
  INVx5_ASAP7_75t_SL U33780 ( .A(n24001), .Y(n24002) );
  MAJIxp5_ASAP7_75t_SL U33781 ( .A(n22842), .B(mult_x_1196_n1891), .C(n22326), 
        .Y(mult_x_1196_n1868) );
  INVx2_ASAP7_75t_SL U33782 ( .A(mult_x_1196_n2558), .Y(n23724) );
  XNOR2xp5_ASAP7_75t_SL U33783 ( .A(mult_x_1196_n2045), .B(mult_x_1196_n2057), 
        .Y(n24116) );
  XNOR2xp5_ASAP7_75t_SL U33784 ( .A(n24073), .B(add_x_735_A_10_), .Y(
        mult_x_1196_n3140) );
  INVx1_ASAP7_75t_SL U33785 ( .A(mult_x_1196_n2388), .Y(n22844) );
  BUFx3_ASAP7_75t_SL U33786 ( .A(n24006), .Y(n23637) );
  XOR2xp5_ASAP7_75t_SL U33787 ( .A(mult_x_1196_n1672), .B(mult_x_1196_n1678), 
        .Y(n22846) );
  MAJIxp5_ASAP7_75t_SL U33788 ( .A(mult_x_1196_n1200), .B(n18931), .C(
        mult_x_1196_n1173), .Y(mult_x_1196_n1167) );
  OAI21xp5_ASAP7_75t_SL U33789 ( .A1(mult_x_1196_n1197), .A2(mult_x_1196_n1168), .B(n22341), .Y(n22847) );
  NAND2xp5_ASAP7_75t_SL U33790 ( .A(mult_x_1196_n1197), .B(mult_x_1196_n1168), 
        .Y(n22848) );
  XNOR2xp5_ASAP7_75t_SL U33791 ( .A(n22850), .B(mult_x_1196_n1200), .Y(n22849)
         );
  INVx1_ASAP7_75t_SL U33792 ( .A(mult_x_1196_n1203), .Y(n22850) );
  INVx1_ASAP7_75t_SL U33793 ( .A(mult_x_1196_n2679), .Y(n22852) );
  XNOR2xp5_ASAP7_75t_SL U33794 ( .A(n23015), .B(n23016), .Y(mult_x_1196_n1525)
         );
  XNOR2xp5_ASAP7_75t_SL U33795 ( .A(n22853), .B(n22475), .Y(mult_x_1196_n1802)
         );
  XNOR2xp5_ASAP7_75t_SL U33796 ( .A(n24110), .B(mult_x_1196_n1801), .Y(n24111)
         );
  XNOR2xp5_ASAP7_75t_SL U33797 ( .A(n22854), .B(n22678), .Y(n23124) );
  XOR2xp5_ASAP7_75t_SL U33798 ( .A(n23411), .B(n23122), .Y(n23123) );
  INVx1_ASAP7_75t_SL U33799 ( .A(mult_x_1196_n1438), .Y(n22854) );
  NAND2xp5_ASAP7_75t_SL U33800 ( .A(mult_x_1196_n1597), .B(mult_x_1196_n1627), 
        .Y(n22856) );
  XOR2xp5_ASAP7_75t_SL U33801 ( .A(mult_x_1196_n2470), .B(mult_x_1196_n2658), 
        .Y(n22858) );
  OAI22xp5_ASAP7_75t_SL U33802 ( .A1(mult_x_1196_n3188), .A2(n23072), .B1(
        mult_x_1196_n3187), .B2(n22248), .Y(n23931) );
  XNOR2xp5_ASAP7_75t_SL U33803 ( .A(n22859), .B(n22861), .Y(mult_x_1196_n2037)
         );
  XNOR2xp5_ASAP7_75t_SL U33804 ( .A(mult_x_1196_n2565), .B(n22860), .Y(n22859)
         );
  XNOR2xp5_ASAP7_75t_SL U33805 ( .A(mult_x_1196_n2693), .B(n23597), .Y(n22861)
         );
  MAJIxp5_ASAP7_75t_SL U33806 ( .A(n22862), .B(mult_x_1196_n2068), .C(
        mult_x_1196_n2080), .Y(mult_x_1196_n2069) );
  XNOR2xp5_ASAP7_75t_SL U33807 ( .A(mult_x_1196_n2068), .B(mult_x_1196_n2080), 
        .Y(n22863) );
  INVx1_ASAP7_75t_SL U33808 ( .A(mult_x_1196_n1554), .Y(n22865) );
  XNOR2xp5_ASAP7_75t_SL U33809 ( .A(mult_x_1196_n1703), .B(mult_x_1196_n1705), 
        .Y(n22866) );
  INVx1_ASAP7_75t_SL U33810 ( .A(mult_x_1196_n1676), .Y(n22867) );
  INVx1_ASAP7_75t_SL U33811 ( .A(n22870), .Y(n22868) );
  INVx1_ASAP7_75t_SL U33812 ( .A(mult_x_1196_n2520), .Y(n22871) );
  INVx1_ASAP7_75t_SL U33813 ( .A(n22874), .Y(n22872) );
  XNOR2xp5_ASAP7_75t_SL U33814 ( .A(n22874), .B(mult_x_1196_n2206), .Y(n22873)
         );
  NOR2x1_ASAP7_75t_SL U33815 ( .A(n22876), .B(n22875), .Y(n22874) );
  NOR2x1_ASAP7_75t_SL U33816 ( .A(mult_x_1196_n3217), .B(n24082), .Y(n22875)
         );
  NOR2x1_ASAP7_75t_SL U33817 ( .A(n23984), .B(mult_x_1196_n3216), .Y(n22876)
         );
  MAJIxp5_ASAP7_75t_SL U33818 ( .A(n22878), .B(mult_x_1196_n2312), .C(
        mult_x_1196_n2158), .Y(mult_x_1196_n1054) );
  XNOR2xp5_ASAP7_75t_SL U33819 ( .A(mult_x_1196_n2312), .B(n22877), .Y(
        mult_x_1196_n1055) );
  OAI22xp5_ASAP7_75t_SL U33820 ( .A1(mult_x_1196_n2945), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2944), .Y(n22878) );
  A2O1A1Ixp33_ASAP7_75t_SL U33821 ( .A1(n22881), .A2(n22880), .B(n24281), .C(
        n22879), .Y(mult_x_1196_n1294) );
  INVx1_ASAP7_75t_SL U33822 ( .A(n22883), .Y(n22880) );
  INVx1_ASAP7_75t_SL U33823 ( .A(n22884), .Y(n22881) );
  XNOR2xp5_ASAP7_75t_SL U33824 ( .A(n24281), .B(n22882), .Y(mult_x_1196_n1295)
         );
  XOR2xp5_ASAP7_75t_SL U33825 ( .A(n22884), .B(n22883), .Y(n22882) );
  MAJIxp5_ASAP7_75t_SL U33826 ( .A(mult_x_1196_n1834), .B(n18303), .C(
        mult_x_1196_n1852), .Y(mult_x_1196_n1825) );
  INVx1_ASAP7_75t_SL U33827 ( .A(n22887), .Y(n22885) );
  XNOR2xp5_ASAP7_75t_SL U33828 ( .A(n22887), .B(mult_x_1196_n1846), .Y(n22886)
         );
  XOR2xp5_ASAP7_75t_SL U33829 ( .A(n22889), .B(n22888), .Y(n22887) );
  INVx1_ASAP7_75t_SL U33830 ( .A(mult_x_1196_n1852), .Y(n22889) );
  MAJIxp5_ASAP7_75t_SL U33831 ( .A(n22890), .B(mult_x_1196_n2627), .C(
        mult_x_1196_n2595), .Y(mult_x_1196_n2012) );
  XNOR2xp5_ASAP7_75t_SL U33832 ( .A(n22893), .B(n22891), .Y(mult_x_1196_n2013)
         );
  XOR2xp5_ASAP7_75t_SL U33833 ( .A(mult_x_1196_n2595), .B(n22892), .Y(n22891)
         );
  INVx1_ASAP7_75t_SL U33834 ( .A(mult_x_1196_n2627), .Y(n22892) );
  INVx1_ASAP7_75t_SL U33835 ( .A(n23541), .Y(n22895) );
  XNOR2x2_ASAP7_75t_SL U33836 ( .A(n23367), .B(n23368), .Y(mult_x_1196_n1887)
         );
  INVx1_ASAP7_75t_SL U33837 ( .A(mult_x_1196_n1351), .Y(n22896) );
  XNOR2xp5_ASAP7_75t_SL U33838 ( .A(mult_x_1196_n1416), .B(mult_x_1196_n1418), 
        .Y(n22898) );
  INVx1_ASAP7_75t_SL U33839 ( .A(mult_x_1196_n1424), .Y(n22899) );
  BUFx5_ASAP7_75t_SL U33840 ( .A(n23444), .Y(n23442) );
  MAJIxp5_ASAP7_75t_SL U33841 ( .A(n22901), .B(mult_x_1196_n1802), .C(n22550), 
        .Y(mult_x_1196_n1796) );
  XOR2xp5_ASAP7_75t_SL U33842 ( .A(mult_x_1196_n1822), .B(mult_x_1196_n1802), 
        .Y(n22900) );
  MAJIxp5_ASAP7_75t_SL U33843 ( .A(n24090), .B(n22521), .C(n22528), .Y(
        mult_x_1196_n1083) );
  XNOR2xp5_ASAP7_75t_SL U33844 ( .A(n22904), .B(n22339), .Y(n22903) );
  INVx1_ASAP7_75t_SL U33845 ( .A(mult_x_1196_n1089), .Y(n22904) );
  NOR2x1_ASAP7_75t_SL U33846 ( .A(n22983), .B(mult_x_1196_n2900), .Y(n24159)
         );
  MAJIxp5_ASAP7_75t_SL U33847 ( .A(mult_x_1196_n1362), .B(n24260), .C(n22905), 
        .Y(mult_x_1196_n1327) );
  XNOR2x2_ASAP7_75t_SL U33848 ( .A(mult_x_1196_n2251), .B(n24093), .Y(
        mult_x_1196_n1057) );
  INVx1_ASAP7_75t_SL U33849 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__31_), .Y(
        n25237) );
  INVx2_ASAP7_75t_SL U33850 ( .A(u0_0_leon3x0_p0_muli[42]), .Y(n23956) );
  HB1xp67_ASAP7_75t_SL U33851 ( .A(n23482), .Y(n22906) );
  XNOR2xp5_ASAP7_75t_SL U33852 ( .A(mult_x_1196_n2040), .B(n22907), .Y(
        mult_x_1196_n2029) );
  XOR2xp5_ASAP7_75t_SL U33853 ( .A(mult_x_1196_n2692), .B(n23500), .Y(n22907)
         );
  MAJIxp5_ASAP7_75t_SL U33854 ( .A(mult_x_1196_n1361), .B(mult_x_1196_n1372), 
        .C(mult_x_1196_n1400), .Y(mult_x_1196_n1362) );
  NAND2xp5_ASAP7_75t_SL U33855 ( .A(n22910), .B(n22908), .Y(mult_x_1196_n893)
         );
  NAND2xp5_ASAP7_75t_SL U33856 ( .A(n22909), .B(mult_x_1196_n910), .Y(n22908)
         );
  NAND2xp5_ASAP7_75t_SL U33857 ( .A(mult_x_1196_n912), .B(mult_x_1196_n899), 
        .Y(n22909) );
  NAND2xp5_ASAP7_75t_SL U33858 ( .A(n22911), .B(n22913), .Y(n22910) );
  XNOR2xp5_ASAP7_75t_SL U33859 ( .A(mult_x_1196_n910), .B(n22912), .Y(
        mult_x_1196_n894) );
  XOR2xp5_ASAP7_75t_SL U33860 ( .A(mult_x_1196_n912), .B(n22913), .Y(n22912)
         );
  INVx1_ASAP7_75t_SL U33861 ( .A(mult_x_1196_n899), .Y(n22913) );
  XNOR2xp5_ASAP7_75t_SL U33862 ( .A(n22914), .B(n22916), .Y(mult_x_1196_n1374)
         );
  XNOR2xp5_ASAP7_75t_SL U33863 ( .A(n22915), .B(mult_x_1196_n1420), .Y(n22914)
         );
  INVx1_ASAP7_75t_SL U33864 ( .A(mult_x_1196_n1422), .Y(n22915) );
  OAI21x1_ASAP7_75t_SL U33865 ( .A1(n23100), .A2(mult_x_1196_n3098), .B(n22917), .Y(n23125) );
  XOR2xp5_ASAP7_75t_SL U33866 ( .A(add_x_735_A_15_), .B(add_x_735_A_16_), .Y(
        mult_x_1196_n3323) );
  MAJIxp5_ASAP7_75t_SL U33867 ( .A(mult_x_1196_n2457), .B(mult_x_1196_n2361), 
        .C(n23679), .Y(mult_x_1196_n1703) );
  OAI22xp5_ASAP7_75t_SL U33868 ( .A1(mult_x_1196_n3029), .A2(n22563), .B1(
        mult_x_1196_n3028), .B2(n22540), .Y(mult_x_1196_n2457) );
  NAND2x1_ASAP7_75t_SL U33869 ( .A(n24193), .B(n24195), .Y(mult_x_1196_n1262)
         );
  XNOR2xp5_ASAP7_75t_SL U33870 ( .A(mult_x_1196_n1443), .B(n23615), .Y(n23614)
         );
  MAJIxp5_ASAP7_75t_SL U33871 ( .A(mult_x_1196_n1522), .B(mult_x_1196_n1488), 
        .C(mult_x_1196_n1524), .Y(n23615) );
  NAND2xp5_ASAP7_75t_SL U33872 ( .A(n22921), .B(n22920), .Y(mult_x_1196_n1312)
         );
  OAI21xp5_ASAP7_75t_SL U33873 ( .A1(n22924), .A2(n22923), .B(n22925), .Y(
        n22920) );
  OR2x2_ASAP7_75t_SL U33874 ( .A(mult_x_1196_n2446), .B(mult_x_1196_n2538), 
        .Y(n22921) );
  XNOR2xp5_ASAP7_75t_SL U33875 ( .A(n22924), .B(n22923), .Y(n22922) );
  INVx1_ASAP7_75t_SL U33876 ( .A(mult_x_1196_n2446), .Y(n22924) );
  INVx1_ASAP7_75t_SL U33877 ( .A(n23306), .Y(n23308) );
  BUFx12f_ASAP7_75t_SL U33878 ( .A(add_x_735_A_32_), .Y(n22926) );
  MAJIxp5_ASAP7_75t_SL U33879 ( .A(mult_x_1196_n1086), .B(mult_x_1196_n1064), 
        .C(mult_x_1196_n1062), .Y(mult_x_1196_n1058) );
  XNOR2xp5_ASAP7_75t_SL U33880 ( .A(mult_x_1196_n1062), .B(n22927), .Y(
        mult_x_1196_n1059) );
  INVx3_ASAP7_75t_SL U33881 ( .A(n23974), .Y(n23976) );
  INVx1_ASAP7_75t_SL U33882 ( .A(mult_x_1196_n1237), .Y(n24238) );
  OAI22x1_ASAP7_75t_SL U33883 ( .A1(mult_x_1196_n2989), .A2(n23311), .B1(
        mult_x_1196_n2988), .B2(n24012), .Y(mult_x_1196_n2417) );
  NOR2x1_ASAP7_75t_SL U33884 ( .A(mult_x_1196_n2730), .B(n24043), .Y(
        mult_x_1196_n2168) );
  OAI21x1_ASAP7_75t_SL U33885 ( .A1(mult_x_1196_n2991), .A2(n23311), .B(n22300), .Y(mult_x_1196_n2419) );
  XNOR2xp5_ASAP7_75t_SL U33886 ( .A(n23664), .B(mult_x_1196_n2035), .Y(
        mult_x_1196_n2030) );
  MAJIxp5_ASAP7_75t_SL U33887 ( .A(mult_x_1196_n1477), .B(mult_x_1196_n1479), 
        .C(mult_x_1196_n1471), .Y(mult_x_1196_n1472) );
  XOR2xp5_ASAP7_75t_SL U33888 ( .A(mult_x_1196_n1477), .B(mult_x_1196_n1479), 
        .Y(n22934) );
  OAI22x1_ASAP7_75t_SL U33889 ( .A1(mult_x_1196_n3120), .A2(n23999), .B1(
        n23997), .B2(mult_x_1196_n3119), .Y(mult_x_1196_n2544) );
  OAI21x1_ASAP7_75t_SL U33890 ( .A1(n25138), .A2(n24686), .B(n25137), .Y(
        add_x_735_A_12_) );
  NAND2x1_ASAP7_75t_SL U33891 ( .A(n22218), .B(n23041), .Y(n24285) );
  XOR2xp5_ASAP7_75t_SL U33892 ( .A(n22937), .B(n24111), .Y(mult_x_1196_n1775)
         );
  INVx1_ASAP7_75t_SL U33893 ( .A(n24077), .Y(n22937) );
  AOI21xp5_ASAP7_75t_SL U33894 ( .A1(n23107), .A2(n23782), .B(n23488), .Y(
        n22938) );
  XOR2xp5_ASAP7_75t_SL U33895 ( .A(mult_x_1196_n1459), .B(mult_x_1196_n1425), 
        .Y(n24108) );
  BUFx6f_ASAP7_75t_SL U33896 ( .A(mult_x_1196_n126), .Y(n24035) );
  INVx1_ASAP7_75t_SL U33897 ( .A(n23107), .Y(n22940) );
  INVx1_ASAP7_75t_SL U33898 ( .A(n23782), .Y(n22941) );
  NAND2x1_ASAP7_75t_SL U33899 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__4_), .B(n24686), .Y(n25087) );
  XOR2xp5_ASAP7_75t_SL U33900 ( .A(n22943), .B(n23924), .Y(n22942) );
  XNOR2xp5_ASAP7_75t_SL U33901 ( .A(n22310), .B(n24199), .Y(n22943) );
  MAJIxp5_ASAP7_75t_SL U33902 ( .A(mult_x_1196_n1204), .B(mult_x_1196_n1196), 
        .C(n22944), .Y(mult_x_1196_n1197) );
  MAJIxp5_ASAP7_75t_SL U33903 ( .A(mult_x_1196_n1237), .B(mult_x_1196_n1240), 
        .C(mult_x_1196_n1270), .Y(n22944) );
  MAJIxp5_ASAP7_75t_SL U33904 ( .A(mult_x_1196_n2054), .B(mult_x_1196_n2139), 
        .C(mult_x_1196_n2060), .Y(mult_x_1196_n2055) );
  OAI21xp5_ASAP7_75t_SL U33905 ( .A1(mult_x_1196_n2065), .A2(mult_x_1196_n2058), .B(n22945), .Y(mult_x_1196_n2052) );
  NAND2xp5_ASAP7_75t_SL U33906 ( .A(n22948), .B(n22946), .Y(n22945) );
  NAND2xp5_ASAP7_75t_SL U33907 ( .A(mult_x_1196_n2065), .B(mult_x_1196_n2058), 
        .Y(n22946) );
  XNOR2xp5_ASAP7_75t_SL U33908 ( .A(n22948), .B(n22947), .Y(mult_x_1196_n2053)
         );
  XOR2xp5_ASAP7_75t_SL U33909 ( .A(mult_x_1196_n2054), .B(n22949), .Y(n22948)
         );
  XOR2xp5_ASAP7_75t_SL U33910 ( .A(mult_x_1196_n2139), .B(mult_x_1196_n2060), 
        .Y(n22949) );
  MAJx2_ASAP7_75t_SL U33911 ( .A(n22439), .B(mult_x_1196_n1318), .C(
        mult_x_1196_n1286), .Y(mult_x_1196_n1235) );
  NOR2xp33_ASAP7_75t_SL U33912 ( .A(mult_x_1196_n3034), .B(n24009), .Y(n22951)
         );
  OAI22x1_ASAP7_75t_SL U33913 ( .A1(mult_x_1196_n2990), .A2(n23311), .B1(
        mult_x_1196_n2989), .B2(n24012), .Y(mult_x_1196_n2418) );
  MAJIxp5_ASAP7_75t_SL U33914 ( .A(mult_x_1196_n2662), .B(mult_x_1196_n2534), 
        .C(n22954), .Y(mult_x_1196_n2048) );
  INVx1_ASAP7_75t_SL U33915 ( .A(n22956), .Y(n22954) );
  XNOR2xp5_ASAP7_75t_SL U33916 ( .A(n22956), .B(n22955), .Y(mult_x_1196_n2049)
         );
  NOR2x1_ASAP7_75t_SL U33917 ( .A(n22958), .B(n22957), .Y(n22956) );
  INVx1_ASAP7_75t_SL U33918 ( .A(mult_x_1196_n2136), .Y(n22959) );
  INVx1_ASAP7_75t_SL U33919 ( .A(mult_x_1196_n1981), .Y(n22960) );
  NAND2xp5_ASAP7_75t_SL U33920 ( .A(n18365), .B(n23359), .Y(n23751) );
  XNOR2xp5_ASAP7_75t_SL U33921 ( .A(mult_x_1196_n1297), .B(n22963), .Y(
        mult_x_1196_n1263) );
  XNOR2xp5_ASAP7_75t_SL U33922 ( .A(n22964), .B(n24191), .Y(n22963) );
  INVx1_ASAP7_75t_SL U33923 ( .A(mult_x_1196_n1299), .Y(n22964) );
  XNOR2xp5_ASAP7_75t_SL U33924 ( .A(mult_x_1196_n1620), .B(n23813), .Y(
        mult_x_1196_n1613) );
  XNOR2xp5_ASAP7_75t_SL U33925 ( .A(n22967), .B(mult_x_1196_n1474), .Y(n22966)
         );
  BUFx5_ASAP7_75t_SL U33926 ( .A(n22285), .Y(n22968) );
  MAJIxp5_ASAP7_75t_SL U33927 ( .A(mult_x_1196_n2252), .B(n22970), .C(
        mult_x_1196_n2406), .Y(mult_x_1196_n1077) );
  XNOR2xp5_ASAP7_75t_SL U33928 ( .A(n22971), .B(n22969), .Y(mult_x_1196_n1078)
         );
  XNOR2xp5_ASAP7_75t_SL U33929 ( .A(n22970), .B(mult_x_1196_n2406), .Y(n22969)
         );
  OAI22xp5_ASAP7_75t_SL U33930 ( .A1(mult_x_1196_n3010), .A2(n22815), .B1(
        n23442), .B2(mult_x_1196_n3009), .Y(n22970) );
  XOR2xp5_ASAP7_75t_SL U33931 ( .A(mult_x_1196_n1113), .B(n22972), .Y(n24090)
         );
  NOR2x1p5_ASAP7_75t_SL U33932 ( .A(mult_x_1196_n526), .B(mult_x_1196_n519), 
        .Y(mult_x_1196_n517) );
  INVx1_ASAP7_75t_SL U33933 ( .A(n23593), .Y(n22973) );
  INVx1_ASAP7_75t_SL U33934 ( .A(mult_x_1196_n2161), .Y(n24117) );
  NOR2x1_ASAP7_75t_SL U33935 ( .A(mult_x_1196_n3094), .B(n18654), .Y(n23109)
         );
  MAJIxp5_ASAP7_75t_SL U33936 ( .A(mult_x_1196_n2160), .B(n22976), .C(
        mult_x_1196_n2313), .Y(mult_x_1196_n1101) );
  XOR2xp5_ASAP7_75t_SL U33937 ( .A(mult_x_1196_n2313), .B(n22975), .Y(
        mult_x_1196_n1102) );
  XNOR2xp5_ASAP7_75t_SL U33938 ( .A(n22976), .B(mult_x_1196_n2160), .Y(n22975)
         );
  OAI22xp5_ASAP7_75t_SL U33939 ( .A1(mult_x_1196_n2851), .A2(n24031), .B1(
        n22743), .B2(mult_x_1196_n2850), .Y(n22976) );
  MAJIxp5_ASAP7_75t_SL U33940 ( .A(n22259), .B(n22211), .C(n22977), .Y(
        mult_x_1196_n1889) );
  INVx1_ASAP7_75t_SL U33941 ( .A(n22978), .Y(n22977) );
  INVx1_ASAP7_75t_SL U33942 ( .A(mult_x_1196_n1916), .Y(n22979) );
  XNOR2xp5_ASAP7_75t_SL U33943 ( .A(mult_x_1196_n2390), .B(n22981), .Y(n22980)
         );
  OAI22xp5_ASAP7_75t_SL U33944 ( .A1(mult_x_1196_n2802), .A2(n24039), .B1(
        mult_x_1196_n2801), .B2(n22391), .Y(n22981) );
  INVx1_ASAP7_75t_SL U33945 ( .A(mult_x_1196_n2300), .Y(n22982) );
  MAJIxp5_ASAP7_75t_SL U33946 ( .A(n22984), .B(n22337), .C(mult_x_1196_n1159), 
        .Y(mult_x_1196_n1147) );
  MAJIxp5_ASAP7_75t_SL U33947 ( .A(mult_x_1196_n1636), .B(n22985), .C(
        mult_x_1196_n1612), .Y(mult_x_1196_n1593) );
  INVx1_ASAP7_75t_SL U33948 ( .A(mult_x_1196_n1078), .Y(n22987) );
  XNOR2xp5_ASAP7_75t_SL U33949 ( .A(n22989), .B(n22988), .Y(mult_x_1196_n1009)
         );
  MAJIxp5_ASAP7_75t_SL U33950 ( .A(n23082), .B(mult_x_1196_n2340), .C(
        mult_x_1196_n2282), .Y(n22988) );
  XNOR2xp5_ASAP7_75t_SL U33951 ( .A(n22990), .B(mult_x_1196_n1028), .Y(n22989)
         );
  INVx1_ASAP7_75t_SL U33952 ( .A(n24253), .Y(n22990) );
  XNOR2xp5_ASAP7_75t_SL U33953 ( .A(mult_x_1196_n1825), .B(n22992), .Y(n22991)
         );
  INVx1_ASAP7_75t_SL U33954 ( .A(mult_x_1196_n1807), .Y(n22992) );
  MAJIxp5_ASAP7_75t_SL U33955 ( .A(mult_x_1196_n1527), .B(n22299), .C(n22994), 
        .Y(mult_x_1196_n1516) );
  XNOR2xp5_ASAP7_75t_SL U33956 ( .A(n22299), .B(n22994), .Y(n22993) );
  MAJx2_ASAP7_75t_SL U33957 ( .A(n23352), .B(mult_x_1196_n1317), .C(n18400), 
        .Y(mult_x_1196_n1269) );
  MAJIxp5_ASAP7_75t_SL U33958 ( .A(mult_x_1196_n2281), .B(n22995), .C(
        mult_x_1196_n2339), .Y(mult_x_1196_n1010) );
  OAI21xp5_ASAP7_75t_SL U33959 ( .A1(mult_x_1196_n2783), .A2(n22412), .B(
        n22996), .Y(n22995) );
  NAND2xp5_ASAP7_75t_SL U33960 ( .A(n22998), .B(n22997), .Y(n22996) );
  INVx1_ASAP7_75t_SL U33961 ( .A(n22936), .Y(n22998) );
  XOR2xp5_ASAP7_75t_SL U33962 ( .A(mult_x_1196_n1559), .B(mult_x_1196_n1557), 
        .Y(n23000) );
  XNOR2xp5_ASAP7_75t_SL U33963 ( .A(mult_x_1196_n1493), .B(n23001), .Y(
        mult_x_1196_n1484) );
  XOR2xp5_ASAP7_75t_SL U33964 ( .A(mult_x_1196_n1497), .B(mult_x_1196_n1501), 
        .Y(n23001) );
  MAJIxp5_ASAP7_75t_SL U33965 ( .A(n23123), .B(mult_x_1196_n1438), .C(
        mult_x_1196_n1483), .Y(mult_x_1196_n1439) );
  NAND2xp5_ASAP7_75t_SL U33966 ( .A(n24192), .B(n22261), .Y(n24193) );
  XOR2xp5_ASAP7_75t_SL U33967 ( .A(mult_x_1196_n1473), .B(n23242), .Y(
        mult_x_1196_n1467) );
  AOI21x1_ASAP7_75t_SL U33968 ( .A1(n24272), .A2(mult_x_1196_n753), .B(
        mult_x_1196_n750), .Y(mult_x_1196_n748) );
  MAJIxp5_ASAP7_75t_SL U33969 ( .A(n23003), .B(n22354), .C(mult_x_1196_n1334), 
        .Y(mult_x_1196_n1297) );
  XNOR2xp5_ASAP7_75t_SL U33970 ( .A(n22595), .B(n23004), .Y(mult_x_1196_n1298)
         );
  XNOR2xp5_ASAP7_75t_SL U33971 ( .A(n22354), .B(mult_x_1196_n1334), .Y(n23004)
         );
  MAJIxp5_ASAP7_75t_SL U33972 ( .A(n24152), .B(n24153), .C(n22350), .Y(n23005)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U33973 ( .A1(mult_x_1196_n2666), .A2(
        mult_x_1196_n2602), .B(mult_x_1196_n2077), .C(n23006), .Y(
        mult_x_1196_n2078) );
  NAND2xp5_ASAP7_75t_SL U33974 ( .A(n23007), .B(n23009), .Y(n23006) );
  INVx1_ASAP7_75t_SL U33975 ( .A(mult_x_1196_n2602), .Y(n23007) );
  NAND2xp5_ASAP7_75t_SL U33976 ( .A(n22222), .B(mult_x_1196_n2075), .Y(
        mult_x_1196_n752) );
  XNOR2xp5_ASAP7_75t_SL U33977 ( .A(n23008), .B(mult_x_1196_n2077), .Y(
        mult_x_1196_n2075) );
  XOR2xp5_ASAP7_75t_SL U33978 ( .A(mult_x_1196_n2602), .B(n23009), .Y(n23008)
         );
  MAJIxp5_ASAP7_75t_SL U33979 ( .A(n24309), .B(n23011), .C(n23010), .Y(
        mult_x_1196_n1822) );
  INVx1_ASAP7_75t_SL U33980 ( .A(n23013), .Y(n23010) );
  MAJIxp5_ASAP7_75t_SL U33981 ( .A(mult_x_1196_n1858), .B(mult_x_1196_n1862), 
        .C(n23088), .Y(n23011) );
  XOR2xp5_ASAP7_75t_SL U33982 ( .A(n23013), .B(n24309), .Y(n23012) );
  XNOR2xp5_ASAP7_75t_SL U33983 ( .A(n23090), .B(n23514), .Y(n23013) );
  MAJIxp5_ASAP7_75t_SL U33984 ( .A(mult_x_1196_n1571), .B(n22651), .C(n23014), 
        .Y(mult_x_1196_n1524) );
  INVx1_ASAP7_75t_SL U33985 ( .A(n23016), .Y(n23014) );
  MAJIxp5_ASAP7_75t_SL U33986 ( .A(n23018), .B(mult_x_1196_n1792), .C(
        mult_x_1196_n1788), .Y(mult_x_1196_n1756) );
  XOR2xp5_ASAP7_75t_SL U33987 ( .A(mult_x_1196_n1792), .B(mult_x_1196_n1788), 
        .Y(n23017) );
  XNOR2xp5_ASAP7_75t_SL U33988 ( .A(mult_x_1196_n2647), .B(n24204), .Y(n23018)
         );
  XNOR2xp5_ASAP7_75t_SL U33989 ( .A(n23019), .B(n23020), .Y(mult_x_1196_n1932)
         );
  XNOR2xp5_ASAP7_75t_SL U33990 ( .A(n23022), .B(n23021), .Y(n23020) );
  XOR2xp5_ASAP7_75t_SL U33991 ( .A(mult_x_1196_n1957), .B(n22307), .Y(n23021)
         );
  INVx1_ASAP7_75t_SL U33992 ( .A(mult_x_1196_n1940), .Y(n23022) );
  XNOR2xp5_ASAP7_75t_SL U33993 ( .A(mult_x_1196_n2284), .B(mult_x_1196_n2220), 
        .Y(n23023) );
  XNOR2xp5_ASAP7_75t_SL U33994 ( .A(mult_x_1196_n1912), .B(mult_x_1196_n1937), 
        .Y(n23025) );
  MAJIxp5_ASAP7_75t_SL U33995 ( .A(n24292), .B(mult_x_1196_n1188), .C(n23028), 
        .Y(mult_x_1196_n1175) );
  INVx1_ASAP7_75t_SL U33996 ( .A(n23030), .Y(n23028) );
  XOR2xp5_ASAP7_75t_SL U33997 ( .A(mult_x_1196_n2378), .B(n24178), .Y(n23030)
         );
  MAJIxp5_ASAP7_75t_SL U33998 ( .A(mult_x_1196_n960), .B(mult_x_1196_n2245), 
        .C(n23032), .Y(mult_x_1196_n944) );
  XNOR2xp5_ASAP7_75t_SL U33999 ( .A(n23032), .B(n23031), .Y(mult_x_1196_n945)
         );
  XOR2xp5_ASAP7_75t_SL U34000 ( .A(mult_x_1196_n2245), .B(mult_x_1196_n960), 
        .Y(n23031) );
  OAI22xp5_ASAP7_75t_SL U34001 ( .A1(n24040), .A2(mult_x_1196_n2746), .B1(
        n18364), .B2(mult_x_1196_n2747), .Y(n23032) );
  XNOR2xp5_ASAP7_75t_SL U34002 ( .A(n24060), .B(n23955), .Y(mult_x_1196_n3229)
         );
  MAJIxp5_ASAP7_75t_SL U34003 ( .A(mult_x_1196_n1433), .B(n22358), .C(n23033), 
        .Y(mult_x_1196_n1394) );
  INVx1_ASAP7_75t_SL U34004 ( .A(n23035), .Y(n23033) );
  XNOR2xp5_ASAP7_75t_SL U34005 ( .A(n23036), .B(n23034), .Y(mult_x_1196_n1395)
         );
  XOR2xp5_ASAP7_75t_SL U34006 ( .A(mult_x_1196_n1433), .B(n23035), .Y(n23034)
         );
  INVx1_ASAP7_75t_SL U34007 ( .A(n22358), .Y(n23036) );
  NAND2x1_ASAP7_75t_SL U34008 ( .A(n23505), .B(n23507), .Y(mult_x_1196_n1113)
         );
  XNOR2xp5_ASAP7_75t_SL U34009 ( .A(n23038), .B(mult_x_1196_n2005), .Y(n23037)
         );
  INVx1_ASAP7_75t_SL U34010 ( .A(mult_x_1196_n1994), .Y(n23038) );
  NAND2xp5_ASAP7_75t_SL U34011 ( .A(n24285), .B(n23040), .Y(mult_x_1196_n540)
         );
  NAND2xp5_ASAP7_75t_SL U34012 ( .A(mult_x_1196_n1295), .B(n23786), .Y(n23041)
         );
  MAJIxp5_ASAP7_75t_SL U34013 ( .A(mult_x_1196_n2562), .B(n23043), .C(
        mult_x_1196_n2594), .Y(mult_x_1196_n1995) );
  XNOR2xp5_ASAP7_75t_SL U34014 ( .A(n23043), .B(mult_x_1196_n2594), .Y(n23042)
         );
  OAI22xp5_ASAP7_75t_SL U34015 ( .A1(mult_x_1196_n3074), .A2(n24007), .B1(
        n24005), .B2(mult_x_1196_n3073), .Y(n23043) );
  INVx1_ASAP7_75t_SL U34016 ( .A(mult_x_1196_n2562), .Y(n23044) );
  OAI21x1_ASAP7_75t_SL U34017 ( .A1(mult_x_1196_n3155), .A2(n24230), .B(n24267), .Y(n24123) );
  MAJIxp5_ASAP7_75t_SL U34018 ( .A(mult_x_1196_n2064), .B(n23045), .C(
        mult_x_1196_n2071), .Y(mult_x_1196_n2061) );
  XOR2xp5_ASAP7_75t_SL U34019 ( .A(n22331), .B(n23047), .Y(n23046) );
  XOR2xp5_ASAP7_75t_SL U34020 ( .A(n23585), .B(n23048), .Y(n23584) );
  INVx1_ASAP7_75t_SL U34021 ( .A(mult_x_1196_n2573), .Y(n23048) );
  OAI22xp5_ASAP7_75t_SL U34022 ( .A1(n24287), .A2(mult_x_1196_n3149), .B1(
        mult_x_1196_n3148), .B2(n23992), .Y(mult_x_1196_n2573) );
  NAND2xp5_ASAP7_75t_SL U34023 ( .A(mult_x_1196_n2686), .B(mult_x_1196_n2526), 
        .Y(n24219) );
  OAI21x1_ASAP7_75t_SL U34024 ( .A1(n23550), .A2(n24686), .B(n25145), .Y(
        add_x_735_A_24_) );
  INVx1_ASAP7_75t_SL U34025 ( .A(mult_x_1196_n1959), .Y(n23051) );
  MAJIxp5_ASAP7_75t_SL U34026 ( .A(mult_x_1196_n2561), .B(n23625), .C(
        mult_x_1196_n2501), .Y(n23052) );
  OAI21x1_ASAP7_75t_SL U34027 ( .A1(mult_x_1196_n387), .A2(mult_x_1196_n434), 
        .B(mult_x_1196_n390), .Y(mult_x_1196_n386) );
  NAND2xp5_ASAP7_75t_SL U34028 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__7_), .B(
        n18911), .Y(n25144) );
  XNOR2x1_ASAP7_75t_SL U34029 ( .A(n23125), .B(n23288), .Y(n24234) );
  INVx1_ASAP7_75t_SL U34030 ( .A(mult_x_1196_n2566), .Y(mult_x_1196_n2045) );
  MAJIxp5_ASAP7_75t_SL U34031 ( .A(mult_x_1196_n1305), .B(n23053), .C(n18934), 
        .Y(mult_x_1196_n1267) );
  INVx1_ASAP7_75t_SL U34032 ( .A(n23055), .Y(n23053) );
  XNOR2xp5_ASAP7_75t_SL U34033 ( .A(n23055), .B(mult_x_1196_n1305), .Y(n23054)
         );
  XOR2xp5_ASAP7_75t_SL U34034 ( .A(mult_x_1196_n1320), .B(n24164), .Y(n23055)
         );
  MAJIxp5_ASAP7_75t_SL U34035 ( .A(n23056), .B(mult_x_1196_n2324), .C(
        mult_x_1196_n2266), .Y(mult_x_1196_n1536) );
  OAI22xp5_ASAP7_75t_SL U34036 ( .A1(mult_x_1196_n3248), .A2(n23981), .B1(
        n22389), .B2(mult_x_1196_n3247), .Y(n23056) );
  MAJIxp5_ASAP7_75t_SL U34037 ( .A(mult_x_1196_n1371), .B(mult_x_1196_n1345), 
        .C(mult_x_1196_n1373), .Y(mult_x_1196_n1334) );
  OAI21x1_ASAP7_75t_SL U34038 ( .A1(mult_x_1196_n3037), .A2(n22815), .B(n22291), .Y(mult_x_1196_n2465) );
  XNOR2xp5_ASAP7_75t_SL U34039 ( .A(n23059), .B(n23058), .Y(mult_x_1196_n1369)
         );
  INVx1_ASAP7_75t_SL U34040 ( .A(n23369), .Y(n23059) );
  MAJIxp5_ASAP7_75t_SL U34041 ( .A(mult_x_1196_n2642), .B(mult_x_1196_n2207), 
        .C(mult_x_1196_n2326), .Y(mult_x_1196_n1609) );
  XNOR2xp5_ASAP7_75t_SL U34042 ( .A(mult_x_1196_n2207), .B(mult_x_1196_n2642), 
        .Y(n23062) );
  INVx1_ASAP7_75t_SL U34043 ( .A(mult_x_1196_n2326), .Y(n23063) );
  OAI21xp5_ASAP7_75t_SL U34044 ( .A1(mult_x_1196_n2335), .A2(mult_x_1196_n2213), .B(n23064), .Y(mult_x_1196_n940) );
  MAJIxp5_ASAP7_75t_SL U34045 ( .A(n23346), .B(mult_x_1196_n2153), .C(
        mult_x_1196_n2278), .Y(n23066) );
  XOR2xp5_ASAP7_75t_SL U34046 ( .A(mult_x_1196_n2335), .B(n23068), .Y(n23067)
         );
  MAJIxp5_ASAP7_75t_SL U34047 ( .A(mult_x_1196_n2512), .B(n23069), .C(
        mult_x_1196_n2640), .Y(mult_x_1196_n1538) );
  XNOR2xp5_ASAP7_75t_SL U34048 ( .A(n23656), .B(mult_x_1196_n2633), .Y(
        mult_x_1196_n2068) );
  MAJIxp5_ASAP7_75t_SL U34049 ( .A(mult_x_1196_n2137), .B(mult_x_1196_n2563), 
        .C(mult_x_1196_n2503), .Y(mult_x_1196_n2010) );
  XNOR2x1_ASAP7_75t_SL U34050 ( .A(n22423), .B(add_x_735_A_26_), .Y(n24033) );
  OAI22x1_ASAP7_75t_SL U34051 ( .A1(mult_x_1196_n3023), .A2(n24009), .B1(
        mult_x_1196_n3022), .B2(n23442), .Y(mult_x_1196_n2451) );
  INVx1_ASAP7_75t_SL U34052 ( .A(mult_x_1196_n1158), .Y(n23074) );
  XOR2xp5_ASAP7_75t_SL U34053 ( .A(mult_x_1196_n2086), .B(n23078), .Y(n23077)
         );
  NAND2xp5_ASAP7_75t_SL U34054 ( .A(n23159), .B(n23080), .Y(n23079) );
  INVx1_ASAP7_75t_SL U34055 ( .A(mult_x_1196_n3209), .Y(n23080) );
  INVx1_ASAP7_75t_SL U34056 ( .A(mult_x_1196_n1034), .Y(n23082) );
  XOR2xp5_ASAP7_75t_SL U34057 ( .A(mult_x_1196_n1034), .B(mult_x_1196_n2340), 
        .Y(n23083) );
  OAI21xp5_ASAP7_75t_SL U34058 ( .A1(mult_x_1196_n2880), .A2(n22464), .B(
        n23084), .Y(mult_x_1196_n1034) );
  NAND2xp5_ASAP7_75t_SL U34059 ( .A(n18536), .B(n23085), .Y(n23084) );
  INVx1_ASAP7_75t_SL U34060 ( .A(mult_x_1196_n2282), .Y(n23086) );
  XOR2xp5_ASAP7_75t_SL U34061 ( .A(n23087), .B(mult_x_1196_n995), .Y(n23668)
         );
  INVx1_ASAP7_75t_SL U34062 ( .A(mult_x_1196_n2338), .Y(n23087) );
  OAI22xp5_ASAP7_75t_SL U34063 ( .A1(mult_x_1196_n2910), .A2(n24022), .B1(
        mult_x_1196_n2909), .B2(n24020), .Y(mult_x_1196_n2338) );
  MAJx2_ASAP7_75t_SL U34064 ( .A(n23504), .B(mult_x_1196_n1510), .C(
        mult_x_1196_n1553), .Y(mult_x_1196_n1471) );
  XNOR2xp5_ASAP7_75t_SL U34065 ( .A(n18982), .B(n23720), .Y(n23088) );
  MAJIxp5_ASAP7_75t_SL U34066 ( .A(mult_x_1196_n2478), .B(mult_x_1196_n1323), 
        .C(n23874), .Y(mult_x_1196_n1318) );
  INVx1_ASAP7_75t_SL U34067 ( .A(mult_x_1196_n1840), .Y(n23090) );
  MAJIxp5_ASAP7_75t_SL U34068 ( .A(n23093), .B(mult_x_1196_n1579), .C(n22652), 
        .Y(mult_x_1196_n1580) );
  XNOR2xp5_ASAP7_75t_SL U34069 ( .A(n23092), .B(n23093), .Y(mult_x_1196_n1581)
         );
  XOR2xp5_ASAP7_75t_SL U34070 ( .A(n23466), .B(n23937), .Y(n23094) );
  MAJIxp5_ASAP7_75t_SL U34071 ( .A(mult_x_1196_n1554), .B(mult_x_1196_n1586), 
        .C(n23752), .Y(n23937) );
  NAND2xp5_ASAP7_75t_SL U34072 ( .A(n23099), .B(n23098), .Y(n23097) );
  INVx1_ASAP7_75t_SL U34073 ( .A(n24002), .Y(n23099) );
  OAI22xp5_ASAP7_75t_SL U34074 ( .A1(n18654), .A2(mult_x_1196_n3085), .B1(
        n22756), .B2(mult_x_1196_n3084), .Y(mult_x_1196_n2510) );
  OAI22xp5_ASAP7_75t_SL U34075 ( .A1(n23100), .A2(mult_x_1196_n3088), .B1(
        n22756), .B2(mult_x_1196_n3087), .Y(mult_x_1196_n2512) );
  OAI22xp5_ASAP7_75t_SL U34076 ( .A1(n18920), .A2(mult_x_1196_n3105), .B1(
        n24002), .B2(mult_x_1196_n3104), .Y(mult_x_1196_n2529) );
  OAI22xp5_ASAP7_75t_SL U34077 ( .A1(n18919), .A2(mult_x_1196_n3103), .B1(
        n22756), .B2(mult_x_1196_n3102), .Y(mult_x_1196_n2527) );
  OAI22xp5_ASAP7_75t_SL U34078 ( .A1(n23100), .A2(mult_x_1196_n3104), .B1(
        n24002), .B2(mult_x_1196_n3103), .Y(mult_x_1196_n2528) );
  OAI22xp5_ASAP7_75t_SL U34079 ( .A1(n18654), .A2(mult_x_1196_n3106), .B1(
        n22756), .B2(mult_x_1196_n3105), .Y(n23544) );
  XNOR2xp5_ASAP7_75t_SL U34080 ( .A(mult_x_1196_n1142), .B(mult_x_1196_n1167), 
        .Y(n23101) );
  INVx1_ASAP7_75t_SL U34081 ( .A(n23533), .Y(n23106) );
  MAJIxp5_ASAP7_75t_SL U34082 ( .A(mult_x_1196_n1129), .B(mult_x_1196_n1127), 
        .C(n23111), .Y(mult_x_1196_n1119) );
  INVx1_ASAP7_75t_SL U34083 ( .A(mult_x_1196_n1152), .Y(n23111) );
  OAI22xp33_ASAP7_75t_SL U34084 ( .A1(n22493), .A2(n24026), .B1(n24025), .B2(
        mult_x_1196_n2906), .Y(mult_x_1196_n2132) );
  INVx1_ASAP7_75t_SL U34085 ( .A(n23119), .Y(n23117) );
  XNOR2xp5_ASAP7_75t_SL U34086 ( .A(mult_x_1196_n2516), .B(n23119), .Y(n23118)
         );
  NOR2x1_ASAP7_75t_SL U34087 ( .A(n23121), .B(n23120), .Y(n23119) );
  NOR2x1_ASAP7_75t_SL U34088 ( .A(n22389), .B(mult_x_1196_n3251), .Y(n23121)
         );
  XNOR2xp5_ASAP7_75t_SL U34089 ( .A(mult_x_1196_n1496), .B(mult_x_1196_n1500), 
        .Y(n23122) );
  MAJIxp5_ASAP7_75t_SL U34090 ( .A(mult_x_1196_n2233), .B(mult_x_1196_n2172), 
        .C(n24227), .Y(mult_x_1196_n1496) );
  INVx1_ASAP7_75t_SL U34091 ( .A(n23129), .Y(n23128) );
  NOR2xp33_ASAP7_75t_SL U34092 ( .A(mult_x_1196_n3034), .B(n24008), .Y(n23131)
         );
  INVx1_ASAP7_75t_SL U34093 ( .A(mult_x_1196_n1805), .Y(n23132) );
  OAI21xp5_ASAP7_75t_SL U34094 ( .A1(mult_x_1196_n2765), .A2(n24041), .B(
        n22282), .Y(n23322) );
  MAJIxp5_ASAP7_75t_SL U34095 ( .A(mult_x_1196_n2398), .B(n23136), .C(
        mult_x_1196_n2554), .Y(mult_x_1196_n1835) );
  XNOR2xp5_ASAP7_75t_SL U34096 ( .A(n23136), .B(mult_x_1196_n2398), .Y(n23135)
         );
  XNOR2xp5_ASAP7_75t_SL U34097 ( .A(n23139), .B(n23138), .Y(mult_x_1196_n1353)
         );
  NOR2x1_ASAP7_75t_SL U34098 ( .A(n24030), .B(mult_x_1196_n2858), .Y(n23140)
         );
  XNOR2x1_ASAP7_75t_SL U34099 ( .A(n23144), .B(add_x_735_A_20_), .Y(n23143) );
  INVx1_ASAP7_75t_SL U34100 ( .A(u0_0_leon3x0_p0_muli[46]), .Y(n23144) );
  OAI21xp5_ASAP7_75t_SL U34101 ( .A1(n24168), .A2(n24206), .B(n23146), .Y(
        n23145) );
  OAI21xp5_ASAP7_75t_SL U34102 ( .A1(n24168), .A2(n24167), .B(n23147), .Y(
        n23146) );
  INVx1_ASAP7_75t_SL U34103 ( .A(mult_x_1196_n2154), .Y(n23147) );
  NOR2x1_ASAP7_75t_SL U34104 ( .A(n24025), .B(mult_x_1196_n2876), .Y(n24167)
         );
  NOR2x1_ASAP7_75t_SL U34105 ( .A(mult_x_1196_n2877), .B(n23708), .Y(n24168)
         );
  MAJIxp5_ASAP7_75t_SL U34106 ( .A(mult_x_1196_n1484), .B(mult_x_1196_n1486), 
        .C(n23918), .Y(mult_x_1196_n1476) );
  MAJIxp5_ASAP7_75t_SL U34107 ( .A(n22589), .B(mult_x_1196_n1535), .C(
        mult_x_1196_n1537), .Y(n23918) );
  XNOR2xp5_ASAP7_75t_SL U34108 ( .A(mult_x_1196_n1534), .B(mult_x_1196_n1536), 
        .Y(n23149) );
  MAJIxp5_ASAP7_75t_SL U34109 ( .A(n23150), .B(mult_x_1196_n2257), .C(
        mult_x_1196_n2196), .Y(mult_x_1196_n1222) );
  INVx1_ASAP7_75t_SL U34110 ( .A(mult_x_1196_n1255), .Y(n23150) );
  NOR2x1_ASAP7_75t_SL U34111 ( .A(n24002), .B(mult_x_1196_n3079), .Y(n23151)
         );
  NOR2x1_ASAP7_75t_SL U34112 ( .A(n18920), .B(mult_x_1196_n3080), .Y(n23152)
         );
  OAI21xp5_ASAP7_75t_SL U34113 ( .A1(mult_x_1196_n3193), .A2(n23522), .B(
        n23157), .Y(n23156) );
  INVx1_ASAP7_75t_SL U34114 ( .A(mult_x_1196_n905), .Y(mult_x_1196_n902) );
  NOR2xp33_ASAP7_75t_SL U34115 ( .A(n22999), .B(n23161), .Y(n31671) );
  XOR2xp5_ASAP7_75t_SL U34116 ( .A(n23968), .B(n28848), .Y(mult_x_1196_n3320)
         );
  NAND2xp5_ASAP7_75t_SL U34117 ( .A(n23161), .B(u0_0_leon3x0_p0_divi[19]), .Y(
        add_x_735_n142) );
  NOR2x1p5_ASAP7_75t_SL U34118 ( .A(n23569), .B(n23568), .Y(n28848) );
  XNOR2xp5_ASAP7_75t_SL U34119 ( .A(mult_x_1196_n2686), .B(mult_x_1196_n2526), 
        .Y(n24218) );
  AND2x2_ASAP7_75t_SL U34120 ( .A(n22278), .B(n25109), .Y(n25491) );
  NAND2xp5_ASAP7_75t_SL U34121 ( .A(n22556), .B(u0_0_leon3x0_p0_divi[25]), .Y(
        add_x_735_n86) );
  O2A1O1Ixp33_ASAP7_75t_SL U34122 ( .A1(n23164), .A2(n25198), .B(n25197), .C(
        n28850), .Y(n25202) );
  AOI21x1_ASAP7_75t_SL U34123 ( .A1(mult_x_1196_n815), .A2(mult_x_1196_n664), 
        .B(mult_x_1196_n657), .Y(mult_x_1196_n655) );
  OR2x2_ASAP7_75t_SL U34124 ( .A(n23260), .B(mult_x_1196_n1581), .Y(n23166) );
  OAI21x1_ASAP7_75t_SL U34125 ( .A1(mult_x_1196_n602), .A2(n23166), .B(
        mult_x_1196_n603), .Y(mult_x_1196_n597) );
  NAND2xp5_ASAP7_75t_SL U34126 ( .A(n23165), .B(mult_x_1196_n807), .Y(
        mult_x_1196_n257) );
  MAJIxp5_ASAP7_75t_SL U34127 ( .A(mult_x_1196_n2059), .B(n18863), .C(n23168), 
        .Y(mult_x_1196_n2050) );
  OAI22xp5_ASAP7_75t_SL U34128 ( .A1(mult_x_1196_n3270), .A2(n23982), .B1(
        n22389), .B2(mult_x_1196_n3269), .Y(n23168) );
  MAJIxp5_ASAP7_75t_SL U34129 ( .A(n22289), .B(mult_x_1196_n2155), .C(n23170), 
        .Y(mult_x_1196_n989) );
  INVx1_ASAP7_75t_SL U34130 ( .A(n23172), .Y(n23170) );
  XNOR2xp5_ASAP7_75t_SL U34131 ( .A(n23171), .B(n22289), .Y(mult_x_1196_n990)
         );
  XNOR2xp5_ASAP7_75t_SL U34132 ( .A(mult_x_1196_n2155), .B(n23172), .Y(n23171)
         );
  INVx1_ASAP7_75t_SL U34133 ( .A(mult_x_1196_n1161), .Y(n23175) );
  MAJIxp5_ASAP7_75t_SL U34134 ( .A(n23500), .B(mult_x_1196_n2692), .C(
        mult_x_1196_n2040), .Y(n23182) );
  NOR2x1_ASAP7_75t_SL U34135 ( .A(n23176), .B(n23597), .Y(mult_x_1196_n2040)
         );
  INVx1_ASAP7_75t_SL U34136 ( .A(mult_x_1196_n2693), .Y(n23176) );
  MAJIxp5_ASAP7_75t_SL U34137 ( .A(n23182), .B(n24265), .C(n23177), .Y(
        mult_x_1196_n2008) );
  INVx1_ASAP7_75t_SL U34138 ( .A(n23179), .Y(n23177) );
  AOI21x1_ASAP7_75t_SL U34139 ( .A1(n24241), .A2(n23181), .B(n23180), .Y(
        n23179) );
  NOR2x1p5_ASAP7_75t_SL U34140 ( .A(mult_x_1196_n2628), .B(mult_x_1196_n2504), 
        .Y(n23180) );
  OAI22x1_ASAP7_75t_SL U34141 ( .A1(mult_x_1196_n3203), .A2(n22248), .B1(
        n23072), .B2(mult_x_1196_n3204), .Y(mult_x_1196_n2628) );
  NAND2x2_ASAP7_75t_SL U34142 ( .A(n23571), .B(n23570), .Y(n24107) );
  INVx3_ASAP7_75t_SL U34143 ( .A(n23757), .Y(n23987) );
  MAJIxp5_ASAP7_75t_SL U34144 ( .A(mult_x_1196_n1637), .B(mult_x_1196_n1641), 
        .C(n22344), .Y(mult_x_1196_n1627) );
  XOR2xp5_ASAP7_75t_SL U34145 ( .A(mult_x_1196_n1641), .B(n22344), .Y(n23184)
         );
  OAI22x1_ASAP7_75t_SL U34146 ( .A1(mult_x_1196_n2894), .A2(n24026), .B1(
        n24025), .B2(mult_x_1196_n2893), .Y(n23185) );
  MAJIxp5_ASAP7_75t_SL U34147 ( .A(mult_x_1196_n2624), .B(mult_x_1196_n2436), 
        .C(n23186), .Y(mult_x_1196_n1964) );
  INVx1_ASAP7_75t_SL U34148 ( .A(n23188), .Y(n23186) );
  XNOR2xp5_ASAP7_75t_SL U34149 ( .A(mult_x_1196_n2624), .B(n23187), .Y(
        mult_x_1196_n1965) );
  XOR2xp5_ASAP7_75t_SL U34150 ( .A(n23190), .B(mult_x_1196_n1168), .Y(
        mult_x_1196_n1166) );
  XNOR2xp5_ASAP7_75t_SL U34151 ( .A(n22341), .B(mult_x_1196_n1197), .Y(n23190)
         );
  MAJIxp5_ASAP7_75t_SL U34152 ( .A(mult_x_1196_n1870), .B(n18937), .C(
        mult_x_1196_n1847), .Y(mult_x_1196_n1844) );
  XOR2xp5_ASAP7_75t_SL U34153 ( .A(mult_x_1196_n1847), .B(n23191), .Y(
        mult_x_1196_n1845) );
  XNOR2xp5_ASAP7_75t_SL U34154 ( .A(n22335), .B(mult_x_1196_n1870), .Y(n23191)
         );
  OAI21xp33_ASAP7_75t_SL U34155 ( .A1(mult_x_1196_n3254), .A2(n23981), .B(
        n23193), .Y(n23192) );
  INVxp67_ASAP7_75t_SL U34156 ( .A(mult_x_1196_n3253), .Y(n23194) );
  XNOR2xp5_ASAP7_75t_SL U34157 ( .A(mult_x_1196_n2635), .B(n23198), .Y(
        mult_x_1196_n2087) );
  INVx1_ASAP7_75t_SL U34158 ( .A(mult_x_1196_n2699), .Y(n23198) );
  XNOR2xp5_ASAP7_75t_SL U34159 ( .A(n23199), .B(n23580), .Y(n23579) );
  XNOR2xp5_ASAP7_75t_SL U34160 ( .A(n23200), .B(mult_x_1196_n2253), .Y(
        mult_x_1196_n1104) );
  OAI21xp5_ASAP7_75t_SL U34161 ( .A1(mult_x_1196_n2755), .A2(n24041), .B(
        n22281), .Y(n23201) );
  XNOR2xp5_ASAP7_75t_SL U34162 ( .A(mult_x_1196_n1222), .B(n23203), .Y(n23202)
         );
  INVx1_ASAP7_75t_SL U34163 ( .A(mult_x_1196_n1216), .Y(n23203) );
  MAJIxp5_ASAP7_75t_SL U34164 ( .A(mult_x_1196_n1877), .B(mult_x_1196_n1879), 
        .C(n23204), .Y(mult_x_1196_n1870) );
  INVx1_ASAP7_75t_SL U34165 ( .A(n23271), .Y(n23205) );
  NOR2x1_ASAP7_75t_SL U34166 ( .A(n23207), .B(n23206), .Y(n23271) );
  NAND3xp33_ASAP7_75t_SL U34167 ( .A(mult_x_1196_n359), .B(n18437), .C(n22584), 
        .Y(n23208) );
  AOI21xp5_ASAP7_75t_SL U34168 ( .A1(mult_x_1196_n360), .A2(n18437), .B(n23210), .Y(n23209) );
  NAND4xp25_ASAP7_75t_SL U34169 ( .A(n23230), .B(mult_x_1196_n359), .C(n18437), 
        .D(n23215), .Y(n23214) );
  MAJIxp5_ASAP7_75t_SL U34170 ( .A(n24295), .B(mult_x_1196_n1684), .C(
        mult_x_1196_n1721), .Y(mult_x_1196_n1685) );
  XNOR2xp5_ASAP7_75t_SL U34171 ( .A(n22827), .B(n23216), .Y(mult_x_1196_n1686)
         );
  XOR2xp5_ASAP7_75t_SL U34172 ( .A(mult_x_1196_n1684), .B(n24295), .Y(n23216)
         );
  INVx1_ASAP7_75t_SL U34173 ( .A(mult_x_1196_n2677), .Y(n23217) );
  OAI22xp5_ASAP7_75t_SL U34174 ( .A1(mult_x_1196_n3253), .A2(n23981), .B1(
        n22389), .B2(mult_x_1196_n3252), .Y(mult_x_1196_n2677) );
  NAND2xp5_ASAP7_75t_SL U34175 ( .A(n25305), .B(n23220), .Y(n23219) );
  NAND2xp5_ASAP7_75t_SL U34176 ( .A(n23225), .B(n23228), .Y(n23220) );
  INVx1_ASAP7_75t_SL U34177 ( .A(n23226), .Y(n23221) );
  NAND3xp33_ASAP7_75t_SL U34178 ( .A(n23230), .B(mult_x_1196_n411), .C(n23228), 
        .Y(n23227) );
  AND2x2_ASAP7_75t_SL U34179 ( .A(n23229), .B(n22367), .Y(n23228) );
  NAND2xp5_ASAP7_75t_SL U34180 ( .A(n23235), .B(n23232), .Y(n23237) );
  AOI31xp33_ASAP7_75t_SL U34181 ( .A1(n23232), .A2(n23235), .A3(n23231), .B(
        n25318), .Y(n23233) );
  NAND3xp33_ASAP7_75t_SL U34182 ( .A(n22361), .B(n23682), .C(n23681), .Y(
        n23232) );
  OAI211xp5_ASAP7_75t_SL U34183 ( .A1(n23600), .A2(n23601), .B(n23234), .C(
        n23233), .Y(n4189) );
  NAND2xp5_ASAP7_75t_SL U34184 ( .A(mult_x_1196_n323), .B(mult_x_1196_n324), 
        .Y(n23235) );
  MAJIxp5_ASAP7_75t_SL U34185 ( .A(n23542), .B(mult_x_1196_n1860), .C(
        mult_x_1196_n1864), .Y(mult_x_1196_n1852) );
  OAI21xp5_ASAP7_75t_SL U34186 ( .A1(n23936), .A2(n23141), .B(n22290), .Y(
        mult_x_1196_n2134) );
  AND2x2_ASAP7_75t_SL U34187 ( .A(mult_x_1196_n1868), .B(mult_x_1196_n1845), 
        .Y(mult_x_1196_n664) );
  MAJIxp5_ASAP7_75t_SL U34188 ( .A(n23342), .B(n23512), .C(n23339), .Y(n23238)
         );
  MAJIxp5_ASAP7_75t_SL U34189 ( .A(n23241), .B(n18915), .C(n23240), .Y(
        mult_x_1196_n1447) );
  XNOR2xp5_ASAP7_75t_SL U34190 ( .A(n23241), .B(n23239), .Y(mult_x_1196_n1448)
         );
  XOR2xp5_ASAP7_75t_SL U34191 ( .A(mult_x_1196_n1475), .B(n23243), .Y(n23242)
         );
  MAJIxp5_ASAP7_75t_SL U34192 ( .A(mult_x_1196_n1548), .B(mult_x_1196_n1517), 
        .C(n23471), .Y(n23243) );
  MAJIxp5_ASAP7_75t_SL U34193 ( .A(n23244), .B(mult_x_1196_n2368), .C(
        mult_x_1196_n2652), .Y(mult_x_1196_n1884) );
  XNOR2xp5_ASAP7_75t_SL U34194 ( .A(mult_x_1196_n881), .B(n23245), .Y(
        mult_x_1196_n870) );
  NAND2xp5_ASAP7_75t_SL U34195 ( .A(mult_x_1196_n2142), .B(n23247), .Y(
        mult_x_1196_n765) );
  INVx1_ASAP7_75t_SL U34196 ( .A(mult_x_1196_n770), .Y(n23246) );
  NAND2xp5_ASAP7_75t_SL U34197 ( .A(mult_x_1196_n2670), .B(mult_x_1196_n2702), 
        .Y(mult_x_1196_n770) );
  AND2x2_ASAP7_75t_SL U34198 ( .A(mult_x_1196_n2703), .B(mult_x_1196_n2143), 
        .Y(mult_x_1196_n771) );
  NOR2x1_ASAP7_75t_SL U34199 ( .A(mult_x_1196_n2142), .B(n23247), .Y(
        mult_x_1196_n764) );
  XNOR2xp5_ASAP7_75t_SL U34200 ( .A(n23248), .B(mult_x_1196_n2669), .Y(n23247)
         );
  OAI22xp5_ASAP7_75t_SL U34201 ( .A1(n24080), .A2(mult_x_1196_n3245), .B1(
        mult_x_1196_n3244), .B2(n23984), .Y(mult_x_1196_n2669) );
  INVx1_ASAP7_75t_SL U34202 ( .A(mult_x_1196_n2701), .Y(n23248) );
  OAI22xp5_ASAP7_75t_SL U34203 ( .A1(mult_x_1196_n3277), .A2(n23982), .B1(
        n23980), .B2(mult_x_1196_n3276), .Y(mult_x_1196_n2701) );
  INVx1_ASAP7_75t_SL U34204 ( .A(n23666), .Y(n23665) );
  XNOR2x1_ASAP7_75t_SL U34205 ( .A(n26683), .B(n23966), .Y(n24237) );
  INVx1_ASAP7_75t_SL U34206 ( .A(n23249), .Y(mult_x_1196_n335) );
  OAI21xp5_ASAP7_75t_SL U34207 ( .A1(n22214), .A2(n22407), .B(mult_x_1196_n339), .Y(n23249) );
  NAND2xp5_ASAP7_75t_SL U34208 ( .A(n22313), .B(mult_x_1196_n877), .Y(
        mult_x_1196_n348) );
  INVx1_ASAP7_75t_SL U34209 ( .A(mult_x_1196_n890), .Y(mult_x_1196_n877) );
  OR2x2_ASAP7_75t_SL U34210 ( .A(mult_x_1196_n904), .B(mult_x_1196_n891), .Y(
        mult_x_1196_n355) );
  A2O1A1Ixp33_ASAP7_75t_SL U34211 ( .A1(n24136), .A2(mult_x_1196_n2141), .B(
        mult_x_1196_n2087), .C(n23252), .Y(mult_x_1196_n2084) );
  NAND2xp5_ASAP7_75t_SL U34212 ( .A(n23253), .B(n24135), .Y(n23252) );
  OAI21xp5_ASAP7_75t_SL U34213 ( .A1(n23522), .A2(n18314), .B(n22316), .Y(
        mult_x_1196_n2141) );
  XOR2xp5_ASAP7_75t_SL U34214 ( .A(n23254), .B(mult_x_1196_n2342), .Y(
        mult_x_1196_n1074) );
  XNOR2xp5_ASAP7_75t_SL U34215 ( .A(n23255), .B(mult_x_1196_n2374), .Y(n23254)
         );
  OAI21xp5_ASAP7_75t_SL U34216 ( .A1(mult_x_1196_n2754), .A2(n24041), .B(
        n22280), .Y(n23255) );
  XNOR2xp5_ASAP7_75t_SL U34217 ( .A(n23257), .B(mult_x_1196_n2631), .Y(
        mult_x_1196_n2060) );
  NOR2xp33_ASAP7_75t_SL U34218 ( .A(mult_x_1196_n3271), .B(n23981), .Y(n23258)
         );
  INVx1_ASAP7_75t_SL U34219 ( .A(mult_x_1196_n1581), .Y(mult_x_1196_n1577) );
  INVx1_ASAP7_75t_SL U34220 ( .A(mult_x_1196_n1578), .Y(n23260) );
  AO21x1_ASAP7_75t_SL U34221 ( .A1(n22355), .A2(mult_x_1196_n1620), .B(n23801), 
        .Y(mult_x_1196_n1578) );
  XNOR2xp5_ASAP7_75t_SL U34222 ( .A(n23864), .B(mult_x_1196_n1152), .Y(n23261)
         );
  OR2x2_ASAP7_75t_SL U34223 ( .A(mult_x_1196_n1058), .B(mult_x_1196_n1037), 
        .Y(n23574) );
  INVx1_ASAP7_75t_SL U34224 ( .A(n23574), .Y(mult_x_1196_n457) );
  INVx1_ASAP7_75t_SL U34225 ( .A(n24121), .Y(n23262) );
  NAND2xp5_ASAP7_75t_SL U34226 ( .A(n22663), .B(n18514), .Y(mult_x_1196_n495)
         );
  XOR2xp5_ASAP7_75t_SL U34227 ( .A(mult_x_1196_n2506), .B(n23265), .Y(n23655)
         );
  AO21x1_ASAP7_75t_SL U34228 ( .A1(n23266), .A2(mult_x_1196_n1520), .B(n22329), 
        .Y(n23269) );
  AND2x2_ASAP7_75t_SL U34229 ( .A(n23747), .B(n24109), .Y(n24001) );
  INVx1_ASAP7_75t_SL U34230 ( .A(mult_x_1196_n2465), .Y(n23270) );
  XOR2xp5_ASAP7_75t_SL U34231 ( .A(n23274), .B(mult_x_1196_n2277), .Y(
        mult_x_1196_n943) );
  XNOR2xp5_ASAP7_75t_SL U34232 ( .A(n23275), .B(mult_x_1196_n2152), .Y(n23274)
         );
  OAI22xp5_ASAP7_75t_SL U34233 ( .A1(mult_x_1196_n2875), .A2(n22464), .B1(
        mult_x_1196_n2874), .B2(n18305), .Y(n23275) );
  MAJIxp5_ASAP7_75t_SL U34234 ( .A(n23793), .B(mult_x_1196_n2468), .C(n23276), 
        .Y(mult_x_1196_n1962) );
  INVx1_ASAP7_75t_SL U34235 ( .A(n23792), .Y(n23276) );
  MAJIxp5_ASAP7_75t_SL U34236 ( .A(n23278), .B(mult_x_1196_n1190), .C(
        mult_x_1196_n2288), .Y(mult_x_1196_n1185) );
  INVx1_ASAP7_75t_SL U34237 ( .A(n23280), .Y(n23278) );
  XNOR2xp5_ASAP7_75t_SL U34238 ( .A(mult_x_1196_n2288), .B(n23279), .Y(
        mult_x_1196_n1186) );
  XNOR2xp5_ASAP7_75t_SL U34239 ( .A(n23280), .B(mult_x_1196_n1190), .Y(n23279)
         );
  NOR2x1_ASAP7_75t_SL U34240 ( .A(n23282), .B(n23281), .Y(n23280) );
  NOR2x1_ASAP7_75t_SL U34241 ( .A(mult_x_1196_n2790), .B(n24039), .Y(n23281)
         );
  NOR2x1_ASAP7_75t_SL U34242 ( .A(mult_x_1196_n2789), .B(n22391), .Y(n23282)
         );
  MAJIxp5_ASAP7_75t_SL U34243 ( .A(n23633), .B(n23632), .C(n23631), .Y(
        mult_x_1196_n1552) );
  MAJIxp5_ASAP7_75t_SL U34244 ( .A(n24094), .B(mult_x_1196_n2190), .C(
        mult_x_1196_n2251), .Y(n23284) );
  OAI21x1_ASAP7_75t_SL U34245 ( .A1(mult_x_1196_n3255), .A2(n23981), .B(n22295), .Y(mult_x_1196_n2679) );
  MAJIxp5_ASAP7_75t_SL U34246 ( .A(n23286), .B(mult_x_1196_n2344), .C(
        mult_x_1196_n2286), .Y(mult_x_1196_n1126) );
  XNOR2xp5_ASAP7_75t_SL U34247 ( .A(n23286), .B(mult_x_1196_n2344), .Y(n23285)
         );
  INVx1_ASAP7_75t_SL U34248 ( .A(mult_x_1196_n2286), .Y(n23287) );
  NAND2xp5_ASAP7_75t_SL U34249 ( .A(n23291), .B(n23290), .Y(n23289) );
  MAJIxp5_ASAP7_75t_SL U34250 ( .A(mult_x_1196_n1753), .B(n22342), .C(n23292), 
        .Y(mult_x_1196_n1747) );
  XOR2xp5_ASAP7_75t_SL U34251 ( .A(n18924), .B(n23293), .Y(mult_x_1196_n1748)
         );
  MAJIxp5_ASAP7_75t_SL U34252 ( .A(n23860), .B(n18916), .C(n23859), .Y(n23292)
         );
  MAJIxp5_ASAP7_75t_SL U34253 ( .A(mult_x_1196_n1247), .B(mult_x_1196_n1251), 
        .C(n24274), .Y(mult_x_1196_n1239) );
  MAJx2_ASAP7_75t_SL U34254 ( .A(mult_x_1196_n1316), .B(n18547), .C(
        mult_x_1196_n1320), .Y(n24274) );
  INVx1_ASAP7_75t_SL U34255 ( .A(mult_x_1196_n2318), .Y(n23295) );
  MAJIxp5_ASAP7_75t_SL U34256 ( .A(n23297), .B(mult_x_1196_n1442), .C(
        mult_x_1196_n1439), .Y(mult_x_1196_n1400) );
  INVx1_ASAP7_75t_SL U34257 ( .A(mult_x_1196_n1423), .Y(n23299) );
  MAJIxp5_ASAP7_75t_SL U34258 ( .A(mult_x_1196_n2370), .B(n23414), .C(n23300), 
        .Y(mult_x_1196_n993) );
  INVx1_ASAP7_75t_SL U34259 ( .A(n23301), .Y(n23300) );
  XOR2xp5_ASAP7_75t_SL U34260 ( .A(n23301), .B(n23412), .Y(mult_x_1196_n994)
         );
  MAJIxp5_ASAP7_75t_SL U34261 ( .A(mult_x_1196_n1983), .B(mult_x_1196_n1995), 
        .C(n23303), .Y(mult_x_1196_n1975) );
  XNOR2xp5_ASAP7_75t_SL U34262 ( .A(n18391), .B(n23302), .Y(mult_x_1196_n1976)
         );
  XOR2xp5_ASAP7_75t_SL U34263 ( .A(mult_x_1196_n1995), .B(mult_x_1196_n1983), 
        .Y(n23302) );
  MAJIxp5_ASAP7_75t_SL U34264 ( .A(n22297), .B(n23544), .C(mult_x_1196_n2690), 
        .Y(n23303) );
  AOI21xp5_ASAP7_75t_SL U34265 ( .A1(n18319), .A2(n22389), .B(
        mult_x_1196_n3247), .Y(n24255) );
  INVx1_ASAP7_75t_SL U34266 ( .A(n23799), .Y(n23305) );
  XNOR2xp5_ASAP7_75t_SL U34267 ( .A(mult_x_1196_n1385), .B(mult_x_1196_n1379), 
        .Y(n23307) );
  OAI22x1_ASAP7_75t_SL U34268 ( .A1(mult_x_1196_n3115), .A2(n23997), .B1(
        mult_x_1196_n3116), .B2(n23999), .Y(mult_x_1196_n2540) );
  XNOR2xp5_ASAP7_75t_SL U34269 ( .A(n23954), .B(n23310), .Y(mult_x_1196_n3228)
         );
  INVx1_ASAP7_75t_SL U34270 ( .A(n24059), .Y(n23310) );
  BUFx12f_ASAP7_75t_SL U34271 ( .A(n24013), .Y(n23311) );
  OAI22xp5_ASAP7_75t_SL U34272 ( .A1(mult_x_1196_n2980), .A2(n24012), .B1(
        n24014), .B2(mult_x_1196_n2981), .Y(mult_x_1196_n2409) );
  OAI22xp5_ASAP7_75t_SL U34273 ( .A1(mult_x_1196_n2979), .A2(n24012), .B1(
        n24014), .B2(mult_x_1196_n2980), .Y(mult_x_1196_n2408) );
  OAI22xp5_ASAP7_75t_SL U34274 ( .A1(mult_x_1196_n3008), .A2(n18308), .B1(
        n18442), .B2(n22216), .Y(mult_x_1196_n2135) );
  OAI22xp5_ASAP7_75t_SL U34275 ( .A1(mult_x_1196_n2978), .A2(n24012), .B1(
        n24014), .B2(mult_x_1196_n2979), .Y(mult_x_1196_n2407) );
  AOI21xp5_ASAP7_75t_SL U34276 ( .A1(n18308), .A2(n18442), .B(
        mult_x_1196_n2975), .Y(n24253) );
  OAI22xp5_ASAP7_75t_SL U34277 ( .A1(mult_x_1196_n2975), .A2(n18308), .B1(
        n18442), .B2(mult_x_1196_n2976), .Y(mult_x_1196_n2404) );
  OAI22xp5_ASAP7_75t_SL U34278 ( .A1(mult_x_1196_n2977), .A2(n24012), .B1(
        n24014), .B2(mult_x_1196_n2978), .Y(mult_x_1196_n2406) );
  OAI21xp5_ASAP7_75t_SL U34279 ( .A1(mult_x_1196_n3000), .A2(n24014), .B(
        n22302), .Y(n23562) );
  OAI21xp5_ASAP7_75t_SL U34280 ( .A1(n24014), .A2(mult_x_1196_n2984), .B(
        n22303), .Y(n23718) );
  OAI21xp5_ASAP7_75t_SL U34281 ( .A1(n24014), .A2(mult_x_1196_n3003), .B(
        n24277), .Y(n23517) );
  NOR2x1_ASAP7_75t_SL U34282 ( .A(mult_x_1196_n2824), .B(n22251), .Y(n23313)
         );
  NAND2xp5_ASAP7_75t_SL U34283 ( .A(n23315), .B(n23314), .Y(n23317) );
  OAI21xp5_ASAP7_75t_SL U34284 ( .A1(n23316), .A2(n23318), .B(
        mult_x_1196_n1487), .Y(n23314) );
  NAND2xp5_ASAP7_75t_SL U34285 ( .A(n23316), .B(n23318), .Y(n23315) );
  INVx1_ASAP7_75t_SL U34286 ( .A(mult_x_1196_n1455), .Y(n23316) );
  INVx1_ASAP7_75t_SL U34287 ( .A(mult_x_1196_n1460), .Y(n23318) );
  MAJIxp5_ASAP7_75t_SL U34288 ( .A(n24211), .B(n23688), .C(n23322), .Y(
        mult_x_1196_n1424) );
  XOR2xp5_ASAP7_75t_SL U34289 ( .A(n23324), .B(mult_x_1196_n2564), .Y(n23323)
         );
  INVx1_ASAP7_75t_SL U34290 ( .A(mult_x_1196_n2596), .Y(n23324) );
  INVx1_ASAP7_75t_SL U34291 ( .A(mult_x_1196_n1757), .Y(n23326) );
  OR3x1_ASAP7_75t_SL U34292 ( .A(n22366), .B(mult_x_1196_n405), .C(n24646), 
        .Y(n23329) );
  XOR2xp5_ASAP7_75t_SL U34293 ( .A(mult_x_1196_n2268), .B(n23330), .Y(n24229)
         );
  XNOR2xp5_ASAP7_75t_SL U34294 ( .A(n23931), .B(n23331), .Y(mult_x_1196_n1674)
         );
  MAJIxp5_ASAP7_75t_SL U34295 ( .A(mult_x_1196_n2369), .B(n23334), .C(
        mult_x_1196_n2337), .Y(mult_x_1196_n971) );
  XNOR2xp5_ASAP7_75t_SL U34296 ( .A(n23334), .B(n23333), .Y(mult_x_1196_n972)
         );
  XOR2xp5_ASAP7_75t_SL U34297 ( .A(mult_x_1196_n2369), .B(mult_x_1196_n2337), 
        .Y(n23333) );
  NAND2xp5_ASAP7_75t_SL U34298 ( .A(mult_x_1196_n1610), .B(mult_x_1196_n1604), 
        .Y(n23335) );
  INVx3_ASAP7_75t_SL U34299 ( .A(n24001), .Y(n24003) );
  XNOR2x1_ASAP7_75t_SL U34300 ( .A(n24052), .B(n22394), .Y(mult_x_1196_n3085)
         );
  MAJIxp5_ASAP7_75t_SL U34301 ( .A(n23337), .B(mult_x_1196_n1441), .C(
        mult_x_1196_n1490), .Y(mult_x_1196_n1442) );
  NAND2xp5_ASAP7_75t_SL U34302 ( .A(mult_x_1196_n1357), .B(n23338), .Y(
        mult_x_1196_n558) );
  NOR2x1_ASAP7_75t_SL U34303 ( .A(n23338), .B(mult_x_1196_n1357), .Y(
        mult_x_1196_n557) );
  INVx1_ASAP7_75t_SL U34304 ( .A(mult_x_1196_n1754), .Y(n23339) );
  MAJIxp5_ASAP7_75t_SL U34305 ( .A(mult_x_1196_n1766), .B(mult_x_1196_n1762), 
        .C(n22253), .Y(mult_x_1196_n1754) );
  INVx1_ASAP7_75t_SL U34306 ( .A(mult_x_1196_n1756), .Y(n23342) );
  XOR2x2_ASAP7_75t_SL U34307 ( .A(n23343), .B(n23398), .Y(mult_x_1196_n1745)
         );
  XNOR2x1_ASAP7_75t_SL U34308 ( .A(n23344), .B(n23345), .Y(n24220) );
  INVx1_ASAP7_75t_SL U34309 ( .A(mult_x_1196_n1397), .Y(n23345) );
  INVx1_ASAP7_75t_SL U34310 ( .A(mult_x_1196_n960), .Y(n23346) );
  XNOR2xp5_ASAP7_75t_SL U34311 ( .A(mult_x_1196_n960), .B(n23347), .Y(
        mult_x_1196_n957) );
  MAJIxp5_ASAP7_75t_SL U34312 ( .A(mult_x_1196_n1611), .B(n24266), .C(n23350), 
        .Y(mult_x_1196_n1563) );
  XNOR2xp5_ASAP7_75t_SL U34313 ( .A(n24266), .B(mult_x_1196_n1611), .Y(n23348)
         );
  INVx1_ASAP7_75t_SL U34314 ( .A(n23350), .Y(n23349) );
  NAND2xp5_ASAP7_75t_SL U34315 ( .A(mult_x_1196_n2154), .B(n23353), .Y(n24206)
         );
  NAND2xp5_ASAP7_75t_SL U34316 ( .A(n23353), .B(n24207), .Y(n24169) );
  INVx1_ASAP7_75t_SL U34317 ( .A(n24167), .Y(n23353) );
  INVx1_ASAP7_75t_SL U34318 ( .A(n23355), .Y(n23354) );
  NAND2xp5_ASAP7_75t_SL U34319 ( .A(n23365), .B(u0_0_leon3x0_p0_divi[29]), .Y(
        add_x_735_n48) );
  NAND2xp5_ASAP7_75t_SL U34320 ( .A(n23360), .B(n29149), .Y(n29151) );
  NOR3xp33_ASAP7_75t_SL U34321 ( .A(n23365), .B(n29148), .C(n24631), .Y(n23361) );
  NOR3xp33_ASAP7_75t_SL U34322 ( .A(n25477), .B(n26155), .C(n23362), .Y(n25908) );
  NAND2xp5_ASAP7_75t_SL U34323 ( .A(n23363), .B(n29145), .Y(n29152) );
  INVx1_ASAP7_75t_SL U34324 ( .A(n18388), .Y(n23365) );
  INVx1_ASAP7_75t_SL U34325 ( .A(mult_x_1196_n1380), .Y(n23369) );
  NAND2xp5_ASAP7_75t_SL U34326 ( .A(mult_x_1196_n1531), .B(n24312), .Y(n23371)
         );
  XNOR2xp5_ASAP7_75t_SL U34327 ( .A(n24312), .B(mult_x_1196_n1531), .Y(n23372)
         );
  XNOR2xp5_ASAP7_75t_SL U34328 ( .A(mult_x_1196_n2133), .B(mult_x_1196_n1866), 
        .Y(n23602) );
  INVx2_ASAP7_75t_SL U34329 ( .A(mult_x_1196_n3327), .Y(n23374) );
  XNOR2x1_ASAP7_75t_SL U34330 ( .A(n23959), .B(n23375), .Y(mult_x_1196_n3327)
         );
  OAI22xp5_ASAP7_75t_SL U34331 ( .A1(n24691), .A2(n24031), .B1(n24029), .B2(
        mult_x_1196_n2872), .Y(n23380) );
  NAND2x1p5_ASAP7_75t_SL U34332 ( .A(n24120), .B(mult_x_1196_n3329), .Y(n23985) );
  XNOR2x1_ASAP7_75t_SL U34333 ( .A(add_x_735_A_4_), .B(n23381), .Y(
        mult_x_1196_n3329) );
  XNOR2x2_ASAP7_75t_SL U34334 ( .A(n23951), .B(u0_0_leon3x0_p0_muli[40]), .Y(
        n23983) );
  INVx1_ASAP7_75t_SL U34335 ( .A(u0_0_leon3x0_p0_muli[40]), .Y(n23381) );
  INVx1_ASAP7_75t_SL U34336 ( .A(mult_x_1196_n2577), .Y(n23382) );
  OAI22xp5_ASAP7_75t_SL U34337 ( .A1(n24035), .A2(mult_x_1196_n2833), .B1(
        n22251), .B2(mult_x_1196_n2832), .Y(n23384) );
  OAI21xp5_ASAP7_75t_SL U34338 ( .A1(mult_x_1196_n312), .A2(mult_x_1196_n390), 
        .B(mult_x_1196_n313), .Y(n23389) );
  NAND2xp5_ASAP7_75t_SL U34339 ( .A(n22409), .B(n23389), .Y(n23388) );
  NOR2x1_ASAP7_75t_SL U34340 ( .A(mult_x_1196_n301), .B(mult_x_1196_n387), .Y(
        n23391) );
  AOI21xp5_ASAP7_75t_SL U34341 ( .A1(n18932), .A2(mult_x_1196_n299), .B(n23392), .Y(mult_x_1196_n298) );
  NOR2x1_ASAP7_75t_SL U34342 ( .A(mult_x_1196_n301), .B(mult_x_1196_n308), .Y(
        mult_x_1196_n299) );
  XNOR2xp5_ASAP7_75t_SL U34343 ( .A(n22425), .B(n22961), .Y(mult_x_1196_n3050)
         );
  XNOR2xp5_ASAP7_75t_SL U34344 ( .A(n22961), .B(n23395), .Y(mult_x_1196_n3061)
         );
  INVx1_ASAP7_75t_SL U34345 ( .A(n24062), .Y(n23395) );
  XOR2xp5_ASAP7_75t_SL U34346 ( .A(n22961), .B(n24065), .Y(mult_x_1196_n3064)
         );
  XOR2xp5_ASAP7_75t_SL U34347 ( .A(n22961), .B(n24075), .Y(mult_x_1196_n3074)
         );
  XOR2xp5_ASAP7_75t_SL U34348 ( .A(n24045), .B(n22961), .Y(mult_x_1196_n3044)
         );
  XOR2xp5_ASAP7_75t_SL U34349 ( .A(n24070), .B(n22961), .Y(mult_x_1196_n3069)
         );
  XNOR2xp5_ASAP7_75t_SL U34350 ( .A(n24064), .B(n23396), .Y(mult_x_1196_n3063)
         );
  XNOR2xp5_ASAP7_75t_SL U34351 ( .A(n24057), .B(n23396), .Y(mult_x_1196_n3056)
         );
  BUFx6f_ASAP7_75t_SL U34352 ( .A(n23959), .Y(n23397) );
  XOR2xp5_ASAP7_75t_SL U34353 ( .A(n23397), .B(n24065), .Y(mult_x_1196_n3166)
         );
  XOR2xp5_ASAP7_75t_SL U34354 ( .A(n23397), .B(n24061), .Y(mult_x_1196_n3162)
         );
  XOR2xp5_ASAP7_75t_SL U34355 ( .A(u0_0_leon3x0_p0_muli[26]), .B(n23397), .Y(
        mult_x_1196_n3159) );
  XNOR2xp5_ASAP7_75t_SL U34356 ( .A(n24057), .B(n23960), .Y(mult_x_1196_n3158)
         );
  XNOR2xp5_ASAP7_75t_SL U34357 ( .A(n24060), .B(n18394), .Y(mult_x_1196_n3161)
         );
  INVx1_ASAP7_75t_SL U34358 ( .A(mult_x_1196_n1750), .Y(n23487) );
  NOR2x1_ASAP7_75t_SL U34359 ( .A(n18928), .B(mult_x_1196_n1745), .Y(n23927)
         );
  INVx1_ASAP7_75t_SL U34360 ( .A(n23402), .Y(n23400) );
  INVx1_ASAP7_75t_SL U34361 ( .A(mult_x_1196_n2599), .Y(n23401) );
  OAI21xp5_ASAP7_75t_SL U34362 ( .A1(mult_x_1196_n3143), .A2(n18397), .B(
        n22287), .Y(n23402) );
  INVx1_ASAP7_75t_SL U34363 ( .A(n23814), .Y(n23403) );
  MAJIxp5_ASAP7_75t_SL U34364 ( .A(mult_x_1196_n2170), .B(n23405), .C(
        mult_x_1196_n2510), .Y(mult_x_1196_n1422) );
  INVx1_ASAP7_75t_SL U34365 ( .A(mult_x_1196_n2510), .Y(n23406) );
  INVx1_ASAP7_75t_SL U34366 ( .A(mult_x_1196_n2343), .Y(n23407) );
  NAND2xp5_ASAP7_75t_SL U34367 ( .A(n22998), .B(n23410), .Y(n23409) );
  MAJIxp5_ASAP7_75t_SL U34368 ( .A(n24280), .B(mult_x_1196_n2451), .C(n22411), 
        .Y(n23411) );
  XNOR2xp5_ASAP7_75t_SL U34369 ( .A(n23414), .B(n23413), .Y(n23412) );
  NOR2x1_ASAP7_75t_SL U34370 ( .A(n24043), .B(mult_x_1196_n2736), .Y(
        mult_x_1196_n2127) );
  OA21x2_ASAP7_75t_SL U34371 ( .A1(n25207), .A2(n18910), .B(n23923), .Y(n23415) );
  NAND2xp5_ASAP7_75t_SL U34372 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__31_), .B(
        n18911), .Y(n23923) );
  INVx1_ASAP7_75t_SL U34373 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__31_), .Y(n25207)
         );
  OAI22xp5_ASAP7_75t_SL U34374 ( .A1(n24000), .A2(mult_x_1196_n3123), .B1(
        n23996), .B2(mult_x_1196_n3122), .Y(mult_x_1196_n2547) );
  OAI22xp5_ASAP7_75t_SL U34375 ( .A1(mult_x_1196_n3128), .A2(n24000), .B1(
        n23996), .B2(mult_x_1196_n3127), .Y(mult_x_1196_n2552) );
  OAI22xp5_ASAP7_75t_SL U34376 ( .A1(mult_x_1196_n3124), .A2(n23999), .B1(
        n23996), .B2(mult_x_1196_n3123), .Y(mult_x_1196_n2548) );
  OAI22xp5_ASAP7_75t_SL U34377 ( .A1(mult_x_1196_n3125), .A2(n18397), .B1(
        n23997), .B2(mult_x_1196_n3124), .Y(mult_x_1196_n2549) );
  MAJIxp5_ASAP7_75t_SL U34378 ( .A(n23817), .B(n23416), .C(mult_x_1196_n2301), 
        .Y(mult_x_1196_n1640) );
  INVx1_ASAP7_75t_SL U34379 ( .A(n23816), .Y(n23416) );
  NOR2x1_ASAP7_75t_SL U34380 ( .A(n23418), .B(n23417), .Y(n23816) );
  NOR2x1_ASAP7_75t_SL U34381 ( .A(mult_x_1196_n3059), .B(n24007), .Y(n23417)
         );
  NOR2x1_ASAP7_75t_SL U34382 ( .A(mult_x_1196_n3058), .B(n24005), .Y(n23418)
         );
  OAI22x1_ASAP7_75t_SL U34383 ( .A1(n23081), .A2(mult_x_1196_n3165), .B1(
        n23992), .B2(n23421), .Y(mult_x_1196_n2589) );
  INVx2_ASAP7_75t_SL U34384 ( .A(n25087), .Y(n23422) );
  NOR2xp67_ASAP7_75t_SL U34385 ( .A(n31475), .B(n24686), .Y(n23423) );
  XNOR2xp5_ASAP7_75t_SL U34386 ( .A(n23426), .B(n23425), .Y(mult_x_1196_n1245)
         );
  XOR2xp5_ASAP7_75t_SL U34387 ( .A(mult_x_1196_n1243), .B(mult_x_1196_n1285), 
        .Y(n23425) );
  OAI21xp5_ASAP7_75t_SL U34388 ( .A1(mult_x_1196_n1323), .A2(n24181), .B(
        n23428), .Y(n23427) );
  NAND2xp5_ASAP7_75t_SL U34389 ( .A(mult_x_1196_n1323), .B(n24181), .Y(n23429)
         );
  NOR2x1_ASAP7_75t_SL U34390 ( .A(n23855), .B(n23854), .Y(n24181) );
  NAND2x2_ASAP7_75t_SL U34391 ( .A(n23991), .B(n23431), .Y(n24287) );
  INVx2_ASAP7_75t_SL U34392 ( .A(n23374), .Y(n23431) );
  OAI21xp5_ASAP7_75t_SL U34393 ( .A1(mult_x_1196_n2000), .A2(n23437), .B(
        n23436), .Y(mult_x_1196_n1991) );
  NAND2xp5_ASAP7_75t_SL U34394 ( .A(n22320), .B(mult_x_1196_n2008), .Y(n23436)
         );
  XOR2xp5_ASAP7_75t_SL U34395 ( .A(n22320), .B(mult_x_1196_n2008), .Y(n23438)
         );
  XOR2xp5_ASAP7_75t_SL U34396 ( .A(n23440), .B(n22565), .Y(mult_x_1196_n1633)
         );
  XNOR2xp5_ASAP7_75t_SL U34397 ( .A(n24130), .B(n24129), .Y(n23439) );
  XNOR2xp5_ASAP7_75t_SL U34398 ( .A(mult_x_1196_n878), .B(mult_x_1196_n893), 
        .Y(n23441) );
  XNOR2x1_ASAP7_75t_SL U34399 ( .A(add_x_735_A_14_), .B(add_x_735_A_15_), .Y(
        n23444) );
  INVx1_ASAP7_75t_SL U34400 ( .A(n23444), .Y(n23443) );
  OAI22xp5_ASAP7_75t_SL U34401 ( .A1(mult_x_1196_n3028), .A2(n22815), .B1(
        mult_x_1196_n3027), .B2(n23442), .Y(mult_x_1196_n2456) );
  OAI22xp5_ASAP7_75t_SL U34402 ( .A1(mult_x_1196_n3021), .A2(n24009), .B1(
        mult_x_1196_n3020), .B2(n23442), .Y(mult_x_1196_n2449) );
  OAI22xp5_ASAP7_75t_SL U34403 ( .A1(mult_x_1196_n3022), .A2(n24009), .B1(
        mult_x_1196_n3021), .B2(n23442), .Y(mult_x_1196_n2450) );
  OAI22xp5_ASAP7_75t_SL U34404 ( .A1(mult_x_1196_n3024), .A2(n24009), .B1(
        mult_x_1196_n3023), .B2(n23442), .Y(mult_x_1196_n2452) );
  OAI22xp5_ASAP7_75t_SL U34405 ( .A1(mult_x_1196_n3027), .A2(n24009), .B1(
        mult_x_1196_n3026), .B2(n23442), .Y(mult_x_1196_n2455) );
  OAI22xp5_ASAP7_75t_SL U34406 ( .A1(mult_x_1196_n3026), .A2(n22815), .B1(
        mult_x_1196_n3025), .B2(n23442), .Y(mult_x_1196_n2454) );
  XNOR2xp5_ASAP7_75t_SL U34407 ( .A(n23446), .B(n23445), .Y(mult_x_1196_n1697)
         );
  XOR2xp5_ASAP7_75t_SL U34408 ( .A(mult_x_1196_n1735), .B(mult_x_1196_n1708), 
        .Y(n23445) );
  XNOR2xp5_ASAP7_75t_SL U34409 ( .A(n24162), .B(n24161), .Y(n23446) );
  XOR2x1_ASAP7_75t_SL U34410 ( .A(n24550), .B(n24693), .Y(n23990) );
  AND2x2_ASAP7_75t_SL U34411 ( .A(n25112), .B(n25113), .Y(n24550) );
  NAND2xp5_ASAP7_75t_SL U34412 ( .A(n23375), .B(u0_0_leon3x0_p0_divi[5]), .Y(
        add_x_735_n248) );
  NAND2xp5_ASAP7_75t_SL U34413 ( .A(mult_x_1196_n2061), .B(mult_x_1196_n2053), 
        .Y(mult_x_1196_n734) );
  INVx1_ASAP7_75t_SL U34414 ( .A(mult_x_1196_n1689), .Y(mult_x_1196_n1681) );
  INVxp33_ASAP7_75t_SL U34415 ( .A(mult_x_1196_n308), .Y(mult_x_1196_n306) );
  NAND2x2_ASAP7_75t_SL U34416 ( .A(n23474), .B(n23683), .Y(mult_x_1196_n312)
         );
  OAI22xp5_ASAP7_75t_SL U34417 ( .A1(mult_x_1196_n2862), .A2(n24031), .B1(
        n24030), .B2(mult_x_1196_n2861), .Y(n23814) );
  OAI22xp5_ASAP7_75t_SL U34418 ( .A1(mult_x_1196_n2850), .A2(n23449), .B1(
        mult_x_1196_n2849), .B2(n18390), .Y(mult_x_1196_n2284) );
  OAI22xp5_ASAP7_75t_SL U34419 ( .A1(mult_x_1196_n2867), .A2(n23449), .B1(
        n24030), .B2(mult_x_1196_n2866), .Y(mult_x_1196_n2301) );
  OAI22xp5_ASAP7_75t_SL U34420 ( .A1(mult_x_1196_n2848), .A2(n22780), .B1(
        n22743), .B2(mult_x_1196_n2847), .Y(mult_x_1196_n2282) );
  OAI22xp5_ASAP7_75t_SL U34421 ( .A1(mult_x_1196_n2847), .A2(n22780), .B1(
        n24030), .B2(mult_x_1196_n2846), .Y(mult_x_1196_n2281) );
  OAI22xp5_ASAP7_75t_SL U34422 ( .A1(mult_x_1196_n2846), .A2(n22780), .B1(
        n18346), .B2(mult_x_1196_n2845), .Y(mult_x_1196_n2280) );
  OAI22x1_ASAP7_75t_SL U34423 ( .A1(n18920), .A2(mult_x_1196_n3084), .B1(
        n22756), .B2(mult_x_1196_n3083), .Y(mult_x_1196_n1387) );
  OAI22x1_ASAP7_75t_SL U34424 ( .A1(n18920), .A2(mult_x_1196_n3089), .B1(
        mult_x_1196_n3088), .B2(n24002), .Y(mult_x_1196_n2513) );
  NOR2x1p5_ASAP7_75t_SL U34425 ( .A(mult_x_1196_n3119), .B(n23999), .Y(n23811)
         );
  OAI21x1_ASAP7_75t_SL U34426 ( .A1(mult_x_1196_n3036), .A2(n24009), .B(n24258), .Y(n24100) );
  INVx2_ASAP7_75t_SL U34427 ( .A(n24027), .Y(n23704) );
  NAND2x1p5_ASAP7_75t_SL U34428 ( .A(n24033), .B(mult_x_1196_n3317), .Y(
        mult_x_1196_n126) );
  BUFx6f_ASAP7_75t_SL U34429 ( .A(n24107), .Y(n23989) );
  AOI21xp5_ASAP7_75t_SL U34430 ( .A1(mult_x_1196_n386), .A2(n23769), .B(n23768), .Y(n23676) );
  NAND2x1_ASAP7_75t_SL U34431 ( .A(n23676), .B(n23675), .Y(mult_x_1196_n360)
         );
  AOI21x1_ASAP7_75t_SL U34432 ( .A1(mult_x_1196_n626), .A2(n24086), .B(n24289), 
        .Y(mult_x_1196_n617) );
  NOR2x1_ASAP7_75t_SL U34433 ( .A(mult_x_1196_n2734), .B(n24043), .Y(
        mult_x_1196_n2172) );
  OR2x6_ASAP7_75t_SL U34434 ( .A(n24028), .B(n24113), .Y(n24031) );
  NAND2xp5_ASAP7_75t_SL U34435 ( .A(n18910), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__5_), .Y(n25193) );
  BUFx6f_ASAP7_75t_SL U34436 ( .A(n24013), .Y(n24014) );
  NAND2xp5_ASAP7_75t_SL U34437 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__23_), .B(
        n22434), .Y(n25145) );
  BUFx6f_ASAP7_75t_SL U34438 ( .A(n23998), .Y(n23999) );
  AOI21x1_ASAP7_75t_SL U34439 ( .A1(mult_x_1196_n611), .A2(n23700), .B(
        mult_x_1196_n612), .Y(n23745) );
  OAI22x1_ASAP7_75t_SL U34440 ( .A1(n23717), .A2(n24038), .B1(n22936), .B2(
        mult_x_1196_n2798), .Y(mult_x_1196_n2233) );
  NAND2x1p5_ASAP7_75t_SL U34441 ( .A(mult_x_1196_n3316), .B(n24037), .Y(
        mult_x_1196_n135) );
  NOR2x1p5_ASAP7_75t_SL U34442 ( .A(mult_x_1196_n507), .B(n22894), .Y(n23730)
         );
  INVx4_ASAP7_75t_SL U34443 ( .A(n24551), .Y(add_x_735_A_4_) );
  XNOR2x1_ASAP7_75t_SL U34444 ( .A(n23973), .B(n23483), .Y(mult_x_1196_n3316)
         );
  OAI22xp5_ASAP7_75t_SL U34445 ( .A1(n24080), .A2(mult_x_1196_n3219), .B1(
        n23984), .B2(mult_x_1196_n3218), .Y(n24130) );
  XNOR2xp5_ASAP7_75t_SL U34446 ( .A(n22426), .B(n23954), .Y(mult_x_1196_n3218)
         );
  OAI21x1_ASAP7_75t_SL U34447 ( .A1(n23927), .A2(mult_x_1196_n646), .B(
        mult_x_1196_n641), .Y(mult_x_1196_n639) );
  OAI21x1_ASAP7_75t_SL U34448 ( .A1(n23453), .A2(n23454), .B(n23452), .Y(
        mult_x_1196_n668) );
  AOI21x1_ASAP7_75t_SL U34449 ( .A1(mult_x_1196_n677), .A2(n24298), .B(
        mult_x_1196_n672), .Y(n23452) );
  NAND2x1_ASAP7_75t_SL U34450 ( .A(n24298), .B(mult_x_1196_n676), .Y(n23453)
         );
  NAND2x1_ASAP7_75t_SL U34451 ( .A(n24304), .B(mult_x_1196_n638), .Y(n23455)
         );
  AOI21xp5_ASAP7_75t_SL U34452 ( .A1(mult_x_1196_n829), .A2(mult_x_1196_n744), 
        .B(n24197), .Y(n24198) );
  AND2x2_ASAP7_75t_SL U34453 ( .A(mult_x_1196_n2069), .B(mult_x_1196_n2062), 
        .Y(n24197) );
  OR2x2_ASAP7_75t_SL U34454 ( .A(mult_x_1196_n978), .B(mult_x_1196_n964), .Y(
        n23576) );
  MAJIxp5_ASAP7_75t_SL U34455 ( .A(mult_x_1196_n1538), .B(n23458), .C(
        mult_x_1196_n1532), .Y(mult_x_1196_n1487) );
  XNOR2xp5_ASAP7_75t_SL U34456 ( .A(mult_x_1196_n1532), .B(mult_x_1196_n1538), 
        .Y(n23456) );
  INVx1_ASAP7_75t_SL U34457 ( .A(n23458), .Y(n23457) );
  MAJIxp5_ASAP7_75t_SL U34458 ( .A(n23459), .B(mult_x_1196_n2613), .C(
        mult_x_1196_n2581), .Y(mult_x_1196_n1707) );
  INVx1_ASAP7_75t_SL U34459 ( .A(n23461), .Y(n23459) );
  XNOR2xp5_ASAP7_75t_SL U34460 ( .A(mult_x_1196_n2613), .B(n23461), .Y(n23460)
         );
  NOR2x1_ASAP7_75t_SL U34461 ( .A(n18390), .B(mult_x_1196_n2868), .Y(n23463)
         );
  MAJx2_ASAP7_75t_SL U34462 ( .A(mult_x_1196_n1112), .B(n22810), .C(n22338), 
        .Y(mult_x_1196_n1081) );
  OAI22xp5_ASAP7_75t_SL U34463 ( .A1(n23994), .A2(mult_x_1196_n3162), .B1(
        n23991), .B2(mult_x_1196_n3161), .Y(n23465) );
  XNOR2x1_ASAP7_75t_SL U34464 ( .A(u0_0_leon3x0_p0_muli[43]), .B(n22206), .Y(
        n23516) );
  OAI21xp5_ASAP7_75t_SL U34465 ( .A1(n23469), .A2(n23468), .B(n23467), .Y(
        n24292) );
  OAI21xp5_ASAP7_75t_SL U34466 ( .A1(mult_x_1196_n1250), .A2(mult_x_1196_n1252), .B(mult_x_1196_n1246), .Y(n23467) );
  INVx1_ASAP7_75t_SL U34467 ( .A(mult_x_1196_n1250), .Y(n23468) );
  INVx1_ASAP7_75t_SL U34468 ( .A(mult_x_1196_n1252), .Y(n23469) );
  MAJIxp5_ASAP7_75t_SL U34469 ( .A(n23699), .B(n23921), .C(mult_x_1196_n2258), 
        .Y(mult_x_1196_n1252) );
  OAI22xp5_ASAP7_75t_SL U34470 ( .A1(mult_x_1196_n2888), .A2(n24026), .B1(
        mult_x_1196_n2887), .B2(n22983), .Y(n23921) );
  INVx1_ASAP7_75t_SL U34471 ( .A(n23471), .Y(n23470) );
  XNOR2xp5_ASAP7_75t_SL U34472 ( .A(mult_x_1196_n1452), .B(n23473), .Y(n23472)
         );
  INVx1_ASAP7_75t_SL U34473 ( .A(mult_x_1196_n1419), .Y(n23473) );
  NAND2x2_ASAP7_75t_SL U34474 ( .A(mult_x_1196_n784), .B(mult_x_1196_n785), 
        .Y(mult_x_1196_n393) );
  NAND4xp75_ASAP7_75t_SL U34475 ( .A(n24252), .B(n24305), .C(n24279), .D(
        mult_x_1196_n343), .Y(mult_x_1196_n330) );
  NAND2xp5_ASAP7_75t_SL U34476 ( .A(n23576), .B(mult_x_1196_n787), .Y(n23475)
         );
  XOR2xp5_ASAP7_75t_SL U34477 ( .A(n23711), .B(n23477), .Y(n23476) );
  INVx1_ASAP7_75t_SL U34478 ( .A(mult_x_1196_n2480), .Y(n23477) );
  INVx1_ASAP7_75t_SL U34479 ( .A(mult_x_1196_n952), .Y(mult_x_1196_n946) );
  INVx1_ASAP7_75t_SL U34480 ( .A(n24251), .Y(n23478) );
  XOR2xp5_ASAP7_75t_SL U34481 ( .A(n23076), .B(n24072), .Y(n23717) );
  XOR2xp5_ASAP7_75t_SL U34482 ( .A(n23479), .B(n24066), .Y(mult_x_1196_n2793)
         );
  XOR2xp5_ASAP7_75t_SL U34483 ( .A(n23479), .B(n24067), .Y(mult_x_1196_n2794)
         );
  XOR2xp5_ASAP7_75t_SL U34484 ( .A(n23479), .B(n24061), .Y(mult_x_1196_n2788)
         );
  XOR2xp5_ASAP7_75t_SL U34485 ( .A(n23479), .B(n24062), .Y(mult_x_1196_n2789)
         );
  XOR2xp5_ASAP7_75t_SL U34486 ( .A(n23479), .B(n24075), .Y(mult_x_1196_n2802)
         );
  XOR2xp5_ASAP7_75t_SL U34487 ( .A(n18556), .B(n23479), .Y(mult_x_1196_n2779)
         );
  XOR2xp5_ASAP7_75t_SL U34488 ( .A(n24063), .B(n23479), .Y(mult_x_1196_n2790)
         );
  XOR2xp5_ASAP7_75t_SL U34489 ( .A(n23479), .B(n24065), .Y(mult_x_1196_n2792)
         );
  XOR2xp5_ASAP7_75t_SL U34490 ( .A(n24058), .B(n23479), .Y(mult_x_1196_n2785)
         );
  XOR2xp5_ASAP7_75t_SL U34491 ( .A(n24069), .B(n23479), .Y(mult_x_1196_n2796)
         );
  XOR2xp5_ASAP7_75t_SL U34492 ( .A(n24064), .B(n23479), .Y(mult_x_1196_n2791)
         );
  XOR2xp5_ASAP7_75t_SL U34493 ( .A(n23479), .B(n24068), .Y(mult_x_1196_n2795)
         );
  XOR2xp5_ASAP7_75t_SL U34494 ( .A(n22227), .B(n23479), .Y(mult_x_1196_n2803)
         );
  XOR2xp5_ASAP7_75t_SL U34495 ( .A(n24060), .B(n23076), .Y(mult_x_1196_n2787)
         );
  XOR2xp5_ASAP7_75t_SL U34496 ( .A(n23479), .B(n24074), .Y(mult_x_1196_n2801)
         );
  XOR2xp5_ASAP7_75t_SL U34497 ( .A(n23479), .B(n24073), .Y(mult_x_1196_n2800)
         );
  MAJIxp5_ASAP7_75t_SL U34498 ( .A(n24300), .B(mult_x_1196_n2450), .C(n23481), 
        .Y(mult_x_1196_n1452) );
  INVx1_ASAP7_75t_SL U34499 ( .A(mult_x_1196_n2450), .Y(n23480) );
  OAI22xp5_ASAP7_75t_SL U34500 ( .A1(mult_x_1196_n3118), .A2(n23999), .B1(
        n23996), .B2(mult_x_1196_n3117), .Y(n23481) );
  INVx1_ASAP7_75t_SL U34501 ( .A(n24278), .Y(n23485) );
  NAND2xp5_ASAP7_75t_SL U34502 ( .A(n23487), .B(n22806), .Y(n23486) );
  XNOR2xp5_ASAP7_75t_SL U34503 ( .A(n23490), .B(mult_x_1196_n39), .Y(n23489)
         );
  INVx1_ASAP7_75t_SL U34504 ( .A(u0_0_leon3x0_p0_muli[43]), .Y(n23490) );
  INVx3_ASAP7_75t_SL U34505 ( .A(mult_x_1196_n60), .Y(n24004) );
  XNOR2x1_ASAP7_75t_SL U34506 ( .A(n23491), .B(n23961), .Y(mult_x_1196_n60) );
  AND2x2_ASAP7_75t_SL U34507 ( .A(n25099), .B(n25100), .Y(n23491) );
  MAJIxp5_ASAP7_75t_SL U34508 ( .A(n24163), .B(n23492), .C(mult_x_1196_n2645), 
        .Y(mult_x_1196_n1709) );
  INVx1_ASAP7_75t_SL U34509 ( .A(n23521), .Y(n23492) );
  NOR2x1_ASAP7_75t_SL U34510 ( .A(n23494), .B(n23493), .Y(n23521) );
  MAJIxp5_ASAP7_75t_SL U34511 ( .A(n23495), .B(n18445), .C(n22372), .Y(
        mult_x_1196_n1036) );
  XNOR2xp5_ASAP7_75t_SL U34512 ( .A(mult_x_1196_n1063), .B(n24248), .Y(n23495)
         );
  INVx1_ASAP7_75t_SL U34513 ( .A(mult_x_1196_n788), .Y(n23496) );
  OAI21xp5_ASAP7_75t_SL U34514 ( .A1(mult_x_1196_n460), .A2(n23499), .B(n23497), .Y(mult_x_1196_n432) );
  NAND2xp5_ASAP7_75t_SL U34515 ( .A(mult_x_1196_n788), .B(n23498), .Y(n23497)
         );
  NAND2xp5_ASAP7_75t_SL U34516 ( .A(mult_x_1196_n451), .B(mult_x_1196_n442), 
        .Y(n23498) );
  INVx1_ASAP7_75t_SL U34517 ( .A(n23502), .Y(n23501) );
  MAJIxp5_ASAP7_75t_SL U34518 ( .A(mult_x_1196_n1591), .B(mult_x_1196_n1561), 
        .C(mult_x_1196_n1596), .Y(n23504) );
  NAND2xp5_ASAP7_75t_SL U34519 ( .A(n23506), .B(n23511), .Y(n23505) );
  NAND2xp5_ASAP7_75t_SL U34520 ( .A(mult_x_1196_n1147), .B(mult_x_1196_n1122), 
        .Y(n23506) );
  NAND2xp5_ASAP7_75t_SL U34521 ( .A(n23508), .B(n23510), .Y(n23507) );
  INVx1_ASAP7_75t_SL U34522 ( .A(mult_x_1196_n1122), .Y(n23510) );
  INVx1_ASAP7_75t_SL U34523 ( .A(n23606), .Y(n23513) );
  XOR2xp5_ASAP7_75t_SL U34524 ( .A(mult_x_1196_n1859), .B(mult_x_1196_n1838), 
        .Y(n23514) );
  XNOR2xp5_ASAP7_75t_SL U34525 ( .A(mult_x_1196_n1074), .B(mult_x_1196_n1095), 
        .Y(n23515) );
  OAI21xp5_ASAP7_75t_SL U34526 ( .A1(mult_x_1196_n689), .A2(mult_x_1196_n693), 
        .B(mult_x_1196_n690), .Y(mult_x_1196_n688) );
  NOR2x1_ASAP7_75t_SL U34527 ( .A(mult_x_1196_n689), .B(mult_x_1196_n692), .Y(
        mult_x_1196_n687) );
  NOR2x1_ASAP7_75t_SL U34528 ( .A(mult_x_1196_n683), .B(mult_x_1196_n678), .Y(
        mult_x_1196_n676) );
  OR2x2_ASAP7_75t_SL U34529 ( .A(mult_x_1196_n1889), .B(mult_x_1196_n1869), 
        .Y(n24298) );
  OR2x2_ASAP7_75t_SL U34530 ( .A(n23996), .B(mult_x_1196_n3128), .Y(n24257) );
  XOR2xp5_ASAP7_75t_SL U34531 ( .A(n23517), .B(mult_x_1196_n2587), .Y(n24225)
         );
  INVx1_ASAP7_75t_SL U34532 ( .A(mult_x_1196_n2134), .Y(n23520) );
  XOR2xp5_ASAP7_75t_SL U34533 ( .A(n23521), .B(n24163), .Y(n24161) );
  BUFx6f_ASAP7_75t_SL U34534 ( .A(n24107), .Y(n23522) );
  AOI21xp5_ASAP7_75t_SL U34535 ( .A1(n24106), .A2(n18528), .B(
        mult_x_1196_n3179), .Y(n23523) );
  OAI22xp5_ASAP7_75t_SL U34536 ( .A1(n23522), .A2(mult_x_1196_n3184), .B1(
        n23987), .B2(mult_x_1196_n3183), .Y(mult_x_1196_n2608) );
  OAI22xp5_ASAP7_75t_SL U34537 ( .A1(n23522), .A2(mult_x_1196_n3181), .B1(
        n22248), .B2(mult_x_1196_n3180), .Y(mult_x_1196_n2605) );
  MAJIxp5_ASAP7_75t_SL U34538 ( .A(n23541), .B(n18913), .C(mult_x_1196_n1660), 
        .Y(n23525) );
  XOR2xp5_ASAP7_75t_SL U34539 ( .A(mult_x_1196_n1674), .B(n23527), .Y(n23526)
         );
  INVx1_ASAP7_75t_SL U34540 ( .A(mult_x_1196_n1625), .Y(n23528) );
  NAND2xp5_ASAP7_75t_SL U34541 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__19_), .B(
        n22434), .Y(n23530) );
  NOR2x1_ASAP7_75t_SL U34542 ( .A(mult_x_1196_n354), .B(mult_x_1196_n347), .Y(
        mult_x_1196_n343) );
  OR2x2_ASAP7_75t_SL U34543 ( .A(mult_x_1196_n918), .B(mult_x_1196_n902), .Y(
        n24279) );
  NAND2xp5_ASAP7_75t_SL U34544 ( .A(n24279), .B(n24305), .Y(mult_x_1196_n361)
         );
  NAND2xp5_ASAP7_75t_SL U34545 ( .A(n24252), .B(mult_x_1196_n343), .Y(
        mult_x_1196_n334) );
  OAI22xp5_ASAP7_75t_SL U34546 ( .A1(n24041), .A2(mult_x_1196_n2749), .B1(
        n24040), .B2(n23534), .Y(mult_x_1196_n2186) );
  XOR2xp5_ASAP7_75t_SL U34547 ( .A(mult_x_1196_n1321), .B(n22720), .Y(n23535)
         );
  INVx1_ASAP7_75t_SL U34548 ( .A(mult_x_1196_n1315), .Y(n23536) );
  INVx1_ASAP7_75t_SL U34549 ( .A(mult_x_1196_n1022), .Y(n23537) );
  INVx1_ASAP7_75t_SL U34550 ( .A(n22363), .Y(n23538) );
  NAND2xp5_ASAP7_75t_SL U34551 ( .A(mult_x_1196_n1016), .B(mult_x_1196_n998), 
        .Y(mult_x_1196_n442) );
  INVx1_ASAP7_75t_SL U34552 ( .A(mult_x_1196_n1098), .Y(n23539) );
  XOR2xp5_ASAP7_75t_SL U34553 ( .A(mult_x_1196_n1124), .B(mult_x_1196_n1102), 
        .Y(n23540) );
  XNOR2xp5_ASAP7_75t_SL U34554 ( .A(n24140), .B(n24139), .Y(mult_x_1196_n1184)
         );
  OR2x2_ASAP7_75t_SL U34555 ( .A(n24137), .B(n24138), .Y(n24140) );
  XNOR2xp5_ASAP7_75t_SL U34556 ( .A(n22297), .B(n23543), .Y(mult_x_1196_n2000)
         );
  XNOR2xp5_ASAP7_75t_SL U34557 ( .A(n23545), .B(n23546), .Y(n23888) );
  INVx1_ASAP7_75t_SL U34558 ( .A(mult_x_1196_n2022), .Y(n23545) );
  XNOR2xp5_ASAP7_75t_SL U34559 ( .A(n23547), .B(mult_x_1196_n2018), .Y(n23546)
         );
  INVx1_ASAP7_75t_SL U34560 ( .A(mult_x_1196_n2034), .Y(n23547) );
  NOR2x1_ASAP7_75t_SL U34561 ( .A(n28956), .B(n23831), .Y(n30604) );
  INVx1_ASAP7_75t_SL U34562 ( .A(u0_0_leon3x0_p0_iu_r_E__INVOP2_), .Y(n23548)
         );
  NOR2xp33_ASAP7_75t_SL U34563 ( .A(n30817), .B(n18884), .Y(n25086) );
  OAI22xp5_ASAP7_75t_SL U34564 ( .A1(n28715), .A2(n23559), .B1(n24689), .B2(
        n23549), .Y(u0_0_leon3x0_p0_muli[20]) );
  OAI22xp5_ASAP7_75t_SL U34565 ( .A1(n28472), .A2(n23831), .B1(n24689), .B2(
        n23550), .Y(u0_0_leon3x0_p0_muli[31]) );
  INVx1_ASAP7_75t_SL U34566 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__23_), .Y(
        n23550) );
  NAND2xp5_ASAP7_75t_SL U34567 ( .A(n23552), .B(n28676), .Y(
        u0_0_leon3x0_p0_muli[21]) );
  NAND2xp5_ASAP7_75t_SL U34568 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__11_), .B(
        n24689), .Y(n23552) );
  NAND2xp5_ASAP7_75t_SL U34569 ( .A(n23553), .B(n28478), .Y(
        u0_0_leon3x0_p0_muli[30]) );
  NAND2xp5_ASAP7_75t_SL U34570 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__22_), .B(
        n24689), .Y(n23553) );
  NAND2xp5_ASAP7_75t_SL U34571 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__14_), .B(
        n24689), .Y(n23554) );
  NAND2xp5_ASAP7_75t_SL U34572 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__31_), .B(
        n23849), .Y(n23555) );
  NAND2xp5_ASAP7_75t_SL U34573 ( .A(n23556), .B(n26987), .Y(
        u0_0_leon3x0_p0_muli[28]) );
  NAND2xp5_ASAP7_75t_SL U34574 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__20_), .B(
        n24689), .Y(n23556) );
  NAND2xp5_ASAP7_75t_SL U34575 ( .A(n23557), .B(n26301), .Y(
        u0_0_leon3x0_p0_muli[16]) );
  NAND2xp5_ASAP7_75t_SL U34576 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__5_), .B(
        n24689), .Y(n23557) );
  NAND2xp5_ASAP7_75t_SL U34577 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__29_), .B(
        n24689), .Y(n23558) );
  OAI21xp5_ASAP7_75t_SL U34578 ( .A1(n30487), .A2(n18884), .B(n26739), .Y(
        n28992) );
  NAND2xp5_ASAP7_75t_SL U34579 ( .A(n18884), .B(n25121), .Y(n26739) );
  XNOR2xp5_ASAP7_75t_SL U34580 ( .A(n23050), .B(n24056), .Y(mult_x_1196_n2987)
         );
  MAJIxp5_ASAP7_75t_SL U34581 ( .A(mult_x_1196_n2396), .B(mult_x_1196_n2552), 
        .C(n23562), .Y(mult_x_1196_n1788) );
  XOR2xp5_ASAP7_75t_SL U34582 ( .A(n23562), .B(n23561), .Y(n23560) );
  INVx1_ASAP7_75t_SL U34583 ( .A(mult_x_1196_n2552), .Y(n23561) );
  MAJIxp5_ASAP7_75t_SL U34584 ( .A(mult_x_1196_n2140), .B(n23564), .C(
        mult_x_1196_n2665), .Y(mult_x_1196_n2071) );
  MAJIxp5_ASAP7_75t_SL U34585 ( .A(mult_x_1196_n1979), .B(mult_x_1196_n1981), 
        .C(mult_x_1196_n1972), .Y(mult_x_1196_n1973) );
  NOR2xp33_ASAP7_75t_SL U34586 ( .A(n27088), .B(n18910), .Y(n23569) );
  INVx2_ASAP7_75t_SL U34587 ( .A(n23986), .Y(n23570) );
  NAND3xp33_ASAP7_75t_SL U34588 ( .A(n23574), .B(n18416), .C(n23573), .Y(
        n23572) );
  XOR2xp5_ASAP7_75t_SL U34589 ( .A(mult_x_1196_n2163), .B(n24179), .Y(n24178)
         );
  OR2x2_ASAP7_75t_SL U34590 ( .A(n24176), .B(n24177), .Y(n24179) );
  INVx2_ASAP7_75t_SL U34591 ( .A(n22929), .Y(mult_x_1196_n580) );
  INVx1_ASAP7_75t_SL U34592 ( .A(n23580), .Y(n23578) );
  MAJIxp5_ASAP7_75t_SL U34593 ( .A(mult_x_1196_n2481), .B(n23585), .C(
        mult_x_1196_n2573), .Y(mult_x_1196_n1420) );
  XNOR2xp5_ASAP7_75t_SL U34594 ( .A(n23586), .B(n23584), .Y(mult_x_1196_n1421)
         );
  INVx1_ASAP7_75t_SL U34595 ( .A(mult_x_1196_n2481), .Y(n23586) );
  OAI21xp5_ASAP7_75t_SL U34596 ( .A1(mult_x_1196_n1964), .A2(mult_x_1196_n1962), .B(mult_x_1196_n1966), .Y(n23592) );
  MAJIxp5_ASAP7_75t_SL U34597 ( .A(mult_x_1196_n2362), .B(n23595), .C(
        mult_x_1196_n2394), .Y(mult_x_1196_n1733) );
  INVx1_ASAP7_75t_SL U34598 ( .A(mult_x_1196_n2394), .Y(n23593) );
  XOR2xp5_ASAP7_75t_SL U34599 ( .A(n23595), .B(mult_x_1196_n2362), .Y(n23594)
         );
  OAI22xp5_ASAP7_75t_SL U34600 ( .A1(mult_x_1196_n3030), .A2(n24009), .B1(
        mult_x_1196_n3029), .B2(n23442), .Y(n23595) );
  AND2x2_ASAP7_75t_SL U34601 ( .A(mult_x_1196_n2519), .B(mult_x_1196_n2679), 
        .Y(n23606) );
  OR2x2_ASAP7_75t_SL U34602 ( .A(n22428), .B(mult_x_1196_n227), .Y(n23600) );
  OAI21xp5_ASAP7_75t_SL U34603 ( .A1(n18423), .A2(n22487), .B(n23603), .Y(
        mult_x_1196_n2133) );
  NAND2xp5_ASAP7_75t_SL U34604 ( .A(n22267), .B(n18563), .Y(n23603) );
  NAND2xp33_ASAP7_75t_SL U34605 ( .A(mult_x_1196_n859), .B(mult_x_1196_n852), 
        .Y(mult_x_1196_n317) );
  MAJIxp5_ASAP7_75t_SL U34606 ( .A(mult_x_1196_n2615), .B(mult_x_1196_n2491), 
        .C(mult_x_1196_n2583), .Y(mult_x_1196_n1765) );
  INVx1_ASAP7_75t_SL U34607 ( .A(mult_x_1196_n2491), .Y(n23604) );
  NAND2xp5_ASAP7_75t_SL U34608 ( .A(mult_x_1196_n1964), .B(mult_x_1196_n1962), 
        .Y(n23605) );
  NAND2xp5_ASAP7_75t_SL U34609 ( .A(n23607), .B(mult_x_1196_n1989), .Y(n24273)
         );
  XNOR2xp5_ASAP7_75t_SL U34610 ( .A(mult_x_1196_n2130), .B(mult_x_1196_n1739), 
        .Y(n23608) );
  XNOR2xp5_ASAP7_75t_SL U34611 ( .A(n23613), .B(n23609), .Y(mult_x_1196_n1544)
         );
  XNOR2xp5_ASAP7_75t_SL U34612 ( .A(mult_x_1196_n1542), .B(mult_x_1196_n1583), 
        .Y(n23609) );
  INVx1_ASAP7_75t_SL U34613 ( .A(mult_x_1196_n1542), .Y(n23610) );
  INVx1_ASAP7_75t_SL U34614 ( .A(mult_x_1196_n1583), .Y(n23611) );
  INVx1_ASAP7_75t_SL U34615 ( .A(mult_x_1196_n1586), .Y(n23612) );
  MAJIxp5_ASAP7_75t_SL U34616 ( .A(n23615), .B(mult_x_1196_n1443), .C(
        mult_x_1196_n1476), .Y(mult_x_1196_n1433) );
  XNOR2xp5_ASAP7_75t_SL U34617 ( .A(n23618), .B(mult_x_1196_n1387), .Y(n23617)
         );
  NOR2xp33_ASAP7_75t_SL U34618 ( .A(n24046), .B(n28769), .Y(n28381) );
  INVx1_ASAP7_75t_SL U34619 ( .A(mult_x_1196_n2004), .Y(mult_x_1196_n2001) );
  INVx1_ASAP7_75t_SL U34620 ( .A(mult_x_1196_n2002), .Y(n23624) );
  MAJx2_ASAP7_75t_SL U34621 ( .A(mult_x_1196_n2022), .B(mult_x_1196_n2034), 
        .C(mult_x_1196_n2018), .Y(mult_x_1196_n2002) );
  XOR2x2_ASAP7_75t_SL U34622 ( .A(u0_0_leon3x0_p0_muli[47]), .B(n24421), .Y(
        n24024) );
  INVx1_ASAP7_75t_SL U34623 ( .A(n23628), .Y(n23625) );
  XOR2xp5_ASAP7_75t_SL U34624 ( .A(n23627), .B(n23626), .Y(mult_x_1196_n1981)
         );
  INVx1_ASAP7_75t_SL U34625 ( .A(mult_x_1196_n2561), .Y(n23626) );
  XNOR2xp5_ASAP7_75t_SL U34626 ( .A(n23628), .B(mult_x_1196_n2501), .Y(n23627)
         );
  NOR2x1_ASAP7_75t_SL U34627 ( .A(n23630), .B(n23629), .Y(n23628) );
  NOR2x1_ASAP7_75t_SL U34628 ( .A(mult_x_1196_n3041), .B(n24009), .Y(n23630)
         );
  INVx1_ASAP7_75t_SL U34629 ( .A(mult_x_1196_n2358), .Y(n23631) );
  INVx1_ASAP7_75t_SL U34630 ( .A(mult_x_1196_n2454), .Y(n23633) );
  MAJIxp5_ASAP7_75t_SL U34631 ( .A(n23634), .B(mult_x_1196_n2305), .C(
        mult_x_1196_n2647), .Y(mult_x_1196_n1767) );
  INVx1_ASAP7_75t_SL U34632 ( .A(n24203), .Y(n23634) );
  NOR2x1_ASAP7_75t_SL U34633 ( .A(mult_x_1196_n2903), .B(n23708), .Y(n23635)
         );
  INVx1_ASAP7_75t_SL U34634 ( .A(n23636), .Y(mult_x_1196_n1331) );
  XNOR2x1_ASAP7_75t_SL U34635 ( .A(u0_0_leon3x0_p0_muli[45]), .B(n23962), .Y(
        n23638) );
  BUFx6f_ASAP7_75t_SL U34636 ( .A(mult_x_1196_n39), .Y(n23639) );
  NAND2xp5_ASAP7_75t_SL U34637 ( .A(n23641), .B(n25404), .Y(n28404) );
  OAI21xp5_ASAP7_75t_SL U34638 ( .A1(n22578), .A2(n28868), .B(n26259), .Y(
        n28966) );
  NAND2xp5_ASAP7_75t_SL U34639 ( .A(n23642), .B(n25787), .Y(n27091) );
  NAND2x2_ASAP7_75t_SL U34640 ( .A(n24237), .B(n23644), .Y(n24013) );
  INVx2_ASAP7_75t_SL U34641 ( .A(n24010), .Y(n23644) );
  XNOR2x1_ASAP7_75t_SL U34642 ( .A(add_x_735_A_16_), .B(n26683), .Y(n24010) );
  BUFx6f_ASAP7_75t_SL U34643 ( .A(n24010), .Y(n23645) );
  INVx1_ASAP7_75t_SL U34644 ( .A(mult_x_1196_n968), .Y(mult_x_1196_n962) );
  OR2x2_ASAP7_75t_SL U34645 ( .A(mult_x_1196_n1194), .B(mult_x_1196_n1166), 
        .Y(mult_x_1196_n507) );
  NOR2x1_ASAP7_75t_SL U34646 ( .A(mult_x_1196_n1929), .B(mult_x_1196_n1932), 
        .Y(mult_x_1196_n689) );
  NOR2x1_ASAP7_75t_SL U34647 ( .A(n22328), .B(n22327), .Y(mult_x_1196_n1929)
         );
  NAND2xp5_ASAP7_75t_SL U34648 ( .A(n23649), .B(n25146), .Y(n25910) );
  INVx1_ASAP7_75t_SL U34649 ( .A(n23960), .Y(n23651) );
  XNOR2xp5_ASAP7_75t_SL U34650 ( .A(n23655), .B(n23654), .Y(mult_x_1196_n1188)
         );
  NAND2xp5_ASAP7_75t_SL U34651 ( .A(mult_x_1196_n963), .B(mult_x_1196_n948), 
        .Y(mult_x_1196_n407) );
  OAI22xp5_ASAP7_75t_SL U34652 ( .A1(mult_x_1196_n3273), .A2(n23981), .B1(
        n23980), .B2(mult_x_1196_n3272), .Y(n23656) );
  XNOR2xp5_ASAP7_75t_SL U34653 ( .A(n22425), .B(n24076), .Y(mult_x_1196_n3118)
         );
  XNOR2xp5_ASAP7_75t_SL U34654 ( .A(n24076), .B(n22426), .Y(mult_x_1196_n3116)
         );
  INVx1_ASAP7_75t_SL U34655 ( .A(n24050), .Y(n23657) );
  XOR2xp5_ASAP7_75t_SL U34656 ( .A(n23643), .B(n24045), .Y(mult_x_1196_n3112)
         );
  XOR2xp5_ASAP7_75t_SL U34657 ( .A(n24076), .B(n24055), .Y(mult_x_1196_n3122)
         );
  XNOR2xp5_ASAP7_75t_SL U34658 ( .A(n23658), .B(n24054), .Y(mult_x_1196_n3121)
         );
  XNOR2xp5_ASAP7_75t_SL U34659 ( .A(n23658), .B(n24046), .Y(mult_x_1196_n3113)
         );
  XOR2xp5_ASAP7_75t_SL U34660 ( .A(n24044), .B(n22578), .Y(mult_x_1196_n3111)
         );
  XNOR2xp5_ASAP7_75t_SL U34661 ( .A(n22448), .B(n24047), .Y(mult_x_1196_n3114)
         );
  XOR2xp5_ASAP7_75t_SL U34662 ( .A(n24076), .B(n24053), .Y(mult_x_1196_n3120)
         );
  XNOR2xp5_ASAP7_75t_SL U34663 ( .A(n23658), .B(n24056), .Y(mult_x_1196_n3123)
         );
  XNOR2x1_ASAP7_75t_SL U34664 ( .A(n23661), .B(mult_x_1196_n1818), .Y(n23660)
         );
  NOR2xp33_ASAP7_75t_SL U34665 ( .A(n23981), .B(mult_x_1196_n3256), .Y(n23662)
         );
  XNOR2xp5_ASAP7_75t_SL U34666 ( .A(mult_x_1196_n2031), .B(mult_x_1196_n2046), 
        .Y(n23664) );
  AND2x2_ASAP7_75t_SL U34667 ( .A(n25093), .B(n25094), .Y(n26683) );
  NAND2xp5_ASAP7_75t_SL U34668 ( .A(n23665), .B(u0_0_leon3x0_p0_divi[15]), .Y(
        add_x_735_n174) );
  NOR2x1_ASAP7_75t_SL U34669 ( .A(n23665), .B(u0_0_leon3x0_p0_divi[15]), .Y(
        add_x_735_n173) );
  MAJIxp5_ASAP7_75t_SL U34670 ( .A(mult_x_1196_n2280), .B(n23667), .C(
        mult_x_1196_n2338), .Y(mult_x_1196_n991) );
  INVx1_ASAP7_75t_SL U34671 ( .A(mult_x_1196_n995), .Y(n23667) );
  XNOR2xp5_ASAP7_75t_SL U34672 ( .A(n23668), .B(mult_x_1196_n2280), .Y(
        mult_x_1196_n992) );
  INVx1_ASAP7_75t_SL U34673 ( .A(mult_x_1196_n357), .Y(mult_x_1196_n359) );
  AOI21xp33_ASAP7_75t_SL U34674 ( .A1(n22254), .A2(n18995), .B(n22252), .Y(
        mult_x_1196_n637) );
  XOR2xp5_ASAP7_75t_SL U34675 ( .A(n22254), .B(mult_x_1196_n263), .Y(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N27) );
  AOI21xp5_ASAP7_75t_SL U34676 ( .A1(mult_x_1196_n386), .A2(n23672), .B(n23671), .Y(n23670) );
  NAND3xp33_ASAP7_75t_SL U34677 ( .A(n23674), .B(n18932), .C(mult_x_1196_n781), 
        .Y(n23673) );
  XNOR2xp5_ASAP7_75t_SL U34678 ( .A(n23678), .B(n23677), .Y(mult_x_1196_n1704)
         );
  INVx1_ASAP7_75t_SL U34679 ( .A(mult_x_1196_n2457), .Y(n23677) );
  OAI21xp5_ASAP7_75t_SL U34680 ( .A1(mult_x_1196_n3061), .A2(n24007), .B(
        n22275), .Y(n23679) );
  NAND2xp5_ASAP7_75t_SL U34681 ( .A(n23683), .B(mult_x_1196_n386), .Y(n23681)
         );
  NAND3xp33_ASAP7_75t_SL U34682 ( .A(mult_x_1196_n465), .B(mult_x_1196_n385), 
        .C(n23683), .Y(n23682) );
  AO21x1_ASAP7_75t_SL U34683 ( .A1(mult_x_1196_n385), .A2(n18932), .B(
        mult_x_1196_n386), .Y(n23765) );
  OAI21xp5_ASAP7_75t_SL U34684 ( .A1(mult_x_1196_n379), .A2(n22533), .B(n23684), .Y(mult_x_1196_n378) );
  INVx1_ASAP7_75t_SL U34685 ( .A(n23765), .Y(n23684) );
  OAI21xp5_ASAP7_75t_SL U34686 ( .A1(mult_x_1196_n1376), .A2(mult_x_1196_n1409), .B(mult_x_1196_n1374), .Y(n23685) );
  NAND2xp5_ASAP7_75t_SL U34687 ( .A(mult_x_1196_n1376), .B(mult_x_1196_n1409), 
        .Y(n23686) );
  XOR2xp5_ASAP7_75t_SL U34688 ( .A(n22363), .B(mult_x_1196_n1006), .Y(n23687)
         );
  INVx1_ASAP7_75t_SL U34689 ( .A(n24210), .Y(n23688) );
  XNOR2xp5_ASAP7_75t_SL U34690 ( .A(n23690), .B(mult_x_1196_n1733), .Y(n23689)
         );
  INVx1_ASAP7_75t_SL U34691 ( .A(mult_x_1196_n1737), .Y(n23690) );
  OAI21xp5_ASAP7_75t_SL U34692 ( .A1(mult_x_1196_n1093), .A2(mult_x_1196_n1067), .B(n23692), .Y(mult_x_1196_n1061) );
  NAND2xp5_ASAP7_75t_SL U34693 ( .A(mult_x_1196_n1088), .B(n23693), .Y(n23692)
         );
  XOR2xp5_ASAP7_75t_SL U34694 ( .A(mult_x_1196_n1093), .B(mult_x_1196_n1067), 
        .Y(n23694) );
  OAI22xp5_ASAP7_75t_SL U34695 ( .A1(n24030), .A2(mult_x_1196_n2859), .B1(
        n24031), .B2(n23695), .Y(mult_x_1196_n2294) );
  INVx1_ASAP7_75t_SL U34696 ( .A(n23697), .Y(n23695) );
  XOR2xp5_ASAP7_75t_SL U34697 ( .A(n23971), .B(n24065), .Y(n23697) );
  INVx1_ASAP7_75t_SL U34698 ( .A(n18416), .Y(n24175) );
  NAND2xp5_ASAP7_75t_SL U34699 ( .A(mult_x_1196_n464), .B(mult_x_1196_n420), 
        .Y(mult_x_1196_n418) );
  AND2x2_ASAP7_75t_SL U34700 ( .A(n18416), .B(n23669), .Y(mult_x_1196_n420) );
  XOR2xp5_ASAP7_75t_SL U34701 ( .A(n23698), .B(n23921), .Y(mult_x_1196_n1253)
         );
  XNOR2xp5_ASAP7_75t_SL U34702 ( .A(n23699), .B(mult_x_1196_n2258), .Y(n23698)
         );
  OAI22xp5_ASAP7_75t_SL U34703 ( .A1(mult_x_1196_n3112), .A2(n23999), .B1(
        n23997), .B2(mult_x_1196_n3111), .Y(n23699) );
  INVx1_ASAP7_75t_SL U34704 ( .A(n23700), .Y(mult_x_1196_n629) );
  XOR2xp5_ASAP7_75t_SL U34705 ( .A(mult_x_1196_n1318), .B(mult_x_1196_n1288), 
        .Y(n23703) );
  INVx1_ASAP7_75t_SL U34706 ( .A(mult_x_1196_n1825), .Y(n23709) );
  MAJIxp5_ASAP7_75t_SL U34707 ( .A(n23712), .B(mult_x_1196_n1074), .C(
        mult_x_1196_n1078), .Y(mult_x_1196_n1066) );
  INVx1_ASAP7_75t_SL U34708 ( .A(mult_x_1196_n1095), .Y(n23712) );
  MAJIxp5_ASAP7_75t_SL U34709 ( .A(n23714), .B(mult_x_1196_n2657), .C(
        mult_x_1196_n2625), .Y(mult_x_1196_n1982) );
  XNOR2xp5_ASAP7_75t_SL U34710 ( .A(mult_x_1196_n2657), .B(n23713), .Y(
        mult_x_1196_n1983) );
  XOR2xp5_ASAP7_75t_SL U34711 ( .A(mult_x_1196_n2625), .B(n23714), .Y(n23713)
         );
  OAI22xp5_ASAP7_75t_SL U34712 ( .A1(mult_x_1196_n3168), .A2(n23992), .B1(
        mult_x_1196_n3169), .B2(n23081), .Y(n23714) );
  INVx1_ASAP7_75t_SL U34713 ( .A(mult_x_1196_n1964), .Y(n23715) );
  MAJIxp5_ASAP7_75t_SL U34714 ( .A(mult_x_1196_n2223), .B(n23716), .C(
        mult_x_1196_n2345), .Y(mult_x_1196_n1154) );
  OAI22xp5_ASAP7_75t_SL U34715 ( .A1(mult_x_1196_n3013), .A2(n22563), .B1(
        mult_x_1196_n3012), .B2(n23442), .Y(n23716) );
  OAI22xp5_ASAP7_75t_SL U34716 ( .A1(mult_x_1196_n2800), .A2(n24038), .B1(
        n22391), .B2(n23717), .Y(n24212) );
  NOR2x1_ASAP7_75t_SL U34717 ( .A(mult_x_1196_n877), .B(n22313), .Y(
        mult_x_1196_n347) );
  MAJIxp5_ASAP7_75t_SL U34718 ( .A(mult_x_1196_n2476), .B(mult_x_1196_n1255), 
        .C(n23718), .Y(mult_x_1196_n1250) );
  OAI21xp5_ASAP7_75t_SL U34719 ( .A1(n23722), .A2(n23724), .B(
        mult_x_1196_n1945), .Y(n23721) );
  XNOR2xp5_ASAP7_75t_SL U34720 ( .A(n23723), .B(mult_x_1196_n1945), .Y(
        mult_x_1196_n1922) );
  XOR2xp5_ASAP7_75t_SL U34721 ( .A(mult_x_1196_n2466), .B(n23724), .Y(n23723)
         );
  MAJIxp5_ASAP7_75t_SL U34722 ( .A(mult_x_1196_n1672), .B(mult_x_1196_n1678), 
        .C(n23725), .Y(mult_x_1196_n1659) );
  INVx1_ASAP7_75t_SL U34723 ( .A(n23726), .Y(n23725) );
  NOR2x1_ASAP7_75t_SL U34724 ( .A(n23729), .B(n23727), .Y(n23726) );
  INVx1_ASAP7_75t_SL U34725 ( .A(mult_x_1196_n1739), .Y(n23728) );
  NOR2x1_ASAP7_75t_SL U34726 ( .A(mult_x_1196_n1712), .B(mult_x_1196_n2130), 
        .Y(n23729) );
  OAI21xp33_ASAP7_75t_SL U34727 ( .A1(mult_x_1196_n496), .A2(mult_x_1196_n488), 
        .B(n18422), .Y(mult_x_1196_n487) );
  INVx1_ASAP7_75t_SL U34728 ( .A(mult_x_1196_n504), .Y(n23731) );
  NAND2xp5_ASAP7_75t_SL U34729 ( .A(mult_x_1196_n1135), .B(mult_x_1196_n1134), 
        .Y(mult_x_1196_n504) );
  MAJIxp5_ASAP7_75t_SL U34730 ( .A(n23913), .B(mult_x_1196_n2162), .C(n23733), 
        .Y(mult_x_1196_n1158) );
  INVx1_ASAP7_75t_SL U34731 ( .A(n24158), .Y(n23733) );
  NOR2x1_ASAP7_75t_SL U34732 ( .A(n24157), .B(n23734), .Y(n24158) );
  AOI21xp33_ASAP7_75t_SL U34733 ( .A1(n18932), .A2(mult_x_1196_n306), .B(
        n22219), .Y(n23736) );
  NAND2xp33_ASAP7_75t_SL U34734 ( .A(mult_x_1196_n464), .B(mult_x_1196_n306), 
        .Y(n23737) );
  XNOR2xp5_ASAP7_75t_SL U34735 ( .A(mult_x_1196_n2535), .B(n23739), .Y(n23738)
         );
  NAND2x2_ASAP7_75t_SL U34736 ( .A(n23741), .B(n22268), .Y(add_x_735_A_25_) );
  NOR2x1_ASAP7_75t_SL U34737 ( .A(mult_x_1196_n330), .B(mult_x_1196_n379), .Y(
        mult_x_1196_n328) );
  OAI21xp5_ASAP7_75t_SL U34738 ( .A1(mult_x_1196_n586), .A2(mult_x_1196_n594), 
        .B(mult_x_1196_n587), .Y(n23744) );
  NAND2xp5_ASAP7_75t_SL U34739 ( .A(mult_x_1196_n1467), .B(n22349), .Y(
        mult_x_1196_n587) );
  NAND2xp5_ASAP7_75t_SL U34740 ( .A(n22345), .B(mult_x_1196_n1504), .Y(
        mult_x_1196_n594) );
  NOR2x1_ASAP7_75t_SL U34741 ( .A(mult_x_1196_n586), .B(mult_x_1196_n591), .Y(
        mult_x_1196_n584) );
  NOR2x1_ASAP7_75t_SL U34742 ( .A(n22349), .B(mult_x_1196_n1467), .Y(
        mult_x_1196_n586) );
  NOR2x1_ASAP7_75t_SL U34743 ( .A(n24222), .B(n24223), .Y(n24224) );
  OAI21xp5_ASAP7_75t_SL U34744 ( .A1(mult_x_1196_n2905), .A2(n23708), .B(
        n22270), .Y(mult_x_1196_n2333) );
  OAI21xp5_ASAP7_75t_SL U34745 ( .A1(n24121), .A2(mult_x_1196_n3225), .B(
        n23751), .Y(mult_x_1196_n2649) );
  NAND2xp5_ASAP7_75t_SL U34746 ( .A(n23756), .B(n23755), .Y(n23754) );
  INVx1_ASAP7_75t_SL U34747 ( .A(mult_x_1196_n1610), .Y(n23755) );
  INVx1_ASAP7_75t_SL U34748 ( .A(mult_x_1196_n1604), .Y(n23756) );
  BUFx6f_ASAP7_75t_SL U34749 ( .A(n23986), .Y(n23757) );
  MAJIxp5_ASAP7_75t_SL U34750 ( .A(mult_x_1196_n1674), .B(mult_x_1196_n1661), 
        .C(mult_x_1196_n1670), .Y(mult_x_1196_n1662) );
  INVx1_ASAP7_75t_SL U34751 ( .A(mult_x_1196_n2588), .Y(n23758) );
  XOR2xp5_ASAP7_75t_SL U34752 ( .A(mult_x_1196_n2400), .B(n23760), .Y(n23759)
         );
  OAI21xp5_ASAP7_75t_SL U34753 ( .A1(n23766), .A2(n22258), .B(n23764), .Y(
        n23763) );
  AOI21xp5_ASAP7_75t_SL U34754 ( .A1(n23765), .A2(n24305), .B(mult_x_1196_n375), .Y(n23764) );
  NAND2xp5_ASAP7_75t_SL U34755 ( .A(n24305), .B(n23767), .Y(n23766) );
  INVx1_ASAP7_75t_SL U34756 ( .A(mult_x_1196_n379), .Y(n23767) );
  INVx1_ASAP7_75t_SL U34757 ( .A(mult_x_1196_n364), .Y(n23768) );
  INVx1_ASAP7_75t_SL U34758 ( .A(mult_x_1196_n361), .Y(n23769) );
  INVx1_ASAP7_75t_SL U34759 ( .A(mult_x_1196_n1015), .Y(mult_x_1196_n1002) );
  INVx1_ASAP7_75t_SL U34760 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__17_), .Y(n23771)
         );
  INVx1_ASAP7_75t_SL U34761 ( .A(n24029), .Y(n23775) );
  NAND2xp5_ASAP7_75t_SL U34762 ( .A(n23779), .B(n23777), .Y(n23776) );
  INVx1_ASAP7_75t_SL U34763 ( .A(mult_x_1196_n2319), .Y(n23777) );
  NOR2x1_ASAP7_75t_SL U34764 ( .A(n23637), .B(mult_x_1196_n3051), .Y(n23780)
         );
  NOR2x1_ASAP7_75t_SL U34765 ( .A(mult_x_1196_n3050), .B(n24005), .Y(n23781)
         );
  XNOR2xp5_ASAP7_75t_SL U34766 ( .A(n23783), .B(mult_x_1196_n1487), .Y(
        mult_x_1196_n1446) );
  XNOR2xp5_ASAP7_75t_SL U34767 ( .A(mult_x_1196_n1991), .B(mult_x_1196_n1976), 
        .Y(n23784) );
  INVxp67_ASAP7_75t_SL U34768 ( .A(mult_x_1196_n1298), .Y(n23785) );
  NOR2x1_ASAP7_75t_SL U34769 ( .A(n24303), .B(n24286), .Y(mult_x_1196_n546) );
  INVx1_ASAP7_75t_SL U34770 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__24_), .Y(
        n26514) );
  AND2x2_ASAP7_75t_SL U34771 ( .A(n24042), .B(n22279), .Y(mult_x_1196_n2154)
         );
  OAI21xp5_ASAP7_75t_SL U34772 ( .A1(mult_x_1196_n3072), .A2(n18561), .B(
        n22277), .Y(n23793) );
  XNOR2xp5_ASAP7_75t_SL U34773 ( .A(n23794), .B(mult_x_1196_n1316), .Y(n24164)
         );
  INVx1_ASAP7_75t_SL U34774 ( .A(mult_x_1196_n1973), .Y(n23796) );
  XOR2xp5_ASAP7_75t_SL U34775 ( .A(mult_x_1196_n1973), .B(n23798), .Y(n23797)
         );
  NAND2xp5_ASAP7_75t_SL U34776 ( .A(mult_x_1196_n902), .B(mult_x_1196_n918), 
        .Y(mult_x_1196_n368) );
  AND2x2_ASAP7_75t_SL U34777 ( .A(mult_x_1196_n1580), .B(mult_x_1196_n1544), 
        .Y(mult_x_1196_n602) );
  NOR2x1_ASAP7_75t_SL U34778 ( .A(n23802), .B(n23803), .Y(n23801) );
  INVx1_ASAP7_75t_SL U34779 ( .A(n22212), .Y(n23802) );
  NOR2x1_ASAP7_75t_SL U34780 ( .A(n22644), .B(mult_x_1196_n1577), .Y(
        mult_x_1196_n607) );
  INVx1_ASAP7_75t_SL U34781 ( .A(mult_x_1196_n1653), .Y(n23803) );
  MAJIxp5_ASAP7_75t_SL U34782 ( .A(mult_x_1196_n1184), .B(mult_x_1196_n1220), 
        .C(mult_x_1196_n1186), .Y(mult_x_1196_n1177) );
  XNOR2xp5_ASAP7_75t_SL U34783 ( .A(n23805), .B(mult_x_1196_n1184), .Y(n23804)
         );
  INVx1_ASAP7_75t_SL U34784 ( .A(mult_x_1196_n1220), .Y(n23805) );
  INVx1_ASAP7_75t_SL U34785 ( .A(mult_x_1196_n1091), .Y(n24096) );
  OR2x2_ASAP7_75t_SL U34786 ( .A(n24159), .B(n24160), .Y(n24163) );
  XNOR2xp5_ASAP7_75t_SL U34787 ( .A(mult_x_1196_n1936), .B(n23807), .Y(n23806)
         );
  NOR2x1_ASAP7_75t_SL U34788 ( .A(n23997), .B(mult_x_1196_n3118), .Y(n23812)
         );
  XNOR2xp5_ASAP7_75t_SL U34789 ( .A(n22212), .B(mult_x_1196_n1653), .Y(n23813)
         );
  XNOR2xp5_ASAP7_75t_SL U34790 ( .A(n23818), .B(n23815), .Y(mult_x_1196_n1641)
         );
  XOR2xp5_ASAP7_75t_SL U34791 ( .A(n23817), .B(n22735), .Y(n23815) );
  OAI21xp5_ASAP7_75t_SL U34792 ( .A1(mult_x_1196_n2995), .A2(n24014), .B(
        n22215), .Y(n23817) );
  INVx1_ASAP7_75t_SL U34793 ( .A(mult_x_1196_n2301), .Y(n23818) );
  XNOR2xp5_ASAP7_75t_SL U34794 ( .A(mult_x_1196_n1434), .B(mult_x_1196_n1472), 
        .Y(n23819) );
  XOR2xp5_ASAP7_75t_SL U34795 ( .A(n23821), .B(n23820), .Y(mult_x_1196_n1706)
         );
  INVx1_ASAP7_75t_SL U34796 ( .A(mult_x_1196_n2549), .Y(n23821) );
  MAJIxp5_ASAP7_75t_SL U34797 ( .A(n23822), .B(mult_x_1196_n2393), .C(
        mult_x_1196_n2549), .Y(mult_x_1196_n1705) );
  MAJIxp5_ASAP7_75t_SL U34798 ( .A(mult_x_1196_n2157), .B(n23824), .C(
        mult_x_1196_n2372), .Y(mult_x_1196_n1028) );
  XNOR2xp5_ASAP7_75t_SL U34799 ( .A(n23825), .B(n23823), .Y(mult_x_1196_n1029)
         );
  INVx1_ASAP7_75t_SL U34800 ( .A(mult_x_1196_n2372), .Y(n23825) );
  XOR2xp5_ASAP7_75t_SL U34801 ( .A(n23827), .B(n23826), .Y(mult_x_1196_n1217)
         );
  INVx1_ASAP7_75t_SL U34802 ( .A(mult_x_1196_n2443), .Y(n23826) );
  BUFx6f_ASAP7_75t_SL U34803 ( .A(n23849), .Y(n23830) );
  INVx3_ASAP7_75t_SL U34804 ( .A(n24688), .Y(n23849) );
  BUFx6f_ASAP7_75t_SL U34805 ( .A(n24688), .Y(n23831) );
  INVx1_ASAP7_75t_SL U34806 ( .A(u0_0_leon3x0_p0_iu_r_E__SHCNT__1_), .Y(n23835) );
  OAI22xp5_ASAP7_75t_SL U34807 ( .A1(n26514), .A2(n23830), .B1(n23831), .B2(
        n23836), .Y(u0_0_leon3x0_p0_muli[32]) );
  OR2x2_ASAP7_75t_SL U34808 ( .A(n23837), .B(n23831), .Y(n30603) );
  INVx1_ASAP7_75t_SL U34809 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__4_), .Y(n23837)
         );
  NAND2xp5_ASAP7_75t_SL U34810 ( .A(n23831), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__4_), .Y(n23838) );
  OAI22xp5_ASAP7_75t_SL U34811 ( .A1(n26562), .A2(n24689), .B1(n23831), .B2(
        n23840), .Y(u0_0_leon3x0_p0_muli[24]) );
  OAI22xp5_ASAP7_75t_SL U34812 ( .A1(n28425), .A2(n23849), .B1(n24688), .B2(
        n23842), .Y(u0_0_leon3x0_p0_muli[33]) );
  INVx1_ASAP7_75t_SL U34813 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__18_), .Y(n23844)
         );
  OAI21xp5_ASAP7_75t_SL U34814 ( .A1(n28720), .A2(n23849), .B(n28719), .Y(
        u0_0_leon3x0_p0_muli[18]) );
  OAI21xp5_ASAP7_75t_SL U34815 ( .A1(n30606), .A2(n23829), .B(n30605), .Y(
        u0_0_leon3x0_p0_muli[12]) );
  NOR2xp67_ASAP7_75t_SL U34816 ( .A(n24686), .B(n30574), .Y(n23850) );
  OAI22xp5_ASAP7_75t_SL U34817 ( .A1(n18537), .A2(mult_x_1196_n2992), .B1(
        mult_x_1196_n2991), .B2(n24012), .Y(n23851) );
  XNOR2xp5_ASAP7_75t_SL U34818 ( .A(n18916), .B(n23862), .Y(n23861) );
  INVx1_ASAP7_75t_SL U34819 ( .A(mult_x_1196_n1814), .Y(n23863) );
  NAND2x1_ASAP7_75t_SL U34820 ( .A(mult_x_1196_n2515), .B(mult_x_1196_n2675), 
        .Y(n24189) );
  OAI22x1_ASAP7_75t_SL U34821 ( .A1(n24002), .A2(mult_x_1196_n3090), .B1(
        n18920), .B2(mult_x_1196_n3091), .Y(mult_x_1196_n2515) );
  XNOR2x1_ASAP7_75t_SL U34822 ( .A(n28848), .B(n23529), .Y(mult_x_1196_n96) );
  MAJIxp5_ASAP7_75t_SL U34823 ( .A(mult_x_1196_n2294), .B(n23865), .C(
        mult_x_1196_n2230), .Y(mult_x_1196_n1381) );
  OAI22xp5_ASAP7_75t_SL U34824 ( .A1(mult_x_1196_n2764), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2763), .Y(n23865) );
  INVx1_ASAP7_75t_SL U34825 ( .A(n23870), .Y(n23867) );
  INVx1_ASAP7_75t_SL U34826 ( .A(mult_x_1196_n2548), .Y(n23868) );
  XNOR2xp5_ASAP7_75t_SL U34827 ( .A(mult_x_1196_n2580), .B(n23870), .Y(n23869)
         );
  NOR2x1_ASAP7_75t_SL U34828 ( .A(n24012), .B(mult_x_1196_n2995), .Y(n23872)
         );
  MAJIxp5_ASAP7_75t_SL U34829 ( .A(mult_x_1196_n2299), .B(mult_x_1196_n2485), 
        .C(n23876), .Y(mult_x_1196_n1569) );
  XNOR2xp5_ASAP7_75t_SL U34830 ( .A(n23922), .B(n23875), .Y(mult_x_1196_n1570)
         );
  XOR2xp5_ASAP7_75t_SL U34831 ( .A(n23876), .B(mult_x_1196_n2299), .Y(n23875)
         );
  OAI22xp5_ASAP7_75t_SL U34832 ( .A1(mult_x_1196_n2993), .A2(n23311), .B1(
        mult_x_1196_n2992), .B2(n24012), .Y(n23876) );
  MAJIxp5_ASAP7_75t_SL U34833 ( .A(mult_x_1196_n2395), .B(mult_x_1196_n2551), 
        .C(n23877), .Y(mult_x_1196_n1763) );
  INVx1_ASAP7_75t_SL U34834 ( .A(n23878), .Y(n23877) );
  OAI21xp5_ASAP7_75t_SL U34835 ( .A1(n28975), .A2(n28976), .B(n28853), .Y(
        n30631) );
  OAI21xp5_ASAP7_75t_SL U34836 ( .A1(uart1_uarto_SCALER__0_), .A2(n28174), .B(
        n28173), .Y(n28175) );
  NAND2xp5_ASAP7_75t_SL U34837 ( .A(n30177), .B(n30176), .Y(n3048) );
  AO21x1_ASAP7_75t_SL U34838 ( .A1(n22421), .A2(n23881), .B(n29099), .Y(n4285)
         );
  INVx1_ASAP7_75t_SL U34839 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUSEL__1_), .Y(
        n28965) );
  NAND2xp5_ASAP7_75t_SL U34840 ( .A(n31307), .B(n23885), .Y(n31311) );
  OA21x2_ASAP7_75t_SL U34841 ( .A1(n32258), .A2(n30182), .B(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__1_), .Y(n23882) );
  NAND2xp5_ASAP7_75t_SL U34842 ( .A(n30177), .B(n30171), .Y(n3049) );
  INVx1_ASAP7_75t_SL U34843 ( .A(n32811), .Y(n32815) );
  NOR2x1_ASAP7_75t_SL U34844 ( .A(timer0_N69), .B(n24354), .Y(n24358) );
  INVx1_ASAP7_75t_SL U34845 ( .A(n28981), .Y(n27108) );
  AO21x1_ASAP7_75t_SL U34846 ( .A1(n23229), .A2(n23883), .B(n29097), .Y(n4281)
         );
  NOR2x1_ASAP7_75t_SL U34847 ( .A(uart1_r_TRADDR__4_), .B(n27390), .Y(n27997)
         );
  NAND2xp5_ASAP7_75t_SL U34848 ( .A(n32564), .B(n32123), .Y(n31934) );
  OAI21xp5_ASAP7_75t_SL U34849 ( .A1(n25068), .A2(n25067), .B(n25066), .Y(
        n29912) );
  NAND2xp5_ASAP7_75t_SL U34850 ( .A(n30015), .B(n31034), .Y(n25066) );
  NAND2xp5_ASAP7_75t_SL U34851 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_), 
        .B(n18806), .Y(n30652) );
  INVx1_ASAP7_75t_SL U34852 ( .A(n26139), .Y(n25092) );
  NAND2xp5_ASAP7_75t_SL U34853 ( .A(add_x_735_n135), .B(add_x_735_n121), .Y(
        add_x_735_n115) );
  OAI21xp5_ASAP7_75t_SL U34854 ( .A1(n22228), .A2(add_x_735_n50), .B(
        add_x_735_n51), .Y(add_x_735_n49) );
  NAND2xp5_ASAP7_75t_SL U34855 ( .A(n31706), .B(n31734), .Y(n31743) );
  NAND2xp5_ASAP7_75t_SL U34856 ( .A(n32825), .B(n32824), .Y(n32831) );
  OAI21xp5_ASAP7_75t_SL U34857 ( .A1(add_x_735_n263), .A2(add_x_735_n259), .B(
        add_x_735_n260), .Y(add_x_735_n258) );
  NAND2xp5_ASAP7_75t_SL U34858 ( .A(add_x_735_n260), .B(add_x_735_n301), .Y(
        add_x_735_n32) );
  NAND2xp5_ASAP7_75t_SL U34859 ( .A(u0_0_leon3x0_p0_divi[2]), .B(n22449), .Y(
        add_x_735_n260) );
  NAND2xp5_ASAP7_75t_SL U34860 ( .A(DP_OP_5187J1_124_3275_n91), .B(
        DP_OP_5187J1_124_3275_n107), .Y(DP_OP_5187J1_124_3275_n6) );
  OAI21xp5_ASAP7_75t_SL U34861 ( .A1(n22225), .A2(DP_OP_5187J1_124_3275_n85), 
        .B(DP_OP_5187J1_124_3275_n86), .Y(DP_OP_5187J1_124_3275_n84) );
  OAI21xp5_ASAP7_75t_SL U34862 ( .A1(DP_OP_5187J1_124_3275_n190), .A2(n22225), 
        .B(DP_OP_5187J1_124_3275_n191), .Y(DP_OP_5187J1_124_3275_n189) );
  AOI21xp5_ASAP7_75t_SL U34863 ( .A1(add_x_735_n151), .A2(add_x_735_n168), .B(
        add_x_735_n152), .Y(add_x_735_n150) );
  NAND2xp5_ASAP7_75t_SL U34864 ( .A(n18909), .B(add_x_735_A_2_), .Y(
        add_x_735_n267) );
  NAND2xp5_ASAP7_75t_SL U34865 ( .A(add_x_735_n167), .B(add_x_735_n185), .Y(
        add_x_735_n165) );
  AOI21xp5_ASAP7_75t_SL U34866 ( .A1(n31845), .A2(timer0_res_19_), .B(n26545), 
        .Y(n26546) );
  AOI21xp5_ASAP7_75t_SL U34867 ( .A1(n31845), .A2(timer0_res_24_), .B(n26518), 
        .Y(n26519) );
  AOI21xp5_ASAP7_75t_SL U34868 ( .A1(n31845), .A2(timer0_res_26_), .B(n26499), 
        .Y(n26500) );
  AOI21xp5_ASAP7_75t_SL U34869 ( .A1(n31845), .A2(timer0_res_29_), .B(n26493), 
        .Y(n26494) );
  AOI21xp5_ASAP7_75t_SL U34870 ( .A1(n31845), .A2(timer0_res_23_), .B(n26531), 
        .Y(n26532) );
  AOI21xp5_ASAP7_75t_SL U34871 ( .A1(n31845), .A2(timer0_res_30_), .B(n26480), 
        .Y(n26481) );
  NAND2xp5_ASAP7_75t_SL U34872 ( .A(n29307), .B(n31352), .Y(n29239) );
  NAND2xp5_ASAP7_75t_SL U34873 ( .A(u0_0_leon3x0_p0_divi[0]), .B(n22999), .Y(
        add_x_735_n272) );
  INVx1_ASAP7_75t_SL U34874 ( .A(timer0_N82), .Y(n24408) );
  NAND2xp5_ASAP7_75t_SL U34875 ( .A(n29894), .B(n29893), .Y(n32575) );
  NAND2xp5_ASAP7_75t_SL U34876 ( .A(n28705), .B(n28704), .Y(n32587) );
  NAND2x1p5_ASAP7_75t_SL U34877 ( .A(n24120), .B(mult_x_1196_n3329), .Y(n24121) );
  OAI22xp5_ASAP7_75t_SL U34878 ( .A1(mult_x_1196_n3237), .A2(n23985), .B1(
        mult_x_1196_n3236), .B2(n24120), .Y(n24243) );
  OAI22xp5_ASAP7_75t_SL U34879 ( .A1(n24082), .A2(mult_x_1196_n3216), .B1(
        mult_x_1196_n3215), .B2(n22538), .Y(mult_x_1196_n2640) );
  NOR2xp33_ASAP7_75t_SL U34880 ( .A(mult_x_1196_n3243), .B(n23985), .Y(n24134)
         );
  OAI21xp5_ASAP7_75t_SL U34881 ( .A1(add_x_735_n108), .A2(n22228), .B(
        add_x_735_n109), .Y(add_x_735_n107) );
  NAND2xp5_ASAP7_75t_SL U34882 ( .A(n30713), .B(n30712), .Y(n32578) );
  AOI21x1_ASAP7_75t_SL U34883 ( .A1(n22274), .A2(
        u0_0_leon3x0_p0_iu_r_E__ALUCIN_), .B(add_x_735_n270), .Y(
        add_x_735_n268) );
  NAND2xp5_ASAP7_75t_SL U34884 ( .A(n22379), .B(n22431), .Y(n26188) );
  NAND2xp5_ASAP7_75t_SL U34885 ( .A(n26757), .B(n22379), .Y(n26354) );
  NAND2xp5_ASAP7_75t_SL U34886 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__7_), .B(
        n28769), .Y(n28768) );
  OAI21xp5_ASAP7_75t_SL U34887 ( .A1(add_x_735_n115), .A2(n22228), .B(
        add_x_735_n116), .Y(add_x_735_n114) );
  AO21x1_ASAP7_75t_SL U34888 ( .A1(n23229), .A2(n23884), .B(n27225), .Y(n4277)
         );
  XNOR2xp5_ASAP7_75t_SL U34889 ( .A(mult_x_1196_n271), .B(n22401), .Y(n23884)
         );
  OAI21xp5_ASAP7_75t_SL U34890 ( .A1(add_x_735_n213), .A2(add_x_735_n209), .B(
        add_x_735_n210), .Y(add_x_735_n204) );
  OAI21xp5_ASAP7_75t_SL U34891 ( .A1(add_x_735_n126), .A2(n22228), .B(
        add_x_735_n127), .Y(add_x_735_n125) );
  OAI21xp5_ASAP7_75t_SL U34892 ( .A1(n22228), .A2(add_x_735_n70), .B(
        add_x_735_n71), .Y(add_x_735_n69) );
  INVx1_ASAP7_75t_SL U34893 ( .A(add_x_735_n272), .Y(add_x_735_n270) );
  OAI21xp5_ASAP7_75t_SL U34894 ( .A1(n29816), .A2(n29815), .B(n29814), .Y(
        n30944) );
  NAND2xp5_ASAP7_75t_SL U34895 ( .A(n26484), .B(n25917), .Y(n29867) );
  NAND2xp5_ASAP7_75t_SL U34896 ( .A(n24716), .B(n24715), .Y(n24723) );
  NOR2x1_ASAP7_75t_SL U34897 ( .A(n24460), .B(n26302), .Y(
        u0_0_leon3x0_p0_divi[4]) );
  AOI21xp5_ASAP7_75t_SL U34898 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__12_), .A2(n22400), .B(
        n25427), .Y(n4756) );
  AOI21xp5_ASAP7_75t_SL U34899 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__6_), .A2(n22400), .B(n25856), .Y(n4713) );
  AOI21x1_ASAP7_75t_SL U34900 ( .A1(n29114), .A2(n24423), .B(n28378), .Y(
        n29017) );
  INVx1_ASAP7_75t_SL U34901 ( .A(n29017), .Y(n29019) );
  AOI21xp5_ASAP7_75t_SL U34902 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__9_), .A2(n22400), .B(n25411), .Y(n4558) );
  AOI21xp5_ASAP7_75t_SL U34903 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__27_), .A2(n22400), .B(
        n26343), .Y(n4529) );
  AOI21xp5_ASAP7_75t_SL U34904 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__0_), .A2(n22400), .B(n28101), .Y(n4367) );
  AOI21xp5_ASAP7_75t_SL U34905 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__28_), .A2(n22400), .B(
        n25434), .Y(n4595) );
  AOI21xp5_ASAP7_75t_SL U34906 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__13_), .A2(n22400), .B(
        n29994), .Y(n4661) );
  AOI21xp5_ASAP7_75t_SL U34907 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__21_), .A2(n22400), .B(
        n26330), .Y(n4383) );
  AOI21xp5_ASAP7_75t_SL U34908 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__5_), .A2(n22400), .B(n30011), .Y(n4745) );
  AOI21xp5_ASAP7_75t_SL U34909 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__24_), .A2(n22400), .B(
        n26510), .Y(n4512) );
  AOI21xp5_ASAP7_75t_SL U34910 ( .A1(n32739), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__1_), .B(n32738), .Y(n2970) );
  HB1xp67_ASAP7_75t_SL U34911 ( .A(n18883), .Y(n23885) );
  INVx1_ASAP7_75t_SL U34912 ( .A(n30190), .Y(n32121) );
  AOI21xp5_ASAP7_75t_SL U34913 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__31_), .A2(n22400), .B(
        n31041), .Y(n4773) );
  AOI21xp5_ASAP7_75t_SL U34914 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__10_), .A2(n22400), .B(
        n30994), .Y(n4454) );
  AOI21xp5_ASAP7_75t_SL U34915 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__31_), .B(n31689), .Y(n4485) );
  AOI21xp5_ASAP7_75t_SL U34916 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__24_), .B(n31777), .Y(n2978) );
  AOI21xp5_ASAP7_75t_SL U34917 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__25_), .B(n31785), .Y(n2977) );
  AOI21xp5_ASAP7_75t_SL U34918 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__26_), .B(n31781), .Y(n2976) );
  AOI21xp5_ASAP7_75t_SL U34919 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__28_), .B(n31773), .Y(n2974) );
  AOI21xp5_ASAP7_75t_SL U34920 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__25_), .A2(n22400), .B(
        n28407), .Y(n4622) );
  AOI21xp5_ASAP7_75t_SL U34921 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__16_), .B(n30535), .Y(n2985) );
  AOI21xp5_ASAP7_75t_SL U34922 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__17_), .B(n30542), .Y(n2984) );
  AOI21xp5_ASAP7_75t_SL U34923 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__19_), .B(n30830), .Y(n2983) );
  AOI21xp5_ASAP7_75t_SL U34924 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__14_), .B(n30512), .Y(n4651) );
  AOI21xp5_ASAP7_75t_SL U34925 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__15_), .B(n30519), .Y(n2986) );
  AOI21xp5_ASAP7_75t_SL U34926 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__14_), .A2(n22400), .B(
        n30558), .Y(n4430) );
  AOI21xp5_ASAP7_75t_SL U34927 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__2_), .A2(n22400), .B(n29565), .Y(n4673) );
  AOI21xp5_ASAP7_75t_SL U34928 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__13_), .B(n30528), .Y(n2987) );
  AOI21xp5_ASAP7_75t_SL U34929 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__20_), .B(n31771), .Y(n2982) );
  AOI21xp5_ASAP7_75t_SL U34930 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__23_), .B(n31764), .Y(n2979) );
  AOI21xp5_ASAP7_75t_SL U34931 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__3_), .A2(n22400), .B(n29506), .Y(n4693) );
  AOI21xp5_ASAP7_75t_SL U34932 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__21_), .B(n31767), .Y(n2981) );
  AOI21xp5_ASAP7_75t_SL U34933 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__29_), .B(n31692), .Y(n2973) );
  AOI21xp5_ASAP7_75t_SL U34934 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__20_), .A2(n22400), .B(
        n26963), .Y(n4500) );
  AOI21xp5_ASAP7_75t_SL U34935 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__23_), .A2(n22400), .B(
        n29908), .Y(n4417) );
  AOI21xp5_ASAP7_75t_SL U34936 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__19_), .A2(n22400), .B(
        n26538), .Y(n4361) );
  AO21x1_ASAP7_75t_SL U34937 ( .A1(mult_x_1196_n687), .A2(n22592), .B(
        mult_x_1196_n688), .Y(n23886) );
  AOI21xp5_ASAP7_75t_SL U34938 ( .A1(n32739), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__0_), .B(n32715), .Y(n2705) );
  OA21x2_ASAP7_75t_SL U34939 ( .A1(DP_OP_5187J1_124_3275_n262), .A2(
        DP_OP_5187J1_124_3275_n290), .B(DP_OP_5187J1_124_3275_n263), .Y(n23887) );
  AOI21xp5_ASAP7_75t_SL U34940 ( .A1(DP_OP_5187J1_124_3275_n264), .A2(
        DP_OP_5187J1_124_3275_n277), .B(DP_OP_5187J1_124_3275_n265), .Y(
        DP_OP_5187J1_124_3275_n263) );
  INVx1_ASAP7_75t_SL U34941 ( .A(n31988), .Y(n30499) );
  AND2x2_ASAP7_75t_SL U34942 ( .A(n25515), .B(n18883), .Y(n31637) );
  AOI21xp5_ASAP7_75t_SL U34943 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__22_), .B(n31775), .Y(n2980) );
  NAND2xp5_ASAP7_75t_SL U34944 ( .A(n18911), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__1_), .Y(n25188) );
  NAND2xp5_ASAP7_75t_SL U34945 ( .A(u0_0_leon3x0_p0_iu_fe_pc_3_), .B(
        u0_0_leon3x0_p0_iu_fe_pc_2_), .Y(add_x_746_n153) );
  NOR2x1_ASAP7_75t_SL U34946 ( .A(n26482), .B(n25130), .Y(n28821) );
  OR2x2_ASAP7_75t_SL U34947 ( .A(n23892), .B(n25517), .Y(n23890) );
  AND2x4_ASAP7_75t_SL U34948 ( .A(n23891), .B(n23890), .Y(n31632) );
  OR2x2_ASAP7_75t_SL U34949 ( .A(n22380), .B(n30916), .Y(n23891) );
  OR2x2_ASAP7_75t_SL U34950 ( .A(n25518), .B(n22380), .Y(n23892) );
  AOI21xp5_ASAP7_75t_SL U34951 ( .A1(n28878), .A2(n26341), .B(n28482), .Y(
        n28692) );
  OAI21xp5_ASAP7_75t_SL U34952 ( .A1(n23954), .A2(n22392), .B(n25763), .Y(
        n28878) );
  OAI21x1_ASAP7_75t_SL U34953 ( .A1(n31460), .A2(n32274), .B(n25410), .Y(
        n23893) );
  NOR2x1_ASAP7_75t_SL U34954 ( .A(n30509), .B(n24515), .Y(n25410) );
  INVx1_ASAP7_75t_SL U34955 ( .A(n25518), .Y(n31460) );
  AOI21xp5_ASAP7_75t_SL U34956 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__26_), .A2(n22400), .B(
        n26232), .Y(n4612) );
  AOI21xp5_ASAP7_75t_SL U34957 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__15_), .A2(n22400), .B(
        n31033), .Y(n4638) );
  AOI21xp5_ASAP7_75t_SL U34958 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__7_), .A2(n22400), .B(n29911), .Y(n4778) );
  AOI21xp5_ASAP7_75t_SL U34959 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__22_), .A2(n22400), .B(
        n26220), .Y(n4576) );
  AOI21xp5_ASAP7_75t_SL U34960 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__1_), .A2(n22400), .B(n27490), .Y(n4535) );
  AOI21xp5_ASAP7_75t_SL U34961 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__30_), .A2(n22400), .B(
        n30572), .Y(n4739) );
  AOI21xp5_ASAP7_75t_SL U34962 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__8_), .A2(n22400), .B(n29758), .Y(n4687) );
  AOI21xp5_ASAP7_75t_SL U34963 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__11_), .A2(n22400), .B(
        n28134), .Y(n4523) );
  AOI21xp5_ASAP7_75t_SL U34964 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__29_), .A2(n22400), .B(
        n26488), .Y(n4667) );
  AOI21xp5_ASAP7_75t_SL U34965 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__16_), .A2(n22400), .B(
        n26663), .Y(n4642) );
  AND3x2_ASAP7_75t_SL U34966 ( .A(n18883), .B(n24684), .C(n25521), .Y(n23894)
         );
  AOI21xp5_ASAP7_75t_SL U34967 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__4_), .A2(n22400), .B(n25870), .Y(n4767) );
  NAND2xp5_ASAP7_75t_SL U34968 ( .A(add_x_746_n36), .B(add_x_746_n58), .Y(
        add_x_746_n2) );
  NAND2xp5_ASAP7_75t_SL U34969 ( .A(add_x_746_n34), .B(n18880), .Y(
        add_x_746_n33) );
  NOR2x1_ASAP7_75t_SL U34970 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__2_), .B(
        n26732), .Y(n31868) );
  NOR2x1_ASAP7_75t_SL U34971 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[36]), .Y(
        n25125) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U34972 ( .A1(u0_0_leon3x0_p0_divi[30]), .A2(
        n28931), .B(n25131), .C(n18530), .Y(n25132) );
  NAND2xp5_ASAP7_75t_SL U34973 ( .A(n26207), .B(n26206), .Y(n32581) );
  NAND2xp5_ASAP7_75t_SL U34974 ( .A(u0_0_leon3x0_p0_div0_vaddin1[10]), .B(
        u0_0_leon3x0_p0_div0_b[10]), .Y(DP_OP_5187J1_124_3275_n245) );
  NAND2xp5_ASAP7_75t_SL U34975 ( .A(n28696), .B(n28695), .Y(n30972) );
  AOI21xp5_ASAP7_75t_SL U34976 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__18_), .B(n31836), .Y(n2569) );
  AOI21xp5_ASAP7_75t_SL U34977 ( .A1(n22381), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__27_), .B(n31788), .Y(n2975) );
  NAND2xp5_ASAP7_75t_SL U34978 ( .A(n32001), .B(n32000), .Y(n18045) );
  NAND2xp5_ASAP7_75t_SL U34979 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__30_), 
        .B(n22381), .Y(n32000) );
  AOI21xp5_ASAP7_75t_SL U34980 ( .A1(DP_OP_1196_128_7433_n345), .A2(
        DP_OP_1196_128_7433_n353), .B(DP_OP_1196_128_7433_n346), .Y(
        DP_OP_1196_128_7433_n2) );
  NAND2xp5_ASAP7_75t_SL U34981 ( .A(n30958), .B(n30962), .Y(n28536) );
  OAI21xp5_ASAP7_75t_SL U34982 ( .A1(DP_OP_5187J1_124_3275_n191), .A2(
        DP_OP_5187J1_124_3275_n187), .B(DP_OP_5187J1_124_3275_n188), .Y(
        DP_OP_5187J1_124_3275_n182) );
  NAND2xp5_ASAP7_75t_SL U34983 ( .A(u0_0_leon3x0_p0_div0_vaddin1[16]), .B(
        u0_0_leon3x0_p0_div0_b[16]), .Y(DP_OP_5187J1_124_3275_n191) );
  AO21x1_ASAP7_75t_SL U34984 ( .A1(n22421), .A2(n23895), .B(n27038), .Y(n4267)
         );
  OAI21xp5_ASAP7_75t_SL U34985 ( .A1(add_x_735_n165), .A2(add_x_735_n214), .B(
        add_x_735_n166), .Y(add_x_735_n164) );
  AOI21xp5_ASAP7_75t_SL U34986 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__18_), .A2(n22400), .B(
        n25714), .Y(n4357) );
  AOI21xp5_ASAP7_75t_SL U34987 ( .A1(n31637), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__0_), .B(n28107), .Y(n4366)
         );
  INVx1_ASAP7_75t_SL U34988 ( .A(DP_OP_5187J1_124_3275_n299), .Y(
        DP_OP_5187J1_124_3275_n298) );
  OAI21xp5_ASAP7_75t_SL U34989 ( .A1(n24317), .A2(DP_OP_5187J1_124_3275_n300), 
        .B(DP_OP_5187J1_124_3275_n301), .Y(DP_OP_5187J1_124_3275_n299) );
  AOI21xp5_ASAP7_75t_SL U34990 ( .A1(DP_OP_5187J1_124_3275_n129), .A2(
        DP_OP_5187J1_124_3275_n146), .B(DP_OP_5187J1_124_3275_n130), .Y(
        DP_OP_5187J1_124_3275_n128) );
  NAND2xp5_ASAP7_75t_SL U34991 ( .A(DP_OP_5187J1_124_3275_n227), .B(
        DP_OP_5187J1_124_3275_n327), .Y(DP_OP_5187J1_124_3275_n27) );
  NAND2xp5_ASAP7_75t_SL U34992 ( .A(u0_0_leon3x0_p0_div0_vaddin1[12]), .B(
        u0_0_leon3x0_p0_div0_b[12]), .Y(DP_OP_5187J1_124_3275_n227) );
  NAND2xp5_ASAP7_75t_SL U34993 ( .A(n32824), .B(n32789), .Y(n32821) );
  HB1xp67_ASAP7_75t_SL U34994 ( .A(n24381), .Y(n23896) );
  NOR2x1_ASAP7_75t_SL U34995 ( .A(DP_OP_5187J1_124_3275_n127), .B(
        DP_OP_5187J1_124_3275_n161), .Y(DP_OP_5187J1_124_3275_n4) );
  NOR2x1_ASAP7_75t_SL U34996 ( .A(n28987), .B(n30635), .Y(n29605) );
  OAI21xp5_ASAP7_75t_SL U34997 ( .A1(n22380), .A2(n32246), .B(n25401), .Y(
        n31042) );
  AOI21xp5_ASAP7_75t_SL U34998 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__17_), .A2(n22400), .B(
        n27248), .Y(n4035) );
  OAI21xp5_ASAP7_75t_SL U34999 ( .A1(DP_OP_5187J1_124_3275_n288), .A2(
        DP_OP_5187J1_124_3275_n282), .B(DP_OP_5187J1_124_3275_n283), .Y(
        DP_OP_5187J1_124_3275_n277) );
  NAND2xp5_ASAP7_75t_SL U35000 ( .A(u0_0_leon3x0_p0_div0_vaddin1[4]), .B(
        u0_0_leon3x0_p0_div0_b[4]), .Y(DP_OP_5187J1_124_3275_n288) );
  OAI21xp5_ASAP7_75t_SL U35001 ( .A1(DP_OP_5187J1_124_3275_n179), .A2(n22225), 
        .B(DP_OP_5187J1_124_3275_n180), .Y(DP_OP_5187J1_124_3275_n178) );
  INVx1_ASAP7_75t_SL U35002 ( .A(timer0_N85), .Y(n24411) );
  OAI21xp5_ASAP7_75t_SL U35003 ( .A1(n32642), .A2(n18851), .B(n31546), .Y(
        n30160) );
  NOR2x1_ASAP7_75t_SL U35004 ( .A(n24547), .B(n30160), .Y(n30189) );
  NOR2x1_ASAP7_75t_SL U35005 ( .A(n28987), .B(n29609), .Y(n28742) );
  INVx1_ASAP7_75t_SL U35006 ( .A(n28921), .Y(n28764) );
  OAI21xp5_ASAP7_75t_SL U35007 ( .A1(n22428), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N25), .B(n29080), .Y(n4265) );
  AOI21xp5_ASAP7_75t_SL U35008 ( .A1(n31637), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__7_), .B(n29941), .Y(n4777)
         );
  AOI21xp5_ASAP7_75t_SL U35009 ( .A1(n31637), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__4_), .B(n25876), .Y(n4766)
         );
  NAND2xp5_ASAP7_75t_SL U35010 ( .A(n32764), .B(n32763), .Y(n32782) );
  NAND2xp5_ASAP7_75t_SL U35011 ( .A(n32816), .B(n32803), .Y(n32810) );
  INVx1_ASAP7_75t_SL U35012 ( .A(n32816), .Y(n32808) );
  AOI21xp5_ASAP7_75t_SL U35013 ( .A1(n31637), .A2(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__6_), .B(n25862), .Y(n4712)
         );
  NAND2xp5_ASAP7_75t_SL U35014 ( .A(add_x_735_n203), .B(add_x_735_n189), .Y(
        add_x_735_n183) );
  OAI21xp5_ASAP7_75t_SL U35015 ( .A1(add_x_735_n181), .A2(add_x_735_n173), .B(
        add_x_735_n174), .Y(add_x_735_n168) );
  OAI21xp5_ASAP7_75t_SL U35016 ( .A1(add_x_735_n97), .A2(n22228), .B(
        add_x_735_n98), .Y(add_x_735_n96) );
  OAI21xp5_ASAP7_75t_SL U35017 ( .A1(n25234), .A2(n18838), .B(n24794), .Y(
        n32179) );
  NAND2xp5_ASAP7_75t_SL U35018 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_), 
        .B(n24796), .Y(n24794) );
  INVx1_ASAP7_75t_SL U35019 ( .A(mult_x_1196_n2456), .Y(mult_x_1196_n1666) );
  OAI21xp5_ASAP7_75t_SL U35020 ( .A1(mult_x_1196_n692), .A2(n22401), .B(
        mult_x_1196_n693), .Y(mult_x_1196_n691) );
  AOI21xp5_ASAP7_75t_SL U35021 ( .A1(DP_OP_5187J1_124_3275_n235), .A2(
        DP_OP_5187J1_124_3275_n250), .B(DP_OP_5187J1_124_3275_n236), .Y(
        DP_OP_5187J1_124_3275_n230) );
  NAND2xp5_ASAP7_75t_SL U35022 ( .A(n26322), .B(n26321), .Y(n31947) );
  AO21x1_ASAP7_75t_SL U35023 ( .A1(n23229), .A2(n23897), .B(n26913), .Y(n4255)
         );
  NAND2xp5_ASAP7_75t_SL U35024 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__2_), .B(
        n24809), .Y(n24810) );
  NAND2xp5_ASAP7_75t_SL U35025 ( .A(n25005), .B(n26854), .Y(n24748) );
  NAND2xp5_ASAP7_75t_SL U35026 ( .A(n24373), .B(n24414), .Y(n24378) );
  NOR3xp33_ASAP7_75t_SL U35027 ( .A(n24333), .B(timer0_N77), .C(timer0_N78), 
        .Y(n24339) );
  INVx5_ASAP7_75t_SL U35028 ( .A(n22933), .Y(n23952) );
  OAI21xp5_ASAP7_75t_SL U35029 ( .A1(mult_x_1196_n718), .A2(mult_x_1196_n730), 
        .B(mult_x_1196_n719), .Y(mult_x_1196_n717) );
  NAND2xp5_ASAP7_75t_SL U35030 ( .A(mult_x_1196_n2002), .B(mult_x_1196_n2001), 
        .Y(mult_x_1196_n712) );
  NAND2xp5_ASAP7_75t_SL U35031 ( .A(n24694), .B(n28119), .Y(n30779) );
  NAND2xp5_ASAP7_75t_SL U35032 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__12_), .B(
        n24689), .Y(n28622) );
  NAND2xp5_ASAP7_75t_SL U35033 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__26_), .B(
        n23849), .Y(n25483) );
  NAND2xp5_ASAP7_75t_SL U35034 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__1_), .B(
        n24689), .Y(n30605) );
  NAND2xp5_ASAP7_75t_SL U35035 ( .A(u0_0_leon3x0_p0_iu_r_E__OP2__8_), .B(
        n23849), .Y(n28719) );
  AOI21xp5_ASAP7_75t_SL U35036 ( .A1(n23886), .A2(mult_x_1196_n819), .B(
        mult_x_1196_n682), .Y(mult_x_1196_n680) );
  O2A1O1Ixp5_ASAP7_75t_SL U35037 ( .A1(n31857), .A2(n26817), .B(n24772), .C(
        n26818), .Y(n23899) );
  AO21x1_ASAP7_75t_SL U35038 ( .A1(n22421), .A2(n23900), .B(n28278), .Y(n4253)
         );
  OAI21xp5_ASAP7_75t_SL U35039 ( .A1(n30339), .A2(n22376), .B(n25166), .Y(
        n28574) );
  AO21x1_ASAP7_75t_SL U35040 ( .A1(n23229), .A2(n23901), .B(n29024), .Y(n4251)
         );
  XOR2xp5_ASAP7_75t_SL U35041 ( .A(mult_x_1196_n258), .B(mult_x_1196_n615), 
        .Y(n23901) );
  NAND2xp5_ASAP7_75t_SL U35042 ( .A(n23002), .B(u0_0_leon3x0_p0_divi[23]), .Y(
        add_x_735_n106) );
  FAx1_ASAP7_75t_SL U35043 ( .A(mult_x_1196_n2668), .B(mult_x_1196_n2700), 
        .CI(mult_x_1196_n2636), .CON(mult_x_1196_n2089), .SN(mult_x_1196_n2090) );
  OAI22xp5_ASAP7_75t_SL U35044 ( .A1(mult_x_1196_n3276), .A2(n23981), .B1(
        n23980), .B2(mult_x_1196_n3275), .Y(mult_x_1196_n2700) );
  INVx1_ASAP7_75t_SL U35045 ( .A(add_x_735_n265), .Y(add_x_735_n264) );
  OAI21xp5_ASAP7_75t_SL U35046 ( .A1(DP_OP_5187J1_124_3275_n258), .A2(n23887), 
        .B(DP_OP_5187J1_124_3275_n259), .Y(DP_OP_5187J1_124_3275_n257) );
  OAI21xp5_ASAP7_75t_SL U35047 ( .A1(n18381), .A2(n25198), .B(n25194), .Y(
        n26377) );
  OAI21xp5_ASAP7_75t_SL U35048 ( .A1(n29561), .A2(n25198), .B(n25107), .Y(
        n26390) );
  AOI21xp5_ASAP7_75t_SL U35049 ( .A1(DP_OP_5187J1_124_3275_n91), .A2(
        DP_OP_5187J1_124_3275_n108), .B(DP_OP_5187J1_124_3275_n92), .Y(
        DP_OP_5187J1_124_3275_n5) );
  INVx1_ASAP7_75t_SL U35050 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__0_), .Y(
        n31961) );
  NAND2xp5_ASAP7_75t_SL U35051 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__CNT__1_), 
        .B(n31961), .Y(n32141) );
  NAND2xp5_ASAP7_75t_SL U35052 ( .A(n18911), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__10_), .Y(n25108) );
  BUFx6f_ASAP7_75t_SL U35053 ( .A(u0_0_leon3x0_p0_iu_r_E__LDBP1_), .Y(n24685)
         );
  NAND2xp5_ASAP7_75t_SL U35054 ( .A(n26074), .B(n27473), .Y(n30872) );
  NAND2xp5_ASAP7_75t_SL U35055 ( .A(n31531), .B(n27316), .Y(n26080) );
  NAND2xp5_ASAP7_75t_SL U35056 ( .A(n26909), .B(n26908), .Y(n26955) );
  AOI22xp5_ASAP7_75t_SL U35057 ( .A1(n27521), .A2(n29746), .B1(
        uart1_r_RCNT__3_), .B2(n27511), .Y(n29982) );
  NAND2xp5_ASAP7_75t_SL U35058 ( .A(n31503), .B(n27503), .Y(n27511) );
  XNOR2x2_ASAP7_75t_SL U35059 ( .A(n24064), .B(n23957), .Y(mult_x_1196_n3199)
         );
  XNOR2xp5_ASAP7_75t_SL U35060 ( .A(mult_x_1196_n253), .B(mult_x_1196_n580), 
        .Y(n23907) );
  NAND2xp5_ASAP7_75t_SL U35061 ( .A(n22436), .B(u0_0_leon3x0_p0_divi[21]), .Y(
        add_x_735_n124) );
  AO21x1_ASAP7_75t_SL U35062 ( .A1(n22421), .A2(n23904), .B(n29093), .Y(n4271)
         );
  XNOR2xp5_ASAP7_75t_SL U35063 ( .A(mult_x_1196_n268), .B(mult_x_1196_n680), 
        .Y(n23904) );
  AO21x1_ASAP7_75t_SL U35064 ( .A1(n22421), .A2(n23905), .B(n27026), .Y(n4269)
         );
  XNOR2xp5_ASAP7_75t_SL U35065 ( .A(mult_x_1196_n267), .B(mult_x_1196_n675), 
        .Y(n23905) );
  AO21x1_ASAP7_75t_SL U35066 ( .A1(n23229), .A2(n23906), .B(n29085), .Y(n4249)
         );
  XOR2xp5_ASAP7_75t_SL U35067 ( .A(mult_x_1196_n257), .B(n18899), .Y(n23906)
         );
  AOI21xp5_ASAP7_75t_SL U35068 ( .A1(n23929), .A2(mult_x_1196_n807), .B(
        mult_x_1196_n606), .Y(mult_x_1196_n604) );
  AOI21xp5_ASAP7_75t_SL U35069 ( .A1(n23929), .A2(n18580), .B(n23919), .Y(
        mult_x_1196_n595) );
  AO21x1_ASAP7_75t_SL U35070 ( .A1(n22421), .A2(n23907), .B(n25272), .Y(n4241)
         );
  OAI21xp5_ASAP7_75t_SL U35071 ( .A1(mult_x_1196_n616), .A2(mult_x_1196_n629), 
        .B(n18535), .Y(mult_x_1196_n615) );
  NAND2xp5_ASAP7_75t_SL U35072 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), 
        .B(n32094), .Y(n24772) );
  INVx1_ASAP7_75t_SL U35073 ( .A(mult_x_1196_n2645), .Y(n24162) );
  INVx1_ASAP7_75t_SL U35074 ( .A(n25574), .Y(n30196) );
  AOI21xp5_ASAP7_75t_SL U35075 ( .A1(n23929), .A2(mult_x_1196_n589), .B(
        mult_x_1196_n590), .Y(mult_x_1196_n588) );
  AND2x2_ASAP7_75t_SL U35076 ( .A(n18516), .B(mult_x_1196_n802), .Y(n23908) );
  NAND2xp5_ASAP7_75t_SL U35077 ( .A(n24789), .B(n24796), .Y(n24790) );
  OAI21xp5_ASAP7_75t_SL U35078 ( .A1(n23902), .A2(mult_x_1196_n654), .B(n22510), .Y(mult_x_1196_n653) );
  OAI21xp5_ASAP7_75t_SL U35079 ( .A1(mult_x_1196_n661), .A2(n23902), .B(n24122), .Y(mult_x_1196_n660) );
  OAI21xp5_ASAP7_75t_SL U35080 ( .A1(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .A2(
        n32186), .B(n24777), .Y(n24779) );
  NAND2xp5_ASAP7_75t_SL U35081 ( .A(n30180), .B(n30162), .Y(n30177) );
  OAI21xp5_ASAP7_75t_SL U35082 ( .A1(n23938), .A2(mult_x_1196_n580), .B(
        mult_x_1196_n568), .Y(mult_x_1196_n566) );
  INVx1_ASAP7_75t_SL U35083 ( .A(n31992), .Y(n30497) );
  NAND2xp5_ASAP7_75t_SL U35084 ( .A(n24681), .B(n31828), .Y(n31992) );
  AO21x1_ASAP7_75t_SL U35085 ( .A1(n22421), .A2(n23909), .B(n26349), .Y(n4243)
         );
  XNOR2xp5_ASAP7_75t_SL U35086 ( .A(mult_x_1196_n254), .B(mult_x_1196_n588), 
        .Y(n23909) );
  AO21x1_ASAP7_75t_SL U35087 ( .A1(n23229), .A2(n23910), .B(n29083), .Y(n4247)
         );
  XNOR2xp5_ASAP7_75t_SL U35088 ( .A(mult_x_1196_n256), .B(mult_x_1196_n604), 
        .Y(n23910) );
  AO21x1_ASAP7_75t_SL U35089 ( .A1(n22421), .A2(n23911), .B(n30608), .Y(n4245)
         );
  XNOR2xp5_ASAP7_75t_SL U35090 ( .A(mult_x_1196_n255), .B(mult_x_1196_n595), 
        .Y(n23911) );
  NAND2xp5_ASAP7_75t_SL U35091 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__16_), .B(
        n24687), .Y(n25093) );
  BUFx2_ASAP7_75t_SL U35092 ( .A(u0_0_leon3x0_p0_muli[43]), .Y(add_x_735_A_9_)
         );
  OAI21xp5_ASAP7_75t_SL U35093 ( .A1(n28720), .A2(n24686), .B(n25098), .Y(
        u0_0_leon3x0_p0_muli[43]) );
  OAI21xp5_ASAP7_75t_SL U35094 ( .A1(mult_x_1196_n578), .A2(mult_x_1196_n580), 
        .B(mult_x_1196_n579), .Y(mult_x_1196_n577) );
  AOI21x1_ASAP7_75t_SL U35095 ( .A1(add_x_735_n257), .A2(add_x_735_n265), .B(
        add_x_735_n258), .Y(add_x_735_n256) );
  INVx1_ASAP7_75t_SL U35096 ( .A(add_x_735_n253), .Y(add_x_735_n252) );
  OAI21xp5_ASAP7_75t_SL U35097 ( .A1(mult_x_1196_n560), .A2(mult_x_1196_n580), 
        .B(mult_x_1196_n561), .Y(mult_x_1196_n559) );
  OAI21xp5_ASAP7_75t_SL U35098 ( .A1(n30905), .A2(n24796), .B(n24795), .Y(
        n32178) );
  NAND2xp5_ASAP7_75t_SL U35099 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__5_), .B(
        n23903), .Y(n25192) );
  NAND2xp5_ASAP7_75t_SL U35100 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__13_), .B(
        n18862), .Y(n25195) );
  NAND2xp5_ASAP7_75t_SL U35101 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__1_), .B(
        n23903), .Y(n25187) );
  NAND2xp5_ASAP7_75t_SL U35102 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__9_), .B(
        n23903), .Y(n25199) );
  NAND2xp5_ASAP7_75t_SL U35103 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__29_), .B(
        n18862), .Y(n24545) );
  NAND2xp5_ASAP7_75t_SL U35104 ( .A(n30603), .B(n28820), .Y(
        u0_0_leon3x0_p0_divi[3]) );
  OAI22xp5_ASAP7_75t_SL U35105 ( .A1(mult_x_1196_n2797), .A2(n24038), .B1(
        mult_x_1196_n2796), .B2(n22391), .Y(mult_x_1196_n2231) );
  OAI22xp5_ASAP7_75t_SL U35106 ( .A1(mult_x_1196_n2927), .A2(n24022), .B1(
        mult_x_1196_n2926), .B2(n24020), .Y(mult_x_1196_n2355) );
  NAND2xp5_ASAP7_75t_SL U35107 ( .A(mult_x_1196_n464), .B(mult_x_1196_n385), 
        .Y(n23915) );
  OR2x2_ASAP7_75t_SL U35108 ( .A(n23915), .B(n23916), .Y(mult_x_1196_n350) );
  OR2x2_ASAP7_75t_SL U35109 ( .A(n22406), .B(mult_x_1196_n361), .Y(n23916) );
  BUFx2_ASAP7_75t_SL U35110 ( .A(mult_x_1196_n1144), .Y(n23917) );
  INVx1_ASAP7_75t_SL U35111 ( .A(DP_OP_5187J1_124_3275_n290), .Y(
        DP_OP_5187J1_124_3275_n289) );
  AOI21xp5_ASAP7_75t_SL U35112 ( .A1(DP_OP_5187J1_124_3275_n291), .A2(
        DP_OP_5187J1_124_3275_n299), .B(DP_OP_5187J1_124_3275_n292), .Y(
        DP_OP_5187J1_124_3275_n290) );
  AOI21xp5_ASAP7_75t_SL U35113 ( .A1(DP_OP_5187J1_124_3275_n289), .A2(
        DP_OP_5187J1_124_3275_n335), .B(DP_OP_5187J1_124_3275_n286), .Y(
        DP_OP_5187J1_124_3275_n284) );
  OAI22xp5_ASAP7_75t_SL U35114 ( .A1(mult_x_1196_n3260), .A2(n23982), .B1(
        n22389), .B2(mult_x_1196_n3259), .Y(mult_x_1196_n2684) );
  OAI22xp5_ASAP7_75t_SL U35115 ( .A1(mult_x_1196_n3073), .A2(n24007), .B1(
        n24005), .B2(mult_x_1196_n3072), .Y(mult_x_1196_n2501) );
  INVx1_ASAP7_75t_SL U35116 ( .A(mult_x_1196_n2560), .Y(mult_x_1196_n1959) );
  OAI22xp5_ASAP7_75t_SL U35117 ( .A1(mult_x_1196_n3048), .A2(n24007), .B1(
        n24005), .B2(mult_x_1196_n3047), .Y(mult_x_1196_n2476) );
  NAND2xp5_ASAP7_75t_SL U35118 ( .A(n24311), .B(mult_x_1196_n1191), .Y(
        mult_x_1196_n520) );
  OAI21xp5_ASAP7_75t_SL U35119 ( .A1(mult_x_1196_n529), .A2(mult_x_1196_n519), 
        .B(mult_x_1196_n520), .Y(mult_x_1196_n518) );
  OAI22xp5_ASAP7_75t_SL U35120 ( .A1(mult_x_1196_n2931), .A2(n22781), .B1(
        mult_x_1196_n2930), .B2(n24020), .Y(mult_x_1196_n2359) );
  NAND2xp5_ASAP7_75t_SL U35121 ( .A(n31405), .B(n22220), .Y(
        u0_0_leon3x0_p0_muli[11]) );
  NOR2x1_ASAP7_75t_SL U35122 ( .A(n24282), .B(mult_x_1196_n1225), .Y(
        mult_x_1196_n526) );
  HB1xp67_ASAP7_75t_SL U35123 ( .A(mult_x_1196_n597), .Y(n23919) );
  OAI22xp5_ASAP7_75t_SL U35124 ( .A1(mult_x_1196_n3171), .A2(n24230), .B1(
        n23992), .B2(mult_x_1196_n3170), .Y(mult_x_1196_n2595) );
  OAI22xp5_ASAP7_75t_SL U35125 ( .A1(mult_x_1196_n2923), .A2(n24022), .B1(
        mult_x_1196_n2922), .B2(n24020), .Y(mult_x_1196_n2351) );
  OAI22xp5_ASAP7_75t_SL U35126 ( .A1(mult_x_1196_n2795), .A2(n24038), .B1(
        mult_x_1196_n2794), .B2(n22391), .Y(mult_x_1196_n2229) );
  OAI22xp5_ASAP7_75t_SL U35127 ( .A1(mult_x_1196_n2786), .A2(n22509), .B1(
        mult_x_1196_n2785), .B2(n22936), .Y(mult_x_1196_n2220) );
  INVx1_ASAP7_75t_SL U35128 ( .A(mult_x_1196_n2444), .Y(mult_x_1196_n1243) );
  OAI22xp5_ASAP7_75t_SL U35129 ( .A1(n23116), .A2(mult_x_1196_n2896), .B1(
        mult_x_1196_n2895), .B2(n24025), .Y(mult_x_1196_n2324) );
  OAI22xp5_ASAP7_75t_SL U35130 ( .A1(mult_x_1196_n2952), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2951), .Y(mult_x_1196_n2380) );
  OAI22xp5_ASAP7_75t_SL U35131 ( .A1(mult_x_1196_n2796), .A2(n24038), .B1(
        mult_x_1196_n2795), .B2(n22391), .Y(mult_x_1196_n2230) );
  OAI22xp5_ASAP7_75t_SL U35132 ( .A1(mult_x_1196_n2852), .A2(n24031), .B1(
        n24030), .B2(mult_x_1196_n2851), .Y(mult_x_1196_n2286) );
  NAND2xp5_ASAP7_75t_SL U35133 ( .A(n22262), .B(n24077), .Y(n24112) );
  OR2x2_ASAP7_75t_SL U35134 ( .A(n24149), .B(n24150), .Y(n23925) );
  INVx1_ASAP7_75t_SL U35135 ( .A(n24270), .Y(n24149) );
  NAND2xp5_ASAP7_75t_SL U35136 ( .A(n23154), .B(u0_0_leon3x0_p0_divi[13]), .Y(
        add_x_735_n192) );
  OAI21xp5_ASAP7_75t_SL U35137 ( .A1(add_x_735_n183), .A2(add_x_735_n214), .B(
        add_x_735_n184), .Y(add_x_735_n182) );
  AOI21xp5_ASAP7_75t_SL U35138 ( .A1(add_x_735_n189), .A2(add_x_735_n204), .B(
        add_x_735_n190), .Y(add_x_735_n184) );
  OAI22xp5_ASAP7_75t_SL U35139 ( .A1(mult_x_1196_n2746), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2745), .Y(mult_x_1196_n2183) );
  NOR2x1_ASAP7_75t_SL U35140 ( .A(mult_x_1196_n1614), .B(mult_x_1196_n1613), 
        .Y(mult_x_1196_n613) );
  NAND2xp5_ASAP7_75t_SL U35141 ( .A(add_x_735_A_10_), .B(n18890), .Y(
        add_x_735_n228) );
  NOR2x1_ASAP7_75t_SL U35142 ( .A(add_x_735_A_10_), .B(n18890), .Y(
        add_x_735_n225) );
  OAI22xp5_ASAP7_75t_SL U35143 ( .A1(mult_x_1196_n2774), .A2(n18341), .B1(
        mult_x_1196_n2773), .B2(n22481), .Y(mult_x_1196_n875) );
  FAx1_ASAP7_75t_SL U35144 ( .A(mult_x_1196_n885), .B(mult_x_1196_n875), .CI(
        mult_x_1196_n883), .CON(mult_x_1196_n871), .SN(mult_x_1196_n872) );
  FAx1_ASAP7_75t_SL U35145 ( .A(mult_x_1196_n2148), .B(mult_x_1196_n2211), 
        .CI(mult_x_1196_n2273), .CON(mult_x_1196_n883), .SN(mult_x_1196_n884)
         );
  OAI22xp5_ASAP7_75t_SL U35146 ( .A1(n24020), .A2(mult_x_1196_n2907), .B1(
        mult_x_1196_n2908), .B2(n24022), .Y(mult_x_1196_n2336) );
  OAI22xp5_ASAP7_75t_SL U35147 ( .A1(mult_x_1196_n2914), .A2(n22781), .B1(
        mult_x_1196_n2913), .B2(n24020), .Y(mult_x_1196_n2342) );
  BUFx6f_ASAP7_75t_SL U35148 ( .A(mult_x_1196_n99), .Y(n24021) );
  OAI22xp5_ASAP7_75t_SL U35149 ( .A1(mult_x_1196_n2946), .A2(n22779), .B1(
        n22694), .B2(mult_x_1196_n2945), .Y(mult_x_1196_n2374) );
  NAND2xp5_ASAP7_75t_SL U35150 ( .A(n24291), .B(mult_x_1196_n829), .Y(n24196)
         );
  NOR2x1_ASAP7_75t_SL U35151 ( .A(n24133), .B(n24134), .Y(n24135) );
  OAI22xp5_ASAP7_75t_SL U35152 ( .A1(mult_x_1196_n2784), .A2(n22412), .B1(
        mult_x_1196_n2783), .B2(n22391), .Y(mult_x_1196_n2218) );
  INVx1_ASAP7_75t_SL U35153 ( .A(mult_x_1196_n1033), .Y(mult_x_1196_n1021) );
  OAI22xp5_ASAP7_75t_SL U35154 ( .A1(mult_x_1196_n2788), .A2(n24038), .B1(
        mult_x_1196_n2787), .B2(n22936), .Y(mult_x_1196_n2222) );
  OAI22xp5_ASAP7_75t_SL U35155 ( .A1(mult_x_1196_n3222), .A2(n23985), .B1(
        mult_x_1196_n3221), .B2(n23984), .Y(mult_x_1196_n2646) );
  OAI22xp5_ASAP7_75t_SL U35156 ( .A1(mult_x_1196_n3039), .A2(n22563), .B1(
        mult_x_1196_n3038), .B2(n22540), .Y(mult_x_1196_n2467) );
  HB1xp67_ASAP7_75t_SL U35157 ( .A(mult_x_1196_n1793), .Y(n23930) );
  OAI22xp5_ASAP7_75t_SL U35158 ( .A1(mult_x_1196_n3275), .A2(n23982), .B1(
        n23980), .B2(mult_x_1196_n3274), .Y(mult_x_1196_n2699) );
  NAND2xp5_ASAP7_75t_SL U35159 ( .A(n31001), .B(n25025), .Y(n25023) );
  NAND2xp5_ASAP7_75t_SL U35160 ( .A(dc_q[31]), .B(n31004), .Y(n25036) );
  AOI21xp5_ASAP7_75t_SL U35161 ( .A1(n25060), .A2(n31001), .B(n25059), .Y(
        n29921) );
  OAI22xp5_ASAP7_75t_SL U35162 ( .A1(mult_x_1196_n3203), .A2(n23072), .B1(
        mult_x_1196_n3202), .B2(n23987), .Y(mult_x_1196_n2627) );
  OAI22xp5_ASAP7_75t_SL U35163 ( .A1(mult_x_1196_n2823), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2822), .Y(mult_x_1196_n2257) );
  OAI22xp5_ASAP7_75t_SL U35164 ( .A1(mult_x_1196_n2871), .A2(n24031), .B1(
        n24030), .B2(mult_x_1196_n2870), .Y(mult_x_1196_n2305) );
  OAI22xp5_ASAP7_75t_SL U35165 ( .A1(mult_x_1196_n2916), .A2(n24021), .B1(
        mult_x_1196_n2915), .B2(n24020), .Y(mult_x_1196_n2344) );
  INVx1_ASAP7_75t_SL U35166 ( .A(mult_x_1196_n706), .Y(mult_x_1196_n704) );
  AOI21xp5_ASAP7_75t_SL U35167 ( .A1(mult_x_1196_n707), .A2(n24273), .B(
        mult_x_1196_n704), .Y(mult_x_1196_n702) );
  BUFx6f_ASAP7_75t_SL U35168 ( .A(mult_x_1196_n72), .Y(n24009) );
  OAI22xp5_ASAP7_75t_SL U35169 ( .A1(n22792), .A2(mult_x_1196_n3064), .B1(
        n24005), .B2(mult_x_1196_n3063), .Y(mult_x_1196_n2492) );
  OAI22xp5_ASAP7_75t_SL U35170 ( .A1(mult_x_1196_n3160), .A2(n24230), .B1(
        n23991), .B2(mult_x_1196_n3159), .Y(mult_x_1196_n2584) );
  OAI22xp5_ASAP7_75t_SL U35171 ( .A1(mult_x_1196_n3187), .A2(n23072), .B1(
        mult_x_1196_n3186), .B2(n23987), .Y(mult_x_1196_n2611) );
  FAx1_ASAP7_75t_SL U35172 ( .A(mult_x_1196_n2528), .B(mult_x_1196_n2688), 
        .CI(mult_x_1196_n1984), .CON(mult_x_1196_n1966), .SN(mult_x_1196_n1967) );
  OAI22xp5_ASAP7_75t_SL U35173 ( .A1(mult_x_1196_n2972), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2971), .Y(mult_x_1196_n2400) );
  FAx1_ASAP7_75t_SL U35174 ( .A(mult_x_1196_n925), .B(n22272), .CI(
        mult_x_1196_n927), .CON(mult_x_1196_n910), .SN(mult_x_1196_n911) );
  OAI22xp5_ASAP7_75t_SL U35175 ( .A1(mult_x_1196_n2919), .A2(n24022), .B1(
        mult_x_1196_n2918), .B2(n24020), .Y(mult_x_1196_n2347) );
  OAI22xp5_ASAP7_75t_SL U35176 ( .A1(n23993), .A2(mult_x_1196_n3159), .B1(
        n23991), .B2(mult_x_1196_n3158), .Y(mult_x_1196_n2583) );
  AOI21xp5_ASAP7_75t_SL U35177 ( .A1(u0_0_leon3x0_p0_dci[8]), .A2(n28902), .B(
        n28901), .Y(n30966) );
  OAI22xp5_ASAP7_75t_SL U35178 ( .A1(mult_x_1196_n3033), .A2(n24009), .B1(
        mult_x_1196_n3032), .B2(n24008), .Y(mult_x_1196_n2461) );
  NAND2xp5_ASAP7_75t_SL U35179 ( .A(n32169), .B(n24765), .Y(n32167) );
  OAI22xp5_ASAP7_75t_SL U35180 ( .A1(mult_x_1196_n3153), .A2(n23992), .B1(
        n23994), .B2(mult_x_1196_n3154), .Y(mult_x_1196_n2578) );
  OAI22xp5_ASAP7_75t_SL U35181 ( .A1(mult_x_1196_n3240), .A2(n23985), .B1(
        mult_x_1196_n3239), .B2(n23984), .Y(mult_x_1196_n2664) );
  OAI22xp5_ASAP7_75t_SL U35182 ( .A1(mult_x_1196_n3062), .A2(n24007), .B1(
        n24005), .B2(mult_x_1196_n3061), .Y(mult_x_1196_n2490) );
  FAx1_ASAP7_75t_SL U35183 ( .A(mult_x_1196_n858), .B(mult_x_1196_n865), .CI(
        mult_x_1196_n863), .CON(mult_x_1196_n859), .SN(mult_x_1196_n860) );
  FAx1_ASAP7_75t_SL U35184 ( .A(mult_x_1196_n2239), .B(mult_x_1196_n2146), 
        .CI(mult_x_1196_n861), .CON(mult_x_1196_n862), .SN(mult_x_1196_n863)
         );
  OAI22xp5_ASAP7_75t_SL U35185 ( .A1(mult_x_1196_n2794), .A2(n24038), .B1(
        mult_x_1196_n2793), .B2(n22936), .Y(mult_x_1196_n2228) );
  OAI22xp5_ASAP7_75t_SL U35186 ( .A1(mult_x_1196_n2792), .A2(n24039), .B1(
        mult_x_1196_n2791), .B2(n22391), .Y(mult_x_1196_n2226) );
  OAI22xp5_ASAP7_75t_SL U35187 ( .A1(mult_x_1196_n3190), .A2(n23989), .B1(
        mult_x_1196_n3189), .B2(n22248), .Y(mult_x_1196_n2614) );
  OAI22xp5_ASAP7_75t_SL U35188 ( .A1(mult_x_1196_n2759), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2758), .Y(mult_x_1196_n2196) );
  OAI22xp5_ASAP7_75t_SL U35189 ( .A1(mult_x_1196_n2964), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2963), .Y(mult_x_1196_n2392) );
  OAI21xp5_ASAP7_75t_SL U35190 ( .A1(n32308), .A2(n22402), .B(n30792), .Y(
        n18209) );
  NAND2xp5_ASAP7_75t_SL U35191 ( .A(mult_x_1196_n1045), .B(mult_x_1196_n1025), 
        .Y(n24146) );
  OAI22xp5_ASAP7_75t_SL U35192 ( .A1(mult_x_1196_n2898), .A2(n23708), .B1(
        mult_x_1196_n2897), .B2(n24025), .Y(mult_x_1196_n2326) );
  OAI22xp5_ASAP7_75t_SL U35193 ( .A1(n24107), .A2(mult_x_1196_n3189), .B1(
        mult_x_1196_n3188), .B2(n23988), .Y(mult_x_1196_n2613) );
  OAI21xp5_ASAP7_75t_SL U35194 ( .A1(n18614), .A2(n22392), .B(n25407), .Y(
        n30619) );
  NAND2xp5_ASAP7_75t_SL U35195 ( .A(n22837), .B(u0_0_leon3x0_p0_divi[9]), .Y(
        add_x_735_n221) );
  INVx1_ASAP7_75t_SL U35196 ( .A(n22837), .Y(n27144) );
  OAI21xp5_ASAP7_75t_SL U35197 ( .A1(n26777), .A2(n24781), .B(n18849), .Y(
        n32184) );
  OAI22xp5_ASAP7_75t_SL U35198 ( .A1(mult_x_1196_n2776), .A2(n22412), .B1(
        mult_x_1196_n2775), .B2(n22481), .Y(mult_x_1196_n900) );
  BUFx6f_ASAP7_75t_SL U35199 ( .A(mult_x_1196_n135), .Y(n24038) );
  INVx1_ASAP7_75t_SL U35200 ( .A(mult_x_1196_n900), .Y(mult_x_1196_n901) );
  AOI21xp5_ASAP7_75t_SL U35201 ( .A1(add_x_735_n121), .A2(add_x_735_n136), .B(
        add_x_735_n122), .Y(add_x_735_n116) );
  FAx1_ASAP7_75t_SL U35202 ( .A(mult_x_1196_n2349), .B(mult_x_1196_n2569), 
        .CI(mult_x_1196_n2227), .CON(mult_x_1196_n1279), .SN(mult_x_1196_n1280) );
  OAI22xp5_ASAP7_75t_SL U35203 ( .A1(mult_x_1196_n2793), .A2(n24039), .B1(
        mult_x_1196_n2792), .B2(n22391), .Y(mult_x_1196_n2227) );
  OAI22xp5_ASAP7_75t_SL U35204 ( .A1(mult_x_1196_n3163), .A2(n23994), .B1(
        n23991), .B2(mult_x_1196_n3162), .Y(mult_x_1196_n2587) );
  OAI22xp5_ASAP7_75t_SL U35205 ( .A1(mult_x_1196_n2854), .A2(n24031), .B1(
        n18390), .B2(mult_x_1196_n2853), .Y(mult_x_1196_n2288) );
  OAI22xp5_ASAP7_75t_SL U35206 ( .A1(n23081), .A2(mult_x_1196_n3157), .B1(
        n23991), .B2(mult_x_1196_n3156), .Y(mult_x_1196_n2581) );
  OR2x2_ASAP7_75t_SL U35207 ( .A(mult_x_1196_n578), .B(n22541), .Y(n23938) );
  NOR2x1_ASAP7_75t_SL U35208 ( .A(mult_x_1196_n1426), .B(mult_x_1196_n1427), 
        .Y(mult_x_1196_n578) );
  INVx1_ASAP7_75t_SL U35209 ( .A(mult_x_1196_n1166), .Y(mult_x_1196_n1162) );
  INVx1_ASAP7_75t_SL U35210 ( .A(mult_x_1196_n1259), .Y(mult_x_1196_n1225) );
  INVx1_ASAP7_75t_SL U35211 ( .A(mult_x_1196_n1295), .Y(n23939) );
  OAI22xp5_ASAP7_75t_SL U35212 ( .A1(mult_x_1196_n2969), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2968), .Y(mult_x_1196_n2397) );
  OAI22xp5_ASAP7_75t_SL U35213 ( .A1(mult_x_1196_n3262), .A2(n23982), .B1(
        n22389), .B2(mult_x_1196_n3261), .Y(mult_x_1196_n2686) );
  XNOR2xp5_ASAP7_75t_SL U35214 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__6_), .B(
        n32185), .Y(n24842) );
  XNOR2xp5_ASAP7_75t_SL U35215 ( .A(n30935), .B(n32185), .Y(n30936) );
  NAND2xp5_ASAP7_75t_SL U35216 ( .A(n30007), .B(n28742), .Y(n28921) );
  NAND2xp5_ASAP7_75t_SL U35217 ( .A(n28877), .B(n28992), .Y(n29609) );
  OAI22xp5_ASAP7_75t_SL U35218 ( .A1(mult_x_1196_n2963), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2962), .Y(mult_x_1196_n2391) );
  INVx1_ASAP7_75t_SL U35219 ( .A(mult_x_1196_n1045), .Y(n24142) );
  OAI22xp5_ASAP7_75t_SL U35220 ( .A1(mult_x_1196_n2965), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2964), .Y(mult_x_1196_n2393) );
  INVx1_ASAP7_75t_SL U35221 ( .A(mult_x_1196_n2037), .Y(mult_x_1196_n2031) );
  NAND2xp5_ASAP7_75t_SL U35222 ( .A(add_x_746_n145), .B(add_x_746_n126), .Y(
        add_x_746_n125) );
  OAI22xp5_ASAP7_75t_SL U35223 ( .A1(mult_x_1196_n3115), .A2(n24000), .B1(
        n23997), .B2(mult_x_1196_n3114), .Y(mult_x_1196_n2539) );
  OAI22xp5_ASAP7_75t_SL U35224 ( .A1(mult_x_1196_n2844), .A2(n18309), .B1(
        n22743), .B2(mult_x_1196_n2843), .Y(mult_x_1196_n2278) );
  NAND2xp5_ASAP7_75t_SL U35225 ( .A(n24897), .B(n24974), .Y(n31627) );
  FAx1_ASAP7_75t_SL U35226 ( .A(mult_x_1196_n2290), .B(mult_x_1196_n2197), 
        .CI(mult_x_1196_n2226), .CON(mult_x_1196_n1248), .SN(mult_x_1196_n1249) );
  NAND2xp5_ASAP7_75t_SL U35227 ( .A(n25410), .B(n32446), .Y(n31040) );
  OAI22xp5_ASAP7_75t_SL U35228 ( .A1(mult_x_1196_n3263), .A2(n23982), .B1(
        n22389), .B2(mult_x_1196_n3262), .Y(mult_x_1196_n2687) );
  OR2x2_ASAP7_75t_SL U35229 ( .A(u0_0_leon3x0_p0_ici[40]), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__10_), .Y(n23945) );
  OR2x2_ASAP7_75t_SL U35230 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__12_), .B(
        u0_0_leon3x0_p0_ici[42]), .Y(n23946) );
  OR2x2_ASAP7_75t_SL U35231 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__16_), .B(
        u0_0_leon3x0_p0_ici[46]), .Y(n23944) );
  OR2x2_ASAP7_75t_SL U35232 ( .A(u0_0_leon3x0_p0_ici[36]), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__6_), .Y(n23949) );
  OR2x2_ASAP7_75t_SL U35233 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__8_), .B(
        u0_0_leon3x0_p0_ici[38]), .Y(n23948) );
  OR2x2_ASAP7_75t_SL U35234 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__5_), .B(
        u0_0_leon3x0_p0_ici[35]), .Y(n23950) );
  OR2x2_ASAP7_75t_SL U35235 ( .A(u0_0_leon3x0_p0_ici[44]), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__14_), .Y(n23943) );
  OR2x2_ASAP7_75t_SL U35236 ( .A(u0_0_leon3x0_p0_ici[51]), .B(n18842), .Y(
        n23942) );
  OR2x2_ASAP7_75t_SL U35237 ( .A(u0_0_leon3x0_p0_ici[48]), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_), .Y(n23947) );
  AND2x2_ASAP7_75t_SL U35238 ( .A(n22227), .B(n24036), .Y(mult_x_1196_n2238)
         );
  AND2x2_ASAP7_75t_SL U35239 ( .A(n18984), .B(n23990), .Y(mult_x_1196_n2602)
         );
  AND2x2_ASAP7_75t_SL U35240 ( .A(n22227), .B(n24010), .Y(mult_x_1196_n2436)
         );
  OR2x2_ASAP7_75t_SL U35241 ( .A(n22227), .B(n22961), .Y(mult_x_1196_n3076) );
  AND2x2_ASAP7_75t_SL U35242 ( .A(n22227), .B(n22265), .Y(mult_x_1196_n2402)
         );
  AND2x2_ASAP7_75t_SL U35243 ( .A(n22227), .B(n18365), .Y(mult_x_1196_n2670)
         );
  AND2x2_ASAP7_75t_SL U35244 ( .A(n22227), .B(n24032), .Y(mult_x_1196_n2272)
         );
  AND2x2_ASAP7_75t_SL U35245 ( .A(n22227), .B(n22962), .Y(mult_x_1196_n2306)
         );
  AND2x2_ASAP7_75t_SL U35246 ( .A(n22227), .B(n23443), .Y(mult_x_1196_n2470)
         );
  AND2x2_ASAP7_75t_SL U35247 ( .A(n22227), .B(n23995), .Y(mult_x_1196_n2568)
         );
  XOR2xp5_ASAP7_75t_SL U35248 ( .A(n24100), .B(mult_x_1196_n2496), .Y(n24101)
         );
  XOR2xp5_ASAP7_75t_SL U35249 ( .A(mult_x_1196_n1486), .B(n23918), .Y(n24102)
         );
  MAJIxp5_ASAP7_75t_SL U35250 ( .A(mult_x_1196_n1349), .B(mult_x_1196_n1355), 
        .C(n22655), .Y(mult_x_1196_n1336) );
  XNOR2xp5_ASAP7_75t_SL U35251 ( .A(mult_x_1196_n1751), .B(mult_x_1196_n1783), 
        .Y(n24104) );
  MAJIxp5_ASAP7_75t_SL U35252 ( .A(mult_x_1196_n2049), .B(mult_x_1196_n2045), 
        .C(mult_x_1196_n2057), .Y(mult_x_1196_n2046) );
  MAJIxp5_ASAP7_75t_SL U35253 ( .A(mult_x_1196_n1793), .B(mult_x_1196_n1814), 
        .C(mult_x_1196_n1812), .Y(mult_x_1196_n1783) );
  XOR2xp5_ASAP7_75t_SL U35254 ( .A(mult_x_1196_n2611), .B(mult_x_1196_n2547), 
        .Y(n24124) );
  MAJIxp5_ASAP7_75t_SL U35255 ( .A(mult_x_1196_n2611), .B(n24123), .C(
        mult_x_1196_n2547), .Y(mult_x_1196_n1642) );
  NOR2xp33_ASAP7_75t_SL U35256 ( .A(n22983), .B(mult_x_1196_n2885), .Y(n24125)
         );
  XOR2xp5_ASAP7_75t_SL U35257 ( .A(mult_x_1196_n2195), .B(mult_x_1196_n2474), 
        .Y(n24139) );
  MAJIxp5_ASAP7_75t_SL U35258 ( .A(mult_x_1196_n2474), .B(mult_x_1196_n2195), 
        .C(n24140), .Y(mult_x_1196_n1183) );
  XNOR2xp5_ASAP7_75t_SL U35259 ( .A(mult_x_1196_n2456), .B(mult_x_1196_n1707), 
        .Y(n24141) );
  XNOR2xp5_ASAP7_75t_SL U35260 ( .A(mult_x_1196_n1042), .B(n24143), .Y(
        mult_x_1196_n1020) );
  XOR2xp5_ASAP7_75t_SL U35261 ( .A(n23963), .B(n24071), .Y(mult_x_1196_n3036)
         );
  XOR2xp5_ASAP7_75t_SL U35262 ( .A(n18299), .B(n24072), .Y(mult_x_1196_n3037)
         );
  XOR2xp5_ASAP7_75t_SL U35263 ( .A(n23963), .B(n24068), .Y(mult_x_1196_n3033)
         );
  XOR2xp5_ASAP7_75t_SL U35264 ( .A(n23963), .B(n24067), .Y(mult_x_1196_n3032)
         );
  XOR2xp5_ASAP7_75t_SL U35265 ( .A(n24069), .B(n23963), .Y(mult_x_1196_n3034)
         );
  XOR2xp5_ASAP7_75t_SL U35266 ( .A(n23963), .B(u0_0_leon3x0_p0_muli[17]), .Y(
        mult_x_1196_n3035) );
  NOR2xp33_ASAP7_75t_SL U35267 ( .A(n24025), .B(mult_x_1196_n2884), .Y(n24157)
         );
  MAJIxp5_ASAP7_75t_SL U35268 ( .A(mult_x_1196_n1406), .B(mult_x_1196_n1417), 
        .C(mult_x_1196_n1421), .Y(mult_x_1196_n1407) );
  OR2x2_ASAP7_75t_SL U35269 ( .A(mult_x_1196_n997), .B(mult_x_1196_n979), .Y(
        mult_x_1196_n787) );
  XNOR2xp5_ASAP7_75t_SL U35270 ( .A(mult_x_1196_n2649), .B(n24182), .Y(n24183)
         );
  XNOR2xp5_ASAP7_75t_SL U35271 ( .A(mult_x_1196_n1262), .B(n24184), .Y(n24185)
         );
  NOR2xp33_ASAP7_75t_SL U35272 ( .A(n22983), .B(mult_x_1196_n2888), .Y(n24186)
         );
  XNOR2xp5_ASAP7_75t_SL U35273 ( .A(mult_x_1196_n1765), .B(mult_x_1196_n1738), 
        .Y(n24190) );
  XOR2xp5_ASAP7_75t_SL U35274 ( .A(n24205), .B(n24071), .Y(mult_x_1196_n3206)
         );
  XOR2xp5_ASAP7_75t_SL U35275 ( .A(n24205), .B(n24073), .Y(mult_x_1196_n3208)
         );
  XOR2xp5_ASAP7_75t_SL U35276 ( .A(n24205), .B(n24072), .Y(mult_x_1196_n3207)
         );
  XNOR2xp5_ASAP7_75t_SL U35277 ( .A(n23957), .B(n24070), .Y(mult_x_1196_n3205)
         );
  XOR2xp5_ASAP7_75t_SL U35278 ( .A(n24205), .B(n24075), .Y(mult_x_1196_n3210)
         );
  MAJIxp5_ASAP7_75t_SL U35279 ( .A(n24220), .B(mult_x_1196_n1363), .C(n18999), 
        .Y(mult_x_1196_n1357) );
  OR2x2_ASAP7_75t_SL U35280 ( .A(n24232), .B(n23983), .Y(n24080) );
  XOR2xp5_ASAP7_75t_SL U35281 ( .A(mult_x_1196_n1246), .B(mult_x_1196_n1252), 
        .Y(n24221) );
  OR2x2_ASAP7_75t_SL U35282 ( .A(mult_x_1196_n1868), .B(mult_x_1196_n1845), 
        .Y(mult_x_1196_n816) );
  XOR2xp5_ASAP7_75t_SL U35283 ( .A(n18423), .B(n24047), .Y(mult_x_1196_n2910)
         );
  XNOR2xp5_ASAP7_75t_SL U35284 ( .A(n23969), .B(n18615), .Y(mult_x_1196_n2912)
         );
  XOR2xp5_ASAP7_75t_SL U35285 ( .A(n23936), .B(n24066), .Y(mult_x_1196_n2963)
         );
  XNOR2xp5_ASAP7_75t_SL U35286 ( .A(n24231), .B(n22227), .Y(mult_x_1196_n2973)
         );
  XNOR2xp5_ASAP7_75t_SL U35287 ( .A(n23967), .B(n24069), .Y(mult_x_1196_n2966)
         );
  XNOR2xp5_ASAP7_75t_SL U35288 ( .A(n24231), .B(n24070), .Y(mult_x_1196_n2967)
         );
  MAJIxp5_ASAP7_75t_SL U35289 ( .A(mult_x_1196_n2514), .B(mult_x_1196_n2674), 
        .C(n24245), .Y(mult_x_1196_n1611) );
  XOR2xp5_ASAP7_75t_SL U35290 ( .A(mult_x_1196_n1048), .B(n24247), .Y(n24248)
         );
  OR2x2_ASAP7_75t_SL U35291 ( .A(mult_x_1196_n839), .B(mult_x_1196_n837), .Y(
        n24250) );
  OR2x2_ASAP7_75t_SL U35292 ( .A(mult_x_1196_n867), .B(mult_x_1196_n866), .Y(
        n24252) );
  OR2x2_ASAP7_75t_SL U35293 ( .A(mult_x_1196_n2702), .B(mult_x_1196_n2670), 
        .Y(n24254) );
  OR2x2_ASAP7_75t_SL U35294 ( .A(mult_x_1196_n3035), .B(n24008), .Y(n24258) );
  OR2x2_ASAP7_75t_SL U35295 ( .A(mult_x_1196_n2083), .B(mult_x_1196_n2082), 
        .Y(n24261) );
  MAJx2_ASAP7_75t_SL U35296 ( .A(mult_x_1196_n1283), .B(mult_x_1196_n1281), 
        .C(mult_x_1196_n1279), .Y(n24263) );
  OR2x2_ASAP7_75t_SL U35297 ( .A(n23997), .B(mult_x_1196_n3121), .Y(n24264) );
  XOR2xp5_ASAP7_75t_SL U35298 ( .A(mult_x_1196_n1719), .B(n24188), .Y(n24269)
         );
  OR2x2_ASAP7_75t_SL U35299 ( .A(mult_x_1196_n3172), .B(n23992), .Y(n24271) );
  OR2x2_ASAP7_75t_SL U35300 ( .A(n22222), .B(mult_x_1196_n2075), .Y(n24272) );
  OR2x2_ASAP7_75t_SL U35301 ( .A(mult_x_1196_n2574), .B(mult_x_1196_n2418), 
        .Y(n24275) );
  OR2x2_ASAP7_75t_SL U35302 ( .A(mult_x_1196_n2052), .B(mult_x_1196_n2044), 
        .Y(n24276) );
  OR2x2_ASAP7_75t_SL U35303 ( .A(mult_x_1196_n3002), .B(n24012), .Y(n24277) );
  MAJx2_ASAP7_75t_SL U35304 ( .A(mult_x_1196_n1364), .B(mult_x_1196_n1329), 
        .C(n22207), .Y(n24281) );
  XOR2xp5_ASAP7_75t_SL U35305 ( .A(n24185), .B(mult_x_1196_n1230), .Y(n24282)
         );
  MAJx2_ASAP7_75t_SL U35306 ( .A(n24244), .B(mult_x_1196_n2470), .C(
        mult_x_1196_n2658), .Y(n24283) );
  MAJx2_ASAP7_75t_SL U35307 ( .A(mult_x_1196_n1640), .B(mult_x_1196_n1642), 
        .C(mult_x_1196_n1638), .Y(n24284) );
  AND2x2_ASAP7_75t_SL U35308 ( .A(n22356), .B(mult_x_1196_n1648), .Y(n24289)
         );
  OR2x2_ASAP7_75t_SL U35309 ( .A(mult_x_1196_n2061), .B(mult_x_1196_n2053), 
        .Y(n24290) );
  MAJx2_ASAP7_75t_SL U35310 ( .A(mult_x_1196_n1242), .B(mult_x_1196_n1245), 
        .C(mult_x_1196_n1273), .Y(n24297) );
  OR2x2_ASAP7_75t_SL U35311 ( .A(mult_x_1196_n3229), .B(n23984), .Y(n24299) );
  MAJx2_ASAP7_75t_SL U35312 ( .A(n18912), .B(mult_x_1196_n1665), .C(
        mult_x_1196_n1668), .Y(n24301) );
  MAJx2_ASAP7_75t_SL U35313 ( .A(mult_x_1196_n1328), .B(mult_x_1196_n1331), 
        .C(n22260), .Y(n24303) );
  OR2x2_ASAP7_75t_SL U35314 ( .A(n24269), .B(mult_x_1196_n1744), .Y(n24304) );
  MAJx2_ASAP7_75t_SL U35315 ( .A(mult_x_1196_n1783), .B(mult_x_1196_n1751), 
        .C(mult_x_1196_n1760), .Y(n24308) );
  MAJx2_ASAP7_75t_SL U35316 ( .A(mult_x_1196_n1230), .B(n18371), .C(
        mult_x_1196_n1262), .Y(n24311) );
  MAJIxp5_ASAP7_75t_SL U35317 ( .A(n24127), .B(mult_x_1196_n2194), .C(
        mult_x_1196_n2255), .Y(mult_x_1196_n1160) );
  XNOR2xp5_ASAP7_75t_SL U35318 ( .A(n24066), .B(n23952), .Y(mult_x_1196_n3269)
         );
  XNOR2xp5_ASAP7_75t_SL U35319 ( .A(n24067), .B(n23952), .Y(mult_x_1196_n3270)
         );
  XNOR2xp5_ASAP7_75t_SL U35320 ( .A(n24068), .B(n23952), .Y(mult_x_1196_n3271)
         );
  NOR2xp33_ASAP7_75t_SL U35321 ( .A(n23984), .B(mult_x_1196_n3235), .Y(n24239)
         );
  NOR2xp33_ASAP7_75t_SL U35322 ( .A(mult_x_1196_n3234), .B(n23984), .Y(n24173)
         );
  NOR2xp33_ASAP7_75t_SL U35323 ( .A(mult_x_1196_n3242), .B(n23984), .Y(n24133)
         );
  XNOR2xp5_ASAP7_75t_SL U35324 ( .A(n24071), .B(n23952), .Y(mult_x_1196_n3274)
         );
  XNOR2xp5_ASAP7_75t_SL U35325 ( .A(n24070), .B(n23952), .Y(mult_x_1196_n3273)
         );
  XNOR2xp5_ASAP7_75t_SL U35326 ( .A(n24069), .B(n23952), .Y(mult_x_1196_n3272)
         );
  INVxp33_ASAP7_75t_SRAM U35327 ( .A(mult_x_1196_n597), .Y(mult_x_1196_n599)
         );
  INVxp33_ASAP7_75t_SRAM U35328 ( .A(mult_x_1196_n547), .Y(mult_x_1196_n545)
         );
  XNOR2xp5_ASAP7_75t_SL U35329 ( .A(n24118), .B(mult_x_1196_n1160), .Y(
        mult_x_1196_n1125) );
  XNOR2xp5_ASAP7_75t_SL U35330 ( .A(n24072), .B(n23952), .Y(mult_x_1196_n3275)
         );
  XNOR2xp5_ASAP7_75t_SL U35331 ( .A(n23957), .B(n24069), .Y(mult_x_1196_n3204)
         );
  XOR2xp5_ASAP7_75t_SL U35332 ( .A(n24205), .B(n24068), .Y(mult_x_1196_n3203)
         );
  XNOR2xp5_ASAP7_75t_SL U35333 ( .A(n24073), .B(n23952), .Y(mult_x_1196_n3276)
         );
  INVxp33_ASAP7_75t_SRAM U35334 ( .A(mult_x_1196_n714), .Y(mult_x_1196_n825)
         );
  INVxp33_ASAP7_75t_SRAM U35335 ( .A(mult_x_1196_n730), .Y(mult_x_1196_n729)
         );
  XNOR2xp5_ASAP7_75t_SL U35336 ( .A(n24225), .B(mult_x_1196_n2555), .Y(
        mult_x_1196_n1862) );
  XNOR2xp5_ASAP7_75t_SL U35337 ( .A(mult_x_1196_n2504), .B(mult_x_1196_n2628), 
        .Y(n24242) );
  XOR2xp5_ASAP7_75t_SL U35338 ( .A(n24205), .B(n24067), .Y(mult_x_1196_n3202)
         );
  NOR2xp33_ASAP7_75t_SL U35339 ( .A(mult_x_1196_n2708), .B(n24043), .Y(
        mult_x_1196_n2146) );
  XNOR2xp5_ASAP7_75t_SL U35340 ( .A(n24231), .B(n24052), .Y(mult_x_1196_n2949)
         );
  XNOR2xp5_ASAP7_75t_SL U35341 ( .A(mult_x_1196_n2513), .B(mult_x_1196_n2673), 
        .Y(n24266) );
  NOR2xp33_ASAP7_75t_SL U35342 ( .A(mult_x_1196_n2710), .B(n24043), .Y(
        mult_x_1196_n2148) );
  INVxp33_ASAP7_75t_SRAM U35343 ( .A(mult_x_1196_n474), .Y(mult_x_1196_n791)
         );
  INVxp33_ASAP7_75t_SRAM U35344 ( .A(mult_x_1196_n613), .Y(mult_x_1196_n808)
         );
  INVxp33_ASAP7_75t_SRAM U35345 ( .A(mult_x_1196_n602), .Y(mult_x_1196_n806)
         );
  NOR2xp33_ASAP7_75t_SL U35346 ( .A(mult_x_1196_n3236), .B(n23985), .Y(n24240)
         );
  INVxp33_ASAP7_75t_SRAM U35347 ( .A(mult_x_1196_n578), .Y(mult_x_1196_n803)
         );
  XOR2xp5_ASAP7_75t_SL U35348 ( .A(n18423), .B(n24046), .Y(mult_x_1196_n2909)
         );
  NOR2xp33_ASAP7_75t_SL U35349 ( .A(mult_x_1196_n2717), .B(n24043), .Y(
        mult_x_1196_n2155) );
  NOR2xp33_ASAP7_75t_SL U35350 ( .A(mult_x_1196_n2718), .B(n24043), .Y(
        mult_x_1196_n2156) );
  XOR2xp5_ASAP7_75t_SL U35351 ( .A(n18423), .B(n24045), .Y(mult_x_1196_n2908)
         );
  XOR2xp5_ASAP7_75t_SL U35352 ( .A(n18423), .B(n24044), .Y(mult_x_1196_n2907)
         );
  XNOR2xp5_ASAP7_75t_SL U35353 ( .A(n23969), .B(n24050), .Y(mult_x_1196_n2913)
         );
  NOR2xp33_ASAP7_75t_SL U35354 ( .A(n24025), .B(mult_x_1196_n2881), .Y(n24091)
         );
  NOR2xp33_ASAP7_75t_SL U35355 ( .A(mult_x_1196_n2882), .B(n23708), .Y(n24092)
         );
  NOR2xp33_ASAP7_75t_SL U35356 ( .A(mult_x_1196_n2722), .B(n24043), .Y(
        mult_x_1196_n2160) );
  XOR2xp5_ASAP7_75t_SL U35357 ( .A(n18423), .B(n24053), .Y(mult_x_1196_n2916)
         );
  NOR2xp33_ASAP7_75t_SL U35358 ( .A(mult_x_1196_n2723), .B(n24043), .Y(
        mult_x_1196_n2161) );
  NOR2xp33_ASAP7_75t_SL U35359 ( .A(mult_x_1196_n2724), .B(n24043), .Y(
        mult_x_1196_n2162) );
  XOR2xp5_ASAP7_75t_SL U35360 ( .A(n23968), .B(n24054), .Y(mult_x_1196_n2917)
         );
  XOR2xp5_ASAP7_75t_SL U35361 ( .A(n18423), .B(n24056), .Y(mult_x_1196_n2919)
         );
  XOR2xp5_ASAP7_75t_SL U35362 ( .A(n23968), .B(n24055), .Y(mult_x_1196_n2918)
         );
  NOR2xp33_ASAP7_75t_SL U35363 ( .A(mult_x_1196_n2917), .B(n24020), .Y(n24137)
         );
  NOR2xp33_ASAP7_75t_SL U35364 ( .A(mult_x_1196_n2918), .B(n24021), .Y(n24138)
         );
  NOR2xp33_ASAP7_75t_SL U35365 ( .A(mult_x_1196_n2725), .B(n24043), .Y(
        mult_x_1196_n2163) );
  NOR2xp33_ASAP7_75t_SL U35366 ( .A(n23442), .B(mult_x_1196_n3013), .Y(n24176)
         );
  NOR2xp33_ASAP7_75t_SL U35367 ( .A(mult_x_1196_n3014), .B(n24009), .Y(n24177)
         );
  XNOR2xp5_ASAP7_75t_SL U35368 ( .A(n24127), .B(n24128), .Y(mult_x_1196_n1161)
         );
  NOR2xp33_ASAP7_75t_SL U35369 ( .A(mult_x_1196_n2727), .B(n24043), .Y(
        mult_x_1196_n2165) );
  XNOR2xp5_ASAP7_75t_SL U35370 ( .A(mult_x_1196_n1250), .B(n24221), .Y(
        mult_x_1196_n1212) );
  NOR2xp33_ASAP7_75t_SL U35371 ( .A(mult_x_1196_n2726), .B(n24043), .Y(
        mult_x_1196_n2164) );
  XNOR2xp5_ASAP7_75t_SL U35372 ( .A(n24052), .B(n23964), .Y(mult_x_1196_n3017)
         );
  XNOR2xp5_ASAP7_75t_SL U35373 ( .A(n24274), .B(n24103), .Y(mult_x_1196_n1240)
         );
  XOR2xp5_ASAP7_75t_SL U35374 ( .A(mult_x_1196_n2537), .B(n24187), .Y(
        mult_x_1196_n1284) );
  NOR2xp33_ASAP7_75t_SL U35375 ( .A(mult_x_1196_n2731), .B(n24043), .Y(
        mult_x_1196_n2169) );
  INVxp33_ASAP7_75t_SRAM U35376 ( .A(mult_x_1196_n1299), .Y(n24192) );
  NAND2xp33_ASAP7_75t_SRAM U35377 ( .A(mult_x_1196_n1299), .B(
        mult_x_1196_n1268), .Y(n24194) );
  NOR2xp33_ASAP7_75t_SL U35378 ( .A(mult_x_1196_n2732), .B(n24043), .Y(
        mult_x_1196_n2170) );
  NOR2xp33_ASAP7_75t_SL U35379 ( .A(mult_x_1196_n3053), .B(mult_x_1196_n60), 
        .Y(n24222) );
  XNOR2xp5_ASAP7_75t_SL U35380 ( .A(mult_x_1196_n1355), .B(n24155), .Y(n24152)
         );
  XOR2xp5_ASAP7_75t_SL U35381 ( .A(n24154), .B(n24152), .Y(n24260) );
  XNOR2xp5_ASAP7_75t_SL U35382 ( .A(n24102), .B(mult_x_1196_n1484), .Y(
        mult_x_1196_n1477) );
  XOR2xp5_ASAP7_75t_SL U35383 ( .A(n23935), .B(n24067), .Y(mult_x_1196_n2964)
         );
  XNOR2xp5_ASAP7_75t_SL U35384 ( .A(n23957), .B(n24052), .Y(mult_x_1196_n3187)
         );
  XNOR2xp5_ASAP7_75t_SL U35385 ( .A(n24115), .B(mult_x_1196_n1574), .Y(
        mult_x_1196_n1559) );
  XOR2xp5_ASAP7_75t_SL U35386 ( .A(n24205), .B(n24055), .Y(mult_x_1196_n3190)
         );
  XOR2xp5_ASAP7_75t_SL U35387 ( .A(n24068), .B(n23935), .Y(mult_x_1196_n2965)
         );
  XOR2xp5_ASAP7_75t_SL U35388 ( .A(n23963), .B(n24066), .Y(mult_x_1196_n3031)
         );
  XOR2xp5_ASAP7_75t_SL U35389 ( .A(n23935), .B(n24072), .Y(mult_x_1196_n2969)
         );
  XOR2xp5_ASAP7_75t_SL U35390 ( .A(n23936), .B(n24071), .Y(mult_x_1196_n2968)
         );
  XNOR2xp5_ASAP7_75t_SL U35391 ( .A(n24203), .B(mult_x_1196_n2305), .Y(n24204)
         );
  XOR2xp5_ASAP7_75t_SL U35392 ( .A(n23936), .B(n24073), .Y(mult_x_1196_n2970)
         );
  XOR2xp5_ASAP7_75t_SL U35393 ( .A(n24183), .B(mult_x_1196_n2333), .Y(
        mult_x_1196_n1817) );
  XOR2xp5_ASAP7_75t_SL U35394 ( .A(n24075), .B(n23936), .Y(mult_x_1196_n2972)
         );
  XOR2xp5_ASAP7_75t_SL U35395 ( .A(n23935), .B(n24074), .Y(mult_x_1196_n2971)
         );
  NOR2xp33_ASAP7_75t_SL U35396 ( .A(mult_x_1196_n2133), .B(mult_x_1196_n1866), 
        .Y(n24132) );
  XOR2xp5_ASAP7_75t_SL U35397 ( .A(n23963), .B(n24074), .Y(mult_x_1196_n3039)
         );
  XOR2xp5_ASAP7_75t_SL U35398 ( .A(n18299), .B(n24073), .Y(mult_x_1196_n3038)
         );
  XNOR2xp5_ASAP7_75t_SL U35399 ( .A(n24241), .B(n24242), .Y(mult_x_1196_n2027)
         );
  INVxp33_ASAP7_75t_SRAM U35400 ( .A(mult_x_1196_n2089), .Y(mult_x_1196_n2083)
         );
  XNOR2xp5_ASAP7_75t_SL U35401 ( .A(n22227), .B(n23952), .Y(mult_x_1196_n3279)
         );
  XNOR2xp5_ASAP7_75t_SL U35402 ( .A(n24075), .B(n23952), .Y(mult_x_1196_n3278)
         );
  XNOR2xp5_ASAP7_75t_SL U35403 ( .A(n24074), .B(n23952), .Y(mult_x_1196_n3277)
         );
  AO21x1_ASAP7_75t_SL U35404 ( .A1(n24261), .A2(mult_x_1196_n759), .B(
        mult_x_1196_n756), .Y(mult_x_1196_n753) );
  INVxp33_ASAP7_75t_SRAM U35405 ( .A(mult_x_1196_n482), .Y(mult_x_1196_n480)
         );
  INVxp33_ASAP7_75t_SRAM U35406 ( .A(mult_x_1196_n333), .Y(mult_x_1196_n331)
         );
  INVxp33_ASAP7_75t_SRAM U35407 ( .A(mult_x_1196_n451), .Y(mult_x_1196_n449)
         );
  INVxp33_ASAP7_75t_SRAM U35408 ( .A(mult_x_1196_n539), .Y(mult_x_1196_n798)
         );
  INVxp33_ASAP7_75t_SRAM U35409 ( .A(mult_x_1196_n546), .Y(mult_x_1196_n799)
         );
  INVxp33_ASAP7_75t_SRAM U35410 ( .A(mult_x_1196_n519), .Y(mult_x_1196_n796)
         );
  INVxp33_ASAP7_75t_SRAM U35411 ( .A(mult_x_1196_n557), .Y(mult_x_1196_n800)
         );
  INVxp33_ASAP7_75t_SRAM U35412 ( .A(n24086), .Y(n24088) );
  INVxp33_ASAP7_75t_SRAM U35413 ( .A(mult_x_1196_n816), .Y(mult_x_1196_n661)
         );
  INVxp33_ASAP7_75t_SRAM U35414 ( .A(mult_x_1196_n668), .Y(mult_x_1196_n667)
         );
  INVxp33_ASAP7_75t_SRAM U35415 ( .A(mult_x_1196_n664), .Y(n24122) );
  INVxp33_ASAP7_75t_SRAM U35416 ( .A(mult_x_1196_n651), .Y(mult_x_1196_n814)
         );
  INVxp33_ASAP7_75t_SRAM U35417 ( .A(mult_x_1196_n591), .Y(mult_x_1196_n805)
         );
  INVxp33_ASAP7_75t_SRAM U35418 ( .A(mult_x_1196_n607), .Y(mult_x_1196_n807)
         );
  INVxp33_ASAP7_75t_SRAM U35419 ( .A(mult_x_1196_n586), .Y(mult_x_1196_n804)
         );
  NAND2xp33_ASAP7_75t_SRAM U35420 ( .A(n24122), .B(mult_x_1196_n816), .Y(
        mult_x_1196_n266) );
  INVxp33_ASAP7_75t_SRAM U35421 ( .A(n24289), .Y(n24083) );
  INVxp33_ASAP7_75t_SRAM U35422 ( .A(mult_x_1196_n640), .Y(mult_x_1196_n812)
         );
  INVxp33_ASAP7_75t_SRAM U35423 ( .A(mult_x_1196_n645), .Y(mult_x_1196_n813)
         );
  INVxp33_ASAP7_75t_SRAM U35424 ( .A(mult_x_1196_n678), .Y(mult_x_1196_n818)
         );
  INVxp33_ASAP7_75t_SRAM U35425 ( .A(mult_x_1196_n684), .Y(mult_x_1196_n682)
         );
  INVxp33_ASAP7_75t_SRAM U35426 ( .A(mult_x_1196_n689), .Y(mult_x_1196_n820)
         );
  INVxp33_ASAP7_75t_SRAM U35427 ( .A(mult_x_1196_n708), .Y(mult_x_1196_n707)
         );
  INVxp33_ASAP7_75t_SRAM U35428 ( .A(n22333), .Y(mult_x_1196_n824) );
  INVxp33_ASAP7_75t_SRAM U35429 ( .A(mult_x_1196_n717), .Y(mult_x_1196_n716)
         );
  FAx1_ASAP7_75t_SL U35430 ( .A(mult_x_1196_n1177), .B(n22306), .CI(
        mult_x_1196_n1153), .CON(mult_x_1196_n1144), .SN(mult_x_1196_n1145) );
  OAI22xp5_ASAP7_75t_SL U35431 ( .A1(mult_x_1196_n2887), .A2(n24026), .B1(
        mult_x_1196_n2886), .B2(n24025), .Y(mult_x_1196_n2315) );
  FAx1_ASAP7_75t_SL U35432 ( .A(mult_x_1196_n2387), .B(mult_x_1196_n2355), 
        .CI(mult_x_1196_n2483), .CON(mult_x_1196_n1494), .SN(mult_x_1196_n1495) );
  INVx11_ASAP7_75t_SL U35433 ( .A(n23968), .Y(n23969) );
  FAx1_ASAP7_75t_SL U35434 ( .A(mult_x_1196_n1294), .B(n22347), .CI(
        mult_x_1196_n1263), .CON(mult_x_1196_n1259), .SN(mult_x_1196_n1260) );
  INVx1_ASAP7_75t_SL U35435 ( .A(mult_x_1196_n1922), .Y(mult_x_1196_n1912) );
  OAI21xp5_ASAP7_75t_SL U35436 ( .A1(mult_x_1196_n444), .A2(n22533), .B(
        mult_x_1196_n445), .Y(mult_x_1196_n443) );
  INVx4_ASAP7_75t_SL U35437 ( .A(n23962), .Y(n24081) );
  FAx1_ASAP7_75t_SL U35438 ( .A(n22357), .B(mult_x_1196_n1706), .CI(
        mult_x_1196_n1704), .CON(mult_x_1196_n1694), .SN(mult_x_1196_n1695) );
  INVx1_ASAP7_75t_SL U35439 ( .A(mult_x_1196_n1695), .Y(mult_x_1196_n1684) );
  INVx2_ASAP7_75t_SL U35440 ( .A(n24024), .Y(n24023) );
  INVx6_ASAP7_75t_SL U35441 ( .A(n24023), .Y(n24025) );
  XNOR2x2_ASAP7_75t_SL U35442 ( .A(n24062), .B(n23957), .Y(mult_x_1196_n3197)
         );
  INVx1_ASAP7_75t_SL U35443 ( .A(mult_x_1196_n674), .Y(mult_x_1196_n672) );
  INVx1_ASAP7_75t_SL U35444 ( .A(mult_x_1196_n377), .Y(mult_x_1196_n375) );
  AOI21xp5_ASAP7_75t_SL U35445 ( .A1(n24279), .A2(mult_x_1196_n375), .B(
        mult_x_1196_n366), .Y(mult_x_1196_n364) );
  OAI22xp5_ASAP7_75t_SL U35446 ( .A1(mult_x_1196_n3047), .A2(n23637), .B1(
        n24005), .B2(mult_x_1196_n3046), .Y(mult_x_1196_n2475) );
  FAx1_ASAP7_75t_SL U35447 ( .A(mult_x_1196_n2475), .B(mult_x_1196_n2507), 
        .CI(mult_x_1196_n2164), .CON(mult_x_1196_n1220), .SN(mult_x_1196_n1221) );
  OAI21xp5_ASAP7_75t_SL U35448 ( .A1(mult_x_1196_n515), .A2(mult_x_1196_n550), 
        .B(mult_x_1196_n516), .Y(mult_x_1196_n514) );
  OAI22xp5_ASAP7_75t_SL U35449 ( .A1(mult_x_1196_n2934), .A2(n22781), .B1(
        mult_x_1196_n2933), .B2(n24020), .Y(mult_x_1196_n2362) );
  NAND2xp5_ASAP7_75t_SL U35450 ( .A(mult_x_1196_n1614), .B(mult_x_1196_n1613), 
        .Y(mult_x_1196_n614) );
  NAND2xp5_ASAP7_75t_SL U35451 ( .A(mult_x_1196_n1225), .B(n24282), .Y(
        mult_x_1196_n529) );
  NAND2xp5_ASAP7_75t_SL U35452 ( .A(n22353), .B(mult_x_1196_n1105), .Y(
        mult_x_1196_n489) );
  OAI22xp5_ASAP7_75t_SL U35453 ( .A1(mult_x_1196_n2815), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2814), .Y(mult_x_1196_n2249) );
  INVx1_ASAP7_75t_SL U35454 ( .A(mult_x_1196_n506), .Y(mult_x_1196_n795) );
  XNOR2x2_ASAP7_75t_SL U35455 ( .A(n24051), .B(n22395), .Y(mult_x_1196_n2812)
         );
  OAI22xp5_ASAP7_75t_SL U35456 ( .A1(mult_x_1196_n2813), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2812), .Y(mult_x_1196_n2247) );
  FAx1_ASAP7_75t_SL U35457 ( .A(mult_x_1196_n2247), .B(mult_x_1196_n995), .CI(
        mult_x_1196_n2186), .CON(mult_x_1196_n975), .SN(mult_x_1196_n976) );
  NAND2xp5_ASAP7_75t_SL U35458 ( .A(mult_x_1196_n997), .B(mult_x_1196_n979), 
        .Y(mult_x_1196_n423) );
  OAI21xp5_ASAP7_75t_SL U35459 ( .A1(mult_x_1196_n531), .A2(mult_x_1196_n580), 
        .B(mult_x_1196_n532), .Y(mult_x_1196_n530) );
  BUFx3_ASAP7_75t_SL U35460 ( .A(n23990), .Y(n24151) );
  INVx6_ASAP7_75t_SL U35461 ( .A(n23977), .Y(n23978) );
  AOI21xp5_ASAP7_75t_SL U35462 ( .A1(mult_x_1196_n534), .A2(mult_x_1196_n517), 
        .B(mult_x_1196_n518), .Y(mult_x_1196_n516) );
  OAI22xp5_ASAP7_75t_SL U35463 ( .A1(mult_x_1196_n2943), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2942), .Y(mult_x_1196_n2371) );
  OAI22xp5_ASAP7_75t_SL U35464 ( .A1(mult_x_1196_n2948), .A2(n22779), .B1(
        n22694), .B2(mult_x_1196_n2947), .Y(mult_x_1196_n2376) );
  INVx1_ASAP7_75t_SL U35465 ( .A(n18921), .Y(mult_x_1196_n552) );
  OAI22xp5_ASAP7_75t_SL U35466 ( .A1(mult_x_1196_n2811), .A2(n24034), .B1(
        n18402), .B2(mult_x_1196_n2810), .Y(mult_x_1196_n2245) );
  NOR2x1_ASAP7_75t_SL U35467 ( .A(mult_x_1196_n515), .B(mult_x_1196_n549), .Y(
        mult_x_1196_n513) );
  XNOR2x2_ASAP7_75t_SL U35468 ( .A(n24058), .B(n23658), .Y(mult_x_1196_n3125)
         );
  FAx1_ASAP7_75t_SL U35469 ( .A(n18906), .B(mult_x_1196_n1057), .CI(
        mult_x_1196_n1044), .CON(mult_x_1196_n1045), .SN(mult_x_1196_n1046) );
  XNOR2x2_ASAP7_75t_SL U35470 ( .A(n24050), .B(n18307), .Y(mult_x_1196_n2811)
         );
  OAI22xp5_ASAP7_75t_SL U35471 ( .A1(mult_x_1196_n2812), .A2(n24034), .B1(
        n18402), .B2(mult_x_1196_n2811), .Y(mult_x_1196_n2246) );
  OAI21xp5_ASAP7_75t_SL U35472 ( .A1(mult_x_1196_n580), .A2(mult_x_1196_n542), 
        .B(mult_x_1196_n543), .Y(mult_x_1196_n541) );
  INVx1_ASAP7_75t_SL U35473 ( .A(mult_x_1196_n1142), .Y(mult_x_1196_n1136) );
  OAI22xp5_ASAP7_75t_SL U35474 ( .A1(mult_x_1196_n2820), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2819), .Y(mult_x_1196_n2254) );
  NAND2xp5_ASAP7_75t_SL U35475 ( .A(mult_x_1196_n1058), .B(mult_x_1196_n1037), 
        .Y(mult_x_1196_n460) );
  XNOR2x2_ASAP7_75t_SL U35476 ( .A(n24047), .B(n22395), .Y(mult_x_1196_n2808)
         );
  FAx1_ASAP7_75t_SL U35477 ( .A(mult_x_1196_n1047), .B(mult_x_1196_n1021), 
        .CI(mult_x_1196_n1027), .CON(mult_x_1196_n1022), .SN(mult_x_1196_n1023) );
  XNOR2x2_ASAP7_75t_SL U35478 ( .A(n24055), .B(n22395), .Y(mult_x_1196_n2816)
         );
  OAI22xp5_ASAP7_75t_SL U35479 ( .A1(mult_x_1196_n2816), .A2(n24034), .B1(
        n22251), .B2(mult_x_1196_n2815), .Y(mult_x_1196_n2250) );
  OAI21xp5_ASAP7_75t_SL U35480 ( .A1(mult_x_1196_n1048), .A2(n18907), .B(
        n24249), .Y(mult_x_1196_n1039) );
  INVx1_ASAP7_75t_SL U35481 ( .A(mult_x_1196_n432), .Y(mult_x_1196_n434) );
  XNOR2x2_ASAP7_75t_SL U35482 ( .A(n24065), .B(n22449), .Y(mult_x_1196_n3234)
         );
  XNOR2x2_ASAP7_75t_SL U35483 ( .A(n24061), .B(n23955), .Y(mult_x_1196_n3230)
         );
  NAND2xp5_ASAP7_75t_SL U35484 ( .A(mult_x_1196_n1820), .B(mult_x_1196_n1797), 
        .Y(mult_x_1196_n652) );
  OAI21xp5_ASAP7_75t_SL U35485 ( .A1(mult_x_1196_n364), .A2(mult_x_1196_n334), 
        .B(mult_x_1196_n335), .Y(mult_x_1196_n333) );
  AOI21xp5_ASAP7_75t_SL U35486 ( .A1(mult_x_1196_n333), .A2(n23474), .B(
        mult_x_1196_n315), .Y(mult_x_1196_n313) );
  FAx1_ASAP7_75t_SL U35487 ( .A(mult_x_1196_n907), .B(mult_x_1196_n889), .CI(
        mult_x_1196_n894), .CON(mult_x_1196_n890), .SN(mult_x_1196_n891) );
  INVx1_ASAP7_75t_SL U35488 ( .A(mult_x_1196_n1117), .Y(mult_x_1196_n1110) );
  FAx1_ASAP7_75t_SL U35489 ( .A(mult_x_1196_n2472), .B(mult_x_1196_n2254), 
        .CI(mult_x_1196_n2408), .CON(mult_x_1196_n1130), .SN(mult_x_1196_n1131) );
  NAND2xp5_ASAP7_75t_SL U35490 ( .A(mult_x_1196_n1083), .B(mult_x_1196_n1059), 
        .Y(mult_x_1196_n475) );
  OAI22xp5_ASAP7_75t_SL U35491 ( .A1(mult_x_1196_n3201), .A2(n23989), .B1(
        mult_x_1196_n3200), .B2(n24106), .Y(mult_x_1196_n2625) );
  NAND2xp5_ASAP7_75t_SL U35492 ( .A(mult_x_1196_n1889), .B(mult_x_1196_n1869), 
        .Y(mult_x_1196_n674) );
  NAND2xp5_ASAP7_75t_SL U35493 ( .A(mult_x_1196_n674), .B(n24298), .Y(
        mult_x_1196_n267) );
  INVx1_ASAP7_75t_SL U35494 ( .A(mult_x_1196_n897), .Y(mult_x_1196_n889) );
  FAx1_ASAP7_75t_SL U35495 ( .A(mult_x_1196_n1077), .B(mult_x_1196_n1075), 
        .CI(mult_x_1196_n1055), .CON(mult_x_1196_n1047), .SN(mult_x_1196_n1048) );
  OAI22xp5_ASAP7_75t_SL U35496 ( .A1(mult_x_1196_n2955), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2954), .Y(mult_x_1196_n2383) );
  OAI22xp5_ASAP7_75t_SL U35497 ( .A1(mult_x_1196_n2959), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2958), .Y(mult_x_1196_n2387) );
  OAI22xp5_ASAP7_75t_SL U35498 ( .A1(mult_x_1196_n2958), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2957), .Y(mult_x_1196_n2386) );
  INVx1_ASAP7_75t_SL U35499 ( .A(n23990), .Y(n24114) );
  NAND2x1p5_ASAP7_75t_SL U35500 ( .A(mult_x_1196_n3327), .B(n24114), .Y(n23993) );
  OAI22xp5_ASAP7_75t_SL U35501 ( .A1(mult_x_1196_n2876), .A2(n22464), .B1(
        mult_x_1196_n2875), .B2(n18305), .Y(mult_x_1196_n960) );
  FAx1_ASAP7_75t_SL U35502 ( .A(mult_x_1196_n1133), .B(mult_x_1196_n2222), 
        .CI(mult_x_1196_n2376), .CON(mult_x_1196_n1128), .SN(mult_x_1196_n1129) );
  AOI21xp5_ASAP7_75t_SL U35503 ( .A1(mult_x_1196_n709), .A2(mult_x_1196_n717), 
        .B(mult_x_1196_n710), .Y(mult_x_1196_n708) );
  OAI22xp5_ASAP7_75t_SL U35504 ( .A1(mult_x_1196_n3226), .A2(n18597), .B1(
        n22538), .B2(mult_x_1196_n3225), .Y(mult_x_1196_n2650) );
  BUFx6f_ASAP7_75t_SL U35505 ( .A(n24027), .Y(n24026) );
  OAI22xp5_ASAP7_75t_SL U35506 ( .A1(mult_x_1196_n3234), .A2(n24121), .B1(
        mult_x_1196_n3233), .B2(n23984), .Y(mult_x_1196_n2658) );
  NAND2xp5_ASAP7_75t_SL U35507 ( .A(mult_x_1196_n1969), .B(mult_x_1196_n1968), 
        .Y(mult_x_1196_n701) );
  INVx1_ASAP7_75t_SL U35508 ( .A(mult_x_1196_n1747), .Y(n24085) );
  INVx2_ASAP7_75t_SL U35509 ( .A(n24037), .Y(n24036) );
  NAND2xp5_ASAP7_75t_SL U35510 ( .A(mult_x_1196_n978), .B(mult_x_1196_n964), 
        .Y(mult_x_1196_n416) );
  OAI21xp5_ASAP7_75t_SL U35511 ( .A1(mult_x_1196_n416), .A2(mult_x_1196_n393), 
        .B(mult_x_1196_n394), .Y(mult_x_1196_n392) );
  INVx1_ASAP7_75t_SL U35512 ( .A(mult_x_1196_n2084), .Y(mult_x_1196_n2077) );
  AOI21xp5_ASAP7_75t_SL U35513 ( .A1(mult_x_1196_n735), .A2(n24290), .B(
        mult_x_1196_n732), .Y(mult_x_1196_n730) );
  NAND2xp5_ASAP7_75t_SL U35514 ( .A(mult_x_1196_n1744), .B(n24269), .Y(
        mult_x_1196_n636) );
  OAI21xp5_ASAP7_75t_SL U35515 ( .A1(n24175), .A2(mult_x_1196_n434), .B(
        mult_x_1196_n423), .Y(mult_x_1196_n421) );
  XNOR2x2_ASAP7_75t_SL U35516 ( .A(n24057), .B(n23089), .Y(mult_x_1196_n2886)
         );
  OAI22xp5_ASAP7_75t_SL U35517 ( .A1(mult_x_1196_n2757), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2756), .Y(mult_x_1196_n2194) );
  FAx1_ASAP7_75t_SL U35518 ( .A(mult_x_1196_n1217), .B(n24263), .CI(
        mult_x_1196_n1221), .CON(mult_x_1196_n1209), .SN(mult_x_1196_n1210) );
  OAI22xp5_ASAP7_75t_SL U35519 ( .A1(mult_x_1196_n3269), .A2(n23982), .B1(
        n23980), .B2(mult_x_1196_n3268), .Y(mult_x_1196_n2693) );
  NAND2xp5_ASAP7_75t_SL U35520 ( .A(n22334), .B(n23888), .Y(mult_x_1196_n715)
         );
  OAI21xp5_ASAP7_75t_SL U35521 ( .A1(mult_x_1196_n715), .A2(n22333), .B(
        mult_x_1196_n712), .Y(mult_x_1196_n710) );
  XNOR2x2_ASAP7_75t_SL U35522 ( .A(n24045), .B(n22897), .Y(mult_x_1196_n2840)
         );
  XNOR2x2_ASAP7_75t_SL U35523 ( .A(n24045), .B(n23964), .Y(mult_x_1196_n3010)
         );
  XNOR2x2_ASAP7_75t_SL U35524 ( .A(n24045), .B(n22394), .Y(mult_x_1196_n3078)
         );
  XNOR2x2_ASAP7_75t_SL U35525 ( .A(n24045), .B(n23960), .Y(mult_x_1196_n3146)
         );
  XNOR2x2_ASAP7_75t_SL U35526 ( .A(n24045), .B(n18307), .Y(mult_x_1196_n2806)
         );
  XNOR2x2_ASAP7_75t_SL U35527 ( .A(n24045), .B(n22968), .Y(mult_x_1196_n2772)
         );
  XNOR2x2_ASAP7_75t_SL U35528 ( .A(n24045), .B(n23976), .Y(mult_x_1196_n2738)
         );
  OAI22xp5_ASAP7_75t_SL U35529 ( .A1(mult_x_1196_n2758), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2757), .Y(mult_x_1196_n2195) );
  OAI22xp5_ASAP7_75t_SL U35530 ( .A1(mult_x_1196_n3045), .A2(n18561), .B1(
        n18550), .B2(mult_x_1196_n3044), .Y(mult_x_1196_n2473) );
  OAI22xp5_ASAP7_75t_SL U35531 ( .A1(mult_x_1196_n3141), .A2(n23999), .B1(
        n23996), .B2(mult_x_1196_n3140), .Y(mult_x_1196_n2565) );
  INVx1_ASAP7_75t_SL U35532 ( .A(mult_x_1196_n728), .Y(mult_x_1196_n726) );
  AOI21xp5_ASAP7_75t_SL U35533 ( .A1(n24307), .A2(mult_x_1196_n726), .B(
        mult_x_1196_n721), .Y(mult_x_1196_n719) );
  INVx1_ASAP7_75t_SL U35534 ( .A(mult_x_1196_n1967), .Y(mult_x_1196_n1954) );
  NAND2xp5_ASAP7_75t_SL U35535 ( .A(mult_x_1196_n1932), .B(mult_x_1196_n1929), 
        .Y(mult_x_1196_n690) );
  OAI22xp5_ASAP7_75t_SL U35536 ( .A1(mult_x_1196_n3012), .A2(n24009), .B1(
        mult_x_1196_n3011), .B2(n23442), .Y(mult_x_1196_n2440) );
  OAI21xp5_ASAP7_75t_SL U35537 ( .A1(mult_x_1196_n482), .A2(mult_x_1196_n474), 
        .B(mult_x_1196_n475), .Y(mult_x_1196_n473) );
  OAI22xp5_ASAP7_75t_SL U35538 ( .A1(mult_x_1196_n2944), .A2(n23141), .B1(
        n24017), .B2(mult_x_1196_n2943), .Y(mult_x_1196_n2372) );
  INVx2_ASAP7_75t_SL U35539 ( .A(mult_x_1196_n1340), .Y(mult_x_1196_n1329) );
  NAND2x1p5_ASAP7_75t_SL U35540 ( .A(mult_x_1196_n517), .B(mult_x_1196_n533), 
        .Y(mult_x_1196_n515) );
  OAI22xp5_ASAP7_75t_SL U35541 ( .A1(mult_x_1196_n2856), .A2(n24031), .B1(
        n24030), .B2(mult_x_1196_n2855), .Y(mult_x_1196_n2290) );
  INVx1_ASAP7_75t_SL U35542 ( .A(n24028), .Y(n24029) );
  OAI22xp5_ASAP7_75t_SL U35543 ( .A1(mult_x_1196_n3207), .A2(n23072), .B1(
        mult_x_1196_n3206), .B2(n24106), .Y(mult_x_1196_n2631) );
  INVx1_ASAP7_75t_SL U35544 ( .A(mult_x_1196_n2063), .Y(mult_x_1196_n2054) );
  FAx1_ASAP7_75t_SL U35545 ( .A(mult_x_1196_n989), .B(mult_x_1196_n976), .CI(
        mult_x_1196_n972), .CON(mult_x_1196_n967), .SN(mult_x_1196_n968) );
  BUFx6f_ASAP7_75t_SL U35546 ( .A(u0_0_leon3x0_p0_muli[14]), .Y(n24073) );
  XNOR2x2_ASAP7_75t_SL U35547 ( .A(n24068), .B(n23091), .Y(mult_x_1196_n3101)
         );
  INVx2_ASAP7_75t_SL U35548 ( .A(n23990), .Y(n23991) );
  OAI21x1_ASAP7_75t_SL U35549 ( .A1(mult_x_1196_n3230), .A2(n18597), .B(n24299), .Y(n24148) );
  XNOR2x2_ASAP7_75t_SL U35550 ( .A(n24063), .B(n24231), .Y(mult_x_1196_n2960)
         );
  FAx1_ASAP7_75t_SL U35551 ( .A(mult_x_1196_n1010), .B(mult_x_1196_n1014), 
        .CI(mult_x_1196_n992), .CON(mult_x_1196_n986), .SN(mult_x_1196_n987)
         );
  NAND2xp5_ASAP7_75t_SL U35552 ( .A(n18983), .B(mult_x_1196_n818), .Y(
        mult_x_1196_n268) );
  OAI22xp5_ASAP7_75t_SL U35553 ( .A1(mult_x_1196_n2994), .A2(n24014), .B1(
        mult_x_1196_n2993), .B2(n24012), .Y(mult_x_1196_n2422) );
  OAI22xp5_ASAP7_75t_SL U35554 ( .A1(mult_x_1196_n3017), .A2(n24009), .B1(
        mult_x_1196_n3016), .B2(n23442), .Y(mult_x_1196_n2445) );
  OAI22xp5_ASAP7_75t_SL U35555 ( .A1(mult_x_1196_n3170), .A2(n23994), .B1(
        n23992), .B2(mult_x_1196_n3169), .Y(mult_x_1196_n2594) );
  AOI21xp5_ASAP7_75t_SL U35556 ( .A1(n24131), .A2(mult_x_1196_n1884), .B(
        n24132), .Y(n24256) );
  NOR2x1_ASAP7_75t_SL U35557 ( .A(n24125), .B(n24126), .Y(mult_x_1196_n1190)
         );
  INVx1_ASAP7_75t_SL U35558 ( .A(mult_x_1196_n1190), .Y(n24127) );
  INVx1_ASAP7_75t_SL U35559 ( .A(mult_x_1196_n1210), .Y(mult_x_1196_n1196) );
  NAND2xp5_ASAP7_75t_SL U35560 ( .A(mult_x_1196_n504), .B(n22663), .Y(
        mult_x_1196_n244) );
  OAI21xp5_ASAP7_75t_SL U35561 ( .A1(mult_x_1196_n623), .A2(mult_x_1196_n629), 
        .B(n23925), .Y(mult_x_1196_n622) );
  FAx1_ASAP7_75t_SL U35562 ( .A(mult_x_1196_n2218), .B(mult_x_1196_n2250), 
        .CI(mult_x_1196_n2404), .CON(mult_x_1196_n1032), .SN(mult_x_1196_n1033) );
  INVx1_ASAP7_75t_SL U35563 ( .A(mult_x_1196_n1322), .Y(mult_x_1196_n1323) );
  BUFx3_ASAP7_75t_SL U35564 ( .A(mult_x_1196_n135), .Y(n24039) );
  INVx1_ASAP7_75t_SL U35565 ( .A(mult_x_1196_n1495), .Y(mult_x_1196_n1480) );
  FAx1_ASAP7_75t_SL U35566 ( .A(mult_x_1196_n2461), .B(mult_x_1196_n2397), 
        .CI(mult_x_1196_n2429), .CON(mult_x_1196_n1812), .SN(mult_x_1196_n1813) );
  INVx6_ASAP7_75t_SL U35567 ( .A(add_x_735_A_4_), .Y(n23954) );
  XNOR2x2_ASAP7_75t_SL U35568 ( .A(n24074), .B(add_x_735_A_4_), .Y(
        mult_x_1196_n3243) );
  XNOR2x2_ASAP7_75t_SL U35569 ( .A(n24075), .B(n22449), .Y(mult_x_1196_n3244)
         );
  XNOR2x2_ASAP7_75t_SL U35570 ( .A(n24073), .B(n18393), .Y(mult_x_1196_n3242)
         );
  INVx1_ASAP7_75t_SL U35571 ( .A(mult_x_1196_n1194), .Y(mult_x_1196_n1163) );
  BUFx6f_ASAP7_75t_SL U35572 ( .A(u0_0_leon3x0_p0_muli[23]), .Y(n24063) );
  BUFx6f_ASAP7_75t_SL U35573 ( .A(n23998), .Y(n24000) );
  OAI22xp5_ASAP7_75t_SL U35574 ( .A1(mult_x_1196_n2962), .A2(n23142), .B1(
        n24017), .B2(mult_x_1196_n2961), .Y(mult_x_1196_n2390) );
  OAI22xp5_ASAP7_75t_SL U35575 ( .A1(mult_x_1196_n2930), .A2(n22781), .B1(
        mult_x_1196_n2929), .B2(n24020), .Y(mult_x_1196_n2358) );
  OAI22xp5_ASAP7_75t_SL U35576 ( .A1(mult_x_1196_n2913), .A2(n24022), .B1(
        mult_x_1196_n2912), .B2(n24020), .Y(mult_x_1196_n2341) );
  INVx1_ASAP7_75t_SL U35577 ( .A(mult_x_1196_n1368), .Y(n24153) );
  NAND2xp5_ASAP7_75t_SL U35578 ( .A(n24194), .B(mult_x_1196_n1297), .Y(n24195)
         );
  NAND2xp5_ASAP7_75t_SL U35579 ( .A(n24146), .B(mult_x_1196_n1042), .Y(n24147)
         );
  OAI22xp5_ASAP7_75t_SL U35580 ( .A1(mult_x_1196_n3220), .A2(n22647), .B1(
        mult_x_1196_n3219), .B2(n23984), .Y(mult_x_1196_n2644) );
  OAI22xp5_ASAP7_75t_SL U35581 ( .A1(mult_x_1196_n3244), .A2(n24121), .B1(
        mult_x_1196_n3243), .B2(n23984), .Y(mult_x_1196_n2668) );
  OAI22xp5_ASAP7_75t_SL U35582 ( .A1(mult_x_1196_n2933), .A2(n24021), .B1(
        mult_x_1196_n2932), .B2(n24020), .Y(mult_x_1196_n2361) );
  BUFx6f_ASAP7_75t_SL U35583 ( .A(n23956), .Y(n24205) );
  BUFx6f_ASAP7_75t_SL U35584 ( .A(mult_x_1196_n99), .Y(n24022) );
  OAI22xp5_ASAP7_75t_SL U35585 ( .A1(mult_x_1196_n2939), .A2(n24022), .B1(
        mult_x_1196_n2938), .B2(n24020), .Y(mult_x_1196_n2367) );
  OAI22xp5_ASAP7_75t_SL U35586 ( .A1(mult_x_1196_n2928), .A2(n24022), .B1(
        mult_x_1196_n2927), .B2(n24020), .Y(mult_x_1196_n2356) );
  OAI22xp5_ASAP7_75t_SL U35587 ( .A1(mult_x_1196_n2921), .A2(n24022), .B1(
        mult_x_1196_n2920), .B2(n24020), .Y(mult_x_1196_n2349) );
  INVx1_ASAP7_75t_SL U35588 ( .A(mult_x_1196_n1145), .Y(n24079) );
  NAND2xp5_ASAP7_75t_SL U35589 ( .A(n24096), .B(n24097), .Y(n24098) );
  OAI22xp5_ASAP7_75t_SL U35590 ( .A1(mult_x_1196_n3065), .A2(n23637), .B1(
        n24005), .B2(mult_x_1196_n3064), .Y(mult_x_1196_n2493) );
  OAI22xp5_ASAP7_75t_SL U35591 ( .A1(mult_x_1196_n2897), .A2(n24026), .B1(
        mult_x_1196_n2896), .B2(n24025), .Y(mult_x_1196_n2325) );
  OAI22xp5_ASAP7_75t_SL U35592 ( .A1(mult_x_1196_n2769), .A2(n24041), .B1(
        n24040), .B2(mult_x_1196_n2768), .Y(mult_x_1196_n2206) );
  OR2x2_ASAP7_75t_SL U35593 ( .A(add_x_735_A_32_), .B(u0_0_leon3x0_p0_divi[30]), .Y(n24313) );
  AO21x1_ASAP7_75t_SL U35594 ( .A1(add_x_735_n62), .A2(add_x_735_n45), .B(
        add_x_735_n46), .Y(n24314) );
  AND2x2_ASAP7_75t_SL U35595 ( .A(add_x_735_n45), .B(add_x_735_n61), .Y(n24315) );
  NOR2xp33_ASAP7_75t_SL U35596 ( .A(n23396), .B(u0_0_leon3x0_p0_divi[12]), .Y(
        add_x_735_n198) );
  NOR2xp33_ASAP7_75t_SL U35597 ( .A(n18908), .B(add_x_735_A_2_), .Y(
        add_x_735_n266) );
  NOR2xp33_ASAP7_75t_SL U35598 ( .A(n23969), .B(u0_0_leon3x0_p0_divi[20]), .Y(
        add_x_735_n130) );
  OAI21xp5_ASAP7_75t_SL U35599 ( .A1(add_x_735_n184), .A2(add_x_735_n149), .B(
        add_x_735_n150), .Y(add_x_735_n148) );
  AOI21x1_ASAP7_75t_SL U35600 ( .A1(add_x_735_n147), .A2(add_x_735_n215), .B(
        add_x_735_n148), .Y(add_x_735_n1) );
  OAI21xp5_ASAP7_75t_SL U35601 ( .A1(add_x_735_n156), .A2(add_x_735_n214), .B(
        add_x_735_n157), .Y(add_x_735_n155) );
  NAND2xp5_ASAP7_75t_SL U35602 ( .A(u0_0_leon3x0_p0_divi[1]), .B(n22939), .Y(
        add_x_735_n263) );
  NAND2xp5_ASAP7_75t_SL U35603 ( .A(n23091), .B(u0_0_leon3x0_p0_divi[10]), .Y(
        add_x_735_n213) );
  OR2x2_ASAP7_75t_SL U35604 ( .A(u0_0_leon3x0_p0_div0_vaddin1[32]), .B(
        u0_0_leon3x0_p0_div0_b[32]), .Y(n24316) );
  OA21x2_ASAP7_75t_SL U35605 ( .A1(DP_OP_5187J1_124_3275_n304), .A2(
        DP_OP_5187J1_124_3275_n306), .B(DP_OP_5187J1_124_3275_n305), .Y(n24317) );
  AOI21xp5_ASAP7_75t_SL U35606 ( .A1(DP_OP_5187J1_124_3275_n167), .A2(
        DP_OP_5187J1_124_3275_n182), .B(DP_OP_5187J1_124_3275_n168), .Y(
        DP_OP_5187J1_124_3275_n162) );
  OAI21x1_ASAP7_75t_SL U35607 ( .A1(DP_OP_5187J1_124_3275_n162), .A2(
        DP_OP_5187J1_124_3275_n127), .B(DP_OP_5187J1_124_3275_n128), .Y(
        DP_OP_5187J1_124_3275_n3) );
  OAI21xp5_ASAP7_75t_SL U35608 ( .A1(n22225), .A2(DP_OP_5187J1_124_3275_n43), 
        .B(DP_OP_5187J1_124_3275_n44), .Y(DP_OP_5187J1_124_3275_n42) );
  XNOR2x2_ASAP7_75t_SL U35609 ( .A(DP_OP_5187J1_124_3275_n7), .B(
        DP_OP_5187J1_124_3275_n42), .Y(u0_0_leon3x0_p0_div0_addout_32_) );
  NAND3xp33_ASAP7_75t_SL U35610 ( .A(n24407), .B(n18871), .C(n24408), .Y(
        n24318) );
  A2O1A1Ixp33_ASAP7_75t_SL U35611 ( .A1(n18871), .A2(n24408), .B(n24407), .C(
        n24318), .Y(timer0_res_10_) );
  NAND3xp33_ASAP7_75t_SL U35612 ( .A(n24406), .B(n24322), .C(n24407), .Y(
        n24321) );
  A2O1A1Ixp33_ASAP7_75t_SL U35613 ( .A1(n24322), .A2(n24407), .B(n24406), .C(
        n24321), .Y(timer0_res_11_) );
  NAND3xp33_ASAP7_75t_SL U35614 ( .A(n24405), .B(n24327), .C(n24406), .Y(
        n24324) );
  A2O1A1Ixp33_ASAP7_75t_SL U35615 ( .A1(n24327), .A2(n24406), .B(n24405), .C(
        n24324), .Y(timer0_res_12_) );
  NAND3xp33_ASAP7_75t_SL U35616 ( .A(n24404), .B(n18874), .C(n24405), .Y(
        n24326) );
  A2O1A1Ixp33_ASAP7_75t_SL U35617 ( .A1(n18874), .A2(n24405), .B(n24404), .C(
        n24326), .Y(timer0_res_13_) );
  NAND3xp33_ASAP7_75t_SL U35618 ( .A(n24403), .B(n24330), .C(n24404), .Y(
        n24329) );
  A2O1A1Ixp33_ASAP7_75t_SL U35619 ( .A1(n24330), .A2(n24404), .B(n24403), .C(
        n24329), .Y(timer0_res_14_) );
  NAND3xp33_ASAP7_75t_SL U35620 ( .A(n24402), .B(n24335), .C(n24403), .Y(
        n24332) );
  A2O1A1Ixp33_ASAP7_75t_SL U35621 ( .A1(n24335), .A2(n24403), .B(n24402), .C(
        n24332), .Y(timer0_res_15_) );
  NAND3xp33_ASAP7_75t_SL U35622 ( .A(n24401), .B(n18868), .C(n24402), .Y(
        n24334) );
  A2O1A1Ixp33_ASAP7_75t_SL U35623 ( .A1(n18868), .A2(n24402), .B(n24401), .C(
        n24334), .Y(timer0_res_16_) );
  NAND3xp33_ASAP7_75t_SL U35624 ( .A(n24400), .B(n24338), .C(n24401), .Y(
        n24337) );
  A2O1A1Ixp33_ASAP7_75t_SL U35625 ( .A1(n24338), .A2(n24401), .B(n24400), .C(
        n24337), .Y(timer0_res_17_) );
  NAND3xp33_ASAP7_75t_SL U35626 ( .A(n24399), .B(n24343), .C(n24400), .Y(
        n24340) );
  A2O1A1Ixp33_ASAP7_75t_SL U35627 ( .A1(n24343), .A2(n24400), .B(n24399), .C(
        n24340), .Y(timer0_res_18_) );
  NAND3xp33_ASAP7_75t_SL U35628 ( .A(n24398), .B(n18881), .C(n24399), .Y(
        n24342) );
  A2O1A1Ixp33_ASAP7_75t_SL U35629 ( .A1(n18881), .A2(n24399), .B(n24398), .C(
        n24342), .Y(timer0_res_19_) );
  NAND3xp33_ASAP7_75t_SL U35630 ( .A(n24397), .B(n24346), .C(n24398), .Y(
        n24345) );
  A2O1A1Ixp33_ASAP7_75t_SL U35631 ( .A1(n24346), .A2(n24398), .B(n24397), .C(
        n24345), .Y(timer0_res_20_) );
  NAND3xp33_ASAP7_75t_SL U35632 ( .A(n24396), .B(n24351), .C(n24397), .Y(
        n24348) );
  A2O1A1Ixp33_ASAP7_75t_SL U35633 ( .A1(n24351), .A2(n24397), .B(n24396), .C(
        n24348), .Y(timer0_res_21_) );
  NAND3xp33_ASAP7_75t_SL U35634 ( .A(n24395), .B(n24396), .C(n24353), .Y(
        n24350) );
  A2O1A1Ixp33_ASAP7_75t_SL U35635 ( .A1(n24353), .A2(n24396), .B(n24395), .C(
        n24350), .Y(timer0_res_22_) );
  NAND3xp33_ASAP7_75t_SL U35636 ( .A(n24394), .B(n24356), .C(n24395), .Y(
        n24352) );
  A2O1A1Ixp33_ASAP7_75t_SL U35637 ( .A1(n24356), .A2(n24395), .B(n24394), .C(
        n24352), .Y(timer0_res_23_) );
  NAND3xp33_ASAP7_75t_SL U35638 ( .A(n24393), .B(n24358), .C(n24394), .Y(
        n24355) );
  A2O1A1Ixp33_ASAP7_75t_SL U35639 ( .A1(n24358), .A2(n24394), .B(n24393), .C(
        n24355), .Y(timer0_res_24_) );
  NAND3xp33_ASAP7_75t_SL U35640 ( .A(n24392), .B(n24361), .C(n24393), .Y(
        n24357) );
  A2O1A1Ixp33_ASAP7_75t_SL U35641 ( .A1(n24361), .A2(n24393), .B(n24392), .C(
        n24357), .Y(timer0_res_25_) );
  NAND3xp33_ASAP7_75t_SL U35642 ( .A(timer0_N65), .B(n24363), .C(n24392), .Y(
        n24360) );
  A2O1A1Ixp33_ASAP7_75t_SL U35643 ( .A1(n24363), .A2(n24392), .B(timer0_N65), 
        .C(n24360), .Y(timer0_res_26_) );
  NAND3xp33_ASAP7_75t_SL U35644 ( .A(n24391), .B(n24366), .C(timer0_N65), .Y(
        n24362) );
  A2O1A1Ixp33_ASAP7_75t_SL U35645 ( .A1(n24366), .A2(timer0_N65), .B(n24391), 
        .C(n24362), .Y(timer0_res_27_) );
  NAND3xp33_ASAP7_75t_SL U35646 ( .A(n24390), .B(n24365), .C(n24391), .Y(
        n24364) );
  A2O1A1Ixp33_ASAP7_75t_SL U35647 ( .A1(n24365), .A2(n24391), .B(n24390), .C(
        n24364), .Y(timer0_res_28_) );
  NAND3xp33_ASAP7_75t_SL U35648 ( .A(n24415), .B(n24416), .C(n22430), .Y(
        n24369) );
  A2O1A1Ixp33_ASAP7_75t_SL U35649 ( .A1(n24416), .A2(n22430), .B(n24415), .C(
        n24369), .Y(timer0_res_2_) );
  NAND3xp33_ASAP7_75t_SL U35650 ( .A(n24388), .B(n24420), .C(n24389), .Y(
        n24370) );
  A2O1A1Ixp33_ASAP7_75t_SL U35651 ( .A1(n24420), .A2(n24389), .B(n24388), .C(
        n24370), .Y(timer0_res_30_) );
  NAND3xp33_ASAP7_75t_SL U35652 ( .A(n24414), .B(n24374), .C(n24415), .Y(
        n24371) );
  A2O1A1Ixp33_ASAP7_75t_SL U35653 ( .A1(n24374), .A2(n24415), .B(n24414), .C(
        n24371), .Y(timer0_res_3_) );
  NAND3xp33_ASAP7_75t_SL U35654 ( .A(n24413), .B(n24373), .C(n24414), .Y(
        n24372) );
  A2O1A1Ixp33_ASAP7_75t_SL U35655 ( .A1(n24373), .A2(n24414), .B(n24413), .C(
        n24372), .Y(timer0_res_4_) );
  NAND3xp33_ASAP7_75t_SL U35656 ( .A(n24412), .B(n24377), .C(n24413), .Y(
        n24376) );
  A2O1A1Ixp33_ASAP7_75t_SL U35657 ( .A1(n24377), .A2(n24413), .B(n24412), .C(
        n24376), .Y(timer0_res_5_) );
  NAND3xp33_ASAP7_75t_SL U35658 ( .A(n24411), .B(n24382), .C(n24412), .Y(
        n24379) );
  A2O1A1Ixp33_ASAP7_75t_SL U35659 ( .A1(n24382), .A2(n24412), .B(n24411), .C(
        n24379), .Y(timer0_res_6_) );
  NAND3xp33_ASAP7_75t_SL U35660 ( .A(n24410), .B(n23896), .C(n24411), .Y(
        n24380) );
  A2O1A1Ixp33_ASAP7_75t_SL U35661 ( .A1(n23896), .A2(n24411), .B(n24410), .C(
        n24380), .Y(timer0_res_7_) );
  NAND3xp33_ASAP7_75t_SL U35662 ( .A(n24409), .B(n24385), .C(n24410), .Y(
        n24384) );
  A2O1A1Ixp33_ASAP7_75t_SL U35663 ( .A1(n24385), .A2(n24410), .B(n24409), .C(
        n24384), .Y(timer0_res_8_) );
  NAND3xp33_ASAP7_75t_SL U35664 ( .A(n24408), .B(n24387), .C(n24409), .Y(
        n24386) );
  A2O1A1Ixp33_ASAP7_75t_SL U35665 ( .A1(n24387), .A2(n24409), .B(n24408), .C(
        n24386), .Y(timer0_res_9_) );
  NOR2xp33_ASAP7_75t_SL U35666 ( .A(timer0_N91), .B(timer0_N90), .Y(n24374) );
  NOR2xp33_ASAP7_75t_SL U35667 ( .A(n18865), .B(n24375), .Y(n24377) );
  NOR2xp33_ASAP7_75t_SL U35668 ( .A(timer0_N87), .B(n24378), .Y(n24382) );
  NOR2xp33_ASAP7_75t_SL U35669 ( .A(timer0_N85), .B(n24383), .Y(n24385) );
  NOR2xp33_ASAP7_75t_SL U35670 ( .A(timer0_N84), .B(n18854), .Y(n24387) );
  NOR2xp33_ASAP7_75t_SL U35671 ( .A(timer0_N82), .B(n24320), .Y(n24322) );
  NOR2xp33_ASAP7_75t_SL U35672 ( .A(timer0_N81), .B(n24325), .Y(n24327) );
  NOR2xp33_ASAP7_75t_SL U35673 ( .A(timer0_N79), .B(n24328), .Y(n24330) );
  NOR2xp33_ASAP7_75t_SL U35674 ( .A(timer0_N78), .B(n18856), .Y(n24335) );
  NOR2xp33_ASAP7_75t_SL U35675 ( .A(timer0_N76), .B(n24336), .Y(n24338) );
  NOR2xp33_ASAP7_75t_SL U35676 ( .A(n24341), .B(timer0_N75), .Y(n24343) );
  NOR2xp33_ASAP7_75t_SL U35677 ( .A(n24367), .B(timer0_N62), .Y(n24368) );
  AOI21xp33_ASAP7_75t_SRAM U35678 ( .A1(timer0_N62), .A2(n24420), .B(n24368), 
        .Y(timer0_res_29_) );
  NOR2xp33_ASAP7_75t_SL U35679 ( .A(timer0_N73), .B(n24344), .Y(n24346) );
  NOR2xp33_ASAP7_75t_SL U35680 ( .A(timer0_N63), .B(timer0_N64), .Y(n24417) );
  NOR3xp33_ASAP7_75t_SL U35681 ( .A(n24378), .B(timer0_N86), .C(timer0_N87), 
        .Y(n24381) );
  NOR3xp33_ASAP7_75t_SL U35682 ( .A(n24319), .B(timer0_N83), .C(timer0_N84), 
        .Y(n24323) );
  INVx1_ASAP7_75t_SL U35683 ( .A(timer0_N88), .Y(n24414) );
  NAND2xp5_ASAP7_75t_SL U35684 ( .A(n24339), .B(n24402), .Y(n24341) );
  NAND2xp5_ASAP7_75t_SL U35685 ( .A(n24323), .B(n24408), .Y(n24325) );
  NAND2xp5_ASAP7_75t_SL U35686 ( .A(n24358), .B(n24394), .Y(n24359) );
  NOR2x1_ASAP7_75t_SL U35687 ( .A(timer0_N67), .B(n24359), .Y(n24363) );
  NOR2x1_ASAP7_75t_SL U35688 ( .A(n18297), .B(n28769), .Y(n28677) );
  NAND2xp5_ASAP7_75t_SL U35689 ( .A(n24832), .B(n26850), .Y(n24866) );
  OAI21xp5_ASAP7_75t_SL U35690 ( .A1(n23980), .A2(n22392), .B(n25520), .Y(
        n29003) );
  NAND2xp5_ASAP7_75t_SL U35691 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__7_), .B(
        n23903), .Y(n25143) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U35692 ( .A1(n29144), .A2(n22449), .B(n28882), 
        .C(n28881), .Y(n28883) );
  INVx1_ASAP7_75t_SL U35693 ( .A(sr1_r_READY_), .Y(n31754) );
  NAND2xp5_ASAP7_75t_SL U35694 ( .A(n32705), .B(n31706), .Y(n32036) );
  INVx1_ASAP7_75t_SL U35695 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__LD_), .Y(n25152) );
  OAI21xp5_ASAP7_75t_SL U35696 ( .A1(n29561), .A2(n22392), .B(n25495), .Y(
        n29564) );
  OAI21xp5_ASAP7_75t_SL U35697 ( .A1(u0_0_leon3x0_p0_mul0_m3232_dwm_N48), .A2(
        n22378), .B(n25291), .Y(n4219) );
  OAI21xp5_ASAP7_75t_SL U35698 ( .A1(n22378), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N49), .B(n25293), .Y(n4217) );
  OAI21xp5_ASAP7_75t_SL U35699 ( .A1(n22378), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N53), .B(n25301), .Y(n4209) );
  OAI21xp5_ASAP7_75t_SL U35700 ( .A1(u0_0_leon3x0_p0_mul0_m3232_dwm_N46), .A2(
        n22378), .B(n25287), .Y(n4223) );
  OAI21xp5_ASAP7_75t_SL U35701 ( .A1(u0_0_leon3x0_p0_mul0_m3232_dwm_N47), .A2(
        n22378), .B(n25289), .Y(n4221) );
  OAI21xp5_ASAP7_75t_SL U35702 ( .A1(n22378), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N57), .B(n25308), .Y(n4201) );
  OAI21xp5_ASAP7_75t_SL U35703 ( .A1(n22378), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N50), .B(n25295), .Y(n4215) );
  OAI21xp5_ASAP7_75t_SL U35704 ( .A1(n22378), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N54), .B(n25303), .Y(n4207) );
  NAND2x1_ASAP7_75t_SL U35705 ( .A(n32030), .B(u0_0_leon3x0_p0_dci[3]), .Y(
        n31257) );
  OAI21xp5_ASAP7_75t_SL U35706 ( .A1(n31400), .A2(n26452), .B(n25213), .Y(
        n30949) );
  NAND2xp5_ASAP7_75t_SL U35707 ( .A(n26715), .B(n26714), .Y(n27263) );
  OAI21xp5_ASAP7_75t_SL U35708 ( .A1(n30635), .A2(n30634), .B(n30633), .Y(
        n30636) );
  NAND2xp5_ASAP7_75t_SL U35709 ( .A(n28766), .B(n28793), .Y(n30799) );
  INVx1_ASAP7_75t_SL U35710 ( .A(n28941), .Y(n30622) );
  INVx1_ASAP7_75t_SL U35711 ( .A(n29594), .Y(n28782) );
  INVx1_ASAP7_75t_SL U35712 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__4_), .Y(
        n31475) );
  NAND2xp5_ASAP7_75t_SL U35713 ( .A(n30007), .B(n27066), .Y(n28887) );
  NAND2xp5_ASAP7_75t_SL U35714 ( .A(n26441), .B(n26440), .Y(n29807) );
  NAND2xp5_ASAP7_75t_SL U35715 ( .A(n3897), .B(
        u0_0_leon3x0_p0_c0mmu_a0_r_BO__0_), .Y(n31602) );
  NAND2xp5_ASAP7_75t_SL U35716 ( .A(n32187), .B(n32188), .Y(n24815) );
  NAND2xp5_ASAP7_75t_SL U35717 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__12_), .B(
        n24687), .Y(n25099) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U35718 ( .A1(n18299), .A2(n25198), .B(n25147), 
        .C(n28850), .Y(n25149) );
  OAI21xp5_ASAP7_75t_SL U35719 ( .A1(n28254), .A2(n22399), .B(n26642), .Y(
        timer0_v_TIMERS__1__VALUE__3_) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U35720 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), .A2(n23898), .B(n31383), .C(
        n31382), .Y(n31388) );
  NAND2xp5_ASAP7_75t_SL U35721 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__6_), .B(
        n18862), .Y(n25112) );
  INVx1_ASAP7_75t_SL U35722 ( .A(n29592), .Y(n28779) );
  NAND2xp5_ASAP7_75t_SL U35723 ( .A(n24634), .B(n26174), .Y(n29594) );
  NAND2xp5_ASAP7_75t_SL U35724 ( .A(n24634), .B(n28480), .Y(n29592) );
  NAND2xp5_ASAP7_75t_SL U35725 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__28_), .B(
        n24687), .Y(n25101) );
  OAI21xp5_ASAP7_75t_SL U35726 ( .A1(n22428), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N52), .B(n25299), .Y(n4211) );
  NAND2xp5_ASAP7_75t_SL U35727 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__27_), .B(
        n18862), .Y(n25139) );
  OAI21xp5_ASAP7_75t_SL U35728 ( .A1(n22378), .A2(
        u0_0_leon3x0_p0_mul0_m3232_dwm_N51), .B(n25297), .Y(n4213) );
  AOI21x1_ASAP7_75t_SL U35729 ( .A1(n29869), .A2(n22375), .B(n25397), .Y(
        n32030) );
  BUFx6f_ASAP7_75t_SL U35730 ( .A(u0_0_leon3x0_p0_iu_r_E__LDBP2_), .Y(n24688)
         );
  OAI21xp5_ASAP7_75t_SL U35731 ( .A1(n29021), .A2(u0_0_leon3x0_p0_div0_vaddsub), .B(n29020), .Y(u0_0_leon3x0_p0_div0_b[0]) );
  NAND2xp5_ASAP7_75t_SL U35732 ( .A(n29021), .B(n24630), .Y(n29020) );
  INVxp33_ASAP7_75t_SRAM U35733 ( .A(resetn), .Y(n4828) );
  INVxp33_ASAP7_75t_SRAM U35734 ( .A(datain[15]), .Y(n4801) );
  INVxp33_ASAP7_75t_SRAM U35735 ( .A(datain[9]), .Y(n4807) );
  INVxp33_ASAP7_75t_SRAM U35736 ( .A(datain[18]), .Y(n4798) );
  INVxp33_ASAP7_75t_SRAM U35737 ( .A(datain[19]), .Y(n4797) );
  INVxp33_ASAP7_75t_SRAM U35738 ( .A(datain[10]), .Y(n4806) );
  INVxp33_ASAP7_75t_SRAM U35739 ( .A(datain[13]), .Y(n4803) );
  INVxp33_ASAP7_75t_SRAM U35740 ( .A(datain[4]), .Y(n4812) );
  INVxp33_ASAP7_75t_SRAM U35741 ( .A(datain[27]), .Y(n4789) );
  INVxp33_ASAP7_75t_SRAM U35742 ( .A(datain[5]), .Y(n4811) );
  INVxp33_ASAP7_75t_SRAM U35743 ( .A(datain[2]), .Y(n4814) );
  INVxp33_ASAP7_75t_SRAM U35744 ( .A(datain[0]), .Y(n4816) );
  INVxp33_ASAP7_75t_SRAM U35745 ( .A(datain[17]), .Y(n4799) );
  INVxp33_ASAP7_75t_SRAM U35746 ( .A(datain[20]), .Y(n4796) );
  INVxp33_ASAP7_75t_SRAM U35747 ( .A(datain[14]), .Y(n4802) );
  INVxp33_ASAP7_75t_SRAM U35748 ( .A(datain[24]), .Y(n4792) );
  INVxp33_ASAP7_75t_SRAM U35749 ( .A(datain[16]), .Y(n4800) );
  INVxp33_ASAP7_75t_SRAM U35750 ( .A(datain[3]), .Y(n4813) );
  INVxp33_ASAP7_75t_SRAM U35751 ( .A(datain[12]), .Y(n4804) );
  INVxp33_ASAP7_75t_SRAM U35752 ( .A(datain[21]), .Y(n4795) );
  INVxp33_ASAP7_75t_SRAM U35753 ( .A(datain[22]), .Y(n4794) );
  INVxp33_ASAP7_75t_SRAM U35754 ( .A(datain[7]), .Y(n4809) );
  INVxp33_ASAP7_75t_SRAM U35755 ( .A(datain[26]), .Y(n4790) );
  INVxp33_ASAP7_75t_SRAM U35756 ( .A(datain[25]), .Y(n4791) );
  INVxp33_ASAP7_75t_SRAM U35757 ( .A(datain[8]), .Y(n4808) );
  INVxp33_ASAP7_75t_SRAM U35758 ( .A(datain[1]), .Y(n4815) );
  INVxp33_ASAP7_75t_SRAM U35759 ( .A(datain[11]), .Y(n4805) );
  INVxp33_ASAP7_75t_SRAM U35760 ( .A(datain[29]), .Y(n4787) );
  INVxp33_ASAP7_75t_SRAM U35761 ( .A(datain[31]), .Y(n4785) );
  INVxp33_ASAP7_75t_SRAM U35762 ( .A(datain[23]), .Y(n4793) );
  INVxp33_ASAP7_75t_SRAM U35763 ( .A(datain[30]), .Y(n4786) );
  INVxp33_ASAP7_75t_SRAM U35764 ( .A(rxd1), .Y(n4784) );
  INVxp33_ASAP7_75t_SRAM U35765 ( .A(datain[6]), .Y(n4810) );
  INVxp33_ASAP7_75t_SRAM U35766 ( .A(datain[28]), .Y(n4788) );
  OAI21xp33_ASAP7_75t_SRAM U35767 ( .A1(n32398), .A2(n32381), .B(n32370), .Y(
        dc_data[18]) );
  AOI21xp33_ASAP7_75t_SRAM U35768 ( .A1(dc_q[16]), .A2(n32385), .B(n32355), 
        .Y(n32359) );
  AOI21xp33_ASAP7_75t_SRAM U35769 ( .A1(dc_q[19]), .A2(n32385), .B(n32372), 
        .Y(n32374) );
  AOI21xp33_ASAP7_75t_SRAM U35770 ( .A1(dc_q[17]), .A2(n32385), .B(n32362), 
        .Y(n32364) );
  INVxp33_ASAP7_75t_SRAM U35771 ( .A(n32386), .Y(n32381) );
  INVxp33_ASAP7_75t_SRAM U35772 ( .A(u0_0_leon3x0_p0_iu_r_X__NERROR_), .Y(
        errorn) );
  INVxp33_ASAP7_75t_SRAM U35773 ( .A(n32356), .Y(n32357) );
  INVxp33_ASAP7_75t_SRAM U35774 ( .A(n32425), .Y(n32414) );
  INVxp33_ASAP7_75t_SRAM U35775 ( .A(n32434), .Y(n32409) );
  OAI21xp33_ASAP7_75t_SRAM U35776 ( .A1(n32426), .A2(n32425), .B(n32424), .Y(
        dc_data[30]) );
  INVxp33_ASAP7_75t_SRAM U35777 ( .A(n32351), .Y(n32352) );
  AOI22xp33_ASAP7_75t_SRAM U35778 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[3]), .A2(
        n32448), .B1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__3_), .B2(n32447), .Y(
        n32442) );
  AOI22xp33_ASAP7_75t_SRAM U35779 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[4]), .A2(
        n32448), .B1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__4_), .B2(n32447), .Y(
        n32449) );
  AOI22xp33_ASAP7_75t_SRAM U35780 ( .A1(it_q[0]), .A2(n32519), .B1(n32518), 
        .B2(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__0_), .Y(n32466) );
  AOI22xp33_ASAP7_75t_SRAM U35781 ( .A1(it_q[1]), .A2(n32519), .B1(n32518), 
        .B2(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__1_), .Y(n32473) );
  AOI22xp33_ASAP7_75t_SRAM U35782 ( .A1(it_q[2]), .A2(n32519), .B1(n32518), 
        .B2(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__2_), .Y(n32480) );
  AOI22xp33_ASAP7_75t_SRAM U35783 ( .A1(it_q[3]), .A2(n32519), .B1(n32518), 
        .B2(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__3_), .Y(n32488) );
  INVxp33_ASAP7_75t_SRAM U35784 ( .A(n32493), .Y(n32494) );
  AOI22xp33_ASAP7_75t_SRAM U35785 ( .A1(it_q[5]), .A2(n32519), .B1(n32518), 
        .B2(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__5_), .Y(n32502) );
  AOI22xp33_ASAP7_75t_SRAM U35786 ( .A1(it_q[6]), .A2(n32519), .B1(n32518), 
        .B2(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__6_), .Y(n32509) );
  AOI22xp33_ASAP7_75t_SRAM U35787 ( .A1(it_q[7]), .A2(n32519), .B1(n32518), 
        .B2(u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__7_), .Y(n32522) );
  INVxp33_ASAP7_75t_SRAM U35788 ( .A(n32490), .Y(n32519) );
  INVxp33_ASAP7_75t_SRAM U35789 ( .A(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__12_), .Y(n32525) );
  INVxp33_ASAP7_75t_SRAM U35790 ( .A(n3474), .Y(rf_addr_b[0]) );
  INVxp33_ASAP7_75t_SRAM U35791 ( .A(n3540), .Y(rf_addr_b[1]) );
  INVxp33_ASAP7_75t_SRAM U35792 ( .A(n2776), .Y(rf_addr_b[4]) );
  AOI22xp33_ASAP7_75t_SRAM U35793 ( .A1(dc_q[11]), .A2(n32344), .B1(n32619), 
        .B2(n24643), .Y(n32335) );
  AOI22xp33_ASAP7_75t_SRAM U35794 ( .A1(dc_q[10]), .A2(n32344), .B1(n32617), 
        .B2(n24643), .Y(n32331) );
  INVxp33_ASAP7_75t_SRAM U35795 ( .A(n32345), .Y(n32341) );
  AOI22xp33_ASAP7_75t_SRAM U35796 ( .A1(dc_q[8]), .A2(n32344), .B1(n32613), 
        .B2(n24643), .Y(n32324) );
  INVxp33_ASAP7_75t_SRAM U35797 ( .A(n32353), .Y(n24642) );
  OAI21xp33_ASAP7_75t_SRAM U35798 ( .A1(n32319), .A2(n32408), .B(n32312), .Y(
        dc_data[5]) );
  AOI22xp33_ASAP7_75t_SRAM U35799 ( .A1(dc_q[5]), .A2(n32318), .B1(n32607), 
        .B2(n24643), .Y(n32312) );
  OAI21xp33_ASAP7_75t_SRAM U35800 ( .A1(n32319), .A2(n32378), .B(n32309), .Y(
        dc_data[4]) );
  AOI22xp33_ASAP7_75t_SRAM U35801 ( .A1(dc_q[4]), .A2(n32318), .B1(n32605), 
        .B2(n24643), .Y(n32309) );
  INVxp33_ASAP7_75t_SRAM U35802 ( .A(n32406), .Y(n32378) );
  OAI21xp33_ASAP7_75t_SRAM U35803 ( .A1(n32319), .A2(n32398), .B(n32304), .Y(
        dc_data[2]) );
  AOI22xp33_ASAP7_75t_SRAM U35804 ( .A1(dc_q[2]), .A2(n32318), .B1(n32601), 
        .B2(n24643), .Y(n32304) );
  OAI21xp33_ASAP7_75t_SRAM U35805 ( .A1(n32319), .A2(n32299), .B(n32298), .Y(
        dc_data[0]) );
  AOI22xp33_ASAP7_75t_SRAM U35806 ( .A1(dc_q[0]), .A2(n32318), .B1(n32599), 
        .B2(n24643), .Y(n32298) );
  INVxp33_ASAP7_75t_SRAM U35807 ( .A(n32393), .Y(n32299) );
  AOI21xp33_ASAP7_75t_SRAM U35808 ( .A1(n32288), .A2(n32287), .B(n32340), .Y(
        n32319) );
  INVxp33_ASAP7_75t_SRAM U35809 ( .A(n32348), .Y(n32340) );
  INVxp33_ASAP7_75t_SRAM U35810 ( .A(n32349), .Y(n32285) );
  INVxp33_ASAP7_75t_SRAM U35811 ( .A(n32294), .Y(n32390) );
  INVxp33_ASAP7_75t_SRAM U35812 ( .A(n32388), .Y(n32286) );
  INVxp33_ASAP7_75t_SRAM U35813 ( .A(n32295), .Y(n32287) );
  AOI21xp33_ASAP7_75t_SRAM U35814 ( .A1(n32290), .A2(
        u0_0_leon3x0_p0_c0mmu_mmudci[0]), .B(n32149), .Y(n32295) );
  INVxp33_ASAP7_75t_SRAM U35815 ( .A(n32290), .Y(n32428) );
  AOI22xp33_ASAP7_75t_SRAM U35816 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[11]), 
        .A2(n32448), .B1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__11_), .B2(n32447), 
        .Y(n32269) );
  AOI22xp33_ASAP7_75t_SRAM U35817 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[7]), .A2(
        n32448), .B1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__7_), .B2(n32447), .Y(
        n32265) );
  AOI22xp33_ASAP7_75t_SRAM U35818 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__6_), 
        .A2(n32447), .B1(u0_0_leon3x0_p0_c0mmu_mmudci[6]), .B2(n32448), .Y(
        n32262) );
  AOI22xp33_ASAP7_75t_SRAM U35819 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[5]), .A2(
        n32448), .B1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__5_), .B2(n32447), .Y(
        n32260) );
  INVxp33_ASAP7_75t_SRAM U35820 ( .A(n32256), .Y(n32254) );
  O2A1O1Ixp5_ASAP7_75t_SL U35821 ( .A1(n32289), .A2(n32241), .B(n32240), .C(
        n32239), .Y(n32242) );
  INVxp33_ASAP7_75t_SRAM U35822 ( .A(n32231), .Y(n32235) );
  INVxp33_ASAP7_75t_SRAM U35823 ( .A(n32214), .Y(n32218) );
  INVxp33_ASAP7_75t_SRAM U35824 ( .A(n32239), .Y(n32204) );
  INVxp33_ASAP7_75t_SRAM U35825 ( .A(n3160), .Y(rf_addr_a[7]) );
  INVxp33_ASAP7_75t_SRAM U35826 ( .A(n32201), .Y(n32275) );
  INVxp33_ASAP7_75t_SRAM U35827 ( .A(n2706), .Y(rf_ce_a) );
  INVxp33_ASAP7_75t_SRAM U35828 ( .A(n3536), .Y(rf_addr_b[2]) );
  INVxp33_ASAP7_75t_SRAM U35829 ( .A(n24543), .Y(n24643) );
  INVxp33_ASAP7_75t_SRAM U35830 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_READ_), 
        .Y(n32144) );
  O2A1O1Ixp5_ASAP7_75t_SL U35831 ( .A1(n32692), .A2(n32691), .B(n32690), .C(
        n32694), .Y(n32693) );
  INVxp33_ASAP7_75t_SRAM U35832 ( .A(n32687), .Y(n32688) );
  INVxp33_ASAP7_75t_SRAM U35833 ( .A(n32686), .Y(n32691) );
  OAI22xp33_ASAP7_75t_SRAM U35834 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[24]), 
        .A2(n32593), .B1(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__24_), .B2(
        n32565), .Y(n32546) );
  INVxp33_ASAP7_75t_SRAM U35835 ( .A(n32594), .Y(n32585) );
  INVxp33_ASAP7_75t_SRAM U35836 ( .A(n32595), .Y(n32588) );
  OAI22xp33_ASAP7_75t_SRAM U35837 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[26]), 
        .A2(n32593), .B1(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__26_), .B2(
        n32565), .Y(n32552) );
  OAI22xp33_ASAP7_75t_SRAM U35838 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[25]), 
        .A2(n32593), .B1(u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__25_), .B2(
        n32565), .Y(n32549) );
  NAND2xp5_ASAP7_75t_SL U35839 ( .A(n18848), .B(n32584), .Y(n32543) );
  INVxp33_ASAP7_75t_SRAM U35840 ( .A(n32593), .Y(n32584) );
  INVxp33_ASAP7_75t_SRAM U35841 ( .A(n32565), .Y(n32561) );
  NOR2xp33_ASAP7_75t_SL U35842 ( .A(n32888), .B(n31639), .Y(n31494) );
  O2A1O1Ixp5_ASAP7_75t_SL U35843 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__3_), .B(n26826), .C(n26809), .Y(
        n3482) );
  O2A1O1Ixp5_ASAP7_75t_SL U35844 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__2_), .B(n26826), .C(n26825), .Y(
        n3499) );
  O2A1O1Ixp5_ASAP7_75t_SL U35845 ( .A1(n23229), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__1_), .B(n26826), .C(n26822), .Y(
        n3756) );
  O2A1O1Ixp5_ASAP7_75t_SL U35846 ( .A1(n28041), .A2(n28040), .B(n28039), .C(
        n24695), .Y(n17444) );
  NOR2xp33_ASAP7_75t_SL U35847 ( .A(n31716), .B(n31727), .Y(n31726) );
  NOR2xp33_ASAP7_75t_SL U35848 ( .A(n31716), .B(n31728), .Y(n31725) );
  NOR2xp33_ASAP7_75t_SL U35849 ( .A(ahb0_r_HADDR__2_), .B(ahb0_r_HADDR__3_), 
        .Y(n25239) );
  NOR2xp33_ASAP7_75t_SL U35850 ( .A(n29945), .B(n28037), .Y(n28033) );
  INVx1_ASAP7_75t_SL U35851 ( .A(n24681), .Y(n24652) );
  INVx1_ASAP7_75t_SL U35852 ( .A(n24681), .Y(n24657) );
  INVx1_ASAP7_75t_SL U35853 ( .A(n24681), .Y(n24656) );
  INVx1_ASAP7_75t_SL U35854 ( .A(n24681), .Y(n24655) );
  INVx1_ASAP7_75t_SL U35855 ( .A(n24681), .Y(n24650) );
  INVx1_ASAP7_75t_SL U35856 ( .A(n24681), .Y(n24653) );
  INVx1_ASAP7_75t_SL U35857 ( .A(n24681), .Y(n24651) );
  INVx1_ASAP7_75t_SL U35858 ( .A(n24681), .Y(n24654) );
  INVx1_ASAP7_75t_SL U35859 ( .A(n32162), .Y(n24641) );
  O2A1O1Ixp5_ASAP7_75t_SL U35860 ( .A1(n30955), .A2(n25703), .B(n24925), .C(
        n25652), .Y(n24995) );
  AOI21xp33_ASAP7_75t_SRAM U35861 ( .A1(n31951), .A2(uart1_r_RCNT__5_), .B(
        n31950), .Y(n31952) );
  OAI21xp33_ASAP7_75t_SRAM U35862 ( .A1(n29451), .A2(n29450), .B(n29449), .Y(
        n29455) );
  AOI21xp33_ASAP7_75t_SRAM U35863 ( .A1(n29448), .A2(n29447), .B(n29446), .Y(
        n29449) );
  INVxp33_ASAP7_75t_SRAM U35864 ( .A(n29445), .Y(n29446) );
  NOR2xp33_ASAP7_75t_SL U35865 ( .A(n24695), .B(n24633), .Y(n28059) );
  INVx1_ASAP7_75t_SL U35866 ( .A(n30548), .Y(n24633) );
  NOR2xp33_ASAP7_75t_SL U35867 ( .A(n24695), .B(n30548), .Y(n28060) );
  INVxp33_ASAP7_75t_SRAM U35868 ( .A(n3704), .Y(n32072) );
  XNOR2xp5_ASAP7_75t_SL U35869 ( .A(n25990), .B(n27496), .Y(n25991) );
  NOR2xp33_ASAP7_75t_SL U35870 ( .A(u0_0_leon3x0_p0_iu_r_A__WOVF_), .B(n29223), 
        .Y(n29667) );
  O2A1O1Ixp5_ASAP7_75t_SL U35871 ( .A1(sr1_r_MCFG1__ROMWWS__0_), .A2(n24695), 
        .B(n30779), .C(n30778), .Y(n2905) );
  O2A1O1Ixp5_ASAP7_75t_SL U35872 ( .A1(sr1_r_MCFG1__ROMWWS__1_), .A2(n24695), 
        .B(n30779), .C(n30072), .Y(n2904) );
  O2A1O1Ixp5_ASAP7_75t_SL U35873 ( .A1(n24542), .A2(n32075), .B(n25710), .C(
        n32076), .Y(n3389) );
  O2A1O1Ixp5_ASAP7_75t_SL U35874 ( .A1(n30780), .A2(n31190), .B(n30775), .C(
        n31188), .Y(n30776) );
  NOR2xp33_ASAP7_75t_SL U35875 ( .A(n32888), .B(n32904), .Y(n32903) );
  NOR2xp33_ASAP7_75t_SL U35876 ( .A(n32913), .B(n32912), .Y(n32973) );
  NOR2xp33_ASAP7_75t_SL U35877 ( .A(n32888), .B(n32860), .Y(n32871) );
  NOR2xp33_ASAP7_75t_SL U35878 ( .A(n32837), .B(n32836), .Y(n32860) );
  NOR2xp33_ASAP7_75t_SL U35879 ( .A(n2357), .B(n32833), .Y(n32886) );
  NOR2xp33_ASAP7_75t_SL U35880 ( .A(n3897), .B(
        u0_0_leon3x0_p0_c0mmu_a0_r_BO__0_), .Y(n25597) );
  INVxp33_ASAP7_75t_SRAM U35881 ( .A(n27373), .Y(n27305) );
  O2A1O1Ixp5_ASAP7_75t_SL U35882 ( .A1(n30073), .A2(n31190), .B(n30067), .C(
        n30071), .Y(n30069) );
  O2A1O1Ixp5_ASAP7_75t_SL U35883 ( .A1(n29510), .A2(n31190), .B(n28233), .C(
        n31188), .Y(n28234) );
  O2A1O1Ixp5_ASAP7_75t_SL U35884 ( .A1(n31197), .A2(n31190), .B(n31189), .C(
        n31188), .Y(n31191) );
  NOR2xp33_ASAP7_75t_SL U35885 ( .A(n26095), .B(n26094), .Y(n29959) );
  NOR2xp33_ASAP7_75t_SL U35886 ( .A(n26093), .B(n26092), .Y(n29955) );
  INVxp33_ASAP7_75t_SRAM U35887 ( .A(uart1_r_RXSTATE__0_), .Y(n26090) );
  NAND2xp33_ASAP7_75t_SRAM U35888 ( .A(n2867), .B(uart1_r_RXSTATE__1_), .Y(
        n29971) );
  NOR2xp33_ASAP7_75t_SL U35889 ( .A(n25556), .B(n25557), .Y(n26356) );
  NOR2xp33_ASAP7_75t_SL U35890 ( .A(n29670), .B(n31443), .Y(n29699) );
  O2A1O1Ixp5_ASAP7_75t_SL U35891 ( .A1(n25703), .A2(n25702), .B(n25701), .C(
        n30957), .Y(n25704) );
  INVxp33_ASAP7_75t_SRAM U35892 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__28_), 
        .Y(n25690) );
  INVxp33_ASAP7_75t_SRAM U35893 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__27_), 
        .Y(n25691) );
  AOI21xp33_ASAP7_75t_SRAM U35894 ( .A1(n25679), .A2(n25678), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .Y(n25685) );
  NAND2xp33_ASAP7_75t_SRAM U35895 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__8_), 
        .B(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__6_), .Y(n25677) );
  O2A1O1Ixp5_ASAP7_75t_SL U35896 ( .A1(n25671), .A2(n25670), .B(n25669), .C(
        n25668), .Y(n25672) );
  XNOR2xp5_ASAP7_75t_SL U35897 ( .A(n27411), .B(n27316), .Y(n27301) );
  NOR2xp33_ASAP7_75t_SL U35898 ( .A(u0_0_leon3x0_p0_iu_r_D__PV_), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__PV_), .Y(n25722) );
  NOR2xp33_ASAP7_75t_SL U35899 ( .A(n25851), .B(timer0_v_TICK_), .Y(n29521) );
  NOR2xp33_ASAP7_75t_SL U35900 ( .A(n4519), .B(n27540), .Y(n29951) );
  O2A1O1Ixp5_ASAP7_75t_SL U35901 ( .A1(n22421), .A2(
        u0_0_leon3x0_p0_iu_r_E__INVOP2_), .B(n25007), .C(n30651), .Y(n3316) );
  NOR2xp33_ASAP7_75t_SL U35902 ( .A(n24538), .B(n25559), .Y(n31987) );
  NOR2xp33_ASAP7_75t_SL U35903 ( .A(n2386), .B(n25996), .Y(n25997) );
  AOI21xp33_ASAP7_75t_SRAM U35904 ( .A1(n26001), .A2(n26023), .B(n26039), .Y(
        n25974) );
  NOR2xp33_ASAP7_75t_SL U35905 ( .A(n24695), .B(n28046), .Y(n27314) );
  NOR2xp33_ASAP7_75t_SL U35906 ( .A(n24695), .B(n27316), .Y(n27315) );
  O2A1O1Ixp5_ASAP7_75t_SL U35907 ( .A1(n29694), .A2(n29222), .B(n29221), .C(
        n29220), .Y(n3362) );
  AOI22xp33_ASAP7_75t_SRAM U35908 ( .A1(sr1_r_MCFG2__RAMRWS__0_), .A2(n31250), 
        .B1(n31235), .B2(sr1_r_MCFG1__ROMRWS__0_), .Y(n28086) );
  AOI22xp33_ASAP7_75t_SRAM U35909 ( .A1(uart1_uarto_RXEN_), .A2(n31950), .B1(
        n31245), .B2(timer0_r_SCALER__0_), .Y(n28087) );
  AOI22xp33_ASAP7_75t_SRAM U35910 ( .A1(uart1_r_RHOLD__13__0_), .A2(n31220), 
        .B1(n31221), .B2(uart1_r_RHOLD__31__0_), .Y(n28074) );
  AOI22xp33_ASAP7_75t_SRAM U35911 ( .A1(n31219), .A2(uart1_r_RHOLD__11__0_), 
        .B1(uart1_r_RHOLD__23__0_), .B2(n31218), .Y(n28075) );
  AOI22xp33_ASAP7_75t_SRAM U35912 ( .A1(n31217), .A2(uart1_r_RHOLD__29__0_), 
        .B1(uart1_r_RHOLD__3__0_), .B2(n31216), .Y(n28076) );
  AOI22xp33_ASAP7_75t_SRAM U35913 ( .A1(n31215), .A2(uart1_r_RHOLD__28__0_), 
        .B1(uart1_r_RHOLD__1__0_), .B2(n31214), .Y(n28077) );
  AOI22xp33_ASAP7_75t_SRAM U35914 ( .A1(n31229), .A2(uart1_r_RHOLD__22__0_), 
        .B1(uart1_r_RHOLD__27__0_), .B2(n31230), .Y(n28070) );
  AOI22xp33_ASAP7_75t_SRAM U35915 ( .A1(n31228), .A2(uart1_r_RHOLD__18__0_), 
        .B1(uart1_r_RHOLD__8__0_), .B2(n31227), .Y(n28071) );
  AOI22xp33_ASAP7_75t_SRAM U35916 ( .A1(uart1_r_RHOLD__10__0_), .A2(n31225), 
        .B1(n31226), .B2(uart1_r_RHOLD__6__0_), .Y(n28072) );
  AOI22xp33_ASAP7_75t_SRAM U35917 ( .A1(uart1_r_RHOLD__2__0_), .A2(n31223), 
        .B1(n31224), .B2(uart1_r_RHOLD__4__0_), .Y(n28073) );
  AOI22xp33_ASAP7_75t_SRAM U35918 ( .A1(uart1_r_RHOLD__26__0_), .A2(n31212), 
        .B1(uart1_r_RHOLD__15__0_), .B2(n31213), .Y(n28064) );
  AOI22xp33_ASAP7_75t_SRAM U35919 ( .A1(n31211), .A2(uart1_r_RHOLD__20__0_), 
        .B1(uart1_r_RHOLD__21__0_), .B2(n31210), .Y(n28065) );
  AOI22xp33_ASAP7_75t_SRAM U35920 ( .A1(n31209), .A2(uart1_r_RHOLD__25__0_), 
        .B1(uart1_r_RHOLD__19__0_), .B2(n31208), .Y(n28066) );
  AOI22xp33_ASAP7_75t_SRAM U35921 ( .A1(uart1_r_RHOLD__17__0_), .A2(n31206), 
        .B1(n31207), .B2(uart1_r_RHOLD__7__0_), .Y(n28067) );
  AOI22xp33_ASAP7_75t_SRAM U35922 ( .A1(n31205), .A2(uart1_r_RHOLD__16__0_), 
        .B1(uart1_r_RHOLD__9__0_), .B2(n31204), .Y(n28061) );
  AOI22xp33_ASAP7_75t_SRAM U35923 ( .A1(uart1_r_RHOLD__12__0_), .A2(n31202), 
        .B1(n31203), .B2(uart1_r_RHOLD__14__0_), .Y(n28062) );
  AOI22xp33_ASAP7_75t_SRAM U35924 ( .A1(n31201), .A2(uart1_r_RHOLD__30__0_), 
        .B1(uart1_r_RHOLD__5__0_), .B2(n31200), .Y(n28063) );
  AOI22xp33_ASAP7_75t_SRAM U35925 ( .A1(uart1_r_THOLD__3__0_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__7__0_), .Y(n28004) );
  AOI22xp33_ASAP7_75t_SRAM U35926 ( .A1(uart1_r_THOLD__23__0_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__11__0_), .Y(n28005) );
  AOI22xp33_ASAP7_75t_SRAM U35927 ( .A1(uart1_r_THOLD__19__0_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__27__0_), .Y(n28006) );
  AOI22xp33_ASAP7_75t_SRAM U35928 ( .A1(n27997), .A2(uart1_r_THOLD__15__0_), 
        .B1(uart1_r_THOLD__31__0_), .B2(n27996), .Y(n28007) );
  INVxp33_ASAP7_75t_SRAM U35929 ( .A(uart1_r_THOLD__17__0_), .Y(n27984) );
  AOI22xp33_ASAP7_75t_SRAM U35930 ( .A1(uart1_r_THOLD__1__0_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__5__0_), .Y(n27981) );
  AO21x1_ASAP7_75t_SL U35931 ( .A1(n26097), .A2(n31249), .B(n24695), .Y(n29385) );
  AOI22xp33_ASAP7_75t_SRAM U35932 ( .A1(uart1_r_RHOLD__6__6_), .A2(n31226), 
        .B1(n31225), .B2(uart1_r_RHOLD__10__6_), .Y(n31233) );
  AOI22xp33_ASAP7_75t_SRAM U35933 ( .A1(uart1_r_RHOLD__4__6_), .A2(n31224), 
        .B1(n31223), .B2(uart1_r_RHOLD__2__6_), .Y(n31234) );
  AOI22xp33_ASAP7_75t_SRAM U35934 ( .A1(uart1_r_RHOLD__31__6_), .A2(n31221), 
        .B1(n31220), .B2(uart1_r_RHOLD__13__6_), .Y(n31222) );
  AOI22xp33_ASAP7_75t_SRAM U35935 ( .A1(uart1_r_THOLD__3__6_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__7__6_), .Y(n27636) );
  AOI22xp33_ASAP7_75t_SRAM U35936 ( .A1(uart1_r_THOLD__19__6_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__27__6_), .Y(n27638) );
  AOI22xp33_ASAP7_75t_SRAM U35937 ( .A1(n27997), .A2(uart1_r_THOLD__15__6_), 
        .B1(uart1_r_THOLD__31__6_), .B2(n27996), .Y(n27639) );
  INVxp33_ASAP7_75t_SRAM U35938 ( .A(uart1_r_THOLD__17__6_), .Y(n27626) );
  AOI22xp33_ASAP7_75t_SRAM U35939 ( .A1(uart1_r_THOLD__1__6_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__5__6_), .Y(n27623) );
  AOI22xp33_ASAP7_75t_SRAM U35940 ( .A1(n31219), .A2(uart1_r_RHOLD__11__3_), 
        .B1(uart1_r_RHOLD__23__3_), .B2(n31218), .Y(n28250) );
  AOI22xp33_ASAP7_75t_SRAM U35941 ( .A1(n31217), .A2(uart1_r_RHOLD__29__3_), 
        .B1(uart1_r_RHOLD__3__3_), .B2(n31216), .Y(n28251) );
  AOI22xp33_ASAP7_75t_SRAM U35942 ( .A1(n31215), .A2(uart1_r_RHOLD__28__3_), 
        .B1(uart1_r_RHOLD__1__3_), .B2(n31214), .Y(n28252) );
  INVxp33_ASAP7_75t_SRAM U35943 ( .A(uart1_r_THOLD__12__3_), .Y(n27840) );
  NAND2xp33_ASAP7_75t_SRAM U35944 ( .A(uart1_r_TRADDR__0_), .B(n27838), .Y(
        n27846) );
  AOI22xp33_ASAP7_75t_SRAM U35945 ( .A1(uart1_r_THOLD__1__3_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__5__3_), .Y(n27834) );
  AOI22xp33_ASAP7_75t_SRAM U35946 ( .A1(uart1_r_THOLD__21__3_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__9__3_), .Y(n27835) );
  AOI22xp33_ASAP7_75t_SRAM U35947 ( .A1(n27997), .A2(uart1_r_THOLD__13__3_), 
        .B1(uart1_r_THOLD__29__3_), .B2(n27996), .Y(n27836) );
  AOI22xp33_ASAP7_75t_SRAM U35948 ( .A1(uart1_r_THOLD__17__3_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__25__3_), .Y(n27837) );
  O2A1O1Ixp5_ASAP7_75t_SL U35949 ( .A1(apbi[27]), .A2(n27292), .B(n27293), .C(
        n28116), .Y(n25959) );
  AOI22xp33_ASAP7_75t_SRAM U35950 ( .A1(uart1_r_RHOLD__13__4_), .A2(n31220), 
        .B1(n31221), .B2(uart1_r_RHOLD__31__4_), .Y(n30785) );
  AOI22xp33_ASAP7_75t_SRAM U35951 ( .A1(n31219), .A2(uart1_r_RHOLD__11__4_), 
        .B1(uart1_r_RHOLD__23__4_), .B2(n31218), .Y(n30786) );
  AOI22xp33_ASAP7_75t_SRAM U35952 ( .A1(n31217), .A2(uart1_r_RHOLD__29__4_), 
        .B1(uart1_r_RHOLD__3__4_), .B2(n31216), .Y(n30787) );
  AOI22xp33_ASAP7_75t_SRAM U35953 ( .A1(n31215), .A2(uart1_r_RHOLD__28__4_), 
        .B1(uart1_r_RHOLD__1__4_), .B2(n31214), .Y(n30788) );
  AOI22xp33_ASAP7_75t_SRAM U35954 ( .A1(n31228), .A2(uart1_r_RHOLD__18__4_), 
        .B1(uart1_r_RHOLD__8__4_), .B2(n31227), .Y(n30784) );
  AOI22xp33_ASAP7_75t_SRAM U35955 ( .A1(uart1_r_THOLD__3__4_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__7__4_), .Y(n27772) );
  INVxp33_ASAP7_75t_SRAM U35956 ( .A(uart1_r_THOLD__27__4_), .Y(n27770) );
  AOI22xp33_ASAP7_75t_SRAM U35957 ( .A1(uart1_r_THOLD__1__4_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__5__4_), .Y(n27757) );
  INVxp33_ASAP7_75t_SRAM U35958 ( .A(uart1_r_THOLD__25__4_), .Y(n27756) );
  NOR3xp33_ASAP7_75t_SL U35959 ( .A(n24596), .B(uart1_uarto_SCALER__8_), .C(
        uart1_uarto_SCALER__7_), .Y(n24587) );
  NOR3xp33_ASAP7_75t_SL U35960 ( .A(n24593), .B(uart1_uarto_SCALER__5_), .C(
        uart1_uarto_SCALER__4_), .Y(n24594) );
  NOR3xp33_ASAP7_75t_SL U35961 ( .A(uart1_uarto_SCALER__1_), .B(
        uart1_uarto_SCALER__2_), .C(uart1_uarto_SCALER__0_), .Y(n24591) );
  NOR2xp33_ASAP7_75t_SL U35962 ( .A(n27329), .B(n27328), .Y(n27376) );
  O2A1O1Ixp5_ASAP7_75t_SL U35963 ( .A1(n29117), .A2(n29116), .B(
        u0_0_leon3x0_p0_divo[32]), .C(n31672), .Y(n2306) );
  XNOR2xp5_ASAP7_75t_SL U35964 ( .A(u0_0_leon3x0_p0_div0_r_QMSB_), .B(n29114), 
        .Y(n29115) );
  AOI22xp33_ASAP7_75t_SRAM U35965 ( .A1(uart1_r_RHOLD__26__1_), .A2(n31212), 
        .B1(uart1_r_RHOLD__15__1_), .B2(n31213), .Y(n27429) );
  AOI22xp33_ASAP7_75t_SRAM U35966 ( .A1(n31211), .A2(uart1_r_RHOLD__20__1_), 
        .B1(uart1_r_RHOLD__21__1_), .B2(n31210), .Y(n27430) );
  AOI22xp33_ASAP7_75t_SRAM U35967 ( .A1(n31209), .A2(uart1_r_RHOLD__25__1_), 
        .B1(uart1_r_RHOLD__19__1_), .B2(n31208), .Y(n27431) );
  AOI22xp33_ASAP7_75t_SRAM U35968 ( .A1(uart1_r_RHOLD__7__1_), .A2(n31207), 
        .B1(n31206), .B2(uart1_r_RHOLD__17__1_), .Y(n27432) );
  AOI22xp33_ASAP7_75t_SRAM U35969 ( .A1(uart1_r_THOLD__1__1_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__5__1_), .Y(n27401) );
  AOI22xp33_ASAP7_75t_SRAM U35970 ( .A1(n28000), .A2(uart1_r_THOLD__9__1_), 
        .B1(uart1_r_THOLD__21__1_), .B2(n28001), .Y(n27402) );
  AOI22xp33_ASAP7_75t_SRAM U35971 ( .A1(uart1_r_THOLD__17__1_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__25__1_), .Y(n27403) );
  AOI22xp33_ASAP7_75t_SRAM U35972 ( .A1(n27997), .A2(uart1_r_THOLD__13__1_), 
        .B1(uart1_r_THOLD__29__1_), .B2(n27996), .Y(n27404) );
  XNOR2xp5_ASAP7_75t_SL U35973 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(
        n29206), .Y(n25003) );
  O2A1O1Ixp5_ASAP7_75t_SL U35974 ( .A1(apbi[18]), .A2(n29652), .B(n29651), .C(
        n29568), .Y(n29331) );
  NOR2xp33_ASAP7_75t_SL U35975 ( .A(n29329), .B(n29294), .Y(n28243) );
  O2A1O1Ixp5_ASAP7_75t_SL U35976 ( .A1(apbi[19]), .A2(n29652), .B(n29651), .C(
        n29510), .Y(n28239) );
  O2A1O1Ixp5_ASAP7_75t_SL U35977 ( .A1(apbi[20]), .A2(n29652), .B(n29651), .C(
        n30780), .Y(n29318) );
  NOR2xp33_ASAP7_75t_SL U35978 ( .A(n29316), .B(n29294), .Y(n29300) );
  O2A1O1Ixp5_ASAP7_75t_SL U35979 ( .A1(apbi[21]), .A2(n29652), .B(n29651), .C(
        n30073), .Y(n29296) );
  O2A1O1Ixp5_ASAP7_75t_SL U35980 ( .A1(apbi[23]), .A2(n29652), .B(n29651), .C(
        n30833), .Y(n29280) );
  O2A1O1Ixp5_ASAP7_75t_SL U35981 ( .A1(apbi[17]), .A2(n29652), .B(n29651), .C(
        n27493), .Y(n27295) );
  NOR2xp33_ASAP7_75t_SL U35982 ( .A(n29316), .B(n29237), .Y(n29238) );
  O2A1O1Ixp5_ASAP7_75t_SL U35983 ( .A1(apbi[31]), .A2(n29652), .B(n29651), .C(
        n29389), .Y(n29392) );
  AOI22xp33_ASAP7_75t_SRAM U35984 ( .A1(uart1_r_THOLD__1__2_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__5__2_), .Y(n27896) );
  AOI22xp33_ASAP7_75t_SRAM U35985 ( .A1(uart1_r_THOLD__21__2_), .A2(n28001), 
        .B1(n28000), .B2(uart1_r_THOLD__9__2_), .Y(n27897) );
  AOI22xp33_ASAP7_75t_SRAM U35986 ( .A1(n27997), .A2(uart1_r_THOLD__13__2_), 
        .B1(uart1_r_THOLD__29__2_), .B2(n27996), .Y(n27898) );
  AOI22xp33_ASAP7_75t_SRAM U35987 ( .A1(uart1_r_THOLD__17__2_), .A2(n27999), 
        .B1(n27998), .B2(uart1_r_THOLD__25__2_), .Y(n27899) );
  NOR2xp33_ASAP7_75t_SL U35988 ( .A(n29316), .B(n29653), .Y(n29245) );
  O2A1O1Ixp5_ASAP7_75t_SL U35989 ( .A1(apbi[28]), .A2(n29652), .B(n29651), .C(
        n29851), .Y(n29241) );
  NOR2xp33_ASAP7_75t_SL U35990 ( .A(n29329), .B(n29653), .Y(n29267) );
  O2A1O1Ixp5_ASAP7_75t_SL U35991 ( .A1(apbi[26]), .A2(n29652), .B(n29651), .C(
        n30978), .Y(n29263) );
  O2A1O1Ixp5_ASAP7_75t_SL U35992 ( .A1(apbi[25]), .A2(n29652), .B(n29651), .C(
        n30139), .Y(n29252) );
  NOR2xp33_ASAP7_75t_SL U35993 ( .A(n3325), .B(n29646), .Y(n29391) );
  NOR2xp33_ASAP7_75t_SL U35994 ( .A(n27470), .B(n27472), .Y(n31242) );
  AOI22xp33_ASAP7_75t_SRAM U35995 ( .A1(uart1_r_RHOLD__31__5_), .A2(n31221), 
        .B1(n31220), .B2(uart1_r_RHOLD__13__5_), .Y(n30094) );
  AOI22xp33_ASAP7_75t_SRAM U35996 ( .A1(n31219), .A2(uart1_r_RHOLD__11__5_), 
        .B1(uart1_r_RHOLD__23__5_), .B2(n31218), .Y(n30095) );
  AOI22xp33_ASAP7_75t_SRAM U35997 ( .A1(n31217), .A2(uart1_r_RHOLD__29__5_), 
        .B1(uart1_r_RHOLD__3__5_), .B2(n31216), .Y(n30096) );
  AOI22xp33_ASAP7_75t_SRAM U35998 ( .A1(n31215), .A2(uart1_r_RHOLD__28__5_), 
        .B1(uart1_r_RHOLD__1__5_), .B2(n31214), .Y(n30097) );
  AOI22xp33_ASAP7_75t_SRAM U35999 ( .A1(uart1_r_RHOLD__22__5_), .A2(n31229), 
        .B1(uart1_r_RHOLD__27__5_), .B2(n31230), .Y(n30090) );
  AOI22xp33_ASAP7_75t_SRAM U36000 ( .A1(n31228), .A2(uart1_r_RHOLD__18__5_), 
        .B1(uart1_r_RHOLD__8__5_), .B2(n31227), .Y(n30091) );
  AOI22xp33_ASAP7_75t_SRAM U36001 ( .A1(uart1_r_RHOLD__6__5_), .A2(n31226), 
        .B1(n31225), .B2(uart1_r_RHOLD__10__5_), .Y(n30092) );
  AOI22xp33_ASAP7_75t_SRAM U36002 ( .A1(uart1_r_RHOLD__4__5_), .A2(n31224), 
        .B1(n31223), .B2(uart1_r_RHOLD__2__5_), .Y(n30093) );
  AOI22xp33_ASAP7_75t_SRAM U36003 ( .A1(uart1_r_RHOLD__26__5_), .A2(n31212), 
        .B1(n31213), .B2(uart1_r_RHOLD__15__5_), .Y(n30084) );
  AOI22xp33_ASAP7_75t_SRAM U36004 ( .A1(n31211), .A2(uart1_r_RHOLD__20__5_), 
        .B1(uart1_r_RHOLD__21__5_), .B2(n31210), .Y(n30085) );
  AOI22xp33_ASAP7_75t_SRAM U36005 ( .A1(n31209), .A2(uart1_r_RHOLD__25__5_), 
        .B1(uart1_r_RHOLD__19__5_), .B2(n31208), .Y(n30086) );
  AOI22xp33_ASAP7_75t_SRAM U36006 ( .A1(uart1_r_RHOLD__7__5_), .A2(n31207), 
        .B1(n31206), .B2(uart1_r_RHOLD__17__5_), .Y(n30087) );
  AOI22xp33_ASAP7_75t_SRAM U36007 ( .A1(n31205), .A2(uart1_r_RHOLD__16__5_), 
        .B1(uart1_r_RHOLD__9__5_), .B2(n31204), .Y(n30081) );
  AOI22xp33_ASAP7_75t_SRAM U36008 ( .A1(uart1_r_RHOLD__14__5_), .A2(n31203), 
        .B1(n31202), .B2(uart1_r_RHOLD__12__5_), .Y(n30082) );
  AOI22xp33_ASAP7_75t_SRAM U36009 ( .A1(n31201), .A2(uart1_r_RHOLD__30__5_), 
        .B1(uart1_r_RHOLD__5__5_), .B2(n31200), .Y(n30083) );
  NOR2xp33_ASAP7_75t_SL U36010 ( .A(n2992), .B(n25951), .Y(n27290) );
  NOR2xp33_ASAP7_75t_SL U36011 ( .A(n28085), .B(n27464), .Y(n31237) );
  NOR2xp33_ASAP7_75t_SL U36012 ( .A(n2931), .B(n27460), .Y(n31252) );
  INVx1_ASAP7_75t_SL U36013 ( .A(n2931), .Y(n26501) );
  NOR2xp33_ASAP7_75t_SL U36014 ( .A(n26071), .B(n25636), .Y(n31248) );
  AND2x2_ASAP7_75t_SL U36015 ( .A(n2992), .B(n4371), .Y(n25961) );
  INVxp33_ASAP7_75t_SRAM U36016 ( .A(uart1_r_THOLD__14__5_), .Y(n27704) );
  AOI22xp33_ASAP7_75t_SRAM U36017 ( .A1(uart1_r_THOLD__3__5_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__7__5_), .Y(n27698) );
  NOR2xp33_ASAP7_75t_SL U36018 ( .A(uart1_r_TRADDR__0_), .B(n27410), .Y(n28015) );
  NOR2xp33_ASAP7_75t_SL U36019 ( .A(uart1_r_TRADDR__0_), .B(n27409), .Y(n28008) );
  NOR2xp33_ASAP7_75t_SL U36020 ( .A(uart1_r_TRADDR__0_), .B(n27408), .Y(n28009) );
  NOR2xp33_ASAP7_75t_SL U36021 ( .A(uart1_r_TRADDR__0_), .B(n27985), .Y(n28010) );
  NOR2xp33_ASAP7_75t_SL U36022 ( .A(uart1_r_TRADDR__0_), .B(n27407), .Y(n28011) );
  NOR2xp33_ASAP7_75t_SL U36023 ( .A(uart1_r_TRADDR__0_), .B(n27405), .Y(n28018) );
  NOR2xp33_ASAP7_75t_SL U36024 ( .A(uart1_r_TRADDR__0_), .B(n27771), .Y(n28017) );
  AOI22xp33_ASAP7_75t_SRAM U36025 ( .A1(uart1_r_THOLD__1__5_), .A2(n28003), 
        .B1(n28002), .B2(uart1_r_THOLD__5__5_), .Y(n27690) );
  NOR2xp33_ASAP7_75t_SL U36026 ( .A(uart1_r_TRADDR__4_), .B(uart1_r_TRADDR__3_), .Y(n27395) );
  AOI22xp33_ASAP7_75t_SRAM U36027 ( .A1(n27997), .A2(uart1_r_THOLD__13__5_), 
        .B1(uart1_r_THOLD__29__5_), .B2(n27996), .Y(n27692) );
  NOR2xp33_ASAP7_75t_SL U36028 ( .A(uart1_r_TRADDR__2_), .B(n27391), .Y(n27392) );
  NOR2xp33_ASAP7_75t_SL U36029 ( .A(n25999), .B(n26014), .Y(n26043) );
  NOR2xp33_ASAP7_75t_SL U36030 ( .A(n25981), .B(n26014), .Y(n26053) );
  NOR2xp33_ASAP7_75t_SL U36031 ( .A(n26006), .B(n26014), .Y(n26066) );
  NOR2xp33_ASAP7_75t_SL U36032 ( .A(n26016), .B(n26014), .Y(n26060) );
  INVx1_ASAP7_75t_SL U36033 ( .A(n24681), .Y(n24660) );
  O2A1O1Ixp5_ASAP7_75t_SL U36034 ( .A1(n29206), .A2(n29205), .B(n23229), .C(
        n29204), .Y(n31439) );
  O2A1O1Ixp5_ASAP7_75t_SL U36035 ( .A1(n29203), .A2(n29202), .B(n29201), .C(
        n29200), .Y(n29204) );
  O2A1O1Ixp5_ASAP7_75t_SL U36036 ( .A1(u0_0_leon3x0_p0_iu_r_X__RESULT__2_), 
        .A2(n29198), .B(n29197), .C(n24659), .Y(n30472) );
  O2A1O1Ixp5_ASAP7_75t_SL U36037 ( .A1(n29189), .A2(n29202), .B(n29188), .C(
        n29187), .Y(n29205) );
  NOR2xp33_ASAP7_75t_SL U36038 ( .A(n27338), .B(n27383), .Y(n27947) );
  NOR2xp33_ASAP7_75t_SL U36039 ( .A(n27388), .B(n27383), .Y(n27975) );
  NOR2xp33_ASAP7_75t_SL U36040 ( .A(n27364), .B(n27383), .Y(n27950) );
  NOR2xp33_ASAP7_75t_SL U36041 ( .A(n27351), .B(n27383), .Y(n27920) );
  NOR2xp33_ASAP7_75t_SL U36042 ( .A(n27369), .B(n27383), .Y(n27962) );
  NOR2xp33_ASAP7_75t_SL U36043 ( .A(n27385), .B(n27383), .Y(n27967) );
  NOR2xp33_ASAP7_75t_SL U36044 ( .A(n27333), .B(n27383), .Y(n27935) );
  NOR2xp33_ASAP7_75t_SL U36045 ( .A(n27353), .B(n27383), .Y(n27928) );
  NAND2xp5_ASAP7_75t_SL U36046 ( .A(n27322), .B(n27325), .Y(n27383) );
  NOR2xp33_ASAP7_75t_SL U36047 ( .A(n27364), .B(n27381), .Y(n27952) );
  NOR2xp33_ASAP7_75t_SL U36048 ( .A(n27385), .B(n27381), .Y(n27968) );
  NOR2xp33_ASAP7_75t_SL U36049 ( .A(n27338), .B(n27381), .Y(n27946) );
  NOR2xp33_ASAP7_75t_SL U36050 ( .A(n27353), .B(n27381), .Y(n27926) );
  NOR2xp33_ASAP7_75t_SL U36051 ( .A(n27369), .B(n27381), .Y(n27960) );
  NOR2xp33_ASAP7_75t_SL U36052 ( .A(n27388), .B(n27381), .Y(n27973) );
  NOR2xp33_ASAP7_75t_SL U36053 ( .A(n27351), .B(n27381), .Y(n27922) );
  NOR2xp33_ASAP7_75t_SL U36054 ( .A(n27333), .B(n27381), .Y(n27939) );
  NOR2xp33_ASAP7_75t_SL U36055 ( .A(n27338), .B(n27387), .Y(n27933) );
  NOR2xp33_ASAP7_75t_SL U36056 ( .A(n27351), .B(n27387), .Y(n27929) );
  NOR2xp33_ASAP7_75t_SL U36057 ( .A(n27369), .B(n27387), .Y(n27948) );
  NOR2xp33_ASAP7_75t_SL U36058 ( .A(n27385), .B(n27387), .Y(n27977) );
  NOR2xp33_ASAP7_75t_SL U36059 ( .A(n27333), .B(n27387), .Y(n27937) );
  NOR2xp33_ASAP7_75t_SL U36060 ( .A(n27364), .B(n27387), .Y(n27951) );
  NOR2xp33_ASAP7_75t_SL U36061 ( .A(n27353), .B(n27387), .Y(n27931) );
  NOR2xp33_ASAP7_75t_SL U36062 ( .A(n27388), .B(n27387), .Y(n27979) );
  NAND2xp5_ASAP7_75t_SL U36063 ( .A(n27310), .B(n27309), .Y(n27387) );
  XNOR2xp5_ASAP7_75t_SL U36064 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__7_), .B(
        n32186), .Y(n30928) );
  XNOR2xp5_ASAP7_75t_SL U36065 ( .A(n30927), .B(n30939), .Y(n30929) );
  XNOR2xp5_ASAP7_75t_SL U36066 ( .A(n30923), .B(n32179), .Y(n30924) );
  XNOR2xp5_ASAP7_75t_SL U36067 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__2_), .B(
        n32178), .Y(n30922) );
  XNOR2xp5_ASAP7_75t_SL U36068 ( .A(n30920), .B(n32183), .Y(n30931) );
  NOR2xp33_ASAP7_75t_SL U36069 ( .A(n24695), .B(n26014), .Y(n29985) );
  NOR2xp33_ASAP7_75t_SL U36070 ( .A(n24695), .B(n26015), .Y(n29987) );
  AOI31xp33_ASAP7_75t_SL U36071 ( .A1(n31194), .A2(n25972), .A3(n30066), .B(
        n27538), .Y(n26015) );
  NOR2xp33_ASAP7_75t_SL U36072 ( .A(n25971), .B(n28189), .Y(n27538) );
  NOR2xp33_ASAP7_75t_SL U36073 ( .A(n29960), .B(n27535), .Y(n31194) );
  NOR2xp33_ASAP7_75t_SL U36074 ( .A(n27522), .B(n27520), .Y(n29977) );
  NOR2xp33_ASAP7_75t_SL U36075 ( .A(n27523), .B(n29980), .Y(n27520) );
  NOR2xp33_ASAP7_75t_SL U36076 ( .A(n29982), .B(n29981), .Y(n29980) );
  NOR2xp33_ASAP7_75t_SL U36077 ( .A(n27519), .B(n27518), .Y(n27522) );
  NOR2xp33_ASAP7_75t_SL U36078 ( .A(n27500), .B(n27501), .Y(n27517) );
  NOR2xp33_ASAP7_75t_SL U36079 ( .A(n29982), .B(n29975), .Y(n29979) );
  NOR2xp33_ASAP7_75t_SL U36080 ( .A(n27507), .B(n27502), .Y(n27513) );
  NOR2xp33_ASAP7_75t_SL U36081 ( .A(n27498), .B(n27497), .Y(n27502) );
  NAND2xp33_ASAP7_75t_SRAM U36082 ( .A(n27495), .B(n31057), .Y(n27498) );
  NOR2xp33_ASAP7_75t_SL U36083 ( .A(n27495), .B(n31057), .Y(n27507) );
  NOR2xp33_ASAP7_75t_SL U36084 ( .A(n25536), .B(n27328), .Y(n28231) );
  NOR2xp33_ASAP7_75t_SL U36085 ( .A(uart1_r_RCNT__1_), .B(n27506), .Y(n27503)
         );
  NOR2xp33_ASAP7_75t_SL U36086 ( .A(n28050), .B(n28049), .Y(n28055) );
  NOR2xp33_ASAP7_75t_SL U36087 ( .A(n29374), .B(n28042), .Y(n28043) );
  NOR2xp33_ASAP7_75t_SL U36088 ( .A(n26081), .B(n28044), .Y(n29374) );
  NOR2xp33_ASAP7_75t_SL U36089 ( .A(n31851), .B(n26079), .Y(n26081) );
  XNOR2xp5_ASAP7_75t_SL U36090 ( .A(n31645), .B(n28044), .Y(n29351) );
  NOR2xp33_ASAP7_75t_SL U36091 ( .A(uart1_r_TCNT__1_), .B(n26080), .Y(n28044)
         );
  NAND2xp5_ASAP7_75t_SL U36092 ( .A(n27540), .B(n28036), .Y(n29949) );
  NOR2xp33_ASAP7_75t_SL U36093 ( .A(n26078), .B(n26077), .Y(n28036) );
  NAND4xp25_ASAP7_75t_SL U36094 ( .A(n29354), .B(uart1_uarto_TXEN_), .C(n4520), 
        .D(n28032), .Y(n26077) );
  NOR2xp33_ASAP7_75t_SL U36095 ( .A(n26076), .B(n28096), .Y(n26078) );
  NOR2xp33_ASAP7_75t_SL U36096 ( .A(n29746), .B(n27510), .Y(n28096) );
  NOR2xp33_ASAP7_75t_SL U36097 ( .A(uart1_r_TCNT__5_), .B(uart1_r_TCNT__4_), 
        .Y(n30873) );
  NAND2xp33_ASAP7_75t_SRAM U36098 ( .A(n33068), .B(n26072), .Y(n26073) );
  NOR4xp25_ASAP7_75t_SL U36099 ( .A(uart1_r_TCNT__1_), .B(uart1_r_TCNT__0_), 
        .C(uart1_r_TCNT__2_), .D(uart1_r_TCNT__3_), .Y(n28045) );
  O2A1O1Ixp5_ASAP7_75t_SL U36100 ( .A1(n29921), .A2(n30014), .B(n29920), .C(
        n30208), .Y(n29922) );
  NOR2xp33_ASAP7_75t_SL U36101 ( .A(n31015), .B(n31016), .Y(n28807) );
  AOI31xp33_ASAP7_75t_SL U36102 ( .A1(n29688), .A2(n31054), .A3(n29687), .B(
        n29501), .Y(n29502) );
  NOR2xp33_ASAP7_75t_SL U36103 ( .A(n31334), .B(n32110), .Y(n31346) );
  INVxp33_ASAP7_75t_SRAM U36104 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[9]), .Y(n31789) );
  AOI22xp33_ASAP7_75t_SRAM U36105 ( .A1(n28935), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__2_), .B1(u0_0_leon3x0_p0_divi[33]), 
        .B2(n30612), .Y(n28936) );
  NOR2xp33_ASAP7_75t_SL U36106 ( .A(n31340), .B(n30464), .Y(n31334) );
  O2A1O1Ixp5_ASAP7_75t_SL U36107 ( .A1(n29505), .A2(n24427), .B(n28895), .C(
        n29503), .Y(n28896) );
  INVxp33_ASAP7_75t_SRAM U36108 ( .A(u0_0_leon3x0_p0_divi[39]), .Y(n28730) );
  NOR2xp33_ASAP7_75t_SL U36109 ( .A(n28647), .B(n28646), .Y(n29845) );
  AO21x1_ASAP7_75t_SL U36110 ( .A1(n28902), .A2(u0_0_leon3x0_p0_dci[9]), .B(
        n28859), .Y(n29626) );
  NOR2xp33_ASAP7_75t_SL U36111 ( .A(n26252), .B(n26251), .Y(n28854) );
  AOI211xp5_ASAP7_75t_SL U36112 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__4_), 
        .A2(n24582), .B(n28887), .C(n28834), .Y(n28837) );
  NOR2xp33_ASAP7_75t_SL U36113 ( .A(n28833), .B(n29592), .Y(n28834) );
  NAND2xp33_ASAP7_75t_SRAM U36114 ( .A(n30614), .B(n30613), .Y(n30615) );
  AOI22xp33_ASAP7_75t_SRAM U36115 ( .A1(u0_0_leon3x0_p0_divi[32]), .A2(n30612), 
        .B1(u0_0_leon3x0_p0_iu_r_W__S__WIM__1_), .B2(n30611), .Y(n30617) );
  NOR2xp33_ASAP7_75t_SL U36116 ( .A(n22952), .B(n28970), .Y(n28852) );
  AOI22xp33_ASAP7_75t_SRAM U36117 ( .A1(n28835), .A2(n27147), .B1(
        u0_0_leon3x0_p0_divi[41]), .B2(n28782), .Y(n27151) );
  NOR2xp33_ASAP7_75t_SL U36118 ( .A(n31340), .B(n30385), .Y(n31048) );
  NOR2xp33_ASAP7_75t_SL U36119 ( .A(n27105), .B(n27104), .Y(n28666) );
  O2A1O1Ixp5_ASAP7_75t_SL U36120 ( .A1(n24491), .A2(n30703), .B(n30708), .C(
        n29726), .Y(n29886) );
  INVxp33_ASAP7_75t_SRAM U36121 ( .A(u0_0_leon3x0_p0_iu_r_M__NALIGN_), .Y(
        n29720) );
  OAI21xp33_ASAP7_75t_SRAM U36122 ( .A1(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__20_), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_), .B(n29471), .Y(n29473) );
  NOR2xp33_ASAP7_75t_SL U36123 ( .A(n22432), .B(n28802), .Y(n28542) );
  INVxp33_ASAP7_75t_SRAM U36124 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__7_), .Y(
        n25765) );
  NOR2xp33_ASAP7_75t_SL U36125 ( .A(n30812), .B(n30811), .Y(n32174) );
  NOR2xp33_ASAP7_75t_SL U36126 ( .A(n26849), .B(n26848), .Y(n28257) );
  NAND4xp25_ASAP7_75t_SL U36127 ( .A(n26862), .B(n26861), .C(n26860), .D(
        n26859), .Y(n26863) );
  XNOR2xp5_ASAP7_75t_SL U36128 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__2_), .B(
        DP_OP_1196_128_7433_n454), .Y(n26859) );
  XNOR2xp5_ASAP7_75t_SL U36129 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__1_), .B(
        DP_OP_1196_128_7433_n453), .Y(n26860) );
  NOR3xp33_ASAP7_75t_SL U36130 ( .A(n26858), .B(n26857), .C(n26856), .Y(n26861) );
  XNOR2xp5_ASAP7_75t_SL U36131 ( .A(n30923), .B(DP_OP_1196_128_7433_n455), .Y(
        n26857) );
  XNOR2xp5_ASAP7_75t_SL U36132 ( .A(n30927), .B(DP_OP_1196_128_7433_n452), .Y(
        n26858) );
  O2A1O1Ixp5_ASAP7_75t_SL U36133 ( .A1(n30595), .A2(n27016), .B(n27015), .C(
        n27014), .Y(n4049) );
  OAI21xp33_ASAP7_75t_SRAM U36134 ( .A1(n26169), .A2(n25820), .B(n25819), .Y(
        n25832) );
  OAI22xp33_ASAP7_75t_SRAM U36135 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__18_), 
        .A2(n27143), .B1(n25816), .B2(n27141), .Y(n25817) );
  OAI22xp33_ASAP7_75t_SRAM U36136 ( .A1(n26176), .A2(n30312), .B1(n25828), 
        .B2(n25812), .Y(n25833) );
  NOR2xp33_ASAP7_75t_SL U36137 ( .A(n27281), .B(n32110), .Y(n27283) );
  INVxp33_ASAP7_75t_SRAM U36138 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__5_), .Y(
        n26698) );
  O2A1O1Ixp5_ASAP7_75t_SL U36139 ( .A1(n27067), .A2(
        u0_0_leon3x0_p0_iu_r_E__JMPL_), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__15_), .C(n28887), .Y(n26571) );
  INVxp33_ASAP7_75t_SRAM U36140 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__3_), .Y(
        n26572) );
  NOR2xp33_ASAP7_75t_SL U36141 ( .A(n25811), .B(n25810), .Y(n26670) );
  AOI22xp33_ASAP7_75t_SRAM U36142 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__6_), 
        .A2(n31364), .B1(n30573), .B2(n31478), .Y(n30565) );
  AOI22xp33_ASAP7_75t_SRAM U36143 ( .A1(it_q[10]), .A2(n24636), .B1(n32625), 
        .B2(n30130), .Y(n25611) );
  AOI22xp33_ASAP7_75t_SRAM U36144 ( .A1(n30995), .A2(n33067), .B1(ic_q[14]), 
        .B2(n22387), .Y(n25612) );
  O2A1O1Ixp5_ASAP7_75t_SL U36145 ( .A1(u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_), 
        .A2(u0_0_leon3x0_p0_dci[6]), .B(n28993), .C(
        u0_0_leon3x0_p0_iu_r_E__ALUSEL__1_), .Y(n29006) );
  NOR2xp33_ASAP7_75t_SL U36146 ( .A(n28919), .B(n28918), .Y(n30627) );
  AOI22xp33_ASAP7_75t_SRAM U36147 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__0_), 
        .A2(n31364), .B1(n30479), .B2(n31478), .Y(n30480) );
  AOI22xp33_ASAP7_75t_SRAM U36148 ( .A1(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__0_), .A2(n30995), .B1(ic_q[0]), 
        .B2(n22387), .Y(n30474) );
  AOI22xp33_ASAP7_75t_SRAM U36149 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__3_), 
        .A2(n31364), .B1(n30968), .B2(n31478), .Y(n30886) );
  NOR2xp33_ASAP7_75t_SL U36150 ( .A(n29992), .B(n24483), .Y(n30026) );
  NOR2xp33_ASAP7_75t_SL U36151 ( .A(n25437), .B(n24482), .Y(n31484) );
  OAI22xp33_ASAP7_75t_SRAM U36152 ( .A1(n31467), .A2(n31466), .B1(n32602), 
        .B2(n31465), .Y(n31468) );
  AOI22xp33_ASAP7_75t_SRAM U36153 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__2_), 
        .A2(n31364), .B1(n31044), .B2(n31478), .Y(n31006) );
  NOR2xp33_ASAP7_75t_SL U36154 ( .A(n26154), .B(n26153), .Y(n28667) );
  NOR2xp33_ASAP7_75t_SL U36155 ( .A(n26559), .B(n26558), .Y(n27209) );
  NOR2xp33_ASAP7_75t_SL U36156 ( .A(n23551), .B(n30575), .Y(n27254) );
  NOR2xp33_ASAP7_75t_SL U36157 ( .A(n26335), .B(n30575), .Y(n26336) );
  AOI31xp33_ASAP7_75t_SL U36158 ( .A1(n26334), .A2(n26333), .A3(n26332), .B(
        n26331), .Y(n30025) );
  AOI22xp33_ASAP7_75t_SRAM U36159 ( .A1(n30130), .A2(n32639), .B1(dt_q[17]), 
        .B2(n29991), .Y(n26334) );
  NAND4xp25_ASAP7_75t_SL U36160 ( .A(n25037), .B(n25036), .C(n25035), .D(
        n25034), .Y(n31035) );
  INVxp33_ASAP7_75t_SRAM U36161 ( .A(n3135), .Y(n25040) );
  INVxp33_ASAP7_75t_SRAM U36162 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__9_), .Y(
        n27069) );
  O2A1O1Ixp5_ASAP7_75t_SL U36163 ( .A1(n32703), .A2(romsn[0]), .B(n32699), .C(
        n32701), .Y(n1661) );
  O2A1O1Ixp5_ASAP7_75t_SL U36164 ( .A1(n32703), .A2(romsn[1]), .B(n32702), .C(
        n32701), .Y(n1659) );
  NOR2xp33_ASAP7_75t_SL U36165 ( .A(n29918), .B(n29917), .Y(n31479) );
  AOI31xp33_ASAP7_75t_SL U36166 ( .A1(n27253), .A2(n27252), .A3(n27251), .B(
        n27250), .Y(n31356) );
  AND2x2_ASAP7_75t_SL U36167 ( .A(n30023), .B(n30022), .Y(n31478) );
  NOR2xp33_ASAP7_75t_SL U36168 ( .A(n30127), .B(n30126), .Y(n30128) );
  NOR2xp33_ASAP7_75t_SL U36169 ( .A(n30016), .B(n25441), .Y(n29913) );
  NOR2xp33_ASAP7_75t_SL U36170 ( .A(n25440), .B(n29916), .Y(n29914) );
  NOR2xp33_ASAP7_75t_SL U36171 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_ASI__0_), 
        .B(n14803), .Y(n25028) );
  O2A1O1Ixp5_ASAP7_75t_SL U36172 ( .A1(n25021), .A2(n25583), .B(n25027), .C(
        n25026), .Y(n25033) );
  NOR2xp33_ASAP7_75t_SL U36173 ( .A(n31340), .B(n29795), .Y(n29803) );
  O2A1O1Ixp5_ASAP7_75t_SL U36174 ( .A1(n30595), .A2(n28516), .B(n28515), .C(
        n28514), .Y(n2517) );
  INVxp33_ASAP7_75t_SRAM U36175 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__15_), .Y(
        n26896) );
  INVxp33_ASAP7_75t_SRAM U36176 ( .A(u0_0_leon3x0_p0_divi[58]), .Y(n26894) );
  AOI21xp33_ASAP7_75t_SRAM U36177 ( .A1(n30264), .A2(n28835), .B(n26418), .Y(
        n26420) );
  INVxp33_ASAP7_75t_SRAM U36178 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__13_), .Y(
        n28422) );
  NOR2xp33_ASAP7_75t_SL U36179 ( .A(n31340), .B(n29768), .Y(n29790) );
  NOR2xp33_ASAP7_75t_SL U36180 ( .A(n25474), .B(n25473), .Y(n28443) );
  NAND2xp33_ASAP7_75t_SRAM U36181 ( .A(n30257), .B(n28835), .Y(n26396) );
  INVxp33_ASAP7_75t_SRAM U36182 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__12_), .Y(
        n26397) );
  INVxp33_ASAP7_75t_SRAM U36183 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__17_), .Y(
        n25896) );
  AOI211xp5_ASAP7_75t_SL U36184 ( .A1(n31342), .A2(n28275), .B(n26949), .C(
        n26948), .Y(n28279) );
  NOR2xp33_ASAP7_75t_SL U36185 ( .A(n31340), .B(n28273), .Y(n26949) );
  NAND2xp33_ASAP7_75t_SRAM U36186 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__28_), 
        .B(n29589), .Y(n26928) );
  INVxp33_ASAP7_75t_SRAM U36187 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__16_), .Y(
        n26929) );
  INVxp33_ASAP7_75t_SRAM U36188 ( .A(u0_0_leon3x0_p0_divi[59]), .Y(n26927) );
  AOI22xp33_ASAP7_75t_SRAM U36189 ( .A1(n29605), .A2(n26914), .B1(n29603), 
        .B2(n29604), .Y(n26942) );
  O2A1O1Ixp5_ASAP7_75t_SL U36190 ( .A1(n28821), .A2(n22721), .B(n28626), .C(
        n28625), .Y(n28627) );
  O2A1O1Ixp5_ASAP7_75t_SL U36191 ( .A1(n28725), .A2(n24489), .B(n28724), .C(
        n28723), .Y(n30396) );
  O2A1O1Ixp5_ASAP7_75t_SL U36192 ( .A1(u0_0_leon3x0_p0_divi[12]), .A2(n28931), 
        .B(n26163), .C(n23396), .Y(n26164) );
  O2A1O1Ixp5_ASAP7_75t_SL U36193 ( .A1(n28830), .A2(n26168), .B(n26162), .C(
        n27200), .Y(n26166) );
  O2A1O1Ixp5_ASAP7_75t_SL U36194 ( .A1(n24691), .A2(n28436), .B(n28435), .C(
        n28434), .Y(n30250) );
  NOR2xp33_ASAP7_75t_SL U36195 ( .A(n27241), .B(n31870), .Y(n26751) );
  NOR2xp33_ASAP7_75t_SL U36196 ( .A(n26750), .B(n28365), .Y(n31870) );
  AND2x2_ASAP7_75t_SL U36197 ( .A(n26368), .B(n26367), .Y(n24428) );
  OR2x2_ASAP7_75t_SL U36198 ( .A(n26368), .B(n26366), .Y(n24514) );
  NOR2xp33_ASAP7_75t_SL U36199 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__WY_), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__WY_), .Y(n26367) );
  O2A1O1Ixp5_ASAP7_75t_SL U36200 ( .A1(u0_0_leon3x0_p0_divi[0]), .A2(n29150), 
        .B(n26743), .C(n23980), .Y(n26744) );
  NOR2xp33_ASAP7_75t_SL U36201 ( .A(n26738), .B(n30446), .Y(n26750) );
  NOR2xp33_ASAP7_75t_SL U36202 ( .A(n26733), .B(n26732), .Y(n29863) );
  NAND3xp33_ASAP7_75t_SL U36203 ( .A(n26733), .B(
        u0_0_leon3x0_p0_iu_r_A__RSEL2__0_), .C(
        u0_0_leon3x0_p0_iu_r_A__RSEL2__1_), .Y(n29865) );
  OR2x2_ASAP7_75t_SL U36204 ( .A(n26872), .B(n26731), .Y(n24541) );
  NOR2xp33_ASAP7_75t_SL U36205 ( .A(n31760), .B(n31733), .Y(n32704) );
  NOR2xp33_ASAP7_75t_SL U36206 ( .A(n31732), .B(n32709), .Y(n31733) );
  NOR2xp33_ASAP7_75t_SL U36207 ( .A(n2292), .B(n32741), .Y(n32742) );
  INVxp33_ASAP7_75t_SRAM U36208 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__18_), .Y(
        n29593) );
  NOR2xp33_ASAP7_75t_SL U36209 ( .A(n28968), .B(n30635), .Y(n29603) );
  AND2x2_ASAP7_75t_SL U36210 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_), 
        .B(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__30_), .Y(n25705) );
  O2A1O1Ixp5_ASAP7_75t_SL U36211 ( .A1(u0_0_leon3x0_p0_divi[19]), .A2(n29150), 
        .B(n26991), .C(n22952), .Y(n26992) );
  NAND3xp33_ASAP7_75t_SL U36212 ( .A(n25210), .B(
        u0_0_leon3x0_p0_iu_r_A__RSEL1__1_), .C(
        u0_0_leon3x0_p0_iu_r_A__RSEL1__0_), .Y(n31396) );
  NOR2xp33_ASAP7_75t_SL U36213 ( .A(n29870), .B(n29816), .Y(n30666) );
  AOI21xp33_ASAP7_75t_SRAM U36214 ( .A1(n30660), .A2(n22919), .B(n24519), .Y(
        n30661) );
  NAND2xp33_ASAP7_75t_SRAM U36215 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__31_), 
        .B(n24581), .Y(n25179) );
  NOR2xp33_ASAP7_75t_SL U36216 ( .A(n24427), .B(n28481), .Y(n27067) );
  NAND2xp33_ASAP7_75t_SRAM U36217 ( .A(n22919), .B(n32130), .Y(n25178) );
  NOR2xp33_ASAP7_75t_SL U36218 ( .A(n25176), .B(n28934), .Y(n26174) );
  NOR2xp33_ASAP7_75t_SL U36219 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__23_), 
        .B(n25172), .Y(n30664) );
  INVxp33_ASAP7_75t_SRAM U36220 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__19_), .Y(
        n25175) );
  NOR2xp33_ASAP7_75t_SL U36221 ( .A(n29575), .B(n25169), .Y(n25176) );
  OR2x2_ASAP7_75t_SL U36222 ( .A(u0_0_leon3x0_p0_iu_r_E__JMPL_), .B(n29000), 
        .Y(n24427) );
  AND2x2_ASAP7_75t_SL U36223 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUOP__2_), .Y(n29147) );
  NOR2xp33_ASAP7_75t_SL U36224 ( .A(u0_0_leon3x0_p0_iu_r_E__JMPL_), .B(n25120), 
        .Y(n28877) );
  O2A1O1Ixp5_ASAP7_75t_SL U36225 ( .A1(n32131), .A2(n23923), .B(n25090), .C(
        u0_0_leon3x0_p0_iu_r_E__SHLEFT_), .Y(n25783) );
  OR2x2_ASAP7_75t_SL U36226 ( .A(n26140), .B(n25092), .Y(n24469) );
  OR2x2_ASAP7_75t_SL U36227 ( .A(u0_0_leon3x0_p0_iu_r_E__JMPL_), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_), .Y(n25123) );
  NOR4xp25_ASAP7_75t_SL U36228 ( .A(n31959), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__30_), .C(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_), .D(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_), .Y(n30663) );
  NOR2xp33_ASAP7_75t_SL U36229 ( .A(n24984), .B(n24966), .Y(n26736) );
  NAND4xp25_ASAP7_75t_SL U36230 ( .A(n24988), .B(n24986), .C(n24965), .D(
        n24983), .Y(n24966) );
  NOR2xp33_ASAP7_75t_SL U36231 ( .A(n25670), .B(n25650), .Y(n24929) );
  NOR2xp33_ASAP7_75t_SL U36232 ( .A(n25661), .B(n25684), .Y(n24965) );
  NOR2xp33_ASAP7_75t_SL U36233 ( .A(n31980), .B(n25697), .Y(n25684) );
  NOR2xp33_ASAP7_75t_SL U36234 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_), 
        .B(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), .Y(n25661) );
  NOR2xp33_ASAP7_75t_SL U36235 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_), 
        .B(n25655), .Y(n24939) );
  NOR2xp33_ASAP7_75t_SL U36236 ( .A(n25667), .B(n24964), .Y(n24988) );
  NOR2xp33_ASAP7_75t_SL U36237 ( .A(n24937), .B(n24930), .Y(n25676) );
  OAI21xp33_ASAP7_75t_SRAM U36238 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .B(n24963), .Y(n24930) );
  NOR2xp33_ASAP7_75t_SL U36239 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), 
        .B(n24944), .Y(n24937) );
  NOR2xp33_ASAP7_75t_SL U36240 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_), 
        .B(n25693), .Y(n25659) );
  NOR2xp33_ASAP7_75t_SL U36241 ( .A(n24949), .B(n24948), .Y(n24987) );
  NOR2xp33_ASAP7_75t_SL U36242 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_), 
        .B(n25692), .Y(n25667) );
  NOR2xp33_ASAP7_75t_SL U36243 ( .A(n24945), .B(n25700), .Y(n25671) );
  NOR2xp33_ASAP7_75t_SL U36244 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_), 
        .B(n25697), .Y(n25700) );
  NOR2xp33_ASAP7_75t_SL U36245 ( .A(n24944), .B(n25697), .Y(n24945) );
  NOR2xp33_ASAP7_75t_SL U36246 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), 
        .B(n25670), .Y(n25652) );
  OR2x2_ASAP7_75t_SL U36247 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), .Y(n30955) );
  NOR2xp33_ASAP7_75t_SL U36248 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), 
        .B(n25675), .Y(n25680) );
  NOR2xp33_ASAP7_75t_SL U36249 ( .A(n32792), .B(n32791), .Y(n32813) );
  NOR2xp33_ASAP7_75t_SL U36250 ( .A(n31739), .B(n31747), .Y(n32791) );
  NOR2xp33_ASAP7_75t_SL U36251 ( .A(sr1_r_BSTATE__1_), .B(n31738), .Y(n32827)
         );
  NAND3xp33_ASAP7_75t_SL U36252 ( .A(n32790), .B(read), .C(oen), .Y(n32820) );
  NOR2xp33_ASAP7_75t_SL U36253 ( .A(n31749), .B(n31748), .Y(n32790) );
  NOR2xp33_ASAP7_75t_SL U36254 ( .A(n31747), .B(n31759), .Y(n31748) );
  NOR2xp33_ASAP7_75t_SL U36255 ( .A(n31746), .B(n31745), .Y(n31759) );
  NOR2xp33_ASAP7_75t_SL U36256 ( .A(sr1_r_MCFG1__ROMWRITE_), .B(n31744), .Y(
        n31746) );
  NOR2xp33_ASAP7_75t_SL U36257 ( .A(n31751), .B(n31745), .Y(n31747) );
  NOR2xp33_ASAP7_75t_SL U36258 ( .A(n2356), .B(sr1_r_MCFG1__IOEN_), .Y(n31745)
         );
  NOR2xp33_ASAP7_75t_SL U36259 ( .A(sr1_r_BSTATE__1_), .B(sr1_r_BSTATE__0_), 
        .Y(n32832) );
  NOR2xp33_ASAP7_75t_SL U36260 ( .A(n32788), .B(n32787), .Y(n32817) );
  NOR2xp33_ASAP7_75t_SL U36261 ( .A(n31698), .B(n31719), .Y(n31699) );
  NOR2xp33_ASAP7_75t_SL U36262 ( .A(n31712), .B(n31714), .Y(n32717) );
  NOR2xp33_ASAP7_75t_SL U36263 ( .A(sr1_r_READY_), .B(n31753), .Y(n32716) );
  AO21x1_ASAP7_75t_SL U36264 ( .A1(sr1_r_MCFG2__RAMBANKSZ__0_), .A2(n32785), 
        .B(n32769), .Y(n32811) );
  NOR2xp33_ASAP7_75t_SL U36265 ( .A(n2924), .B(sr1_r_MCFG2__RAMBANKSZ__3_), 
        .Y(n32771) );
  AND2x2_ASAP7_75t_SL U36266 ( .A(n2924), .B(sr1_r_MCFG2__RAMBANKSZ__3_), .Y(
        n32772) );
  NOR2xp33_ASAP7_75t_SL U36267 ( .A(n2924), .B(n32762), .Y(n32775) );
  NOR2xp33_ASAP7_75t_SL U36268 ( .A(sr1_r_MCFG2__RAMBANKSZ__3_), .B(n32761), 
        .Y(n32773) );
  NOR2xp33_ASAP7_75t_SL U36269 ( .A(n2924), .B(n32774), .Y(n32753) );
  INVxp33_ASAP7_75t_SRAM U36270 ( .A(n32085), .Y(n32088) );
  NAND2xp33_ASAP7_75t_SRAM U36271 ( .A(n32689), .B(n31897), .Y(n31936) );
  NOR2xp33_ASAP7_75t_SL U36272 ( .A(n32097), .B(n32104), .Y(n31387) );
  NOR2xp33_ASAP7_75t_SL U36273 ( .A(n18819), .B(n18842), .Y(n31379) );
  HB1xp67_ASAP7_75t_SL U36274 ( .A(n31679), .Y(n24639) );
  NOR2xp33_ASAP7_75t_SL U36275 ( .A(n24430), .B(n26187), .Y(n31679) );
  AOI31xp33_ASAP7_75t_SL U36276 ( .A1(n32057), .A2(n32091), .A3(n32056), .B(
        n32104), .Y(n32058) );
  NAND2xp33_ASAP7_75t_SRAM U36277 ( .A(n4318), .B(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_NOMDS_), .Y(n31446) );
  NOR2xp33_ASAP7_75t_SL U36278 ( .A(n31881), .B(n31880), .Y(n31882) );
  NOR2xp33_ASAP7_75t_SL U36279 ( .A(n22380), .B(n32045), .Y(n32129) );
  NOR4xp25_ASAP7_75t_SL U36280 ( .A(n31932), .B(n31931), .C(n31930), .D(n31929), .Y(n32454) );
  NAND4xp25_ASAP7_75t_SL U36281 ( .A(n31928), .B(n31927), .C(n31926), .D(
        n31925), .Y(n31929) );
  XNOR2xp5_ASAP7_75t_SL U36282 ( .A(it_q[18]), .B(u0_0_leon3x0_p0_ici[80]), 
        .Y(n31925) );
  XNOR2xp5_ASAP7_75t_SL U36283 ( .A(it_q[24]), .B(u0_0_leon3x0_p0_ici[86]), 
        .Y(n31926) );
  XNOR2xp5_ASAP7_75t_SL U36284 ( .A(it_q[20]), .B(u0_0_leon3x0_p0_ici[82]), 
        .Y(n31928) );
  NAND4xp25_ASAP7_75t_SL U36285 ( .A(n31924), .B(n31923), .C(n31922), .D(
        n31921), .Y(n31930) );
  NAND4xp25_ASAP7_75t_SL U36286 ( .A(n31920), .B(n31919), .C(n31918), .D(
        n31917), .Y(n31931) );
  AND2x2_ASAP7_75t_SL U36287 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__0_), 
        .B(n3135), .Y(n32482) );
  OAI22xp33_ASAP7_75t_SRAM U36288 ( .A1(n32497), .A2(n32669), .B1(
        u0_0_leon3x0_p0_ici[60]), .B2(n32491), .Y(n31904) );
  NOR2xp33_ASAP7_75t_SL U36289 ( .A(n31901), .B(n31900), .Y(n31906) );
  NAND2xp33_ASAP7_75t_SRAM U36290 ( .A(it_q[3]), .B(u0_0_leon3x0_p0_ici[60]), 
        .Y(n31899) );
  NAND2xp33_ASAP7_75t_SRAM U36291 ( .A(it_q[1]), .B(u0_0_leon3x0_p0_ici[60]), 
        .Y(n31898) );
  NOR2xp33_ASAP7_75t_SL U36292 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_UNDERRUN_), 
        .B(n31879), .Y(n31894) );
  NOR2xp33_ASAP7_75t_SL U36293 ( .A(n31891), .B(n32125), .Y(n32124) );
  OAI21xp33_ASAP7_75t_SRAM U36294 ( .A1(u0_0_leon3x0_p0_c0mmu_mcii[0]), .A2(
        n32662), .B(u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_), .Y(n32125) );
  NOR2xp33_ASAP7_75t_SL U36295 ( .A(u0_0_dbgo_OPTYPE__1_), .B(n29214), .Y(
        n29211) );
  XNOR2xp5_ASAP7_75t_SL U36296 ( .A(n32169), .B(n26805), .Y(n29202) );
  NAND2xp33_ASAP7_75t_SRAM U36297 ( .A(n22379), .B(n26797), .Y(n26798) );
  XNOR2xp5_ASAP7_75t_SL U36298 ( .A(u0_0_leon3x0_p0_iu_r_W__S__CWP__2_), .B(
        n26787), .Y(n26801) );
  NOR2xp33_ASAP7_75t_SL U36299 ( .A(n26783), .B(n31426), .Y(n31429) );
  NAND2xp33_ASAP7_75t_SRAM U36300 ( .A(n22379), .B(n26766), .Y(n26767) );
  INVxp33_ASAP7_75t_SRAM U36301 ( .A(n26791), .Y(n26764) );
  NOR2xp33_ASAP7_75t_SL U36302 ( .A(n25606), .B(n26758), .Y(n25608) );
  NOR2xp33_ASAP7_75t_SL U36303 ( .A(u0_0_dbgo_OPTYPE__0_), .B(n25605), .Y(
        n26791) );
  NOR2xp33_ASAP7_75t_SL U36304 ( .A(n26759), .B(n26758), .Y(n29179) );
  NOR3xp33_ASAP7_75t_SL U36305 ( .A(n31984), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__ANNUL_), .C(u0_0_dbgo_OPTYPE__4_), .Y(
        n25451) );
  NOR2xp33_ASAP7_75t_SL U36306 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__20_), 
        .B(n26756), .Y(n26789) );
  NAND2xp33_ASAP7_75t_SRAM U36307 ( .A(u0_0_dbgo_OPTYPE__1_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__19_), .Y(n26756) );
  NOR2xp33_ASAP7_75t_SL U36308 ( .A(n26755), .B(n26754), .Y(n26761) );
  NAND2xp33_ASAP7_75t_SRAM U36309 ( .A(u0_0_dbgo_OPTYPE__1_), .B(n26753), .Y(
        n26754) );
  NOR2xp33_ASAP7_75t_SL U36310 ( .A(u0_0_leon3x0_p0_iu_r_D__ANNUL_), .B(n24889), .Y(n24872) );
  NOR2xp33_ASAP7_75t_SL U36311 ( .A(n30681), .B(n24735), .Y(n24869) );
  NOR2xp33_ASAP7_75t_SL U36312 ( .A(n29741), .B(n24680), .Y(n31352) );
  NOR2xp33_ASAP7_75t_SL U36313 ( .A(u0_0_leon3x0_p0_iu_r_A__CTRL__ANNUL_), .B(
        u0_0_leon3x0_p0_iu_r_A__CTRL__TT__0_), .Y(n31811) );
  O2A1O1Ixp5_ASAP7_75t_SL U36314 ( .A1(n31450), .A2(n31449), .B(n25014), .C(
        n32443), .Y(n25015) );
  NOR2xp33_ASAP7_75t_SL U36315 ( .A(n30533), .B(n22385), .Y(n32529) );
  NOR2xp33_ASAP7_75t_SL U36316 ( .A(n30540), .B(n22385), .Y(n32530) );
  NOR2xp33_ASAP7_75t_SL U36317 ( .A(n30506), .B(n22385), .Y(n32527) );
  NOR2xp33_ASAP7_75t_SL U36318 ( .A(n30974), .B(n22385), .Y(n32589) );
  NOR2xp33_ASAP7_75t_SL U36319 ( .A(n30526), .B(n22385), .Y(n32526) );
  NOR2xp33_ASAP7_75t_SL U36320 ( .A(n30517), .B(n22385), .Y(n32528) );
  NOR2xp33_ASAP7_75t_SL U36321 ( .A(n30828), .B(n22385), .Y(n32532) );
  NOR2xp33_ASAP7_75t_SL U36322 ( .A(n31687), .B(n22385), .Y(n32558) );
  NOR2xp33_ASAP7_75t_SL U36323 ( .A(n30524), .B(n22385), .Y(n32523) );
  NOR2xp33_ASAP7_75t_SL U36324 ( .A(n32574), .B(n22385), .Y(n32573) );
  NOR2xp33_ASAP7_75t_SL U36325 ( .A(n32580), .B(n22385), .Y(n32579) );
  NOR2xp33_ASAP7_75t_SL U36326 ( .A(n32577), .B(n22385), .Y(n32576) );
  NOR2xp33_ASAP7_75t_SL U36327 ( .A(n31454), .B(n31453), .Y(n31583) );
  NOR2xp33_ASAP7_75t_SL U36328 ( .A(n31018), .B(n22385), .Y(n32569) );
  NOR2xp33_ASAP7_75t_SL U36329 ( .A(n32567), .B(n22385), .Y(n32560) );
  NOR2xp33_ASAP7_75t_SL U36330 ( .A(n31690), .B(n22385), .Y(n32555) );
  NOR2xp33_ASAP7_75t_SL U36331 ( .A(n31834), .B(n22385), .Y(n32531) );
  NOR2xp33_ASAP7_75t_SL U36332 ( .A(n31786), .B(n22385), .Y(n32553) );
  NOR2xp33_ASAP7_75t_SL U36333 ( .A(n31765), .B(n22385), .Y(n32536) );
  NOR2xp33_ASAP7_75t_SL U36334 ( .A(n32586), .B(n22385), .Y(n32582) );
  NOR2xp33_ASAP7_75t_SL U36335 ( .A(n32669), .B(n22385), .Y(n32664) );
  NOR2x1_ASAP7_75t_SL U36336 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_), 
        .B(n31883), .Y(n32564) );
  XNOR2xp5_ASAP7_75t_SL U36337 ( .A(n2933), .B(n32662), .Y(n30913) );
  NOR2xp33_ASAP7_75t_SL U36338 ( .A(n28100), .B(n28105), .Y(n32293) );
  OAI22xp33_ASAP7_75t_SRAM U36339 ( .A1(n32410), .A2(n24637), .B1(n32417), 
        .B2(n22383), .Y(n26488) );
  OAI22xp33_ASAP7_75t_SRAM U36340 ( .A1(n32333), .A2(n24637), .B1(n32332), 
        .B2(n22383), .Y(n28134) );
  OAI22xp33_ASAP7_75t_SRAM U36341 ( .A1(n32315), .A2(n24637), .B1(n32314), 
        .B2(n22383), .Y(n25856) );
  OAI22xp33_ASAP7_75t_SRAM U36342 ( .A1(n31509), .A2(n24637), .B1(n32405), 
        .B2(n22383), .Y(n25434) );
  OAI22xp33_ASAP7_75t_SRAM U36343 ( .A1(n32367), .A2(n24637), .B1(n32366), 
        .B2(n22383), .Y(n25714) );
  OAI22xp33_ASAP7_75t_SRAM U36344 ( .A1(n30155), .A2(n24637), .B1(n32325), 
        .B2(n22383), .Y(n25411) );
  OAI22xp33_ASAP7_75t_SRAM U36345 ( .A1(n32382), .A2(n24637), .B1(n32383), 
        .B2(n22383), .Y(n26220) );
  INVx1_ASAP7_75t_SL U36346 ( .A(n2929), .Y(n31529) );
  NOR2xp33_ASAP7_75t_SL U36347 ( .A(n31577), .B(n31576), .Y(n31590) );
  NAND2xp33_ASAP7_75t_SRAM U36348 ( .A(n31571), .B(n31570), .Y(n31598) );
  NAND2xp33_ASAP7_75t_SRAM U36349 ( .A(n4318), .B(n32274), .Y(n31571) );
  NOR2xp33_ASAP7_75t_SL U36350 ( .A(n3134), .B(n25409), .Y(n32274) );
  NOR2xp33_ASAP7_75t_SL U36351 ( .A(n31455), .B(n32443), .Y(n25402) );
  NOR2xp33_ASAP7_75t_SL U36352 ( .A(u0_0_leon3x0_p0_ico_DIAGRDY_), .B(n13499), 
        .Y(n31564) );
  NOR2xp33_ASAP7_75t_SL U36353 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_), .B(n3134), .Y(n32238) );
  NOR2xp33_ASAP7_75t_SL U36354 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__0_), 
        .B(n30180), .Y(n30164) );
  NOR2xp33_ASAP7_75t_SL U36355 ( .A(n31303), .B(n32193), .Y(n31464) );
  INVxp33_ASAP7_75t_SRAM U36356 ( .A(ahb0_r_DEFSLV_), .Y(n25599) );
  AOI31xp33_ASAP7_75t_SL U36357 ( .A1(n32524), .A2(n3065), .A3(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__6_), .B(n31561), .Y(n3066) );
  NOR2xp33_ASAP7_75t_SL U36358 ( .A(n3054), .B(n30181), .Y(n30183) );
  NOR2xp33_ASAP7_75t_SL U36359 ( .A(n30407), .B(n29736), .Y(n29739) );
  NOR2xp33_ASAP7_75t_SL U36360 ( .A(u0_0_leon3x0_p0_div0_v_ZERO2_), .B(n22421), 
        .Y(n25936) );
  INVxp33_ASAP7_75t_SRAM U36361 ( .A(u0_0_leon3x0_p0_div0_addout_4_), .Y(
        n25923) );
  INVxp33_ASAP7_75t_SRAM U36362 ( .A(u0_0_leon3x0_p0_div0_addout_5_), .Y(
        n25925) );
  AOI31xp33_ASAP7_75t_SL U36363 ( .A1(n32066), .A2(n32010), .A3(
        u0_0_leon3x0_p0_iu_r_A__DIVSTART_), .B(n31678), .Y(n25919) );
  NOR2xp33_ASAP7_75t_SL U36364 ( .A(u0_0_leon3x0_p0_div0_addout_17_), .B(
        u0_0_leon3x0_p0_div0_addout_18_), .Y(n25922) );
  AOI22xp33_ASAP7_75t_SRAM U36365 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__3_), .B1(u0_0_leon3x0_p0_divo[3]), .B2(
        n28371), .Y(n28358) );
  AOI22xp33_ASAP7_75t_SRAM U36366 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__4_), .B1(u0_0_leon3x0_p0_divo[4]), .B2(
        n28371), .Y(n28354) );
  AOI22xp33_ASAP7_75t_SRAM U36367 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__0_), .B1(u0_0_leon3x0_p0_divo[0]), .B2(
        n28371), .Y(n28368) );
  AOI21xp33_ASAP7_75t_SRAM U36368 ( .A1(u0_0_leon3x0_p0_divo[0]), .A2(n31658), 
        .B(n22431), .Y(n28374) );
  INVxp33_ASAP7_75t_SRAM U36369 ( .A(n3727), .Y(n28372) );
  AOI22xp33_ASAP7_75t_SRAM U36370 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__1_), .B1(u0_0_leon3x0_p0_divo[1]), .B2(
        n28371), .Y(n28362) );
  AOI22xp33_ASAP7_75t_SRAM U36371 ( .A1(n22431), .A2(
        u0_0_leon3x0_p0_div0_r_X__2_), .B1(u0_0_leon3x0_p0_divo[2]), .B2(
        n28371), .Y(n28360) );
  NOR2xp33_ASAP7_75t_SL U36372 ( .A(n4949), .B(n28379), .Y(n29109) );
  AND2x2_ASAP7_75t_SL U36373 ( .A(n3725), .B(n3727), .Y(n29112) );
  AND2x2_ASAP7_75t_SL U36374 ( .A(n4325), .B(n3727), .Y(n28291) );
  NOR2xp33_ASAP7_75t_SL U36375 ( .A(u0_0_leon3x0_p0_ici[62]), .B(n22379), .Y(
        n29480) );
  NOR2xp33_ASAP7_75t_SL U36376 ( .A(n25596), .B(n25595), .Y(n2998) );
  INVx2_ASAP7_75t_SL U36377 ( .A(apbi[7]), .Y(n30833) );
  INVx2_ASAP7_75t_SL U36378 ( .A(apbi[4]), .Y(n30780) );
  INVx2_ASAP7_75t_SL U36379 ( .A(apbi[5]), .Y(n30073) );
  INVx2_ASAP7_75t_SL U36380 ( .A(apbi[3]), .Y(n29510) );
  INVx2_ASAP7_75t_SL U36381 ( .A(apbi[6]), .Y(n31197) );
  HB1xp67_ASAP7_75t_SL U36382 ( .A(n31841), .Y(n24640) );
  NOR2xp33_ASAP7_75t_SL U36383 ( .A(timer0_vtimers_1__LOAD_), .B(n26472), .Y(
        n26473) );
  NOR2xp33_ASAP7_75t_SL U36384 ( .A(n26468), .B(n31953), .Y(n26469) );
  OR2x2_ASAP7_75t_SL U36385 ( .A(n27479), .B(n26467), .Y(n31953) );
  NOR2xp33_ASAP7_75t_SL U36386 ( .A(n25984), .B(n25988), .Y(n27463) );
  NAND2xp5_ASAP7_75t_SL U36387 ( .A(apbi[34]), .B(n25941), .Y(n25988) );
  NOR2xp33_ASAP7_75t_SL U36388 ( .A(n25532), .B(n25531), .Y(n25941) );
  NOR2xp33_ASAP7_75t_SL U36389 ( .A(apbi[39]), .B(apbi[38]), .Y(n25528) );
  NOR2xp33_ASAP7_75t_SL U36390 ( .A(apbi[43]), .B(apbi[42]), .Y(n25529) );
  NOR2xp33_ASAP7_75t_SL U36391 ( .A(apbi[44]), .B(apbi[45]), .Y(n25530) );
  NOR2xp33_ASAP7_75t_SL U36392 ( .A(apbi[37]), .B(apbi[36]), .Y(n25527) );
  INVx1_ASAP7_75t_SL U36393 ( .A(apbi[35]), .Y(n25984) );
  NOR2xp33_ASAP7_75t_SL U36394 ( .A(n2925), .B(n1637), .Y(n25846) );
  INVx1_ASAP7_75t_SL U36395 ( .A(apbi[33]), .Y(n25952) );
  NOR2x1_ASAP7_75t_SL U36396 ( .A(n25986), .B(n25985), .Y(n26097) );
  INVx1_ASAP7_75t_SL U36397 ( .A(apbi[32]), .Y(n25985) );
  NOR2xp33_ASAP7_75t_SL U36398 ( .A(n5061), .B(n1752), .Y(timer0_N78) );
  NOR2xp33_ASAP7_75t_SL U36399 ( .A(n5061), .B(n2322), .Y(timer0_N77) );
  NOR2xp33_ASAP7_75t_SL U36400 ( .A(n5061), .B(n1728), .Y(timer0_N85) );
  NOR2xp33_ASAP7_75t_SL U36401 ( .A(n5061), .B(n1630), .Y(timer0_N87) );
  NOR2xp33_ASAP7_75t_SL U36402 ( .A(n5061), .B(n2838), .Y(timer0_N86) );
  NOR2xp33_ASAP7_75t_SL U36403 ( .A(n5061), .B(n2840), .Y(timer0_N88) );
  NOR2xp33_ASAP7_75t_SL U36404 ( .A(n26463), .B(n26462), .Y(n26472) );
  NOR2xp33_ASAP7_75t_SL U36405 ( .A(n4742), .B(timer0_gpto_TICK__1_), .Y(
        n26462) );
  NOR2xp33_ASAP7_75t_SL U36406 ( .A(n24512), .B(n26508), .Y(n32391) );
  O2A1O1Ixp5_ASAP7_75t_SL U36407 ( .A1(n31608), .A2(n31607), .B(n32445), .C(
        n31606), .Y(n31610) );
  NOR2xp33_ASAP7_75t_SL U36408 ( .A(n31603), .B(n32719), .Y(n32451) );
  NOR2xp33_ASAP7_75t_SL U36409 ( .A(n24898), .B(n24974), .Y(n25245) );
  NOR2xp33_ASAP7_75t_SL U36410 ( .A(n4082), .B(n31876), .Y(n24898) );
  AND2x2_ASAP7_75t_SL U36411 ( .A(u0_0_leon3x0_p0_c0mmu_a0_r_NBA_), .B(
        u0_0_leon3x0_p0_c0mmu_a0_r_NBO__1_), .Y(n24479) );
  NOR2xp33_ASAP7_75t_SL U36412 ( .A(n24977), .B(n22393), .Y(n31897) );
  OR2x2_ASAP7_75t_SL U36413 ( .A(n4076), .B(
        u0_0_leon3x0_p0_c0mmu_a0_r_HLOCKEN_), .Y(n31604) );
  NOR2xp33_ASAP7_75t_SL U36414 ( .A(n31589), .B(n31591), .Y(n31601) );
  AND2x2_ASAP7_75t_SL U36415 ( .A(u0_0_leon3x0_p0_dci[4]), .B(
        u0_0_leon3x0_p0_dci[5]), .Y(n31584) );
  NOR2xp33_ASAP7_75t_SL U36416 ( .A(n31297), .B(n32284), .Y(n31463) );
  NOR4xp25_ASAP7_75t_SL U36417 ( .A(n24534), .B(n31295), .C(n31294), .D(n31293), .Y(n31301) );
  NAND4xp25_ASAP7_75t_SL U36418 ( .A(n31292), .B(n31291), .C(n31290), .D(
        n31289), .Y(n31293) );
  XNOR2xp5_ASAP7_75t_SL U36419 ( .A(dt_q[24]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[28]), .Y(n31290) );
  XNOR2xp5_ASAP7_75t_SL U36420 ( .A(dt_q[23]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[27]), .Y(n31291) );
  XNOR2xp5_ASAP7_75t_SL U36421 ( .A(dt_q[21]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[25]), .Y(n31292) );
  NAND4xp25_ASAP7_75t_SL U36422 ( .A(n31288), .B(n31287), .C(n31286), .D(
        n31285), .Y(n31294) );
  NAND4xp25_ASAP7_75t_SL U36423 ( .A(n31284), .B(n31283), .C(n31282), .D(
        n31281), .Y(n31295) );
  XNOR2xp5_ASAP7_75t_SL U36424 ( .A(dt_q[20]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[24]), .Y(n31281) );
  XNOR2xp5_ASAP7_75t_SL U36425 ( .A(dt_q[22]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[26]), .Y(n31282) );
  NOR2xp33_ASAP7_75t_SL U36426 ( .A(n31280), .B(n31279), .Y(n31284) );
  XNOR2xp5_ASAP7_75t_SL U36427 ( .A(n31277), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[30]), .Y(n31280) );
  XNOR2xp5_ASAP7_75t_SL U36428 ( .A(dt_q[8]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[12]), .Y(n31273) );
  XNOR2xp5_ASAP7_75t_SL U36429 ( .A(dt_q[12]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[16]), .Y(n31270) );
  NOR2xp33_ASAP7_75t_SL U36430 ( .A(n31266), .B(n31265), .Y(n31296) );
  NAND2xp33_ASAP7_75t_SRAM U36431 ( .A(u0_0_leon3x0_p0_dci[40]), .B(n31264), 
        .Y(n31297) );
  NOR2xp33_ASAP7_75t_SL U36432 ( .A(n24518), .B(n25421), .Y(n29861) );
  NOR2xp33_ASAP7_75t_SL U36433 ( .A(n24535), .B(n30005), .Y(n32311) );
  NOR2xp33_ASAP7_75t_SL U36434 ( .A(n24537), .B(n25854), .Y(n32315) );
  NOR2xp33_ASAP7_75t_SL U36435 ( .A(n3899), .B(ahb0_r_CFGA11_), .Y(n30001) );
  NOR2xp33_ASAP7_75t_SL U36436 ( .A(n3899), .B(n30975), .Y(n30000) );
  NOR2xp33_ASAP7_75t_SL U36437 ( .A(n3899), .B(n30975), .Y(n24574) );
  NOR2xp33_ASAP7_75t_SL U36438 ( .A(n25571), .B(n32662), .Y(n25572) );
  NOR2xp33_ASAP7_75t_SL U36439 ( .A(n25569), .B(n25568), .Y(n25570) );
  NAND3xp33_ASAP7_75t_SL U36440 ( .A(n32689), .B(
        u0_0_leon3x0_p0_c0mmu_icache0_r_OVERRUN_), .C(n25567), .Y(n25571) );
  INVx1_ASAP7_75t_SL U36441 ( .A(n32676), .Y(n32689) );
  NAND2xp5_ASAP7_75t_SL U36442 ( .A(n3880), .B(
        u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_), .Y(n32676) );
  NOR2xp33_ASAP7_75t_SL U36443 ( .A(u0_0_leon3x0_p0_iu_r_X__MEXC_), .B(n26137), 
        .Y(n29731) );
  OR2x2_ASAP7_75t_SL U36444 ( .A(n25946), .B(n25945), .Y(n26137) );
  NAND4xp25_ASAP7_75t_SL U36445 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__3_), 
        .B(u0_0_leon3x0_p0_iu_r_X__CTRL__TT__5_), .C(
        u0_0_leon3x0_p0_iu_r_X__CTRL__TT__2_), .D(
        u0_0_leon3x0_p0_iu_r_X__CTRL__TT__1_), .Y(n25945) );
  NOR2xp33_ASAP7_75t_SL U36446 ( .A(n31559), .B(n32566), .Y(n31554) );
  NOR2xp33_ASAP7_75t_SL U36447 ( .A(n30174), .B(n30175), .Y(n30179) );
  NAND4xp25_ASAP7_75t_SL U36448 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__0_), .B(u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__3_), .C(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__2_), .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__1_), .Y(n30175) );
  NOR2xp33_ASAP7_75t_SL U36449 ( .A(n32258), .B(n30180), .Y(n30163) );
  NOR2xp33_ASAP7_75t_SL U36450 ( .A(n30202), .B(n31265), .Y(n30915) );
  NOR2xp33_ASAP7_75t_SL U36451 ( .A(n3046), .B(n30201), .Y(n31283) );
  NOR2xp33_ASAP7_75t_SL U36452 ( .A(n30510), .B(n30509), .Y(n32736) );
  NOR2xp33_ASAP7_75t_SL U36453 ( .A(n32243), .B(n32446), .Y(n30507) );
  INVx1_ASAP7_75t_SL U36454 ( .A(n32443), .Y(n32446) );
  NAND2xp33_ASAP7_75t_SRAM U36455 ( .A(n3071), .B(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_RBURST_), .Y(n32712) );
  INVx1_ASAP7_75t_SL U36456 ( .A(n24682), .Y(n24678) );
  NOR4xp25_ASAP7_75t_SL U36457 ( .A(n29996), .B(n29995), .C(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__5_), .D(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__7_), .Y(n29997) );
  NAND4xp25_ASAP7_75t_SL U36458 ( .A(n31260), .B(n32681), .C(n31573), .D(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_CCTRLWR_), .Y(n29996) );
  INVxp33_ASAP7_75t_SRAM U36459 ( .A(n4318), .Y(n31258) );
  NOR2xp33_ASAP7_75t_SL U36460 ( .A(n31263), .B(n31575), .Y(n31458) );
  NOR2xp33_ASAP7_75t_SL U36461 ( .A(n25580), .B(n25579), .Y(n31585) );
  NOR3xp33_ASAP7_75t_SL U36462 ( .A(n25574), .B(u0_0_leon3x0_p0_dci[41]), .C(
        u0_0_leon3x0_p0_dci[40]), .Y(n25580) );
  NOR2xp33_ASAP7_75t_SL U36463 ( .A(n30196), .B(n30193), .Y(n25584) );
  NOR2xp33_ASAP7_75t_SL U36464 ( .A(u0_0_leon3x0_p0_dci[40]), .B(n25585), .Y(
        n30197) );
  NOR2xp33_ASAP7_75t_SL U36465 ( .A(n30119), .B(n25581), .Y(n30192) );
  NOR2xp33_ASAP7_75t_SL U36466 ( .A(u0_0_leon3x0_p0_dci[37]), .B(n25575), .Y(
        n25576) );
  NOR2xp33_ASAP7_75t_SL U36467 ( .A(u0_0_leon3x0_p0_dci[40]), .B(
        u0_0_leon3x0_p0_dci[39]), .Y(n30161) );
  AND2x2_ASAP7_75t_SL U36468 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__3_), 
        .B(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__4_), .Y(n31558) );
  OAI22xp33_ASAP7_75t_SRAM U36469 ( .A1(n26523), .A2(n26522), .B1(n26521), 
        .B2(n30007), .Y(n26525) );
  NOR2xp33_ASAP7_75t_SL U36470 ( .A(n26454), .B(n26216), .Y(n26219) );
  NOR2xp33_ASAP7_75t_SL U36471 ( .A(n25628), .B(n25645), .Y(n27215) );
  NOR2xp33_ASAP7_75t_SL U36472 ( .A(n26231), .B(n26612), .Y(n32401) );
  NOR2xp33_ASAP7_75t_SL U36473 ( .A(n26342), .B(n28133), .Y(n32402) );
  AOI22xp33_ASAP7_75t_SRAM U36474 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__27_), 
        .A2(n22375), .B1(n26950), .B2(n28403), .Y(n26339) );
  NOR2xp33_ASAP7_75t_SL U36475 ( .A(n26613), .B(n26612), .Y(n32329) );
  NOR2xp33_ASAP7_75t_SL U36476 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .B(
        n26230), .Y(n26612) );
  NOR2xp33_ASAP7_75t_SL U36477 ( .A(n22375), .B(n28692), .Y(n28133) );
  NOR2xp33_ASAP7_75t_SL U36478 ( .A(n25408), .B(n28406), .Y(n32325) );
  NAND2xp33_ASAP7_75t_SRAM U36479 ( .A(n30007), .B(n26918), .Y(n25431) );
  NOR2xp33_ASAP7_75t_SL U36480 ( .A(n26169), .B(n28823), .Y(n28825) );
  NOR2xp33_ASAP7_75t_SL U36481 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .B(
        n26447), .Y(n26509) );
  NOR2xp33_ASAP7_75t_SL U36482 ( .A(n22375), .B(n25428), .Y(n28402) );
  NOR2xp33_ASAP7_75t_SL U36483 ( .A(n25855), .B(n28486), .Y(n25428) );
  NOR2xp33_ASAP7_75t_SL U36484 ( .A(n25624), .B(n22392), .Y(n28486) );
  AND2x2_ASAP7_75t_SL U36485 ( .A(n25488), .B(n22392), .Y(n28403) );
  NOR2xp33_ASAP7_75t_SL U36486 ( .A(n26482), .B(n26454), .Y(n28405) );
  NOR2xp33_ASAP7_75t_SL U36487 ( .A(n26454), .B(n30009), .Y(n26483) );
  NOR2xp33_ASAP7_75t_SL U36488 ( .A(n25893), .B(n24481), .Y(n30009) );
  NOR2xp33_ASAP7_75t_SL U36489 ( .A(n22375), .B(n26574), .Y(n28132) );
  NOR2xp33_ASAP7_75t_SL U36490 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .B(
        n28824), .Y(n25488) );
  NOR2xp33_ASAP7_75t_SL U36491 ( .A(n22375), .B(n30620), .Y(n28131) );
  OR2x2_ASAP7_75t_SL U36492 ( .A(n26169), .B(n22375), .Y(n26454) );
  INVx1_ASAP7_75t_SL U36493 ( .A(n24682), .Y(n24677) );
  NOR2xp33_ASAP7_75t_SL U36494 ( .A(n25423), .B(n25422), .Y(n28823) );
  NOR2xp33_ASAP7_75t_SL U36495 ( .A(n28829), .B(n22392), .Y(n25422) );
  AOI21xp33_ASAP7_75t_SRAM U36496 ( .A1(n22375), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__7_), .B(n30006), .Y(n29935) );
  NOR2xp33_ASAP7_75t_SL U36497 ( .A(n30010), .B(n29910), .Y(n29939) );
  NOR2xp33_ASAP7_75t_SL U36498 ( .A(n25168), .B(n24476), .Y(n29910) );
  NOR2xp33_ASAP7_75t_SL U36499 ( .A(n32443), .B(n32024), .Y(n31621) );
  NOR2xp33_ASAP7_75t_SL U36500 ( .A(n29504), .B(n22375), .Y(n30006) );
  NAND3xp33_ASAP7_75t_SL U36501 ( .A(n25177), .B(n26482), .C(
        u0_0_leon3x0_p0_iu_r_E__ALUOP__2_), .Y(n29504) );
  XNOR2xp5_ASAP7_75t_SL U36502 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__6_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__6_), .Y(n25160) );
  XNOR2xp5_ASAP7_75t_SL U36503 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__1_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__1_), .Y(n25161) );
  XNOR2xp5_ASAP7_75t_SL U36504 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__5_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__5_), .Y(n25158) );
  XNOR2xp5_ASAP7_75t_SL U36505 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__7_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__7_), .Y(n25159) );
  NAND4xp25_ASAP7_75t_SL U36506 ( .A(n25157), .B(n25156), .C(n25155), .D(
        n25154), .Y(n25164) );
  XNOR2xp5_ASAP7_75t_SL U36507 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__4_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__4_), .Y(n25154) );
  XNOR2xp5_ASAP7_75t_SL U36508 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__0_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__0_), .Y(n25155) );
  XNOR2xp5_ASAP7_75t_SL U36509 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__2_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__2_), .Y(n25156) );
  XNOR2xp5_ASAP7_75t_SL U36510 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__3_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__RD__3_), .Y(n25157) );
  NAND4xp25_ASAP7_75t_SL U36511 ( .A(n25153), .B(n32141), .C(n22376), .D(
        u0_0_leon3x0_p0_iu_r_X__CTRL__WREG_), .Y(n25165) );
  NOR2xp33_ASAP7_75t_SL U36512 ( .A(n22375), .B(n25855), .Y(n29563) );
  OR2x2_ASAP7_75t_SL U36513 ( .A(n25403), .B(n25901), .Y(n30620) );
  OR2x2_ASAP7_75t_SL U36514 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUOP__2_), .Y(n28824) );
  NOR2xp33_ASAP7_75t_SL U36515 ( .A(n29675), .B(n29638), .Y(n25395) );
  NOR2xp33_ASAP7_75t_SL U36516 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__TRAP_), .B(
        n29883), .Y(n30212) );
  NAND3xp33_ASAP7_75t_SL U36517 ( .A(n25565), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__PV_), .C(n31444), .Y(n25390) );
  NOR2xp33_ASAP7_75t_SL U36518 ( .A(n25389), .B(n27194), .Y(n25565) );
  NOR2xp33_ASAP7_75t_SL U36519 ( .A(u0_0_leon3x0_p0_dco_WERR_), .B(n25388), 
        .Y(n25389) );
  NOR2xp33_ASAP7_75t_SL U36520 ( .A(u0_0_leon3x0_p0_iu_r_M__CTRL__ANNUL_), .B(
        n31813), .Y(n31960) );
  NOR2xp33_ASAP7_75t_SL U36521 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), 
        .B(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_), .Y(n25381) );
  NOR2xp33_ASAP7_75t_SL U36522 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), 
        .B(n29705), .Y(n29701) );
  NOR2xp33_ASAP7_75t_SL U36523 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[2]), .B(
        n29716), .Y(n29715) );
  NOR4xp25_ASAP7_75t_SL U36524 ( .A(n29674), .B(n25378), .C(n25377), .D(n25376), .Y(n25391) );
  NOR2xp33_ASAP7_75t_SL U36525 ( .A(n4752), .B(
        u0_0_leon3x0_p0_iu_r_W__S__PIL__1_), .Y(n25372) );
  NOR3xp33_ASAP7_75t_SL U36526 ( .A(n25370), .B(n4752), .C(n4774), .Y(n25375)
         );
  NOR2xp33_ASAP7_75t_SL U36527 ( .A(n29704), .B(n29472), .Y(n29721) );
  AOI21xp33_ASAP7_75t_SRAM U36528 ( .A1(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__21_), .A2(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_), .B(n25366), .Y(n25368) );
  AND2x2_ASAP7_75t_SL U36529 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), 
        .B(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__21_), .Y(n29706) );
  NOR2xp33_ASAP7_75t_SL U36530 ( .A(n25364), .B(n25363), .Y(n30157) );
  AND2x2_ASAP7_75t_SL U36531 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_), 
        .B(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_), .Y(n25382) );
  NOR2xp33_ASAP7_75t_SL U36532 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__20_), 
        .B(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), .Y(n29702) );
  NOR2xp33_ASAP7_75t_SL U36533 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[3]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[4]), .Y(n29469) );
  NOR2xp33_ASAP7_75t_SL U36534 ( .A(n25361), .B(n25360), .Y(n29884) );
  INVx1_ASAP7_75t_SL U36535 ( .A(u0_0_leon3x0_p0_iu_r_M__CASA_), .Y(n25080) );
  NOR3xp33_ASAP7_75t_SL U36536 ( .A(n25351), .B(u0_0_leon3x0_p0_dci[26]), .C(
        u0_0_leon3x0_p0_dci[32]), .Y(n25352) );
  NOR2xp33_ASAP7_75t_SL U36537 ( .A(n25151), .B(n24705), .Y(n32140) );
  NOR2xp33_ASAP7_75t_SL U36538 ( .A(u0_0_leon3x0_p0_dci[18]), .B(
        u0_0_leon3x0_p0_dci[22]), .Y(n25349) );
  NOR2xp33_ASAP7_75t_SL U36539 ( .A(u0_0_leon3x0_p0_dci[20]), .B(
        u0_0_leon3x0_p0_dci[19]), .Y(n25350) );
  NAND2xp33_ASAP7_75t_SRAM U36540 ( .A(n25106), .B(n25105), .Y(add_x_735_A_19_) );
  NOR2xp33_ASAP7_75t_SL U36541 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[30]), .Y(
        n28479) );
  NOR2xp33_ASAP7_75t_SL U36542 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[29]), .Y(
        n27057) );
  NOR2xp33_ASAP7_75t_SL U36543 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[32]), .Y(
        n26381) );
  NOR2xp33_ASAP7_75t_SL U36544 ( .A(n25338), .B(n31452), .Y(n25513) );
  NOR2xp33_ASAP7_75t_SL U36545 ( .A(n31594), .B(n25399), .Y(n32289) );
  INVx1_ASAP7_75t_SL U36546 ( .A(n3071), .Y(n32250) );
  NOR2xp33_ASAP7_75t_SL U36547 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_STPEND_), 
        .B(n32443), .Y(n31605) );
  NOR2xp33_ASAP7_75t_SL U36548 ( .A(n32237), .B(n31565), .Y(n31462) );
  NOR2xp33_ASAP7_75t_SL U36549 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_), .B(n25512), .Y(n32237) );
  NAND2xp33_ASAP7_75t_SRAM U36550 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_), .B(n3134), .Y(n25511) );
  NOR2xp33_ASAP7_75t_SL U36551 ( .A(n31455), .B(n31452), .Y(n31572) );
  NOR2xp33_ASAP7_75t_SL U36552 ( .A(n32197), .B(n31306), .Y(n31452) );
  INVx1_ASAP7_75t_SL U36553 ( .A(n4082), .Y(n32197) );
  INVx1_ASAP7_75t_SL U36554 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_), 
        .Y(n31594) );
  NOR2xp33_ASAP7_75t_SL U36555 ( .A(n22380), .B(n25521), .Y(n25515) );
  INVx1_ASAP7_75t_SL U36556 ( .A(n3899), .Y(n32037) );
  INVx1_ASAP7_75t_SL U36557 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_STPEND_), .Y(
        n31455) );
  NOR2xp33_ASAP7_75t_SL U36558 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[25]), .Y(
        n26703) );
  NOR2xp33_ASAP7_75t_SL U36559 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[24]), .Y(
        n26563) );
  NOR2xp33_ASAP7_75t_SL U36560 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[19]), .Y(
        n27111) );
  NOR2xp33_ASAP7_75t_SL U36561 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[20]), .Y(
        n27138) );
  XNOR2xp5_ASAP7_75t_SL U36562 ( .A(u0_0_leon3x0_p0_iu_r_E__INVOP2_), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__3_), .Y(n25085) );
  XNOR2xp5_ASAP7_75t_SL U36563 ( .A(u0_0_leon3x0_p0_iu_r_E__INVOP2_), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__2_), .Y(n25083) );
  NOR2xp33_ASAP7_75t_SL U36564 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[16]), .Y(
        n26302) );
  NOR2xp33_ASAP7_75t_SL U36565 ( .A(n31813), .B(n26199), .Y(n31828) );
  AND2x2_ASAP7_75t_SL U36566 ( .A(n23229), .B(n31833), .Y(n31996) );
  NOR2xp33_ASAP7_75t_SL U36567 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), 
        .B(n24879), .Y(n25221) );
  NOR2xp33_ASAP7_75t_SL U36568 ( .A(n24854), .B(n32082), .Y(n32055) );
  NOR2xp33_ASAP7_75t_SL U36569 ( .A(n24847), .B(n29206), .Y(n24848) );
  NOR2xp33_ASAP7_75t_SL U36570 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), 
        .B(n32097), .Y(n24846) );
  NOR2xp33_ASAP7_75t_SL U36571 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__30_), 
        .B(n31958), .Y(n25230) );
  NOR2xp33_ASAP7_75t_SL U36572 ( .A(n31537), .B(n30956), .Y(n25231) );
  NOR2xp33_ASAP7_75t_SL U36573 ( .A(n24843), .B(n24842), .Y(n30940) );
  AOI21xp33_ASAP7_75t_SRAM U36574 ( .A1(n24882), .A2(n32084), .B(n24816), .Y(
        n24833) );
  NOR2xp33_ASAP7_75t_SL U36575 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__5_), .B(
        n32165), .Y(n24828) );
  XNOR2xp5_ASAP7_75t_SL U36576 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_), .Y(n24788) );
  NOR2xp33_ASAP7_75t_SL U36577 ( .A(n24785), .B(n24784), .Y(n32180) );
  XNOR2xp5_ASAP7_75t_SL U36578 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_), .Y(n24785) );
  NOR2xp33_ASAP7_75t_SL U36579 ( .A(n26842), .B(n24782), .Y(n24805) );
  NOR2xp33_ASAP7_75t_SL U36580 ( .A(n24780), .B(n24779), .Y(n24809) );
  NOR2xp33_ASAP7_75t_SL U36581 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__18_), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__17_), .Y(n24776) );
  NOR2xp33_ASAP7_75t_SL U36582 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__28_), .Y(n31380) );
  NOR2xp33_ASAP7_75t_SL U36583 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__1_), .B(
        n24780), .Y(n24778) );
  NOR2xp33_ASAP7_75t_SL U36584 ( .A(n24807), .B(n24774), .Y(n24780) );
  NOR2xp33_ASAP7_75t_SL U36585 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__1_), .B(
        n24763), .Y(n24766) );
  NOR2xp33_ASAP7_75t_SL U36586 ( .A(n24755), .B(n24754), .Y(n24797) );
  NOR2xp33_ASAP7_75t_SL U36587 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(
        n30791), .Y(n26855) );
  AND2x2_ASAP7_75t_SL U36588 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(
        DP_OP_1196_128_7433_n456), .Y(n24763) );
  NOR2xp33_ASAP7_75t_SL U36589 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__1_), .B(
        n32171), .Y(n24747) );
  NOR2xp33_ASAP7_75t_SL U36590 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), 
        .B(n32083), .Y(n24858) );
  NOR2xp33_ASAP7_75t_SL U36591 ( .A(n24887), .B(n25218), .Y(n24888) );
  AOI211xp5_ASAP7_75t_SL U36592 ( .A1(n18799), .A2(n31657), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), .C(n24912), .Y(n25218) );
  NOR2xp33_ASAP7_75t_SL U36593 ( .A(n24845), .B(n32081), .Y(n32050) );
  NOR2xp33_ASAP7_75t_SL U36594 ( .A(u0_0_leon3x0_p0_iu_r_D__ANNUL_), .B(n32097), .Y(n32048) );
  NOR2xp33_ASAP7_75t_SL U36595 ( .A(n24886), .B(n31655), .Y(n31657) );
  NOR2xp33_ASAP7_75t_SL U36596 ( .A(n24885), .B(n24903), .Y(n24906) );
  NOR2xp33_ASAP7_75t_SL U36597 ( .A(n3727), .B(n31658), .Y(n31420) );
  INVx1_ASAP7_75t_SL U36598 ( .A(n4325), .Y(n31656) );
  NOR2xp33_ASAP7_75t_SL U36599 ( .A(u0_0_leon3x0_p0_iu_r_D__ANNUL_), .B(n26818), .Y(n24882) );
  NOR2xp33_ASAP7_75t_SL U36600 ( .A(n31813), .B(n26197), .Y(n26203) );
  NAND4xp25_ASAP7_75t_SL U36601 ( .A(n26196), .B(n32016), .C(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__31_), .D(n31441), .Y(n31884) );
  NOR2xp33_ASAP7_75t_SL U36602 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_), 
        .B(n31964), .Y(n32016) );
  NOR3xp33_ASAP7_75t_SL U36603 ( .A(n26195), .B(
        u0_0_leon3x0_p0_iu_r_E__CTRL__ANNUL_), .C(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__30_), .Y(n26196) );
  INVx1_ASAP7_75t_SL U36604 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__ANNUL_), .Y(
        n30115) );
  AND2x2_ASAP7_75t_SL U36605 ( .A(n3730), .B(n3704), .Y(n26757) );
  OR2x2_ASAP7_75t_SL U36606 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__TRAP_), .B(
        u0_0_leon3x0_p0_iu_r_X__MEXC_), .Y(n26352) );
  NOR2xp33_ASAP7_75t_SL U36607 ( .A(n22380), .B(n25607), .Y(n24736) );
  INVx1_ASAP7_75t_SL U36608 ( .A(n3730), .Y(n25607) );
  NOR2xp33_ASAP7_75t_SL U36609 ( .A(u0_0_leon3x0_p0_iu_r_D__ANNUL_), .B(n32091), .Y(n26192) );
  NOR2xp33_ASAP7_75t_SL U36610 ( .A(n25937), .B(n24739), .Y(n26190) );
  NOR2xp33_ASAP7_75t_SL U36611 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__24_), 
        .B(n18819), .Y(n32052) );
  NOR2xp33_ASAP7_75t_SL U36612 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__25_), 
        .B(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__26_), .Y(n24844) );
  NOR3xp33_ASAP7_75t_SL U36613 ( .A(n24727), .B(u0_0_leon3x0_p0_iu_de_icc_2_), 
        .C(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_), .Y(n24728) );
  NOR2xp33_ASAP7_75t_SL U36614 ( .A(u0_0_leon3x0_p0_iu_r_E__CTRL__ANNUL_), .B(
        n25453), .Y(n24734) );
  NOR2xp33_ASAP7_75t_SL U36615 ( .A(u0_0_leon3x0_p0_iu_de_icc_3_), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__25_), .Y(n24711) );
  NAND2xp33_ASAP7_75t_SRAM U36616 ( .A(n25306), .B(n24672), .Y(n25305) );
  OR2x2_ASAP7_75t_SL U36617 ( .A(n24544), .B(n24431), .Y(
        u0_0_leon3x0_p0_muli[38]) );
  NOR2xp33_ASAP7_75t_SL U36618 ( .A(n25095), .B(n24686), .Y(n24544) );
  NOR2xp33_ASAP7_75t_SL U36619 ( .A(u0_0_leon3x0_p0_iu_r_A__TICC_), .B(
        u0_0_leon3x0_p0_iu_r_A__WUNF_), .Y(n29669) );
  AND2x2_ASAP7_75t_SL U36620 ( .A(n26357), .B(n26356), .Y(n24511) );
  NOR2xp33_ASAP7_75t_SL U36621 ( .A(uart1_r_RCNT__5_), .B(n33065), .Y(n25972)
         );
  INVx1_ASAP7_75t_SL U36622 ( .A(uart1_v_RXDB__1_), .Y(n33065) );
  NAND2xp5_ASAP7_75t_SL U36623 ( .A(n26072), .B(n28231), .Y(n31057) );
  AOI21xp33_ASAP7_75t_SRAM U36624 ( .A1(n24582), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__19_), .B(n28887), .Y(n25764) );
  NOR2xp33_ASAP7_75t_SL U36625 ( .A(n25019), .B(n25020), .Y(n31259) );
  NOR2xp33_ASAP7_75t_SL U36626 ( .A(u0_0_leon3x0_p0_iu_r_M__WCWP_), .B(n31428), 
        .Y(n26775) );
  NOR2xp33_ASAP7_75t_SL U36627 ( .A(n5061), .B(n1626), .Y(timer0_N84) );
  NOR2xp33_ASAP7_75t_SL U36628 ( .A(n5061), .B(n1741), .Y(timer0_N83) );
  NOR2xp33_ASAP7_75t_SL U36629 ( .A(n26465), .B(timer0_N60), .Y(n26466) );
  O2A1O1Ixp5_ASAP7_75t_SL U36630 ( .A1(n31621), .A2(n31610), .B(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_RBURST_), .C(n32273), .Y(n31611) );
  INVxp33_ASAP7_75t_SRAM U36631 ( .A(n26169), .Y(n25626) );
  NAND2xp33_ASAP7_75t_SRAM U36632 ( .A(n25102), .B(n25101), .Y(add_x_735_A_29_) );
  NOR2xp33_ASAP7_75t_SL U36633 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[31]), .Y(
        n26416) );
  INVxp33_ASAP7_75t_SRAM U36634 ( .A(n3550), .Y(rf_addr_b[7]) );
  INVxp33_ASAP7_75t_SRAM U36635 ( .A(n2772), .Y(rf_addr_a[5]) );
  NOR2xp33_ASAP7_75t_SL U36636 ( .A(n29669), .B(n29668), .Y(n29673) );
  INVx1_ASAP7_75t_SL U36637 ( .A(n29949), .Y(n28030) );
  NOR2xp33_ASAP7_75t_SL U36638 ( .A(uart1_r_RCNT__0_), .B(uart1_r_RCNT__3_), 
        .Y(n25983) );
  O2A1O1Ixp5_ASAP7_75t_SL U36639 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__4_), .A2(
        n30007), .B(n28842), .C(n28841), .Y(n28857) );
  AOI22xp33_ASAP7_75t_SRAM U36640 ( .A1(u0_0_leon3x0_p0_iu_de_icc_0_), .A2(
        n30621), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__8_), .B2(n28779), .Y(
        n26995) );
  AOI22xp33_ASAP7_75t_SRAM U36641 ( .A1(n29603), .A2(n28499), .B1(n28742), 
        .B2(n27077), .Y(n27081) );
  OAI22xp33_ASAP7_75t_SRAM U36642 ( .A1(n31353), .A2(n31469), .B1(n32461), 
        .B2(n31466), .Y(n31355) );
  AOI22xp33_ASAP7_75t_SRAM U36643 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__22_), 
        .A2(u0_0_leon3x0_p0_iu_r_E__JMPL_), .B1(u0_0_leon3x0_p0_iu_de_icc_2_), 
        .B2(n30621), .Y(n28492) );
  AOI22xp33_ASAP7_75t_SRAM U36644 ( .A1(u0_0_leon3x0_p0_iu_de_icc_3_), .A2(
        n30621), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__11_), .B2(n28779), .Y(
        n26419) );
  NOR2xp33_ASAP7_75t_SL U36645 ( .A(n26186), .B(n26188), .Y(n24430) );
  NOR2xp33_ASAP7_75t_SL U36646 ( .A(n22427), .B(n31428), .Y(n31427) );
  NOR2xp33_ASAP7_75t_SL U36647 ( .A(n31656), .B(n22422), .Y(n31672) );
  NOR2xp33_ASAP7_75t_SL U36648 ( .A(n5061), .B(n4635), .Y(timer0_N76) );
  INVxp33_ASAP7_75t_SRAM U36649 ( .A(n3552), .Y(rf_addr_b[3]) );
  INVxp33_ASAP7_75t_SRAM U36650 ( .A(n4169), .Y(rf_addr_a[0]) );
  INVxp33_ASAP7_75t_SRAM U36651 ( .A(n3758), .Y(rf_addr_a[1]) );
  INVxp33_ASAP7_75t_SRAM U36652 ( .A(n2774), .Y(rf_addr_a[6]) );
  NOR2xp33_ASAP7_75t_SL U36653 ( .A(n32076), .B(n31987), .Y(n24584) );
  NOR2xp33_ASAP7_75t_SL U36654 ( .A(n32076), .B(n31987), .Y(n31986) );
  AOI22xp33_ASAP7_75t_SRAM U36655 ( .A1(sr1_r_MCFG2__RAMBANKSZ__0_), .A2(
        n31250), .B1(sr1_r_MCFG1__ROMWIDTH__1_), .B2(n31235), .Y(n30142) );
  AOI22xp33_ASAP7_75t_SRAM U36656 ( .A1(sr1_r_MCFG2__RAMRWS__1_), .A2(n31250), 
        .B1(n31235), .B2(sr1_r_MCFG1__ROMRWS__1_), .Y(n27480) );
  AOI22xp33_ASAP7_75t_SRAM U36657 ( .A1(sr1_r_MCFG2__RAMWIDTH__1_), .A2(n31250), .B1(n31235), .B2(sr1_r_MCFG1__ROMWWS__1_), .Y(n30078) );
  NOR2xp33_ASAP7_75t_SL U36658 ( .A(n26073), .B(n29558), .Y(n26074) );
  NOR2xp33_ASAP7_75t_SL U36659 ( .A(n2924), .B(n33049), .Y(n32750) );
  AOI31xp33_ASAP7_75t_SL U36660 ( .A1(n25884), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__29_), .A3(n24855), .B(n31814), .Y(
        n24735) );
  NOR2xp33_ASAP7_75t_SL U36661 ( .A(n32063), .B(n18798), .Y(n31814) );
  INVx1_ASAP7_75t_SL U36662 ( .A(n24681), .Y(n24658) );
  NOR2xp33_ASAP7_75t_SL U36663 ( .A(n28110), .B(n26469), .Y(n26471) );
  NOR2xp33_ASAP7_75t_SL U36664 ( .A(n5061), .B(n4354), .Y(timer0_N73) );
  NOR2xp33_ASAP7_75t_SL U36665 ( .A(n5061), .B(n1771), .Y(timer0_N75) );
  NOR2xp33_ASAP7_75t_SL U36666 ( .A(n5061), .B(n4032), .Y(timer0_N74) );
  NOR2xp33_ASAP7_75t_SL U36667 ( .A(n5061), .B(n1792), .Y(timer0_N82) );
  NAND4xp25_ASAP7_75t_SL U36668 ( .A(n30159), .B(n30158), .C(n30157), .D(
        n30687), .Y(n31546) );
  NOR2xp33_ASAP7_75t_SL U36669 ( .A(n30010), .B(n28823), .Y(n25874) );
  XNOR2xp5_ASAP7_75t_SL U36670 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__3_), .B(
        DP_OP_1196_128_7433_n455), .Y(n24750) );
  NOR2xp33_ASAP7_75t_SL U36671 ( .A(n29340), .B(n29341), .Y(n29344) );
  NOR2xp33_ASAP7_75t_SL U36672 ( .A(n29334), .B(n29335), .Y(n29338) );
  AOI22xp33_ASAP7_75t_SRAM U36673 ( .A1(irqctrl0_r_ILEVEL__12_), .A2(n31248), 
        .B1(irqctrl0_r_IPEND__12_), .B2(n31247), .Y(n29856) );
  AOI22xp33_ASAP7_75t_SRAM U36674 ( .A1(irqctrl0_r_ILEVEL__9_), .A2(n31248), 
        .B1(uart1_r_TFIFOIRQEN_), .B2(n31950), .Y(n30144) );
  NOR2xp33_ASAP7_75t_SL U36675 ( .A(uart1_uarto_TXEN_), .B(uart1_uarto_RXEN_), 
        .Y(n28167) );
  AOI22xp33_ASAP7_75t_SRAM U36676 ( .A1(irqctrl0_r_ILEVEL__1_), .A2(n31248), 
        .B1(irqctrl0_r_IPEND__1_), .B2(n31247), .Y(n27466) );
  AOI22xp33_ASAP7_75t_SRAM U36677 ( .A1(irqctrl0_r_ILEVEL__5_), .A2(n31248), 
        .B1(irqctrl0_r_IPEND__5_), .B2(n31247), .Y(n30076) );
  AOI22xp33_ASAP7_75t_SRAM U36678 ( .A1(u0_0_leon3x0_p0_dci[0]), .A2(n30621), 
        .B1(n29307), .B2(n28779), .Y(n28781) );
  AOI21xp33_ASAP7_75t_SRAM U36679 ( .A1(n29603), .A2(n28763), .B(n26276), .Y(
        n26283) );
  AOI22xp33_ASAP7_75t_SRAM U36680 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__PS_), .A2(
        n30621), .B1(irqo[1]), .B2(n28779), .Y(n26267) );
  AOI211xp5_ASAP7_75t_SL U36681 ( .A1(n28411), .A2(n29919), .B(n26375), .C(
        n30578), .Y(n3011) );
  OAI22xp33_ASAP7_75t_SRAM U36682 ( .A1(n25897), .A2(n29595), .B1(n30230), 
        .B2(n29594), .Y(n25898) );
  NAND2xp33_ASAP7_75t_SRAM U36683 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__29_), 
        .B(n29589), .Y(n25895) );
  NOR2xp33_ASAP7_75t_SL U36684 ( .A(n18860), .B(n4385), .Y(timer0_N70) );
  NOR2xp33_ASAP7_75t_SL U36685 ( .A(n5061), .B(n2233), .Y(timer0_N80) );
  NOR2xp33_ASAP7_75t_SL U36686 ( .A(n28769), .B(u0_0_leon3x0_p0_muli[35]), .Y(
        n25891) );
  NOR2xp33_ASAP7_75t_SL U36687 ( .A(n22380), .B(n3730), .Y(n26198) );
  INVxp33_ASAP7_75t_SRAM U36688 ( .A(n2463), .Y(rf_ce_b) );
  INVxp33_ASAP7_75t_SRAM U36689 ( .A(n3501), .Y(rf_addr_a[2]) );
  INVxp33_ASAP7_75t_SRAM U36690 ( .A(n2567), .Y(rf_addr_a[3]) );
  NOR2xp33_ASAP7_75t_SL U36691 ( .A(n2929), .B(n29743), .Y(n29376) );
  NOR2xp33_ASAP7_75t_SL U36692 ( .A(n28920), .B(n28854), .Y(n31015) );
  AOI211xp5_ASAP7_75t_SL U36693 ( .A1(n28411), .A2(n30024), .B(n25418), .C(
        n30578), .Y(n3004) );
  AOI211xp5_ASAP7_75t_SL U36694 ( .A1(n28411), .A2(n30968), .B(n26347), .C(
        n30578), .Y(n3008) );
  AOI211xp5_ASAP7_75t_SL U36695 ( .A1(n28411), .A2(n30563), .B(n26225), .C(
        n30578), .Y(n3012) );
  AOI211xp5_ASAP7_75t_SL U36696 ( .A1(n28411), .A2(n31005), .B(n25718), .C(
        n30578), .Y(n3017) );
  AOI211xp5_ASAP7_75t_SL U36697 ( .A1(n28411), .A2(n31480), .B(n26968), .C(
        n30578), .Y(n3016) );
  NAND4xp25_ASAP7_75t_SL U36698 ( .A(n22413), .B(n25057), .C(n25056), .D(
        n25055), .Y(n25060) );
  AND2x2_ASAP7_75t_SL U36699 ( .A(n24634), .B(n28995), .Y(n30621) );
  NAND4xp25_ASAP7_75t_SL U36700 ( .A(n25482), .B(n24472), .C(n25481), .D(
        n25480), .Y(n28440) );
  NOR2xp33_ASAP7_75t_SL U36701 ( .A(n18819), .B(n25225), .Y(n26868) );
  INVx1_ASAP7_75t_SL U36702 ( .A(n24681), .Y(n24649) );
  O2A1O1Ixp5_ASAP7_75t_SL U36703 ( .A1(n31388), .A2(n32049), .B(n31387), .C(
        n31386), .Y(n3158) );
  O2A1O1Ixp5_ASAP7_75t_SL U36704 ( .A1(n31598), .A2(n31597), .B(n31596), .C(
        n31595), .Y(n3070) );
  NOR2xp33_ASAP7_75t_SL U36705 ( .A(n18860), .B(n4414), .Y(timer0_N68) );
  NOR2xp33_ASAP7_75t_SL U36706 ( .A(n18860), .B(n4363), .Y(timer0_N72) );
  NOR2xp33_ASAP7_75t_SL U36707 ( .A(n18860), .B(n4497), .Y(timer0_N71) );
  NOR2xp33_ASAP7_75t_SL U36708 ( .A(n18860), .B(n4573), .Y(timer0_N69) );
  NOR2xp33_ASAP7_75t_SL U36709 ( .A(n18860), .B(n2271), .Y(timer0_N67) );
  NOR2xp33_ASAP7_75t_SL U36710 ( .A(n18860), .B(n4624), .Y(timer0_N66) );
  NOR2xp33_ASAP7_75t_SL U36711 ( .A(n18864), .B(n4770), .Y(timer0_N60) );
  NOR3xp33_ASAP7_75t_SL U36712 ( .A(n25380), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__19_), .C(n32713), .Y(n25385) );
  AOI22xp33_ASAP7_75t_SRAM U36713 ( .A1(dc_q[12]), .A2(n32344), .B1(n32621), 
        .B2(n24643), .Y(n32338) );
  AOI22xp33_ASAP7_75t_SRAM U36714 ( .A1(dc_q[9]), .A2(n32344), .B1(n32615), 
        .B2(n24643), .Y(n32327) );
  AOI22xp33_ASAP7_75t_SRAM U36715 ( .A1(n31849), .A2(n31848), .B1(
        sr1_r_MCFG1__IOWS__1_), .B2(n32003), .Y(n31850) );
  OR2x2_ASAP7_75t_SL U36716 ( .A(n25937), .B(n22378), .Y(n24495) );
  INVx1_ASAP7_75t_SL U36717 ( .A(n28180), .Y(n29369) );
  NOR2xp33_ASAP7_75t_SL U36718 ( .A(n27321), .B(n27328), .Y(n27325) );
  NOR2xp33_ASAP7_75t_SL U36719 ( .A(n31038), .B(n31047), .Y(n3022) );
  NOR4xp25_ASAP7_75t_SL U36720 ( .A(n25445), .B(n30018), .C(n29915), .D(n31364), .Y(n31043) );
  O2A1O1Ixp5_ASAP7_75t_SL U36721 ( .A1(n25615), .A2(n24484), .B(n31001), .C(
        n25614), .Y(n30566) );
  NOR2xp33_ASAP7_75t_SL U36722 ( .A(n25438), .B(n25069), .Y(n25070) );
  NOR2xp33_ASAP7_75t_SL U36723 ( .A(n25058), .B(n31001), .Y(n25059) );
  O2A1O1Ixp5_ASAP7_75t_SL U36724 ( .A1(u0_0_leon3x0_p0_iu_r_X__DCI__SIZE__1_), 
        .A2(n30020), .B(n30019), .C(n30018), .Y(n30023) );
  NOR2xp33_ASAP7_75t_SL U36725 ( .A(n25178), .B(n26269), .Y(n28995) );
  O2A1O1Ixp5_ASAP7_75t_SL U36726 ( .A1(n25912), .A2(n28975), .B(n25150), .C(
        n27208), .Y(n25186) );
  NAND2xp33_ASAP7_75t_SRAM U36727 ( .A(n31379), .B(n25221), .Y(n25222) );
  NAND2xp33_ASAP7_75t_SRAM U36728 ( .A(n3880), .B(n24684), .Y(n31891) );
  NOR2xp33_ASAP7_75t_SL U36729 ( .A(n18872), .B(n4741), .Y(timer0_N61) );
  NOR2xp33_ASAP7_75t_SL U36730 ( .A(n18864), .B(n4669), .Y(timer0_N62) );
  NOR2xp33_ASAP7_75t_SL U36731 ( .A(n18864), .B(n4531), .Y(timer0_N64) );
  NOR2xp33_ASAP7_75t_SL U36732 ( .A(n18864), .B(n1775), .Y(timer0_N63) );
  AOI31xp33_ASAP7_75t_SL U36733 ( .A1(n30194), .A2(u0_0_leon3x0_p0_dci[38]), 
        .A3(n30193), .B(n30192), .Y(n30199) );
  INVx1_ASAP7_75t_SL U36734 ( .A(n31813), .Y(n30503) );
  AOI22xp33_ASAP7_75t_SRAM U36735 ( .A1(n32269), .A2(n32268), .B1(n3054), .B2(
        n33067), .Y(dt_address[6]) );
  AOI21xp33_ASAP7_75t_SRAM U36736 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__29_), 
        .A2(n32239), .B(n33067), .Y(n32230) );
  AOI21xp33_ASAP7_75t_SRAM U36737 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__27_), 
        .A2(n32239), .B(n33067), .Y(n32227) );
  AOI21xp33_ASAP7_75t_SRAM U36738 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__26_), 
        .A2(n32239), .B(n33067), .Y(n32225) );
  AOI21xp33_ASAP7_75t_SRAM U36739 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__25_), 
        .A2(n32239), .B(n33067), .Y(n32223) );
  AOI21xp33_ASAP7_75t_SRAM U36740 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__24_), 
        .A2(n32239), .B(n33067), .Y(n32221) );
  INVxp33_ASAP7_75t_SRAM U36741 ( .A(n28189), .Y(n26089) );
  AOI22xp33_ASAP7_75t_SRAM U36742 ( .A1(timer0_vtimers_1__RELOAD__0_), .A2(
        n31956), .B1(n28089), .B2(n30789), .Y(n28090) );
  OR2x2_ASAP7_75t_SL U36743 ( .A(n24695), .B(n27292), .Y(n29652) );
  NOR2xp33_ASAP7_75t_SL U36744 ( .A(n26023), .B(n26021), .Y(n26036) );
  AOI21xp33_ASAP7_75t_SRAM U36745 ( .A1(n30621), .A2(
        u0_0_leon3x0_p0_iu_r_W__S__PIL__1_), .B(n27114), .Y(n27115) );
  O2A1O1Ixp5_ASAP7_75t_SL U36746 ( .A1(n30651), .A2(n30489), .B(n29016), .C(
        n29015), .Y(n2701) );
  AOI22xp33_ASAP7_75t_SRAM U36747 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__26_), 
        .A2(n24582), .B1(u0_0_leon3x0_p0_iu_r_W__S__TBA__14_), .B2(n28779), 
        .Y(n25485) );
  O2A1O1Ixp5_ASAP7_75t_SL U36748 ( .A1(n29790), .A2(n29791), .B(n31054), .C(
        n26443), .Y(n4418) );
  AOI22xp33_ASAP7_75t_SRAM U36749 ( .A1(n28835), .A2(n30249), .B1(
        u0_0_leon3x0_p0_divi[56]), .B2(n28782), .Y(n28428) );
  NOR2xp33_ASAP7_75t_SL U36750 ( .A(n26737), .B(n26736), .Y(n27017) );
  NOR2xp33_ASAP7_75t_SL U36751 ( .A(n32823), .B(n32711), .Y(n32743) );
  NOR2xp33_ASAP7_75t_SL U36752 ( .A(n32710), .B(n32709), .Y(n32823) );
  NOR2xp33_ASAP7_75t_SL U36753 ( .A(n31673), .B(n26188), .Y(n31674) );
  NAND4xp25_ASAP7_75t_SL U36754 ( .A(n31914), .B(n31913), .C(n31912), .D(
        n31911), .Y(n31915) );
  NAND4xp25_ASAP7_75t_SL U36755 ( .A(n31910), .B(n31909), .C(n31908), .D(
        n31907), .Y(n31916) );
  AND2x2_ASAP7_75t_SL U36756 ( .A(n31420), .B(n22379), .Y(n24517) );
  NAND2xp33_ASAP7_75t_SRAM U36757 ( .A(n24231), .B(n28402), .Y(n26537) );
  AOI211xp5_ASAP7_75t_SL U36758 ( .A1(n28402), .A2(n22436), .B(n26219), .C(
        n26218), .Y(n32383) );
  NAND2xp33_ASAP7_75t_SRAM U36759 ( .A(n18530), .B(n28402), .Y(n26457) );
  NOR2xp33_ASAP7_75t_SL U36760 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__5_), .B(
        n32184), .Y(n24841) );
  NAND2xp33_ASAP7_75t_SRAM U36761 ( .A(n24688), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__0_), .Y(n31405) );
  NAND2xp33_ASAP7_75t_SRAM U36762 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__21_), 
        .B(n24688), .Y(n27056) );
  AOI22xp33_ASAP7_75t_SRAM U36763 ( .A1(dc_q[15]), .A2(n32344), .B1(n32627), 
        .B2(n24643), .Y(n32347) );
  AOI22xp33_ASAP7_75t_SRAM U36764 ( .A1(u0_0_leon3x0_p0_c0mmu_mmudci[2]), .A2(
        n32448), .B1(n32437), .B2(n32447), .Y(n32440) );
  OAI22xp33_ASAP7_75t_SRAM U36765 ( .A1(n32494), .A2(n32565), .B1(n32593), 
        .B2(n32606), .Y(it_data[4]) );
  OAI22xp33_ASAP7_75t_SRAM U36766 ( .A1(n32622), .A2(n32543), .B1(n32525), 
        .B2(n32542), .Y(it_data[8]) );
  OAI22xp33_ASAP7_75t_SRAM U36767 ( .A1(n32638), .A2(n32543), .B1(n32542), 
        .B2(n32535), .Y(it_data[16]) );
  INVxp33_ASAP7_75t_SRAM U36768 ( .A(n32273), .Y(n32278) );
  AOI22xp33_ASAP7_75t_SRAM U36769 ( .A1(n32260), .A2(n32259), .B1(n33067), 
        .B2(n32258), .Y(dt_address[0]) );
  INVxp33_ASAP7_75t_SRAM U36770 ( .A(n32292), .Y(n32251) );
  OAI21xp33_ASAP7_75t_SRAM U36771 ( .A1(n32217), .A2(n32628), .B(n32208), .Y(
        dt_data[11]) );
  OAI21xp33_ASAP7_75t_SRAM U36772 ( .A1(n32217), .A2(n32626), .B(n32207), .Y(
        dt_data[10]) );
  OAI21xp33_ASAP7_75t_SRAM U36773 ( .A1(n32217), .A2(n32624), .B(n32206), .Y(
        dt_data[9]) );
  OAI21xp33_ASAP7_75t_SRAM U36774 ( .A1(n32622), .A2(n32217), .B(n32205), .Y(
        dt_data[8]) );
  OAI21xp33_ASAP7_75t_SRAM U36775 ( .A1(n3067), .A2(n14803), .B(n32672), .Y(
        ic_address[0]) );
  INVxp33_ASAP7_75t_SRAM U36776 ( .A(n14803), .Y(n32694) );
  OAI22xp33_ASAP7_75t_SRAM U36777 ( .A1(n32642), .A2(n32543), .B1(n32542), 
        .B2(n32538), .Y(it_data[18]) );
  OAI22xp33_ASAP7_75t_SRAM U36778 ( .A1(n32644), .A2(n32543), .B1(n32542), 
        .B2(n32541), .Y(it_data[19]) );
  OAI22xp33_ASAP7_75t_SRAM U36779 ( .A1(apbi[2]), .A2(n29745), .B1(n29568), 
        .B2(n29376), .Y(n29382) );
  OAI21xp33_ASAP7_75t_SRAM U36780 ( .A1(n30073), .A2(n29516), .B(n24694), .Y(
        n25869) );
  OAI21xp33_ASAP7_75t_SRAM U36781 ( .A1(n31197), .A2(n29516), .B(n24694), .Y(
        n25866) );
  OAI21xp33_ASAP7_75t_SRAM U36782 ( .A1(n27493), .A2(n29516), .B(n24694), .Y(
        n26135) );
  OAI21xp33_ASAP7_75t_SRAM U36783 ( .A1(n30780), .A2(n29516), .B(n24694), .Y(
        n25880) );
  OAI21xp33_ASAP7_75t_SRAM U36784 ( .A1(n29568), .A2(n29516), .B(n24694), .Y(
        n29520) );
  OAI21xp33_ASAP7_75t_SRAM U36785 ( .A1(n29510), .A2(n29516), .B(n24694), .Y(
        n29513) );
  AOI22xp33_ASAP7_75t_SRAM U36786 ( .A1(n31849), .A2(n31529), .B1(
        sr1_r_MCFG1__IOWS__0_), .B2(n32003), .Y(n31530) );
  AOI21xp33_ASAP7_75t_SRAM U36787 ( .A1(timer0_vtimers_1__ENABLE_), .A2(n30790), .B(n28088), .Y(n28091) );
  INVx1_ASAP7_75t_SL U36788 ( .A(apb0_r_CFGSEL_), .Y(n31954) );
  OAI22xp33_ASAP7_75t_SRAM U36789 ( .A1(n31197), .A2(n29652), .B1(n29312), 
        .B2(n29650), .Y(n29310) );
  NOR2xp33_ASAP7_75t_SL U36790 ( .A(n25638), .B(n25954), .Y(n31249) );
  NOR2xp33_ASAP7_75t_SL U36791 ( .A(n31848), .B(n26658), .Y(n27459) );
  INVxp33_ASAP7_75t_SRAM U36792 ( .A(n31057), .Y(n29358) );
  AOI21xp33_ASAP7_75t_SRAM U36793 ( .A1(n28888), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__6_), .B(n28887), .Y(n26266) );
  AOI211xp5_ASAP7_75t_SL U36794 ( .A1(n29881), .A2(n29645), .B(n29644), .C(
        n29643), .Y(n3326) );
  NOR2xp33_ASAP7_75t_SL U36795 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[25]), .B(
        n22379), .Y(n28449) );
  OAI21xp33_ASAP7_75t_SRAM U36796 ( .A1(n28730), .A2(n28934), .B(n30616), .Y(
        n28731) );
  AOI22xp33_ASAP7_75t_SRAM U36797 ( .A1(n28821), .A2(u0_0_leon3x0_p0_divi[3]), 
        .B1(u0_0_leon3x0_p0_iu_r_W__S__WIM__4_), .B2(n30611), .Y(n28822) );
  INVxp33_ASAP7_75t_SRAM U36798 ( .A(n28536), .Y(n28543) );
  NOR2xp33_ASAP7_75t_SL U36799 ( .A(n24677), .B(n28546), .Y(n31821) );
  NOR2xp33_ASAP7_75t_SL U36800 ( .A(n22375), .B(n30637), .Y(n28902) );
  AOI21xp33_ASAP7_75t_SRAM U36801 ( .A1(u0_0_leon3x0_p0_iu_r_E__JMPL_), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__13_), .B(n22375), .Y(n26179) );
  AOI22xp33_ASAP7_75t_SRAM U36802 ( .A1(n28980), .A2(n22449), .B1(n24231), 
        .B2(n28979), .Y(n28870) );
  NOR2xp33_ASAP7_75t_SL U36803 ( .A(n22378), .B(n30488), .Y(n31873) );
  AOI22xp33_ASAP7_75t_SRAM U36804 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__13_), .A2(n30207), .B1(
        ic_q[13]), .B2(n22387), .Y(n29990) );
  AOI22xp33_ASAP7_75t_SRAM U36805 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__12_), .A2(n30207), .B1(
        it_q[8]), .B2(n24636), .Y(n25436) );
  AOI21xp33_ASAP7_75t_SRAM U36806 ( .A1(n24577), .A2(n24231), .B(n26155), .Y(
        n25759) );
  AOI22xp33_ASAP7_75t_SRAM U36807 ( .A1(n28821), .A2(u0_0_leon3x0_p0_divi[13]), 
        .B1(n27195), .B2(n27194), .Y(n27214) );
  AOI22xp33_ASAP7_75t_SRAM U36808 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__22_), .A2(n30207), .B1(
        ic_q[22]), .B2(n22387), .Y(n26222) );
  AOI22xp33_ASAP7_75t_SRAM U36809 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__19_), .A2(n30207), .B1(
        ic_q[19]), .B2(n22387), .Y(n25743) );
  AOI22xp33_ASAP7_75t_SRAM U36810 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__18_), .A2(n30207), .B1(
        ic_q[18]), .B2(n22387), .Y(n25716) );
  AOI22xp33_ASAP7_75t_SRAM U36811 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__20_), .A2(n30207), .B1(
        ic_q[20]), .B2(n22387), .Y(n26965) );
  NOR2xp33_ASAP7_75t_SL U36812 ( .A(n31396), .B(n27086), .Y(n31544) );
  OAI22xp33_ASAP7_75t_SRAM U36813 ( .A1(n30125), .A2(n31469), .B1(n30124), 
        .B2(n31001), .Y(n30129) );
  OAI21xp33_ASAP7_75t_SRAM U36814 ( .A1(n30245), .A2(n28934), .B(n30616), .Y(
        n25498) );
  AOI21xp33_ASAP7_75t_SRAM U36815 ( .A1(n28935), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__22_), .B(n28482), .Y(n28483) );
  NAND2xp33_ASAP7_75t_SRAM U36816 ( .A(n18606), .B(n24578), .Y(n25795) );
  NOR2xp33_ASAP7_75t_SL U36817 ( .A(n26745), .B(n26744), .Y(n28964) );
  NAND2xp33_ASAP7_75t_SRAM U36818 ( .A(n18530), .B(u0_0_leon3x0_p0_divi[30]), 
        .Y(n30656) );
  NOR2xp33_ASAP7_75t_SL U36819 ( .A(n30952), .B(n27020), .Y(n30671) );
  AOI21xp33_ASAP7_75t_SRAM U36820 ( .A1(n22416), .A2(n22436), .B(n18813), .Y(
        n25114) );
  NOR2xp33_ASAP7_75t_SL U36821 ( .A(n28977), .B(n28845), .Y(n28981) );
  AOI21xp33_ASAP7_75t_SRAM U36822 ( .A1(n22416), .A2(add_x_735_A_19_), .B(
        n18813), .Y(n25107) );
  NAND2xp33_ASAP7_75t_SRAM U36823 ( .A(u0_0_leon3x0_p0_iu_r_E__SARI_), .B(
        n18567), .Y(n25090) );
  NOR2xp33_ASAP7_75t_SL U36824 ( .A(n31537), .B(n32010), .Y(n24943) );
  NOR2xp33_ASAP7_75t_SL U36825 ( .A(n31858), .B(n32078), .Y(n32054) );
  NOR2xp33_ASAP7_75t_SL U36826 ( .A(n25513), .B(n30509), .Y(n32246) );
  AOI211xp5_ASAP7_75t_SL U36827 ( .A1(n28402), .A2(n18296), .B(n26525), .C(
        n26524), .Y(n32387) );
  AOI22xp33_ASAP7_75t_SRAM U36828 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__13_), 
        .A2(n22375), .B1(n23396), .B2(n28131), .Y(n26599) );
  NAND2xp33_ASAP7_75t_SRAM U36829 ( .A(n25106), .B(n25105), .Y(n24571) );
  OAI21xp33_ASAP7_75t_SRAM U36830 ( .A1(n25234), .A2(n30909), .B(n30908), .Y(
        DP_OP_1196_128_7433_n480) );
  OAI21xp33_ASAP7_75t_SRAM U36831 ( .A1(n31858), .A2(n30909), .B(n30908), .Y(
        DP_OP_1196_128_7433_n476) );
  OAI21xp33_ASAP7_75t_SRAM U36832 ( .A1(n30906), .A2(n30909), .B(n30908), .Y(
        DP_OP_1196_128_7433_n478) );
  OAI21xp33_ASAP7_75t_SRAM U36833 ( .A1(n30909), .A2(n32079), .B(n30908), .Y(
        DP_OP_1196_128_7433_n474) );
  NOR2xp33_ASAP7_75t_SL U36834 ( .A(n22380), .B(n32153), .Y(n31824) );
  XNOR2xp5_ASAP7_75t_SL U36835 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__1_), .B(
        DP_OP_1196_128_7433_n453), .Y(n24817) );
  OAI22xp33_ASAP7_75t_SRAM U36836 ( .A1(n32367), .A2(n24543), .B1(n32634), 
        .B2(n32429), .Y(n32368) );
  OAI22xp33_ASAP7_75t_SRAM U36837 ( .A1(n32354), .A2(n24543), .B1(n32630), 
        .B2(n32429), .Y(n32355) );
  OAI22xp33_ASAP7_75t_SRAM U36838 ( .A1(n32371), .A2(n24543), .B1(n32636), 
        .B2(n32429), .Y(n32372) );
  OAI22xp33_ASAP7_75t_SRAM U36839 ( .A1(n32361), .A2(n24543), .B1(n32632), 
        .B2(n32429), .Y(n32362) );
  OAI22xp33_ASAP7_75t_SRAM U36840 ( .A1(n32410), .A2(n24543), .B1(n32656), 
        .B2(n32429), .Y(n32411) );
  OAI22xp33_ASAP7_75t_SRAM U36841 ( .A1(n32419), .A2(n24543), .B1(n32658), 
        .B2(n32429), .Y(n32420) );
  NAND2xp33_ASAP7_75t_SRAM U36842 ( .A(n32351), .B(n32353), .Y(n32431) );
  AOI22xp33_ASAP7_75t_SRAM U36843 ( .A1(n32446), .A2(n32445), .B1(n32444), 
        .B2(u0_0_leon3x0_p0_dci[9]), .Y(n32450) );
  AOI21xp33_ASAP7_75t_SRAM U36844 ( .A1(n32317), .A2(n32353), .B(n32316), .Y(
        n32433) );
  AOI21xp33_ASAP7_75t_SRAM U36845 ( .A1(n32314), .A2(n32353), .B(n32313), .Y(
        n32423) );
  NAND2xp33_ASAP7_75t_SRAM U36846 ( .A(n32294), .B(n32296), .Y(n32435) );
  AOI21xp33_ASAP7_75t_SRAM U36847 ( .A1(n18859), .A2(n32280), .B(n32279), .Y(
        n32282) );
  INVxp33_ASAP7_75t_SRAM U36848 ( .A(n32274), .Y(n32277) );
  INVxp33_ASAP7_75t_SRAM U36849 ( .A(n32272), .Y(n32283) );
  AOI21xp33_ASAP7_75t_SRAM U36850 ( .A1(n32444), .A2(u0_0_leon3x0_p0_dci[16]), 
        .B(n32267), .Y(n32268) );
  AOI22xp33_ASAP7_75t_SRAM U36851 ( .A1(n32446), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[40]), .B1(n32444), .B2(
        u0_0_leon3x0_p0_dci[12]), .Y(n32266) );
  AOI22xp33_ASAP7_75t_SRAM U36852 ( .A1(n32446), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[39]), .B1(u0_0_leon3x0_p0_dci[11]), .B2(
        n32444), .Y(n32263) );
  AOI21xp33_ASAP7_75t_SRAM U36853 ( .A1(n32444), .A2(u0_0_leon3x0_p0_dci[10]), 
        .B(n32257), .Y(n32259) );
  OAI21xp33_ASAP7_75t_SRAM U36854 ( .A1(n32254), .A2(n32253), .B(n32252), .Y(
        n32447) );
  AOI21xp33_ASAP7_75t_SRAM U36855 ( .A1(n32183), .A2(n22421), .B(n32182), .Y(
        rf_addr_a[4]) );
  AOI22xp33_ASAP7_75t_SRAM U36856 ( .A1(n32234), .A2(n32343), .B1(n32214), 
        .B2(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__15_), .Y(n32208) );
  AOI22xp33_ASAP7_75t_SRAM U36857 ( .A1(n32234), .A2(n32342), .B1(n32214), 
        .B2(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__14_), .Y(n32207) );
  AOI22xp33_ASAP7_75t_SRAM U36858 ( .A1(n32234), .A2(n32339), .B1(n32214), 
        .B2(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__13_), .Y(n32206) );
  AOI22xp33_ASAP7_75t_SRAM U36859 ( .A1(n32234), .A2(n32336), .B1(
        u0_0_leon3x0_p0_dco_ICDIAG__ADDR__12_), .B2(n32214), .Y(n32205) );
  NAND2xp33_ASAP7_75t_SRAM U36860 ( .A(n3055), .B(n32231), .Y(n32217) );
  NAND2xp33_ASAP7_75t_SRAM U36861 ( .A(n32292), .B(n32443), .Y(n32239) );
  OAI21xp33_ASAP7_75t_SRAM U36862 ( .A1(n32317), .A2(n32232), .B(n32203), .Y(
        dt_data[7]) );
  OAI21xp33_ASAP7_75t_SRAM U36863 ( .A1(n32314), .A2(n32232), .B(n32203), .Y(
        dt_data[6]) );
  OAI21xp33_ASAP7_75t_SRAM U36864 ( .A1(n32310), .A2(n32232), .B(n32203), .Y(
        dt_data[5]) );
  OAI21xp33_ASAP7_75t_SRAM U36865 ( .A1(n32307), .A2(n32232), .B(n32203), .Y(
        dt_data[4]) );
  OAI21xp33_ASAP7_75t_SRAM U36866 ( .A1(n32305), .A2(n32232), .B(n32203), .Y(
        dt_data[3]) );
  OAI21xp33_ASAP7_75t_SRAM U36867 ( .A1(n32302), .A2(n32232), .B(n32203), .Y(
        dt_data[2]) );
  OAI21xp33_ASAP7_75t_SRAM U36868 ( .A1(n32300), .A2(n32232), .B(n32203), .Y(
        dt_data[1]) );
  OAI21xp33_ASAP7_75t_SRAM U36869 ( .A1(n32293), .A2(n32232), .B(n32203), .Y(
        dt_data[0]) );
  OAI21xp33_ASAP7_75t_SRAM U36870 ( .A1(n32197), .A2(n32275), .B(n32202), .Y(
        dt_wren) );
  INVxp33_ASAP7_75t_SRAM U36871 ( .A(n32333), .Y(n32619) );
  INVxp33_ASAP7_75t_SRAM U36872 ( .A(n32328), .Y(n32617) );
  INVxp33_ASAP7_75t_SRAM U36873 ( .A(n32322), .Y(n32613) );
  INVxp33_ASAP7_75t_SRAM U36874 ( .A(n32315), .Y(n32609) );
  INVxp33_ASAP7_75t_SRAM U36875 ( .A(n32311), .Y(n32607) );
  INVxp33_ASAP7_75t_SRAM U36876 ( .A(n32308), .Y(n32605) );
  INVxp33_ASAP7_75t_SRAM U36877 ( .A(n32306), .Y(n32603) );
  INVxp33_ASAP7_75t_SRAM U36878 ( .A(n32303), .Y(n32601) );
  INVxp33_ASAP7_75t_SRAM U36879 ( .A(n32301), .Y(n32600) );
  INVxp33_ASAP7_75t_SRAM U36880 ( .A(n32297), .Y(n32599) );
  OAI22xp33_ASAP7_75t_SRAM U36881 ( .A1(n32687), .A2(n32669), .B1(n32668), 
        .B2(n32676), .Y(n32670) );
  OAI21xp33_ASAP7_75t_SRAM U36882 ( .A1(n32681), .A2(n14803), .B(n32680), .Y(
        ic_address[1]) );
  OAI22xp33_ASAP7_75t_SRAM U36883 ( .A1(n32687), .A2(n32677), .B1(n2935), .B2(
        n32676), .Y(n32678) );
  OAI21xp33_ASAP7_75t_SRAM U36884 ( .A1(n33054), .A2(n32152), .B(n32153), .Y(
        rf_addr_w[0]) );
  AOI22xp33_ASAP7_75t_SRAM U36885 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VADDRESS__4_), .A2(n32689), .B1(
        u0_0_leon3x0_p0_ici[62]), .B2(n32688), .Y(n32690) );
  INVxp33_ASAP7_75t_SRAM U36886 ( .A(n32545), .Y(n32559) );
  NAND2xp33_ASAP7_75t_SRAM U36887 ( .A(n18848), .B(n32561), .Y(n32542) );
  OAI21xp33_ASAP7_75t_SRAM U36888 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_), .A2(n24684), .B(n32562), 
        .Y(n32563) );
  NAND2xp33_ASAP7_75t_SRAM U36889 ( .A(n32561), .B(n32686), .Y(n32595) );
  AOI21xp33_ASAP7_75t_SRAM U36890 ( .A1(n2867), .A2(n29960), .B(n27536), .Y(
        n27526) );
  OAI21xp33_ASAP7_75t_SRAM U36891 ( .A1(u0_0_leon3x0_p0_c0mmu_a0_r_BG_), .A2(
        n32705), .B(n24684), .Y(n4390) );
  OAI21xp33_ASAP7_75t_SRAM U36892 ( .A1(n32705), .A2(ahb0_r_HMASTERD_), .B(
        n22393), .Y(n3901) );
  INVxp33_ASAP7_75t_SRAM U36893 ( .A(n24989), .Y(n24991) );
  AOI21xp33_ASAP7_75t_SRAM U36894 ( .A1(n25693), .A2(n25670), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__1_), .Y(n24994) );
  OAI21xp33_ASAP7_75t_SRAM U36895 ( .A1(n4770), .A2(n31953), .B(n31952), .Y(
        n31955) );
  OAI21xp33_ASAP7_75t_SRAM U36896 ( .A1(n29851), .A2(n29743), .B(
        irqctrl0_r_IPEND__12_), .Y(n29243) );
  OAI21xp33_ASAP7_75t_SRAM U36897 ( .A1(n28116), .A2(n29743), .B(
        irqctrl0_r_IPEND__11_), .Y(n25964) );
  OAI21xp33_ASAP7_75t_SRAM U36898 ( .A1(n29568), .A2(n29743), .B(n29377), .Y(
        n29381) );
  OAI21xp33_ASAP7_75t_SRAM U36899 ( .A1(n30372), .A2(n31404), .B(n22379), .Y(
        n30373) );
  OAI21xp33_ASAP7_75t_SRAM U36900 ( .A1(n30441), .A2(n31404), .B(n22379), .Y(
        n30442) );
  OAI21xp33_ASAP7_75t_SRAM U36901 ( .A1(n30454), .A2(n31404), .B(n22379), .Y(
        n30455) );
  AOI22xp33_ASAP7_75t_SRAM U36902 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .A2(n25700), .B1(n25699), 
        .B2(n25698), .Y(n25701) );
  INVxp33_ASAP7_75t_SRAM U36903 ( .A(n25680), .Y(n25681) );
  OAI21xp33_ASAP7_75t_SRAM U36904 ( .A1(n25695), .A2(n25676), .B(n25675), .Y(
        n25688) );
  OAI21xp33_ASAP7_75t_SRAM U36905 ( .A1(n31678), .A2(n31404), .B(n22379), .Y(
        n30216) );
  OAI21xp33_ASAP7_75t_SRAM U36906 ( .A1(n30287), .A2(n31404), .B(n22379), .Y(
        n30288) );
  NOR2xp33_ASAP7_75t_SL U36907 ( .A(n24678), .B(n26869), .Y(n30813) );
  INVxp33_ASAP7_75t_SRAM U36908 ( .A(n24974), .Y(n24975) );
  AOI22xp33_ASAP7_75t_SRAM U36909 ( .A1(n31325), .A2(n31324), .B1(
        sr1_r_MCFG1__BRDYEN_), .B2(n32003), .Y(n31326) );
  AOI21xp33_ASAP7_75t_SRAM U36910 ( .A1(n30430), .A2(u0_0_leon3x0_p0_divi[56]), 
        .B(n24680), .Y(n30253) );
  OAI21xp33_ASAP7_75t_SRAM U36911 ( .A1(n2925), .A2(n26501), .B(n26658), .Y(
        n30806) );
  AOI22xp33_ASAP7_75t_SRAM U36912 ( .A1(irqctrl0_r_IMASK__0__12_), .A2(n31249), 
        .B1(irqctrl0_r_IFORCE__0__12_), .B2(n31251), .Y(n29852) );
  AOI22xp33_ASAP7_75t_SRAM U36913 ( .A1(irqctrl0_r_IMASK__0__9_), .A2(n31249), 
        .B1(irqctrl0_r_IFORCE__0__9_), .B2(n31251), .Y(n30143) );
  AOI22xp33_ASAP7_75t_SRAM U36914 ( .A1(n31249), .A2(n29412), .B1(
        irqctrl0_r_IFORCE__0__11_), .B2(n31251), .Y(n28122) );
  AOI22xp33_ASAP7_75t_SRAM U36915 ( .A1(timer0_vtimers_1__RESTART_), .A2(
        n30790), .B1(timer0_vtimers_1__RELOAD__1_), .B2(n31956), .Y(n27484) );
  AOI22xp33_ASAP7_75t_SRAM U36916 ( .A1(irqctrl0_r_IMASK__0__1_), .A2(n31249), 
        .B1(irqctrl0_r_IFORCE__0__1_), .B2(n31251), .Y(n27481) );
  AOI22xp33_ASAP7_75t_SRAM U36917 ( .A1(irqctrl0_r_IMASK__0__8_), .A2(n31249), 
        .B1(irqctrl0_r_IFORCE__0__8_), .B2(n31251), .Y(n29750) );
  NOR2xp33_ASAP7_75t_SL U36918 ( .A(apb0_r_CFGSEL_), .B(n31953), .Y(n32008) );
  AOI22xp33_ASAP7_75t_SRAM U36919 ( .A1(irqctrl0_r_IMASK__0__10_), .A2(n31249), 
        .B1(irqctrl0_r_IFORCE__0__10_), .B2(n31251), .Y(n30981) );
  INVxp33_ASAP7_75t_SRAM U36920 ( .A(n31956), .Y(n31243) );
  AOI22xp33_ASAP7_75t_SRAM U36921 ( .A1(irqctrl0_r_IMASK__0__5_), .A2(n31249), 
        .B1(irqctrl0_r_IFORCE__0__5_), .B2(n31251), .Y(n30079) );
  INVxp33_ASAP7_75t_SRAM U36922 ( .A(n27463), .Y(n28085) );
  INVxp33_ASAP7_75t_SRAM U36923 ( .A(n31953), .Y(n30789) );
  AOI22xp33_ASAP7_75t_SRAM U36924 ( .A1(ahb0_r_HADDR__7_), .A2(n22393), .B1(
        n32705), .B2(n32995), .Y(n4758) );
  AOI22xp33_ASAP7_75t_SRAM U36925 ( .A1(ahb0_r_HADDR__6_), .A2(n22393), .B1(
        n32705), .B2(n32994), .Y(n2345) );
  OAI21xp33_ASAP7_75t_SRAM U36926 ( .A1(n31627), .A2(n32035), .B(n24684), .Y(
        n3905) );
  INVxp33_ASAP7_75t_SRAM U36927 ( .A(n32071), .Y(n30689) );
  INVxp33_ASAP7_75t_SRAM U36928 ( .A(n32187), .Y(n32189) );
  INVxp33_ASAP7_75t_SRAM U36929 ( .A(n31960), .Y(n31966) );
  AOI22xp33_ASAP7_75t_SRAM U36930 ( .A1(n30622), .A2(u0_0_leon3x0_p0_divi[5]), 
        .B1(u0_0_leon3x0_p0_iu_r_W__S__WIM__6_), .B2(n28890), .Y(n26271) );
  AOI22xp33_ASAP7_75t_SRAM U36931 ( .A1(n31790), .A2(n22415), .B1(n31789), 
        .B2(n32719), .Y(n31793) );
  AOI21xp33_ASAP7_75t_SRAM U36932 ( .A1(n28821), .A2(n18904), .B(n28731), .Y(
        n28733) );
  INVxp33_ASAP7_75t_SRAM U36933 ( .A(n18316), .Y(n28633) );
  AOI21xp33_ASAP7_75t_SRAM U36934 ( .A1(n29588), .A2(u0_0_leon3x0_p0_divi[10]), 
        .B(n22375), .Y(n28687) );
  AOI21xp33_ASAP7_75t_SRAM U36935 ( .A1(n29721), .A2(n29720), .B(n29719), .Y(
        n29722) );
  INVxp33_ASAP7_75t_SRAM U36936 ( .A(n29716), .Y(n29718) );
  AOI21xp33_ASAP7_75t_SRAM U36937 ( .A1(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__19_), .A2(n29708), .B(n29707), .Y(
        n29709) );
  AOI21xp33_ASAP7_75t_SRAM U36938 ( .A1(n29706), .A2(n29705), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__24_), .Y(n29710) );
  INVxp33_ASAP7_75t_SRAM U36939 ( .A(n29704), .Y(n29711) );
  INVxp33_ASAP7_75t_SRAM U36940 ( .A(n29701), .Y(n29714) );
  AOI22xp33_ASAP7_75t_SRAM U36941 ( .A1(n29583), .A2(n24231), .B1(n28529), 
        .B2(n29598), .Y(n25779) );
  AOI22xp33_ASAP7_75t_SRAM U36942 ( .A1(n18327), .A2(n28631), .B1(n28835), 
        .B2(n30302), .Y(n25769) );
  INVxp33_ASAP7_75t_SRAM U36943 ( .A(n28878), .Y(n25771) );
  AOI21xp33_ASAP7_75t_SRAM U36944 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__31_), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__13_), .B(n24679), .Y(n26870) );
  AOI21xp33_ASAP7_75t_SRAM U36945 ( .A1(n28631), .A2(u0_0_leon3x0_p0_muli[28]), 
        .B(n26997), .Y(n27000) );
  AOI21xp33_ASAP7_75t_SRAM U36946 ( .A1(u0_0_leon3x0_p0_iu_r_E__JMPL_), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__18_), .B(n22375), .Y(n25829) );
  INVxp33_ASAP7_75t_SRAM U36947 ( .A(u0_0_leon3x0_p0_muli[26]), .Y(n25816) );
  OAI21xp33_ASAP7_75t_SRAM U36948 ( .A1(n25813), .A2(n28481), .B(n29504), .Y(
        n25814) );
  INVxp33_ASAP7_75t_SRAM U36949 ( .A(n28486), .Y(n25812) );
  AOI22xp33_ASAP7_75t_SRAM U36950 ( .A1(u0_0_leon3x0_p0_muli[25]), .A2(n28631), 
        .B1(n28835), .B2(n30322), .Y(n26704) );
  AOI22xp33_ASAP7_75t_SRAM U36951 ( .A1(n27065), .A2(n30619), .B1(n28894), 
        .B2(n30326), .Y(n26705) );
  OAI22xp33_ASAP7_75t_SRAM U36952 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__13_), 
        .A2(n27143), .B1(n26171), .B2(n27141), .Y(n26172) );
  INVxp33_ASAP7_75t_SRAM U36953 ( .A(u0_0_leon3x0_p0_muli[23]), .Y(n26171) );
  OAI21xp33_ASAP7_75t_SRAM U36954 ( .A1(n28593), .A2(n28481), .B(n29504), .Y(
        n26170) );
  AO22x1_ASAP7_75t_SL U36955 ( .A1(dc_q[14]), .A2(n31473), .B1(dt_q[10]), .B2(
        n29991), .Y(n24484) );
  INVxp33_ASAP7_75t_SRAM U36956 ( .A(n30557), .Y(n32625) );
  OAI22xp33_ASAP7_75t_SRAM U36957 ( .A1(n23061), .A2(n26294), .B1(n18381), 
        .B2(n28843), .Y(n26295) );
  OAI21xp33_ASAP7_75t_SRAM U36958 ( .A1(n31475), .A2(n31474), .B(n31491), .Y(
        n31476) );
  AOI22xp33_ASAP7_75t_SRAM U36959 ( .A1(n30622), .A2(u0_0_leon3x0_p0_divi[20]), 
        .B1(u0_0_leon3x0_p0_iu_de_icc_1_), .B2(n30621), .Y(n27070) );
  INVxp33_ASAP7_75t_SRAM U36960 ( .A(n30017), .Y(n30020) );
  OAI22xp33_ASAP7_75t_SRAM U36961 ( .A1(n32301), .A2(n31470), .B1(n24426), 
        .B2(n32468), .Y(n31354) );
  AOI21xp33_ASAP7_75t_SRAM U36962 ( .A1(n28486), .A2(n22436), .B(n28485), .Y(
        n28487) );
  AOI21xp33_ASAP7_75t_SRAM U36963 ( .A1(n24581), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__27_), .B(n22375), .Y(n26895) );
  INVxp33_ASAP7_75t_SRAM U36964 ( .A(n29869), .Y(n29176) );
  OAI22xp33_ASAP7_75t_SRAM U36965 ( .A1(n22493), .A2(n27075), .B1(n29910), 
        .B2(n26675), .Y(n26422) );
  AOI22xp33_ASAP7_75t_SRAM U36966 ( .A1(n29583), .A2(n18606), .B1(n29783), 
        .B2(n29598), .Y(n28437) );
  AOI21xp33_ASAP7_75t_SRAM U36967 ( .A1(n28631), .A2(u0_0_leon3x0_p0_muli[33]), 
        .B(n28423), .Y(n28429) );
  AOI21xp33_ASAP7_75t_SRAM U36968 ( .A1(n24581), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__25_), .B(n22375), .Y(n28421) );
  AOI21xp33_ASAP7_75t_SRAM U36969 ( .A1(n29588), .A2(u0_0_leon3x0_p0_divi[23]), 
        .B(n22375), .Y(n26395) );
  INVxp33_ASAP7_75t_SRAM U36970 ( .A(n26915), .Y(n26936) );
  INVxp33_ASAP7_75t_SRAM U36971 ( .A(u0_0_leon3x0_p0_muli[35]), .Y(n25892) );
  AOI21xp33_ASAP7_75t_SRAM U36972 ( .A1(n26565), .A2(n29150), .B(n18299), .Y(
        n26567) );
  INVxp33_ASAP7_75t_SRAM U36973 ( .A(u0_0_leon3x0_p0_divi[18]), .Y(n25773) );
  INVxp33_ASAP7_75t_SRAM U36974 ( .A(n24066), .Y(n27142) );
  AOI22xp33_ASAP7_75t_SRAM U36975 ( .A1(n24937), .A2(n25659), .B1(n25667), 
        .B2(n25652), .Y(n24918) );
  AOI22xp33_ASAP7_75t_SRAM U36976 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__30_), 
        .A2(n29589), .B1(u0_0_leon3x0_p0_divi[29]), .B2(n29588), .Y(n29590) );
  INVxp33_ASAP7_75t_SRAM U36977 ( .A(u0_0_leon3x0_p0_divi[20]), .Y(n27059) );
  INVxp33_ASAP7_75t_SRAM U36978 ( .A(u0_0_leon3x0_p0_divi[0]), .Y(n30660) );
  AOI21xp33_ASAP7_75t_SRAM U36979 ( .A1(n22416), .A2(n22968), .B(n18813), .Y(
        n25197) );
  AOI22xp33_ASAP7_75t_SRAM U36980 ( .A1(n29583), .A2(n18530), .B1(n26725), 
        .B2(n29598), .Y(n25184) );
  AOI21xp33_ASAP7_75t_SRAM U36981 ( .A1(n22416), .A2(n18530), .B(n18813), .Y(
        n25147) );
  AOI21xp33_ASAP7_75t_SRAM U36982 ( .A1(n22416), .A2(n18296), .B(n18813), .Y(
        n25146) );
  AOI21xp33_ASAP7_75t_SRAM U36983 ( .A1(n31418), .A2(n29150), .B(n23974), .Y(
        n25133) );
  AOI21xp33_ASAP7_75t_SRAM U36984 ( .A1(n26278), .A2(add_x_735_A_32_), .B(
        n26155), .Y(n25097) );
  INVxp33_ASAP7_75t_SRAM U36985 ( .A(n31627), .Y(n31628) );
  INVxp33_ASAP7_75t_SRAM U36986 ( .A(n31697), .Y(n31701) );
  OAI21xp33_ASAP7_75t_SRAM U36987 ( .A1(n25226), .A2(n32087), .B(n26868), .Y(
        n25227) );
  AOI21xp33_ASAP7_75t_SRAM U36988 ( .A1(n32087), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), .B(n32079), .Y(n25223) );
  INVxp33_ASAP7_75t_SRAM U36989 ( .A(n32081), .Y(n25220) );
  NAND2xp33_ASAP7_75t_SRAM U36990 ( .A(n32238), .B(n31565), .Y(n32292) );
  INVxp33_ASAP7_75t_SRAM U36991 ( .A(n31452), .Y(n32200) );
  AOI22xp33_ASAP7_75t_SRAM U36992 ( .A1(n29112), .A2(n31417), .B1(n31420), 
        .B2(u0_0_leon3x0_p0_div0_addout_32_), .Y(n28289) );
  INVxp33_ASAP7_75t_SRAM U36993 ( .A(n32022), .Y(n32026) );
  AOI21xp33_ASAP7_75t_SRAM U36994 ( .A1(n2963), .A2(n31306), .B(n31608), .Y(
        n31307) );
  INVxp33_ASAP7_75t_SRAM U36995 ( .A(n31306), .Y(n31302) );
  AOI21xp33_ASAP7_75t_SRAM U36996 ( .A1(u0_0_leon3x0_p0_dci[34]), .A2(n31828), 
        .B(n29026), .Y(n29028) );
  AOI21xp33_ASAP7_75t_SRAM U36997 ( .A1(u0_0_leon3x0_p0_dci[26]), .A2(n31828), 
        .B(n27040), .Y(n27042) );
  AOI21xp33_ASAP7_75t_SRAM U36998 ( .A1(u0_0_leon3x0_p0_dci[20]), .A2(n31828), 
        .B(n28566), .Y(n28568) );
  AOI21xp33_ASAP7_75t_SRAM U36999 ( .A1(u0_0_leon3x0_p0_dci[17]), .A2(n31828), 
        .B(n29820), .Y(n29822) );
  AOI21xp33_ASAP7_75t_SRAM U37000 ( .A1(u0_0_leon3x0_p0_dci[36]), .A2(n31828), 
        .B(n31682), .Y(n31684) );
  AOI21xp33_ASAP7_75t_SRAM U37001 ( .A1(u0_0_leon3x0_p0_dci[24]), .A2(n31828), 
        .B(n30823), .Y(n30825) );
  AOI21xp33_ASAP7_75t_SRAM U37002 ( .A1(u0_0_leon3x0_p0_dci[32]), .A2(n31828), 
        .B(n26874), .Y(n26876) );
  AOI21xp33_ASAP7_75t_SRAM U37003 ( .A1(u0_0_leon3x0_p0_c0mmu_mcdi[0]), .A2(
        n31572), .B(n25588), .Y(n25590) );
  AOI22xp33_ASAP7_75t_SRAM U37004 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__9_), .A2(
        n22375), .B1(add_x_735_A_10_), .B2(n28131), .Y(n25405) );
  AOI22xp33_ASAP7_75t_SRAM U37005 ( .A1(u0_0_leon3x0_p0_iu_r_E__OP1__15_), 
        .A2(n22375), .B1(n23964), .B2(n28131), .Y(n26587) );
  OAI21xp33_ASAP7_75t_SRAM U37006 ( .A1(n30905), .A2(n30909), .B(n30908), .Y(
        DP_OP_1196_128_7433_n479) );
  NOR2xp33_ASAP7_75t_SL U37007 ( .A(n27477), .B(n26467), .Y(n31956) );
  NAND2xp5_ASAP7_75t_SL U37008 ( .A(n25979), .B(n31057), .Y(n26012) );
  NOR2xp33_ASAP7_75t_SL U37009 ( .A(n2925), .B(n27479), .Y(n26072) );
  AOI211xp5_ASAP7_75t_SL U37010 ( .A1(dc_q[18]), .A2(n32385), .B(n32369), .C(
        n32368), .Y(n32370) );
  NOR2xp33_ASAP7_75t_SL U37011 ( .A(n32366), .B(n32431), .Y(n32369) );
  NAND2xp33_ASAP7_75t_SRAM U37012 ( .A(n32393), .B(n32386), .Y(n32358) );
  NAND2xp33_ASAP7_75t_SRAM U37013 ( .A(n32403), .B(n32386), .Y(n32373) );
  NAND2xp33_ASAP7_75t_SRAM U37014 ( .A(n32396), .B(n32386), .Y(n32363) );
  NAND2xp33_ASAP7_75t_SRAM U37015 ( .A(n32345), .B(n32433), .Y(n32346) );
  NOR2xp33_ASAP7_75t_SL U37016 ( .A(n32435), .B(n32357), .Y(n32386) );
  NAND2xp33_ASAP7_75t_SRAM U37017 ( .A(n32350), .B(n32389), .Y(n32385) );
  NAND2xp33_ASAP7_75t_SRAM U37018 ( .A(n32414), .B(n32413), .Y(n32415) );
  AOI211xp5_ASAP7_75t_SL U37019 ( .A1(dc_q[29]), .A2(n33069), .B(n32412), .C(
        n32411), .Y(n32416) );
  NOR2xp33_ASAP7_75t_SL U37020 ( .A(n32409), .B(n32408), .Y(n32412) );
  AOI211xp5_ASAP7_75t_SL U37021 ( .A1(n32423), .A2(n32434), .B(n32422), .C(
        n32421), .Y(n32424) );
  NOR2xp33_ASAP7_75t_SL U37022 ( .A(n32418), .B(n32431), .Y(n32422) );
  OR2x2_ASAP7_75t_SL U37023 ( .A(n32353), .B(n32352), .Y(n32429) );
  NAND2xp33_ASAP7_75t_SRAM U37024 ( .A(n32350), .B(n32321), .Y(n33069) );
  NOR2xp33_ASAP7_75t_SL U37025 ( .A(n24643), .B(n32349), .Y(n32351) );
  NOR2xp33_ASAP7_75t_SL U37026 ( .A(n32390), .B(n32389), .Y(n32434) );
  NAND2xp33_ASAP7_75t_SRAM U37027 ( .A(n32444), .B(n32438), .Y(n32439) );
  NAND2xp33_ASAP7_75t_SRAM U37028 ( .A(n32444), .B(u0_0_leon3x0_p0_dci[8]), 
        .Y(n32441) );
  NAND2xp33_ASAP7_75t_SRAM U37029 ( .A(n32450), .B(n32449), .Y(dc_address[2])
         );
  NAND2xp33_ASAP7_75t_SRAM U37030 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[0]), .B(
        n32584), .Y(n32464) );
  NAND2xp33_ASAP7_75t_SRAM U37031 ( .A(n32584), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[1]), .Y(n32471) );
  NAND2xp33_ASAP7_75t_SRAM U37032 ( .A(n32584), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[2]), .Y(n32478) );
  NAND2xp33_ASAP7_75t_SRAM U37033 ( .A(n32584), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[3]), .Y(n32486) );
  NAND2xp33_ASAP7_75t_SRAM U37034 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[5]), .B(
        n32584), .Y(n32500) );
  NAND2xp33_ASAP7_75t_SRAM U37035 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[6]), .B(
        n32584), .Y(n32507) );
  NAND2xp33_ASAP7_75t_SRAM U37036 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[7]), .B(
        n32584), .Y(n32520) );
  NAND2xp33_ASAP7_75t_SRAM U37037 ( .A(n32345), .B(n32406), .Y(n32337) );
  NAND2xp33_ASAP7_75t_SRAM U37038 ( .A(n32345), .B(n32403), .Y(n32334) );
  NAND2xp33_ASAP7_75t_SRAM U37039 ( .A(n32340), .B(n32400), .Y(n32330) );
  NAND2xp33_ASAP7_75t_SRAM U37040 ( .A(n32345), .B(n32396), .Y(n32326) );
  NAND2xp33_ASAP7_75t_SRAM U37041 ( .A(n32345), .B(n32393), .Y(n32323) );
  NOR2xp33_ASAP7_75t_SL U37042 ( .A(n32356), .B(n32350), .Y(n32345) );
  NAND2xp33_ASAP7_75t_SRAM U37043 ( .A(n32349), .B(n32288), .Y(n32350) );
  NAND2xp33_ASAP7_75t_SRAM U37044 ( .A(n32435), .B(n32321), .Y(n32344) );
  NAND2xp33_ASAP7_75t_SRAM U37045 ( .A(n32296), .B(n32151), .Y(n32321) );
  NOR2xp33_ASAP7_75t_SL U37046 ( .A(n32295), .B(n32286), .Y(n32151) );
  NOR2xp33_ASAP7_75t_SL U37047 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[7]), .B(
        n32353), .Y(n32316) );
  NOR2xp33_ASAP7_75t_SL U37048 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[6]), .B(
        n32353), .Y(n32313) );
  NAND2xp33_ASAP7_75t_SRAM U37049 ( .A(n32435), .B(n32389), .Y(n32318) );
  NAND2xp33_ASAP7_75t_SRAM U37050 ( .A(n32295), .B(n32388), .Y(n32356) );
  NOR2xp33_ASAP7_75t_SL U37051 ( .A(n24643), .B(n32285), .Y(n32296) );
  NOR2xp33_ASAP7_75t_SL U37052 ( .A(n32290), .B(n32289), .Y(n32291) );
  NOR2xp33_ASAP7_75t_SL U37053 ( .A(n32730), .B(n32428), .Y(n32427) );
  NOR2xp33_ASAP7_75t_SL U37054 ( .A(n32148), .B(n32290), .Y(n32149) );
  NOR2xp33_ASAP7_75t_SL U37055 ( .A(n24643), .B(n32294), .Y(n32288) );
  NOR2xp33_ASAP7_75t_SL U37056 ( .A(n32147), .B(n32146), .Y(n32294) );
  NOR2xp33_ASAP7_75t_SL U37057 ( .A(n32734), .B(n32428), .Y(n32146) );
  NOR2xp33_ASAP7_75t_SL U37058 ( .A(n32145), .B(n32290), .Y(n32147) );
  NAND2xp33_ASAP7_75t_SRAM U37059 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_VALID_), 
        .B(u0_0_leon3x0_p0_dco_HIT_), .Y(n32276) );
  NAND2xp33_ASAP7_75t_SRAM U37060 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__2_), .B(n33067), .Y(n32264) );
  NAND2xp33_ASAP7_75t_SRAM U37061 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__1_), .B(n33067), .Y(n32261) );
  OAI31xp33_ASAP7_75t_SL U37062 ( .A1(n3132), .A2(n32250), .A3(n32249), .B(
        n32248), .Y(n32448) );
  NAND2xp33_ASAP7_75t_SRAM U37063 ( .A(n32247), .B(n32246), .Y(n32256) );
  NOR2xp33_ASAP7_75t_SL U37064 ( .A(u0_0_leon3x0_p0_dci[2]), .B(n32236), .Y(
        n32255) );
  NAND2xp33_ASAP7_75t_SRAM U37065 ( .A(n32234), .B(n32228), .Y(n32229) );
  NAND2xp33_ASAP7_75t_SRAM U37066 ( .A(n32231), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[27]), .Y(n32226) );
  NAND2xp33_ASAP7_75t_SRAM U37067 ( .A(n32231), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[26]), .Y(n32224) );
  NAND2xp33_ASAP7_75t_SRAM U37068 ( .A(n32231), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[25]), .Y(n32222) );
  NAND2xp33_ASAP7_75t_SRAM U37069 ( .A(n32231), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[24]), .Y(n32220) );
  NOR2xp33_ASAP7_75t_SL U37070 ( .A(n32204), .B(n33067), .Y(n32214) );
  NOR2xp33_ASAP7_75t_SL U37071 ( .A(n32234), .B(n32239), .Y(n32231) );
  INVx1_ASAP7_75t_SL U37072 ( .A(n32234), .Y(n32232) );
  AND2x2_ASAP7_75t_SL U37073 ( .A(n32196), .B(n18859), .Y(n32234) );
  NOR2xp33_ASAP7_75t_SL U37074 ( .A(n32195), .B(n32194), .Y(n32196) );
  NAND2xp33_ASAP7_75t_SRAM U37075 ( .A(n32458), .B(n14803), .Y(n32597) );
  NAND2xp33_ASAP7_75t_SRAM U37076 ( .A(u0_0_leon3x0_p0_dci[2]), .B(n32290), 
        .Y(n32143) );
  NOR2xp33_ASAP7_75t_SL U37077 ( .A(n32559), .B(n32546), .Y(it_data[20]) );
  NOR2xp33_ASAP7_75t_SL U37078 ( .A(n32559), .B(n32552), .Y(it_data[22]) );
  NOR2xp33_ASAP7_75t_SL U37079 ( .A(n32559), .B(n32549), .Y(it_data[21]) );
  NOR2xp33_ASAP7_75t_SL U37080 ( .A(n32565), .B(n32676), .Y(n32590) );
  OR2x2_ASAP7_75t_SL U37081 ( .A(n32583), .B(n14803), .Y(n32593) );
  NOR2xp33_ASAP7_75t_SL U37082 ( .A(n32687), .B(n32565), .Y(n32594) );
  AOI21xp33_ASAP7_75t_SRAM U37083 ( .A1(n4316), .A2(n32564), .B(n32563), .Y(
        n32687) );
  AOI21xp33_ASAP7_75t_SRAM U37084 ( .A1(n3880), .A2(n4316), .B(
        u0_0_leon3x0_p0_c0mmu_icache0_r_ISTATE__1_), .Y(n32686) );
  NOR2xp33_ASAP7_75t_SL U37085 ( .A(n17251), .B(n17252), .Y(apb0_N1148) );
  NOR2xp33_ASAP7_75t_SL U37086 ( .A(n31020), .B(n31019), .Y(n2333) );
  NOR2xp33_ASAP7_75t_SL U37087 ( .A(n30833), .B(n22397), .Y(n29942) );
  NOR2xp33_ASAP7_75t_SL U37088 ( .A(n31197), .B(n22397), .Y(n25863) );
  NOR2xp33_ASAP7_75t_SL U37089 ( .A(n29568), .B(n22397), .Y(n29569) );
  NOR2xp33_ASAP7_75t_SL U37090 ( .A(n29510), .B(n22397), .Y(n29509) );
  NOR2xp33_ASAP7_75t_SL U37091 ( .A(n30073), .B(n22397), .Y(n30029) );
  NOR2xp33_ASAP7_75t_SL U37092 ( .A(n28108), .B(n22397), .Y(n28109) );
  NOR2xp33_ASAP7_75t_SL U37093 ( .A(n30780), .B(n22397), .Y(n25877) );
  NOR2xp33_ASAP7_75t_SL U37094 ( .A(n27493), .B(n22397), .Y(n27494) );
  NOR2xp33_ASAP7_75t_SL U37095 ( .A(n26544), .B(n22397), .Y(n26542) );
  NOR2xp33_ASAP7_75t_SL U37096 ( .A(n28181), .B(n28182), .Y(n28185) );
  NOR2xp33_ASAP7_75t_SL U37097 ( .A(n30906), .B(n24646), .Y(n26822) );
  NOR2xp33_ASAP7_75t_SL U37098 ( .A(n30147), .B(n30136), .Y(n30135) );
  NOR2xp33_ASAP7_75t_SL U37099 ( .A(n4536), .B(n30134), .Y(n30136) );
  NOR2xp33_ASAP7_75t_SL U37100 ( .A(n2292), .B(n31719), .Y(n31729) );
  NOR2xp33_ASAP7_75t_SL U37101 ( .A(n28032), .B(n29947), .Y(n28041) );
  NOR2xp33_ASAP7_75t_SL U37102 ( .A(n31711), .B(n31710), .Y(n31727) );
  NAND2xp33_ASAP7_75t_SRAM U37103 ( .A(n31751), .B(n32832), .Y(n31728) );
  NOR2xp33_ASAP7_75t_SL U37104 ( .A(sr1_r_WS__2_), .B(n31723), .Y(n31717) );
  NOR2xp33_ASAP7_75t_SL U37105 ( .A(n31713), .B(n32716), .Y(n31722) );
  NOR2xp33_ASAP7_75t_SL U37106 ( .A(n29970), .B(n29969), .Y(n2866) );
  NOR2xp33_ASAP7_75t_SL U37107 ( .A(n29968), .B(n29967), .Y(n29969) );
  NAND2xp33_ASAP7_75t_SRAM U37108 ( .A(uart1_r_RXSTATE__1_), .B(n29960), .Y(
        n29963) );
  NOR2xp33_ASAP7_75t_SL U37109 ( .A(n32136), .B(n32135), .Y(n3584) );
  AOI211xp5_ASAP7_75t_SL U37110 ( .A1(u0_0_leon3x0_p0_muli[8]), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__22_), .C(n32131), .Y(n32133) );
  NOR2xp33_ASAP7_75t_SL U37111 ( .A(n25234), .B(n24646), .Y(n26809) );
  NOR2xp33_ASAP7_75t_SL U37112 ( .A(n30905), .B(n24646), .Y(n26825) );
  NOR2xp33_ASAP7_75t_SL U37113 ( .A(n30119), .B(n22379), .Y(n30122) );
  NOR2xp33_ASAP7_75t_SL U37114 ( .A(u0_0_leon3x0_p0_iu_r_W__S__PS_), .B(n30117), .Y(n30116) );
  NAND2xp33_ASAP7_75t_SRAM U37115 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__RETT_), 
        .B(n30115), .Y(n30117) );
  NOR2xp33_ASAP7_75t_SL U37116 ( .A(n31981), .B(n24646), .Y(n30878) );
  NOR2xp33_ASAP7_75t_SL U37117 ( .A(ahb0_r_HADDR__2_), .B(n17285), .Y(n31020)
         );
  NAND3xp33_ASAP7_75t_SL U37118 ( .A(n25241), .B(n25240), .C(ahb0_r_HADDR__5_), 
        .Y(n17271) );
  NOR2xp33_ASAP7_75t_SL U37119 ( .A(n25238), .B(n30802), .Y(n25242) );
  NOR2xp33_ASAP7_75t_SL U37120 ( .A(ahb0_r_HADDR__8_), .B(ahb0_r_HADDR__10_), 
        .Y(n24982) );
  AOI211xp5_ASAP7_75t_SL U37121 ( .A1(uart1_r_TSEMPTY_), .A2(n29949), .B(
        n24695), .C(n29367), .Y(n2243) );
  NOR2xp33_ASAP7_75t_SL U37122 ( .A(n31395), .B(n24641), .Y(rf_di_w[0]) );
  NOR2xp33_ASAP7_75t_SL U37123 ( .A(n22919), .B(n22427), .Y(n32018) );
  NAND2xp33_ASAP7_75t_SRAM U37124 ( .A(uart1_r_RXSTATE__0_), .B(n29967), .Y(
        n28188) );
  NOR2xp33_ASAP7_75t_SL U37125 ( .A(n28187), .B(n28186), .Y(n29967) );
  NOR2xp33_ASAP7_75t_SL U37126 ( .A(n24921), .B(n24646), .Y(n24927) );
  NAND2xp33_ASAP7_75t_SRAM U37127 ( .A(n18567), .B(n24674), .Y(n25076) );
  NOR2xp33_ASAP7_75t_SL U37128 ( .A(n24695), .B(n31198), .Y(n29523) );
  NOR2xp33_ASAP7_75t_SL U37129 ( .A(n24695), .B(n26136), .Y(n29524) );
  AND2x2_ASAP7_75t_SL U37130 ( .A(n26501), .B(n26130), .Y(n31198) );
  NAND2xp33_ASAP7_75t_SRAM U37131 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__25_), .B(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__29_), .Y(n25558) );
  NOR2xp33_ASAP7_75t_SL U37132 ( .A(n29345), .B(n29359), .Y(n29349) );
  NOR2xp33_ASAP7_75t_SL U37133 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_VALID_), 
        .B(n32270), .Y(n32271) );
  NOR2xp33_ASAP7_75t_SL U37134 ( .A(n26088), .B(n28030), .Y(uart1_v_TXTICK_)
         );
  NAND2xp33_ASAP7_75t_SRAM U37135 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_), .B(n22379), .Y(n24990) );
  NAND2xp33_ASAP7_75t_SRAM U37136 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), .B(n25697), .Y(n24925) );
  NOR2xp33_ASAP7_75t_SL U37137 ( .A(n32135), .B(n24971), .Y(n24981) );
  NOR2xp33_ASAP7_75t_SL U37138 ( .A(n24970), .B(n32014), .Y(n32135) );
  NOR2xp33_ASAP7_75t_SL U37139 ( .A(n25151), .B(n22427), .Y(n32132) );
  NOR2xp33_ASAP7_75t_SL U37140 ( .A(n29399), .B(n29424), .Y(n29630) );
  NOR2xp33_ASAP7_75t_SL U37141 ( .A(n29658), .B(n29659), .Y(n29636) );
  NOR2xp33_ASAP7_75t_SL U37142 ( .A(n4775), .B(n29418), .Y(n29414) );
  NOR2xp33_ASAP7_75t_SL U37143 ( .A(n29628), .B(n29627), .Y(n29664) );
  NOR2xp33_ASAP7_75t_SL U37144 ( .A(n29633), .B(n29635), .Y(n29442) );
  NOR2xp33_ASAP7_75t_SL U37145 ( .A(n29444), .B(n29450), .Y(n29441) );
  NOR2xp33_ASAP7_75t_SL U37146 ( .A(n29461), .B(n29460), .Y(n29436) );
  NOR2xp33_ASAP7_75t_SL U37147 ( .A(n30552), .B(n29631), .Y(n29460) );
  NOR2xp33_ASAP7_75t_SL U37148 ( .A(n29428), .B(n29632), .Y(n29461) );
  NOR2xp33_ASAP7_75t_SL U37149 ( .A(n29427), .B(n29462), .Y(n29435) );
  NOR2xp33_ASAP7_75t_SL U37150 ( .A(n29426), .B(n29629), .Y(n29462) );
  NOR2xp33_ASAP7_75t_SL U37151 ( .A(n29425), .B(n29424), .Y(n29427) );
  NOR2xp33_ASAP7_75t_SL U37152 ( .A(irqctrl0_r_IPEND__12_), .B(
        irqctrl0_r_IFORCE__0__12_), .Y(n29424) );
  NOR2xp33_ASAP7_75t_SL U37153 ( .A(n29456), .B(n29457), .Y(n29438) );
  NOR2xp33_ASAP7_75t_SL U37154 ( .A(n2236), .B(n29433), .Y(n29457) );
  NOR2xp33_ASAP7_75t_SL U37155 ( .A(n30984), .B(n29432), .Y(n29456) );
  AOI31xp33_ASAP7_75t_SL U37156 ( .A1(irqctrl0_r_IMASK__0__8_), .A2(
        irqctrl0_r_ILEVEL__8_), .A3(n29431), .B(n29458), .Y(n29434) );
  NOR2xp33_ASAP7_75t_SL U37157 ( .A(n29430), .B(n29429), .Y(n29458) );
  NOR2xp33_ASAP7_75t_SL U37158 ( .A(n29404), .B(n29403), .Y(n29422) );
  NOR2xp33_ASAP7_75t_SL U37159 ( .A(irqctrl0_r_IPEND__5_), .B(
        irqctrl0_r_IFORCE__0__5_), .Y(n29403) );
  NOR2xp33_ASAP7_75t_SL U37160 ( .A(n29402), .B(n29401), .Y(n29421) );
  NOR2xp33_ASAP7_75t_SL U37161 ( .A(irqctrl0_r_IPEND__4_), .B(
        irqctrl0_r_IFORCE__0__4_), .Y(n29401) );
  NOR2xp33_ASAP7_75t_SL U37162 ( .A(n29453), .B(n29452), .Y(n29423) );
  NOR2xp33_ASAP7_75t_SL U37163 ( .A(n29420), .B(n29419), .Y(n29452) );
  NOR2xp33_ASAP7_75t_SL U37164 ( .A(n29418), .B(n24536), .Y(n29453) );
  NOR2xp33_ASAP7_75t_SL U37165 ( .A(irqctrl0_r_IPEND__7_), .B(
        irqctrl0_r_IFORCE__0__7_), .Y(n29418) );
  NOR2xp33_ASAP7_75t_SL U37166 ( .A(n29416), .B(n29415), .Y(n29447) );
  NOR2xp33_ASAP7_75t_SL U37167 ( .A(n29411), .B(n29410), .Y(n29660) );
  NOR2xp33_ASAP7_75t_SL U37168 ( .A(n29409), .B(n29408), .Y(n29411) );
  NOR2xp33_ASAP7_75t_SL U37169 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__5_), 
        .B(n24646), .Y(n30114) );
  NOR2xp33_ASAP7_75t_SL U37170 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__7_), 
        .B(n24646), .Y(n28759) );
  NOR2xp33_ASAP7_75t_SL U37171 ( .A(n32066), .B(n24510), .Y(n31440) );
  NOR2xp33_ASAP7_75t_SL U37172 ( .A(n24695), .B(n27464), .Y(n25849) );
  NOR2xp33_ASAP7_75t_SL U37173 ( .A(n26131), .B(n28119), .Y(n26132) );
  NOR2xp33_ASAP7_75t_SL U37174 ( .A(n24695), .B(n25991), .Y(n17459) );
  NOR2xp33_ASAP7_75t_SL U37175 ( .A(n30780), .B(n31501), .Y(n30778) );
  NOR2xp33_ASAP7_75t_SL U37176 ( .A(n30073), .B(n31501), .Y(n30072) );
  NOR2xp33_ASAP7_75t_SL U37177 ( .A(n24695), .B(n28030), .Y(n26085) );
  NOR2xp33_ASAP7_75t_SL U37178 ( .A(n5014), .B(n26086), .Y(n26087) );
  NOR2xp33_ASAP7_75t_SL U37179 ( .A(n30777), .B(n30776), .Y(n1734) );
  NOR4xp25_ASAP7_75t_SL U37180 ( .A(n30774), .B(uart1_r_RSEMPTY_), .C(n24695), 
        .D(n30980), .Y(n30777) );
  AOI211xp5_ASAP7_75t_SL U37181 ( .A1(n32983), .A2(n32938), .B(n32937), .C(
        n32936), .Y(n1692) );
  NOR2xp33_ASAP7_75t_SL U37182 ( .A(n32979), .B(n32935), .Y(n32936) );
  AOI211xp5_ASAP7_75t_SL U37183 ( .A1(n32983), .A2(n32946), .B(n32945), .C(
        n32944), .Y(n1691) );
  NOR2xp33_ASAP7_75t_SL U37184 ( .A(n32979), .B(n32943), .Y(n32944) );
  AOI211xp5_ASAP7_75t_SL U37185 ( .A1(n32983), .A2(n32954), .B(n32953), .C(
        n32952), .Y(n1690) );
  NOR2xp33_ASAP7_75t_SL U37186 ( .A(n32979), .B(n32951), .Y(n32952) );
  AOI211xp5_ASAP7_75t_SL U37187 ( .A1(n32983), .A2(n32922), .B(n32921), .C(
        n32920), .Y(n1694) );
  NOR2xp33_ASAP7_75t_SL U37188 ( .A(n32979), .B(n32919), .Y(n32920) );
  AOI211xp5_ASAP7_75t_SL U37189 ( .A1(n32983), .A2(n32930), .B(n32929), .C(
        n32928), .Y(n1693) );
  NOR2xp33_ASAP7_75t_SL U37190 ( .A(n32979), .B(n32927), .Y(n32928) );
  AOI211xp5_ASAP7_75t_SL U37191 ( .A1(n32983), .A2(n32962), .B(n32961), .C(
        n32960), .Y(n1689) );
  NOR2xp33_ASAP7_75t_SL U37192 ( .A(n32979), .B(n32959), .Y(n32960) );
  AOI211xp5_ASAP7_75t_SL U37193 ( .A1(n32983), .A2(n32982), .B(n32981), .C(
        n32980), .Y(n1687) );
  NOR2xp33_ASAP7_75t_SL U37194 ( .A(n32979), .B(n32978), .Y(n32980) );
  AOI211xp5_ASAP7_75t_SL U37195 ( .A1(n32983), .A2(n32970), .B(n32969), .C(
        n32968), .Y(n1688) );
  NOR2xp33_ASAP7_75t_SL U37196 ( .A(n32979), .B(n32967), .Y(n32968) );
  NOR2xp33_ASAP7_75t_SL U37197 ( .A(n1724), .B(address[1]), .Y(n32917) );
  AOI211xp5_ASAP7_75t_SL U37198 ( .A1(address[0]), .A2(n32884), .B(n22433), 
        .C(n32885), .Y(n32972) );
  NOR2xp33_ASAP7_75t_SL U37199 ( .A(n1723), .B(address[0]), .Y(n32837) );
  AND2x2_ASAP7_75t_SL U37200 ( .A(datadir[0]), .B(n32832), .Y(n24527) );
  NOR2xp33_ASAP7_75t_SL U37201 ( .A(u0_0_leon3x0_p0_iu_r_A__RFA1__4_), .B(
        n23229), .Y(n32182) );
  NAND2xp33_ASAP7_75t_SRAM U37202 ( .A(n30066), .B(n30065), .Y(n30070) );
  NOR2xp33_ASAP7_75t_SL U37203 ( .A(n29337), .B(n29336), .Y(n30071) );
  AOI31xp33_ASAP7_75t_SL U37204 ( .A1(n28235), .A2(n31194), .A3(n31193), .B(
        n28234), .Y(n1746) );
  AOI31xp33_ASAP7_75t_SL U37205 ( .A1(n31194), .A2(n31193), .A3(n31192), .B(
        n31191), .Y(n1747) );
  NOR2xp33_ASAP7_75t_SL U37206 ( .A(uart1_v_RXDB__1_), .B(n24695), .Y(n31193)
         );
  NOR2xp33_ASAP7_75t_SL U37207 ( .A(n29243), .B(n29745), .Y(n29247) );
  NOR2xp33_ASAP7_75t_SL U37208 ( .A(n25964), .B(n29745), .Y(n25968) );
  AOI211xp5_ASAP7_75t_SL U37209 ( .A1(uart1_r_RSHIFT__1_), .A2(n29959), .B(
        n29958), .C(n29957), .Y(n2865) );
  NOR2xp33_ASAP7_75t_SL U37210 ( .A(n29956), .B(n29955), .Y(n29957) );
  NOR2xp33_ASAP7_75t_SL U37211 ( .A(n27528), .B(n27539), .Y(n26091) );
  NOR2xp33_ASAP7_75t_SL U37212 ( .A(n26090), .B(n29971), .Y(n27528) );
  NOR2xp33_ASAP7_75t_SL U37213 ( .A(uart1_r_RXTICK_), .B(n26095), .Y(n26093)
         );
  NOR2xp33_ASAP7_75t_SL U37214 ( .A(n29966), .B(n29961), .Y(n26095) );
  NOR2xp33_ASAP7_75t_SL U37215 ( .A(uart1_r_RXSTATE__0_), .B(n29971), .Y(
        n29961) );
  NOR2xp33_ASAP7_75t_SL U37216 ( .A(n24942), .B(n24941), .Y(n24950) );
  NOR2xp33_ASAP7_75t_SL U37217 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__CNT__1_), 
        .B(n24993), .Y(n24936) );
  NOR2xp33_ASAP7_75t_SL U37218 ( .A(irqctrl0_r_IFORCE__0__8_), .B(n29742), .Y(
        n15074) );
  NOR2xp33_ASAP7_75t_SL U37219 ( .A(n24902), .B(n24901), .Y(n24905) );
  AND2x2_ASAP7_75t_SL U37220 ( .A(n24694), .B(n31501), .Y(n31735) );
  NOR2xp33_ASAP7_75t_SL U37221 ( .A(n28583), .B(n30580), .Y(n28584) );
  NOR2xp33_ASAP7_75t_SL U37222 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__14_), .B(
        n22379), .Y(n28583) );
  NOR2xp33_ASAP7_75t_SL U37223 ( .A(n29396), .B(n29395), .Y(n29397) );
  NOR2xp33_ASAP7_75t_SL U37224 ( .A(irqctrl0_r_IPEND__15_), .B(n29745), .Y(
        n29395) );
  NOR2xp33_ASAP7_75t_SL U37225 ( .A(apbi[15]), .B(n29745), .Y(n29398) );
  AOI211xp5_ASAP7_75t_SL U37226 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__12_), .A2(
        n22429), .B(n30374), .C(n30373), .Y(n30375) );
  NOR2xp33_ASAP7_75t_SL U37227 ( .A(n30371), .B(n24638), .Y(n30374) );
  AOI211xp5_ASAP7_75t_SL U37228 ( .A1(u0_0_leon3x0_p0_muli[3]), .A2(n22429), 
        .B(n30443), .C(n30442), .Y(n30444) );
  NOR2xp33_ASAP7_75t_SL U37229 ( .A(n30440), .B(n24638), .Y(n30443) );
  NOR2xp33_ASAP7_75t_SL U37230 ( .A(n22378), .B(n27147), .Y(n30387) );
  NOR2xp33_ASAP7_75t_SL U37231 ( .A(n29876), .B(n29875), .Y(n30702) );
  NAND2xp33_ASAP7_75t_SRAM U37232 ( .A(n25693), .B(n25692), .Y(n25694) );
  NOR4xp25_ASAP7_75t_SL U37233 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__22_), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__5_), .C(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__7_), .D(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__9_), .Y(n25679) );
  AOI211xp5_ASAP7_75t_SL U37234 ( .A1(n25705), .A2(n25674), .B(n25673), .C(
        n25672), .Y(n29225) );
  AOI211xp5_ASAP7_75t_SL U37235 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_), 
        .A2(n30956), .B(n25680), .C(n25665), .Y(n25673) );
  NOR2xp33_ASAP7_75t_SL U37236 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), 
        .B(n25670), .Y(n25682) );
  NAND2xp33_ASAP7_75t_SRAM U37237 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), .B(n25692), .Y(n25664) );
  NOR2xp33_ASAP7_75t_SL U37238 ( .A(n25657), .B(n25656), .Y(n29700) );
  NOR2xp33_ASAP7_75t_SL U37239 ( .A(n25651), .B(n25650), .Y(n25657) );
  NOR2xp33_ASAP7_75t_SL U37240 ( .A(u0_0_leon3x0_p0_iu_r_A__WOVF_), .B(
        u0_0_leon3x0_p0_iu_r_A__WUNF_), .Y(n29873) );
  NOR2xp33_ASAP7_75t_SL U37241 ( .A(n26355), .B(n26354), .Y(n32161) );
  NOR2xp33_ASAP7_75t_SL U37242 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), .B(
        n30701), .Y(n30655) );
  AOI211xp5_ASAP7_75t_SL U37243 ( .A1(n2267), .A2(n27307), .B(n24695), .C(
        n27308), .Y(n17717) );
  NOR2xp33_ASAP7_75t_SL U37244 ( .A(n28613), .B(n30580), .Y(n28614) );
  NOR2xp33_ASAP7_75t_SL U37245 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__12_), .B(
        n22379), .Y(n28613) );
  NOR2xp33_ASAP7_75t_SL U37246 ( .A(n28962), .B(n30814), .Y(n28963) );
  NOR2xp33_ASAP7_75t_SL U37247 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__0_), .B(
        n30813), .Y(n28962) );
  AOI211xp5_ASAP7_75t_SL U37248 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__30_), .A2(
        n22429), .B(n30217), .C(n30216), .Y(n30218) );
  NOR2xp33_ASAP7_75t_SL U37249 ( .A(n30215), .B(n24638), .Y(n30217) );
  AOI211xp5_ASAP7_75t_SL U37250 ( .A1(u0_0_dbgo_SU_), .A2(n24646), .B(n29737), 
        .C(n29217), .Y(n3366) );
  NOR2xp33_ASAP7_75t_SL U37251 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__11_), 
        .B(n24646), .Y(n29207) );
  AOI211xp5_ASAP7_75t_SL U37252 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__20_), .A2(
        n22429), .B(n30289), .C(n30288), .Y(n30290) );
  NOR2xp33_ASAP7_75t_SL U37253 ( .A(n30286), .B(n24638), .Y(n30289) );
  AOI211xp5_ASAP7_75t_SL U37254 ( .A1(n29521), .A2(timer0_scaler_5_), .B(
        n25869), .C(n25868), .Y(n1638) );
  NOR2xp33_ASAP7_75t_SL U37255 ( .A(n25867), .B(n29517), .Y(n25868) );
  AOI211xp5_ASAP7_75t_SL U37256 ( .A1(n29521), .A2(timer0_scaler_6_), .B(
        n25866), .C(n25865), .Y(n1726) );
  NOR2xp33_ASAP7_75t_SL U37257 ( .A(n25864), .B(n29517), .Y(n25865) );
  AOI211xp5_ASAP7_75t_SL U37258 ( .A1(n29521), .A2(timer0_scaler_1_), .B(
        n26135), .C(n26134), .Y(n2230) );
  NOR2xp33_ASAP7_75t_SL U37259 ( .A(n26133), .B(n29517), .Y(n26134) );
  AOI211xp5_ASAP7_75t_SL U37260 ( .A1(n29521), .A2(timer0_scaler_4_), .B(
        n25880), .C(n25879), .Y(n1628) );
  NOR2xp33_ASAP7_75t_SL U37261 ( .A(n25878), .B(n29517), .Y(n25879) );
  AOI211xp5_ASAP7_75t_SL U37262 ( .A1(n29521), .A2(timer0_scaler_2_), .B(
        n29520), .C(n29519), .Y(n1749) );
  NOR2xp33_ASAP7_75t_SL U37263 ( .A(n29518), .B(n29517), .Y(n29519) );
  AOI211xp5_ASAP7_75t_SL U37264 ( .A1(n29521), .A2(timer0_scaler_3_), .B(
        n29513), .C(n29512), .Y(n1739) );
  NOR2xp33_ASAP7_75t_SL U37265 ( .A(n29511), .B(n29517), .Y(n29512) );
  NAND2xp33_ASAP7_75t_SRAM U37266 ( .A(n2929), .B(n30555), .Y(n25850) );
  NOR2xp33_ASAP7_75t_SL U37267 ( .A(n25721), .B(n26354), .Y(n29737) );
  NAND2xp33_ASAP7_75t_SRAM U37268 ( .A(n30115), .B(n26352), .Y(n25721) );
  NOR2xp33_ASAP7_75t_SL U37269 ( .A(n32076), .B(n29738), .Y(n25725) );
  NOR2xp33_ASAP7_75t_SL U37270 ( .A(irqctrl0_r_IPEND__5_), .B(n29745), .Y(
        n29298) );
  NOR2xp33_ASAP7_75t_SL U37271 ( .A(n30073), .B(n29376), .Y(n29302) );
  NOR2xp33_ASAP7_75t_SL U37272 ( .A(irqctrl0_r_IPEND__4_), .B(n29745), .Y(
        n29320) );
  NOR2xp33_ASAP7_75t_SL U37273 ( .A(n30780), .B(n29376), .Y(n29324) );
  NOR2xp33_ASAP7_75t_SL U37274 ( .A(n29284), .B(n29283), .Y(n29285) );
  NOR2xp33_ASAP7_75t_SL U37275 ( .A(irqctrl0_r_IPEND__7_), .B(n29745), .Y(
        n29283) );
  NOR2xp33_ASAP7_75t_SL U37276 ( .A(n30833), .B(n29376), .Y(n29286) );
  NOR2xp33_ASAP7_75t_SL U37277 ( .A(irqctrl0_r_IPEND__6_), .B(n29745), .Y(
        n29311) );
  NOR2xp33_ASAP7_75t_SL U37278 ( .A(n31197), .B(n29376), .Y(n29315) );
  NOR2xp33_ASAP7_75t_SL U37279 ( .A(irqctrl0_r_IPEND__3_), .B(n29745), .Y(
        n28241) );
  NOR2xp33_ASAP7_75t_SL U37280 ( .A(n29510), .B(n29376), .Y(n28245) );
  NOR2xp33_ASAP7_75t_SL U37281 ( .A(irqctrl0_r_IPEND__10_), .B(n29745), .Y(
        n29265) );
  NOR2xp33_ASAP7_75t_SL U37282 ( .A(n30978), .B(n29376), .Y(n29269) );
  NOR2xp33_ASAP7_75t_SL U37283 ( .A(n28588), .B(n30580), .Y(n28589) );
  AND2x2_ASAP7_75t_SL U37284 ( .A(n25938), .B(n30813), .Y(n30580) );
  NOR2xp33_ASAP7_75t_SL U37285 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__13_), .B(
        n22379), .Y(n28588) );
  NOR2xp33_ASAP7_75t_SL U37286 ( .A(n30815), .B(n30814), .Y(n30816) );
  NOR2xp33_ASAP7_75t_SL U37287 ( .A(n24646), .B(n30813), .Y(n30814) );
  NOR2xp33_ASAP7_75t_SL U37288 ( .A(u0_0_leon3x0_p0_iu_r_A__IMM__3_), .B(
        n30813), .Y(n30815) );
  NOR2xp33_ASAP7_75t_SL U37289 ( .A(n24684), .B(n24677), .Y(n32076) );
  AOI211xp5_ASAP7_75t_SL U37290 ( .A1(n2386), .A2(n25996), .B(n24695), .C(
        n25997), .Y(n17456) );
  NOR2xp33_ASAP7_75t_SL U37291 ( .A(n2389), .B(n2388), .Y(n25992) );
  NOR2xp33_ASAP7_75t_SL U37292 ( .A(n30680), .B(n31814), .Y(n32065) );
  NOR2xp33_ASAP7_75t_SL U37293 ( .A(n18800), .B(n32705), .Y(n31625) );
  NOR2xp33_ASAP7_75t_SL U37294 ( .A(n2267), .B(n27307), .Y(n27308) );
  AOI211xp5_ASAP7_75t_SL U37295 ( .A1(n32008), .A2(n31855), .B(n31854), .C(
        n31853), .Y(n4384) );
  NOR2xp33_ASAP7_75t_SL U37296 ( .A(n31852), .B(n32004), .Y(n31853) );
  AOI211xp5_ASAP7_75t_SL U37297 ( .A1(n32008), .A2(n31978), .B(n31977), .C(
        n31976), .Y(n4413) );
  NOR2xp33_ASAP7_75t_SL U37298 ( .A(n31975), .B(n32004), .Y(n31976) );
  AOI211xp5_ASAP7_75t_SL U37299 ( .A1(n32008), .A2(n31535), .B(n31534), .C(
        n31533), .Y(n4496) );
  NOR2xp33_ASAP7_75t_SL U37300 ( .A(n31532), .B(n32004), .Y(n31533) );
  AOI211xp5_ASAP7_75t_SL U37301 ( .A1(n32008), .A2(n26505), .B(n26504), .C(
        n26503), .Y(n4513) );
  NOR2xp33_ASAP7_75t_SL U37302 ( .A(n26520), .B(n32004), .Y(n26503) );
  AOI211xp5_ASAP7_75t_SL U37303 ( .A1(n32008), .A2(n32007), .B(n24540), .C(
        n32006), .Y(n4362) );
  NOR2xp33_ASAP7_75t_SL U37304 ( .A(n32005), .B(n32004), .Y(n32006) );
  AOI211xp5_ASAP7_75t_SL U37305 ( .A1(n32008), .A2(n31376), .B(n31375), .C(
        n31374), .Y(n4623) );
  NOR2xp33_ASAP7_75t_SL U37306 ( .A(n31373), .B(n32004), .Y(n31374) );
  AOI211xp5_ASAP7_75t_SL U37307 ( .A1(n32008), .A2(n31507), .B(n31506), .C(
        n31505), .Y(n4596) );
  NOR2xp33_ASAP7_75t_SL U37308 ( .A(n31504), .B(n32004), .Y(n31505) );
  AOI211xp5_ASAP7_75t_SL U37309 ( .A1(n32008), .A2(n31649), .B(n31648), .C(
        n31647), .Y(n4572) );
  NOR2xp33_ASAP7_75t_SL U37310 ( .A(n31646), .B(n32004), .Y(n31647) );
  AOI211xp5_ASAP7_75t_SL U37311 ( .A1(n32008), .A2(n26662), .B(n26661), .C(
        n26660), .Y(n1770) );
  NOR2xp33_ASAP7_75t_SL U37312 ( .A(n26659), .B(n32004), .Y(n26660) );
  AOI211xp5_ASAP7_75t_SL U37313 ( .A1(n32008), .A2(n31331), .B(n31330), .C(
        n31329), .Y(n4613) );
  NOR2xp33_ASAP7_75t_SL U37314 ( .A(n31328), .B(n32004), .Y(n31329) );
  AOI211xp5_ASAP7_75t_SL U37315 ( .A1(n32008), .A2(n30902), .B(n30901), .C(
        n30900), .Y(n4530) );
  NOR2xp33_ASAP7_75t_SL U37316 ( .A(n30899), .B(n32004), .Y(n30900) );
  NOR2xp33_ASAP7_75t_SL U37317 ( .A(n27390), .B(n27313), .Y(n27317) );
  NOR2xp33_ASAP7_75t_SL U37318 ( .A(n29219), .B(n22379), .Y(n29220) );
  NOR2xp33_ASAP7_75t_SL U37319 ( .A(n30554), .B(n30553), .Y(n17066) );
  NOR2xp33_ASAP7_75t_SL U37320 ( .A(n28079), .B(n28078), .Y(n28081) );
  NOR2xp33_ASAP7_75t_SL U37321 ( .A(n28069), .B(n28068), .Y(n28082) );
  NOR2xp33_ASAP7_75t_SL U37322 ( .A(n28026), .B(n28025), .Y(n28084) );
  AOI211xp5_ASAP7_75t_SL U37323 ( .A1(uart1_r_TRADDR__0_), .A2(n28024), .B(
        n28023), .C(n28022), .Y(n28025) );
  AOI211xp5_ASAP7_75t_SL U37324 ( .A1(uart1_r_THOLD__16__0_), .A2(n28010), .B(
        uart1_r_TRADDR__1_), .C(n27988), .Y(n27992) );
  NOR2xp33_ASAP7_75t_SL U37325 ( .A(n27987), .B(n27986), .Y(n27988) );
  NOR2xp33_ASAP7_75t_SL U37326 ( .A(n25566), .B(n29883), .Y(
        u0_0_leon3x0_p0_iu_v_M__WERR_) );
  NOR2xp33_ASAP7_75t_SL U37327 ( .A(n29261), .B(n29260), .Y(n2822) );
  NOR2xp33_ASAP7_75t_SL U37328 ( .A(n29259), .B(n29385), .Y(n29260) );
  NOR2xp33_ASAP7_75t_SL U37329 ( .A(n30978), .B(n29384), .Y(n29261) );
  NOR2xp33_ASAP7_75t_SL U37330 ( .A(n29290), .B(n29289), .Y(n2823) );
  NOR2xp33_ASAP7_75t_SL U37331 ( .A(n29404), .B(n29385), .Y(n29289) );
  NOR2xp33_ASAP7_75t_SL U37332 ( .A(n30073), .B(n29384), .Y(n29290) );
  NOR2xp33_ASAP7_75t_SL U37333 ( .A(n29327), .B(n29326), .Y(n2825) );
  NOR2xp33_ASAP7_75t_SL U37334 ( .A(n29400), .B(n29385), .Y(n29326) );
  NOR2xp33_ASAP7_75t_SL U37335 ( .A(n29568), .B(n29384), .Y(n29327) );
  NOR2xp33_ASAP7_75t_SL U37336 ( .A(n25642), .B(n25641), .Y(n4432) );
  NOR2xp33_ASAP7_75t_SL U37337 ( .A(n25640), .B(n29385), .Y(n25641) );
  NOR2xp33_ASAP7_75t_SL U37338 ( .A(n30547), .B(n29384), .Y(n25642) );
  NOR2xp33_ASAP7_75t_SL U37339 ( .A(n27300), .B(n27299), .Y(n2826) );
  NOR2xp33_ASAP7_75t_SL U37340 ( .A(n27298), .B(n29385), .Y(n27299) );
  NOR2xp33_ASAP7_75t_SL U37341 ( .A(n27493), .B(n29384), .Y(n27300) );
  NOR2xp33_ASAP7_75t_SL U37342 ( .A(n29251), .B(n29250), .Y(n1795) );
  NOR2xp33_ASAP7_75t_SL U37343 ( .A(n29249), .B(n29385), .Y(n29250) );
  NOR2xp33_ASAP7_75t_SL U37344 ( .A(n30139), .B(n29384), .Y(n29251) );
  NOR2xp33_ASAP7_75t_SL U37345 ( .A(n29235), .B(n29234), .Y(n1754) );
  NOR2xp33_ASAP7_75t_SL U37346 ( .A(n30805), .B(n29385), .Y(n29234) );
  NOR2xp33_ASAP7_75t_SL U37347 ( .A(n29236), .B(n29384), .Y(n29235) );
  NOR2xp33_ASAP7_75t_SL U37348 ( .A(n29388), .B(n29387), .Y(n2321) );
  NOR2xp33_ASAP7_75t_SL U37349 ( .A(n29386), .B(n29385), .Y(n29387) );
  NOR2xp33_ASAP7_75t_SL U37350 ( .A(n29389), .B(n29384), .Y(n29388) );
  NOR2xp33_ASAP7_75t_SL U37351 ( .A(n29273), .B(n29272), .Y(n1743) );
  NOR2xp33_ASAP7_75t_SL U37352 ( .A(n29409), .B(n29385), .Y(n29272) );
  NOR2xp33_ASAP7_75t_SL U37353 ( .A(n29744), .B(n29384), .Y(n29273) );
  NOR2xp33_ASAP7_75t_SL U37354 ( .A(n28248), .B(n28247), .Y(n2824) );
  NOR2xp33_ASAP7_75t_SL U37355 ( .A(n28246), .B(n29385), .Y(n28247) );
  NOR2xp33_ASAP7_75t_SL U37356 ( .A(n29510), .B(n29384), .Y(n28248) );
  NOR2xp33_ASAP7_75t_SL U37357 ( .A(n29306), .B(n29305), .Y(n1730) );
  NOR2xp33_ASAP7_75t_SL U37358 ( .A(n29304), .B(n29385), .Y(n29305) );
  NOR2xp33_ASAP7_75t_SL U37359 ( .A(n31197), .B(n29384), .Y(n29306) );
  NOR2xp33_ASAP7_75t_SL U37360 ( .A(n24695), .B(n26468), .Y(n25639) );
  NOR2xp33_ASAP7_75t_SL U37361 ( .A(n27649), .B(n27648), .Y(n31239) );
  AOI211xp5_ASAP7_75t_SL U37362 ( .A1(uart1_r_TRADDR__0_), .A2(n27647), .B(
        n27646), .C(n27645), .Y(n27648) );
  AOI211xp5_ASAP7_75t_SL U37363 ( .A1(uart1_r_THOLD__16__6_), .A2(n28010), .B(
        uart1_r_TRADDR__1_), .C(n27628), .Y(n27632) );
  NOR2xp33_ASAP7_75t_SL U37364 ( .A(n27627), .B(n27986), .Y(n27628) );
  AOI211xp5_ASAP7_75t_SL U37365 ( .A1(n28018), .A2(uart1_r_THOLD__28__3_), .B(
        n27842), .C(n27841), .Y(n27845) );
  AOI211xp5_ASAP7_75t_SL U37366 ( .A1(n28010), .A2(uart1_r_THOLD__18__3_), .B(
        n28016), .C(n24529), .Y(n27833) );
  NOR2xp33_ASAP7_75t_SL U37367 ( .A(n24695), .B(n25966), .Y(n25958) );
  NOR2xp33_ASAP7_75t_SL U37368 ( .A(n29329), .B(n29237), .Y(n25966) );
  AOI211xp5_ASAP7_75t_SL U37369 ( .A1(n32008), .A2(n29859), .B(n29858), .C(
        n29857), .Y(n1633) );
  NOR2xp33_ASAP7_75t_SL U37370 ( .A(n27459), .B(n31323), .Y(n29858) );
  AOI211xp5_ASAP7_75t_SL U37371 ( .A1(n32008), .A2(n31030), .B(n31029), .C(
        n31028), .Y(n4634) );
  NOR2xp33_ASAP7_75t_SL U37372 ( .A(n31021), .B(n32004), .Y(n31029) );
  NOR2xp33_ASAP7_75t_SL U37373 ( .A(n30153), .B(n30152), .Y(n4559) );
  AOI211xp5_ASAP7_75t_SL U37374 ( .A1(n26813), .A2(n26812), .B(n31510), .C(
        n26811), .Y(n26814) );
  NOR2xp33_ASAP7_75t_SL U37375 ( .A(n27785), .B(n27784), .Y(n30782) );
  AOI211xp5_ASAP7_75t_SL U37376 ( .A1(uart1_r_THOLD__26__4_), .A2(n28017), .B(
        n28016), .C(n27776), .Y(n27780) );
  NOR2xp33_ASAP7_75t_SL U37377 ( .A(n27775), .B(n27774), .Y(n27776) );
  AOI211xp5_ASAP7_75t_SL U37378 ( .A1(uart1_r_THOLD__16__4_), .A2(n28010), .B(
        uart1_r_TRADDR__1_), .C(n27760), .Y(n27764) );
  NOR2xp33_ASAP7_75t_SL U37379 ( .A(n27759), .B(n27986), .Y(n27760) );
  NOR2xp33_ASAP7_75t_SL U37380 ( .A(n28178), .B(n28177), .Y(n2872) );
  OR2x2_ASAP7_75t_SL U37381 ( .A(n28167), .B(n28142), .Y(n28179) );
  NOR2xp33_ASAP7_75t_SL U37382 ( .A(n28108), .B(n28056), .Y(n28178) );
  NAND2xp33_ASAP7_75t_SRAM U37383 ( .A(n27474), .B(n28231), .Y(n28056) );
  AOI211xp5_ASAP7_75t_SL U37384 ( .A1(n32517), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__1_), .B(n32470), .C(n32469), 
        .Y(n2286) );
  NOR2xp33_ASAP7_75t_SL U37385 ( .A(n32468), .B(n32513), .Y(n32469) );
  NOR2xp33_ASAP7_75t_SL U37386 ( .A(n32472), .B(n32512), .Y(n32470) );
  AOI211xp5_ASAP7_75t_SL U37387 ( .A1(n32517), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__6_), .B(n32506), .C(n32505), 
        .Y(n2282) );
  NOR2xp33_ASAP7_75t_SL U37388 ( .A(n32504), .B(n32513), .Y(n32505) );
  NOR2xp33_ASAP7_75t_SL U37389 ( .A(n32508), .B(n32512), .Y(n32506) );
  AOI211xp5_ASAP7_75t_SL U37390 ( .A1(n32517), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__5_), .B(n32499), .C(n32498), 
        .Y(n2283) );
  NOR2xp33_ASAP7_75t_SL U37391 ( .A(n32497), .B(n32513), .Y(n32498) );
  NOR2xp33_ASAP7_75t_SL U37392 ( .A(n32501), .B(n32512), .Y(n32499) );
  NOR2xp33_ASAP7_75t_SL U37393 ( .A(u0_0_leon3x0_p0_c0mmu_mcii[1]), .B(n32510), 
        .Y(n32495) );
  AOI211xp5_ASAP7_75t_SL U37394 ( .A1(n32517), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__3_), .B(n32485), .C(n32484), 
        .Y(n2284) );
  NOR2xp33_ASAP7_75t_SL U37395 ( .A(n32483), .B(n32513), .Y(n32484) );
  NOR2xp33_ASAP7_75t_SL U37396 ( .A(n32487), .B(n32512), .Y(n32485) );
  AOI211xp5_ASAP7_75t_SL U37397 ( .A1(n32517), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__2_), .B(n32477), .C(n32476), 
        .Y(n2285) );
  NOR2xp33_ASAP7_75t_SL U37398 ( .A(n32475), .B(n32513), .Y(n32476) );
  NOR2xp33_ASAP7_75t_SL U37399 ( .A(n32479), .B(n32512), .Y(n32477) );
  NOR2xp33_ASAP7_75t_SL U37400 ( .A(n32496), .B(n32503), .Y(n32474) );
  AOI211xp5_ASAP7_75t_SL U37401 ( .A1(n32517), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_VALID__0__7_), .B(n32516), .C(n32515), 
        .Y(n2281) );
  NOR2xp33_ASAP7_75t_SL U37402 ( .A(n32514), .B(n32513), .Y(n32515) );
  NOR2xp33_ASAP7_75t_SL U37403 ( .A(n32492), .B(n32462), .Y(n32513) );
  NOR2xp33_ASAP7_75t_SL U37404 ( .A(n32490), .B(n32512), .Y(n32462) );
  NOR2xp33_ASAP7_75t_SL U37405 ( .A(n32521), .B(n32512), .Y(n32516) );
  NOR2xp33_ASAP7_75t_SL U37406 ( .A(n32492), .B(n32460), .Y(n32517) );
  NOR2xp33_ASAP7_75t_SL U37407 ( .A(n32518), .B(n32512), .Y(n32460) );
  NOR2xp33_ASAP7_75t_SL U37408 ( .A(n32660), .B(n32458), .Y(n32492) );
  OR2x2_ASAP7_75t_SL U37409 ( .A(n32456), .B(n32662), .Y(n32512) );
  NOR2xp33_ASAP7_75t_SL U37410 ( .A(n28130), .B(n28129), .Y(n4524) );
  AOI211xp5_ASAP7_75t_SL U37411 ( .A1(n31950), .A2(n33068), .B(n28124), .C(
        n28123), .Y(n28128) );
  NOR2xp33_ASAP7_75t_SL U37412 ( .A(n2236), .B(n30983), .Y(n28123) );
  NOR2xp33_ASAP7_75t_SL U37413 ( .A(n26003), .B(n25977), .Y(n25978) );
  AOI211xp5_ASAP7_75t_SL U37414 ( .A1(n31240), .A2(n27915), .B(n27488), .C(
        n27487), .Y(n16969) );
  AOI211xp5_ASAP7_75t_SL U37415 ( .A1(n31246), .A2(uart1_r_BRATE__1_), .B(
        n27483), .C(n27482), .Y(n27485) );
  AOI211xp5_ASAP7_75t_SL U37416 ( .A1(timer0_vtimers_1__RELOAD__8_), .A2(
        n30993), .B(n29757), .C(n29756), .Y(n4688) );
  NAND2xp33_ASAP7_75t_SRAM U37417 ( .A(irqctrl0_r_ILEVEL__8_), .B(n31248), .Y(
        n29749) );
  AND2x2_ASAP7_75t_SL U37418 ( .A(n31954), .B(n31235), .Y(n32003) );
  AOI211xp5_ASAP7_75t_SL U37419 ( .A1(timer0_vtimers_1__RELOAD__10_), .A2(
        n30993), .B(n30992), .C(n30991), .Y(n4455) );
  AOI211xp5_ASAP7_75t_SL U37420 ( .A1(n31950), .A2(uart1_r_RFIFOIRQEN_), .B(
        n30986), .C(n30985), .Y(n30990) );
  NOR2xp33_ASAP7_75t_SL U37421 ( .A(n30984), .B(n30983), .Y(n30985) );
  NOR2xp33_ASAP7_75t_SL U37422 ( .A(n2931), .B(n31323), .Y(n31849) );
  NOR2xp33_ASAP7_75t_SL U37423 ( .A(n26812), .B(n26813), .Y(n26811) );
  NOR2xp33_ASAP7_75t_SL U37424 ( .A(n29329), .B(n29328), .Y(n29379) );
  NOR2xp33_ASAP7_75t_SL U37425 ( .A(n29316), .B(n29328), .Y(n29322) );
  AOI211xp5_ASAP7_75t_SL U37426 ( .A1(n28010), .A2(uart1_r_THOLD__18__2_), .B(
        n28016), .C(n24520), .Y(n27909) );
  AOI211xp5_ASAP7_75t_SL U37427 ( .A1(uart1_r_THOLD__16__2_), .A2(n28010), .B(
        uart1_r_TRADDR__1_), .C(n27901), .Y(n27905) );
  NOR2xp33_ASAP7_75t_SL U37428 ( .A(n27900), .B(n27986), .Y(n27901) );
  NOR2xp33_ASAP7_75t_SL U37429 ( .A(n28833), .B(n29239), .Y(n29390) );
  NOR2xp33_ASAP7_75t_SL U37430 ( .A(n29654), .B(n29328), .Y(n29313) );
  NOR2xp33_ASAP7_75t_SL U37431 ( .A(irqo[1]), .B(n27294), .Y(n29275) );
  AOI211xp5_ASAP7_75t_SL U37432 ( .A1(u0_0_leon3x0_p0_iu_r_X__Y__31_), .A2(
        n22429), .B(n31409), .C(n31408), .Y(n31410) );
  NOR2xp33_ASAP7_75t_SL U37433 ( .A(n31407), .B(n24638), .Y(n31408) );
  NOR2xp33_ASAP7_75t_SL U37434 ( .A(n22378), .B(n31401), .Y(n31411) );
  NOR2xp33_ASAP7_75t_SL U37435 ( .A(n24679), .B(n30453), .Y(n31412) );
  NOR2xp33_ASAP7_75t_SL U37436 ( .A(n29654), .B(n29653), .Y(n29656) );
  OR2x2_ASAP7_75t_SL U37437 ( .A(n24695), .B(n27293), .Y(n29651) );
  NOR2xp33_ASAP7_75t_SL U37438 ( .A(n26468), .B(n25954), .Y(n25963) );
  NOR2xp33_ASAP7_75t_SL U37439 ( .A(n29208), .B(n29211), .Y(n29209) );
  OR2x2_ASAP7_75t_SL U37440 ( .A(n24658), .B(n32153), .Y(n32075) );
  AOI211xp5_ASAP7_75t_SL U37441 ( .A1(n31241), .A2(uart1_r_RHOLD__24__5_), .B(
        n30112), .C(n30111), .Y(n16599) );
  AOI211xp5_ASAP7_75t_SL U37442 ( .A1(n30105), .A2(n30789), .B(n30104), .C(
        n30103), .Y(n30110) );
  AND2x2_ASAP7_75t_SL U37443 ( .A(n28232), .B(n27473), .Y(n31951) );
  AND2x2_ASAP7_75t_SL U37444 ( .A(n27474), .B(n27473), .Y(n31246) );
  NOR2xp33_ASAP7_75t_SL U37445 ( .A(n30099), .B(n30098), .Y(n30101) );
  NOR2xp33_ASAP7_75t_SL U37446 ( .A(n27446), .B(n27439), .Y(n31220) );
  NOR2xp33_ASAP7_75t_SL U37447 ( .A(n27449), .B(n27450), .Y(n31221) );
  NOR2xp33_ASAP7_75t_SL U37448 ( .A(n27449), .B(n27438), .Y(n31218) );
  NOR2xp33_ASAP7_75t_SL U37449 ( .A(n27451), .B(n27439), .Y(n31219) );
  NOR2xp33_ASAP7_75t_SL U37450 ( .A(n27451), .B(n27437), .Y(n31216) );
  NOR2xp33_ASAP7_75t_SL U37451 ( .A(n27446), .B(n27450), .Y(n31217) );
  NOR2xp33_ASAP7_75t_SL U37452 ( .A(n27469), .B(n27437), .Y(n31214) );
  NOR2xp33_ASAP7_75t_SL U37453 ( .A(n27446), .B(n27471), .Y(n31215) );
  NOR2xp33_ASAP7_75t_SL U37454 ( .A(n27451), .B(n27450), .Y(n31230) );
  NOR2xp33_ASAP7_75t_SL U37455 ( .A(n27449), .B(n27448), .Y(n31229) );
  NOR2xp33_ASAP7_75t_SL U37456 ( .A(n27469), .B(n27447), .Y(n31227) );
  NOR2xp33_ASAP7_75t_SL U37457 ( .A(n27448), .B(n27451), .Y(n31228) );
  NOR2xp33_ASAP7_75t_SL U37458 ( .A(n27451), .B(n27447), .Y(n31225) );
  NOR2xp33_ASAP7_75t_SL U37459 ( .A(n27449), .B(n27470), .Y(n31226) );
  NOR2xp33_ASAP7_75t_SL U37460 ( .A(n27451), .B(n27470), .Y(n31223) );
  NOR2xp33_ASAP7_75t_SL U37461 ( .A(n27446), .B(n27470), .Y(n31224) );
  NOR2xp33_ASAP7_75t_SL U37462 ( .A(n30089), .B(n30088), .Y(n30102) );
  NOR2xp33_ASAP7_75t_SL U37463 ( .A(n27449), .B(n27439), .Y(n31213) );
  NOR2xp33_ASAP7_75t_SL U37464 ( .A(n27451), .B(n27471), .Y(n31212) );
  NOR2xp33_ASAP7_75t_SL U37465 ( .A(n27446), .B(n27438), .Y(n31210) );
  NOR2xp33_ASAP7_75t_SL U37466 ( .A(n27446), .B(n27448), .Y(n31211) );
  NOR2xp33_ASAP7_75t_SL U37467 ( .A(n27451), .B(n27438), .Y(n31208) );
  NOR2xp33_ASAP7_75t_SL U37468 ( .A(n27469), .B(n27450), .Y(n31209) );
  NOR2xp33_ASAP7_75t_SL U37469 ( .A(n27469), .B(n27438), .Y(n31206) );
  NOR2xp33_ASAP7_75t_SL U37470 ( .A(n27449), .B(n27437), .Y(n31207) );
  NOR2xp33_ASAP7_75t_SL U37471 ( .A(n27469), .B(n27439), .Y(n31204) );
  NOR2xp33_ASAP7_75t_SL U37472 ( .A(n2389), .B(n2386), .Y(n27427) );
  NOR2xp33_ASAP7_75t_SL U37473 ( .A(n27469), .B(n27448), .Y(n31205) );
  NOR2xp33_ASAP7_75t_SL U37474 ( .A(n27446), .B(n27447), .Y(n31202) );
  NOR2xp33_ASAP7_75t_SL U37475 ( .A(n27449), .B(n27447), .Y(n31203) );
  NOR2xp33_ASAP7_75t_SL U37476 ( .A(n27446), .B(n27437), .Y(n31200) );
  NOR2xp33_ASAP7_75t_SL U37477 ( .A(n2389), .B(n27445), .Y(n27426) );
  NOR2xp33_ASAP7_75t_SL U37478 ( .A(n27449), .B(n27471), .Y(n31201) );
  NOR2xp33_ASAP7_75t_SL U37479 ( .A(n27479), .B(n27478), .Y(n31235) );
  NOR2xp33_ASAP7_75t_SL U37480 ( .A(n27477), .B(n27478), .Y(n31250) );
  NOR2xp33_ASAP7_75t_SL U37481 ( .A(n27476), .B(n27475), .Y(n27478) );
  AND2x2_ASAP7_75t_SL U37482 ( .A(n27459), .B(n27473), .Y(n31950) );
  NOR2xp33_ASAP7_75t_SL U37483 ( .A(n31848), .B(n27477), .Y(n28232) );
  NOR2xp33_ASAP7_75t_SL U37484 ( .A(n25635), .B(n25954), .Y(n27462) );
  NOR2xp33_ASAP7_75t_SL U37485 ( .A(apbi[34]), .B(n25984), .Y(n25634) );
  AOI211xp5_ASAP7_75t_SL U37486 ( .A1(n28018), .A2(uart1_r_THOLD__30__5_), .B(
        n27706), .C(n27705), .Y(n27709) );
  AOI211xp5_ASAP7_75t_SL U37487 ( .A1(n28017), .A2(uart1_r_THOLD__24__5_), .B(
        uart1_r_TRADDR__1_), .C(n24522), .Y(n27697) );
  NOR2xp33_ASAP7_75t_SL U37488 ( .A(n25999), .B(n26015), .Y(n26044) );
  NOR2xp33_ASAP7_75t_SL U37489 ( .A(n2456), .B(n26003), .Y(n25998) );
  NOR2xp33_ASAP7_75t_SL U37490 ( .A(n29369), .B(n26039), .Y(n26038) );
  INVx1_ASAP7_75t_SL U37491 ( .A(n25975), .Y(n26039) );
  NOR2xp33_ASAP7_75t_SL U37492 ( .A(n26068), .B(n29369), .Y(n26065) );
  NOR2xp33_ASAP7_75t_SL U37493 ( .A(uart1_r_RWADDR__2_), .B(n26021), .Y(n26068) );
  NOR2xp33_ASAP7_75t_SL U37494 ( .A(n26032), .B(n29369), .Y(n26031) );
  NOR2xp33_ASAP7_75t_SL U37495 ( .A(uart1_r_RWADDR__2_), .B(n26001), .Y(n26032) );
  NOR2xp33_ASAP7_75t_SL U37496 ( .A(n26062), .B(n29369), .Y(n26059) );
  NOR2xp33_ASAP7_75t_SL U37497 ( .A(n26045), .B(n29369), .Y(n26042) );
  NOR2xp33_ASAP7_75t_SL U37498 ( .A(n25981), .B(n26015), .Y(n26054) );
  NOR2xp33_ASAP7_75t_SL U37499 ( .A(uart1_r_RWADDR__4_), .B(n26004), .Y(n25980) );
  NOR2xp33_ASAP7_75t_SL U37500 ( .A(n26049), .B(n29369), .Y(n26048) );
  NOR2xp33_ASAP7_75t_SL U37501 ( .A(n26006), .B(n26015), .Y(n26067) );
  NOR2xp33_ASAP7_75t_SL U37502 ( .A(n26004), .B(n26003), .Y(n26005) );
  NOR2xp33_ASAP7_75t_SL U37503 ( .A(n26055), .B(n29369), .Y(n26052) );
  NOR2xp33_ASAP7_75t_SL U37504 ( .A(n26016), .B(n26015), .Y(n26061) );
  NOR2xp33_ASAP7_75t_SL U37505 ( .A(n2456), .B(uart1_r_RWADDR__4_), .Y(n26013)
         );
  NOR2xp33_ASAP7_75t_SL U37506 ( .A(n26036), .B(n29369), .Y(n26035) );
  NOR2xp33_ASAP7_75t_SL U37507 ( .A(n30977), .B(n30976), .Y(n4476) );
  NOR2xp33_ASAP7_75t_SL U37508 ( .A(n22393), .B(n33002), .Y(n30976) );
  NOR2xp33_ASAP7_75t_SL U37509 ( .A(n30975), .B(n32705), .Y(n30977) );
  AOI31xp33_ASAP7_75t_SL U37510 ( .A1(n29375), .A2(n29374), .A3(n29373), .B(
        n29372), .Y(n1757) );
  AOI31xp33_ASAP7_75t_SL U37511 ( .A1(n29367), .A2(uart1_r_TSEMPTYIRQEN_), 
        .A3(n29366), .B(n29365), .Y(n29368) );
  NOR2xp33_ASAP7_75t_SL U37512 ( .A(n4519), .B(n27581), .Y(n29367) );
  NOR2xp33_ASAP7_75t_SL U37513 ( .A(n22380), .B(n32705), .Y(n32042) );
  NOR2xp33_ASAP7_75t_SL U37514 ( .A(n29195), .B(n31014), .Y(n29194) );
  NOR2xp33_ASAP7_75t_SL U37515 ( .A(n30429), .B(n29198), .Y(n29192) );
  NOR2xp33_ASAP7_75t_SL U37516 ( .A(n29191), .B(n31437), .Y(n29203) );
  NOR2xp33_ASAP7_75t_SL U37517 ( .A(n31423), .B(n29198), .Y(n29190) );
  NOR2xp33_ASAP7_75t_SL U37518 ( .A(n30439), .B(n29198), .Y(n29185) );
  NOR2xp33_ASAP7_75t_SL U37519 ( .A(n29195), .B(n30796), .Y(n29184) );
  NOR2xp33_ASAP7_75t_SL U37520 ( .A(n30418), .B(n29198), .Y(n29182) );
  NOR2xp33_ASAP7_75t_SL U37521 ( .A(n29191), .B(n31347), .Y(n29189) );
  NOR2xp33_ASAP7_75t_SL U37522 ( .A(n29180), .B(n29198), .Y(n29181) );
  NAND3xp33_ASAP7_75t_SL U37523 ( .A(n29179), .B(n29178), .C(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__20_), .Y(n29198) );
  AOI31xp33_ASAP7_75t_SL U37524 ( .A1(n29983), .A2(n29982), .A3(n29981), .B(
        n29980), .Y(n29984) );
  NOR2xp33_ASAP7_75t_SL U37525 ( .A(uart1_r_TWADDR__0_), .B(uart1_r_TWADDR__1_), .Y(n27320) );
  NOR2xp33_ASAP7_75t_SL U37526 ( .A(uart1_r_TWADDR__4_), .B(n2267), .Y(n27310)
         );
  NOR2xp33_ASAP7_75t_SL U37527 ( .A(n27355), .B(n27373), .Y(n27380) );
  NOR2xp33_ASAP7_75t_SL U37528 ( .A(n30941), .B(n22379), .Y(n30942) );
  AOI31xp33_ASAP7_75t_SL U37529 ( .A1(n32192), .A2(n32191), .A3(n32190), .B(
        n24516), .Y(n2706) );
  NOR2xp33_ASAP7_75t_SL U37530 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__0_), .B(
        n22421), .Y(n32107) );
  NOR2xp33_ASAP7_75t_SL U37531 ( .A(n31333), .B(n30940), .Y(n32192) );
  AOI31xp33_ASAP7_75t_SL U37532 ( .A1(n32139), .A2(n31964), .A3(n32137), .B(
        n31963), .Y(n31965) );
  NOR2xp33_ASAP7_75t_SL U37533 ( .A(uart1_r_RCNT__2_), .B(n30898), .Y(n27504)
         );
  NOR2xp33_ASAP7_75t_SL U37534 ( .A(n27510), .B(n31238), .Y(n27521) );
  NOR2xp33_ASAP7_75t_SL U37535 ( .A(n26071), .B(n27328), .Y(n27309) );
  NOR2xp33_ASAP7_75t_SL U37536 ( .A(n28047), .B(n28046), .Y(n28051) );
  NOR2xp33_ASAP7_75t_SL U37537 ( .A(n28799), .B(n28803), .Y(n28801) );
  NOR2xp33_ASAP7_75t_SL U37538 ( .A(n28815), .B(n22379), .Y(n28816) );
  AOI31xp33_ASAP7_75t_SL U37539 ( .A1(n29686), .A2(n31542), .A3(n29685), .B(
        n26325), .Y(n26326) );
  NOR2xp33_ASAP7_75t_SL U37540 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__5_), .B(
        n23229), .Y(n26325) );
  NOR2xp33_ASAP7_75t_SL U37541 ( .A(n28799), .B(n27135), .Y(n27134) );
  AOI211xp5_ASAP7_75t_SL U37542 ( .A1(n28894), .A2(n30406), .B(n28787), .C(
        n28786), .Y(n28788) );
  NOR2xp33_ASAP7_75t_SL U37543 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__6_), .B(
        n30007), .Y(n26282) );
  AOI211xp5_ASAP7_75t_SL U37544 ( .A1(n28894), .A2(n30416), .B(n26274), .C(
        n26273), .Y(n26275) );
  NAND2xp33_ASAP7_75t_SRAM U37545 ( .A(n26268), .B(n29584), .Y(n26272) );
  NAND2xp33_ASAP7_75t_SRAM U37546 ( .A(n24634), .B(n28879), .Y(n28785) );
  NOR2xp33_ASAP7_75t_SL U37547 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__3_), .B(
        n22379), .Y(n29501) );
  NOR4xp25_ASAP7_75t_SL U37548 ( .A(n33033), .B(n31798), .C(n33040), .D(n32751), .Y(n31800) );
  AOI211xp5_ASAP7_75t_SL U37549 ( .A1(u0_0_leon3x0_p0_iu_r_E__CWP__2_), .A2(
        n30621), .B(n28943), .C(n28942), .Y(n28944) );
  NOR2xp33_ASAP7_75t_SL U37550 ( .A(n28941), .B(n28940), .Y(n28943) );
  AOI211xp5_ASAP7_75t_SL U37551 ( .A1(n28924), .A2(n30631), .B(n28923), .C(
        n28922), .Y(n28950) );
  NOR2xp33_ASAP7_75t_SL U37552 ( .A(n28914), .B(n28913), .Y(n28923) );
  NOR2xp33_ASAP7_75t_SL U37553 ( .A(n31334), .B(n31343), .Y(n30471) );
  AOI211xp5_ASAP7_75t_SL U37554 ( .A1(n28894), .A2(n30449), .B(n28893), .C(
        n28892), .Y(n28895) );
  NOR2xp33_ASAP7_75t_SL U37555 ( .A(n24427), .B(n26308), .Y(n28890) );
  NOR2xp33_ASAP7_75t_SL U37556 ( .A(n28992), .B(n28913), .Y(n28875) );
  NOR2xp33_ASAP7_75t_SL U37557 ( .A(n28992), .B(n28971), .Y(n28874) );
  NOR2xp33_ASAP7_75t_SL U37558 ( .A(n28799), .B(n28757), .Y(n28756) );
  NOR2xp33_ASAP7_75t_SL U37559 ( .A(n22378), .B(n31967), .Y(n29881) );
  NOR2xp33_ASAP7_75t_SL U37560 ( .A(n28799), .B(n28611), .Y(n28610) );
  NOR2xp33_ASAP7_75t_SL U37561 ( .A(n28799), .B(n28581), .Y(n28580) );
  AOI211xp5_ASAP7_75t_SL U37562 ( .A1(u0_0_leon3x0_p0_divi[40]), .A2(n28782), 
        .B(n27117), .C(n27116), .Y(n27118) );
  NAND2xp33_ASAP7_75t_SRAM U37563 ( .A(n30614), .B(n30395), .Y(n28732) );
  NOR2xp33_ASAP7_75t_SL U37564 ( .A(n25284), .B(n22373), .Y(n30395) );
  NOR2xp33_ASAP7_75t_SL U37565 ( .A(n28729), .B(n28728), .Y(n28739) );
  NOR2xp33_ASAP7_75t_SL U37566 ( .A(n28808), .B(n28656), .Y(n28655) );
  AOI211xp5_ASAP7_75t_SL U37567 ( .A1(n28894), .A2(n30380), .B(n28639), .C(
        n28638), .Y(n28640) );
  NOR2xp33_ASAP7_75t_SL U37568 ( .A(n28975), .B(n28917), .Y(n26251) );
  NOR2xp33_ASAP7_75t_SL U37569 ( .A(n28921), .B(n28913), .Y(n28841) );
  NOR2xp33_ASAP7_75t_SL U37570 ( .A(n24526), .B(n24984), .Y(n31872) );
  AOI211xp5_ASAP7_75t_SL U37571 ( .A1(n30632), .A2(n30631), .B(n30630), .C(
        n30629), .Y(n30633) );
  NOR2xp33_ASAP7_75t_SL U37572 ( .A(n30628), .B(n30627), .Y(n30629) );
  AOI211xp5_ASAP7_75t_SL U37573 ( .A1(n28981), .A2(n28978), .B(n28852), .C(
        n28851), .Y(n28853) );
  NOR2xp33_ASAP7_75t_SL U37574 ( .A(n28850), .B(n28849), .Y(n28851) );
  NOR2xp33_ASAP7_75t_SL U37575 ( .A(n28799), .B(n28560), .Y(n28559) );
  NOR2xp33_ASAP7_75t_SL U37576 ( .A(n27153), .B(n27152), .Y(n27157) );
  AOI211xp5_ASAP7_75t_SL U37577 ( .A1(n28924), .A2(n28675), .B(n28674), .C(
        n28673), .Y(n28696) );
  NOR2xp33_ASAP7_75t_SL U37578 ( .A(n29764), .B(n31047), .Y(n3030) );
  NOR2xp33_ASAP7_75t_SL U37579 ( .A(n30971), .B(n31047), .Y(n3027) );
  NOR2xp33_ASAP7_75t_SL U37580 ( .A(n25448), .B(n31047), .Y(n3023) );
  AOI211xp5_ASAP7_75t_SL U37581 ( .A1(n28424), .A2(n26680), .B(n26679), .C(
        n26678), .Y(n26691) );
  AOI211xp5_ASAP7_75t_SL U37582 ( .A1(n28762), .A2(n26709), .B(n26672), .C(
        n26671), .Y(n26696) );
  NOR2xp33_ASAP7_75t_SL U37583 ( .A(n28921), .B(n27209), .Y(n26672) );
  NOR2xp33_ASAP7_75t_SL U37584 ( .A(n22427), .B(n30159), .Y(n29726) );
  NOR2xp33_ASAP7_75t_SL U37585 ( .A(n29470), .B(n30686), .Y(n29719) );
  NOR2xp33_ASAP7_75t_SL U37586 ( .A(n29473), .B(n29472), .Y(n29723) );
  NAND2xp33_ASAP7_75t_SRAM U37587 ( .A(n29705), .B(n29702), .Y(n29471) );
  NAND2xp33_ASAP7_75t_SRAM U37588 ( .A(n29718), .B(n29717), .Y(n29724) );
  NOR2xp33_ASAP7_75t_SL U37589 ( .A(n29638), .B(n30706), .Y(n30708) );
  NOR2xp33_ASAP7_75t_SL U37590 ( .A(n28799), .B(n28534), .Y(n28533) );
  NOR2xp33_ASAP7_75t_SL U37591 ( .A(n27281), .B(n31343), .Y(n25840) );
  NOR2xp33_ASAP7_75t_SL U37592 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__19_), .B(
        n30007), .Y(n25803) );
  AOI211xp5_ASAP7_75t_SL U37593 ( .A1(n29605), .A2(n26709), .B(n25781), .C(
        n25780), .Y(n25804) );
  AOI211xp5_ASAP7_75t_SL U37594 ( .A1(u0_0_leon3x0_p0_divi[50]), .A2(n28782), 
        .B(n25767), .C(n25766), .Y(n25770) );
  NOR2xp33_ASAP7_75t_SL U37595 ( .A(n32173), .B(n32172), .Y(n32175) );
  NOR2xp33_ASAP7_75t_SL U37596 ( .A(n27013), .B(n22379), .Y(n27014) );
  NOR2xp33_ASAP7_75t_SL U37597 ( .A(n30579), .B(n30578), .Y(n3000) );
  AOI211xp5_ASAP7_75t_SL U37598 ( .A1(u0_0_leon3x0_p0_divi[49]), .A2(n26174), 
        .B(n25818), .C(n25817), .Y(n25819) );
  NOR2xp33_ASAP7_75t_SL U37599 ( .A(n31396), .B(n25809), .Y(n27281) );
  AOI211xp5_ASAP7_75t_SL U37600 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__17_), 
        .A2(n24581), .B(n28887), .C(n26699), .Y(n26700) );
  NOR2xp33_ASAP7_75t_SL U37601 ( .A(n26698), .B(n29592), .Y(n26699) );
  AOI211xp5_ASAP7_75t_SL U37602 ( .A1(u0_0_leon3x0_p0_divi[44]), .A2(n26174), 
        .B(n26173), .C(n26172), .Y(n26175) );
  AOI211xp5_ASAP7_75t_SL U37603 ( .A1(n28855), .A2(n28675), .B(n26159), .C(
        n26158), .Y(n26185) );
  AOI31xp33_ASAP7_75t_SL U37604 ( .A1(n24634), .A2(n28737), .A3(n26585), .B(
        n26575), .Y(n26576) );
  AOI211xp5_ASAP7_75t_SL U37605 ( .A1(n28855), .A2(n28615), .B(n26561), .C(
        n26560), .Y(n26583) );
  NOR2xp33_ASAP7_75t_SL U37606 ( .A(n28618), .B(n27209), .Y(n26561) );
  NOR2xp33_ASAP7_75t_SL U37607 ( .A(n32710), .B(n31750), .Y(n31757) );
  NOR2xp33_ASAP7_75t_SL U37608 ( .A(n32040), .B(n31734), .Y(n31803) );
  NOR2xp33_ASAP7_75t_SL U37609 ( .A(n25613), .B(n31001), .Y(n25614) );
  AOI211xp5_ASAP7_75t_SL U37610 ( .A1(it_q[6]), .A2(n24636), .B(n30562), .C(
        n30561), .Y(n30569) );
  NOR2xp33_ASAP7_75t_SL U37611 ( .A(n32315), .B(n31470), .Y(n30561) );
  NAND2xp33_ASAP7_75t_SRAM U37612 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_), .B(n32012), .Y(n26270) );
  NOR2xp33_ASAP7_75t_SL U37613 ( .A(n28977), .B(n28917), .Y(n28918) );
  NOR2xp33_ASAP7_75t_SL U37614 ( .A(n26250), .B(n26249), .Y(n28917) );
  NOR2xp33_ASAP7_75t_SL U37615 ( .A(n26298), .B(n27109), .Y(n26249) );
  NOR2xp33_ASAP7_75t_SL U37616 ( .A(n28977), .B(n28976), .Y(n28990) );
  NAND2xp33_ASAP7_75t_SRAM U37617 ( .A(n18606), .B(n28982), .Y(n26259) );
  AOI211xp5_ASAP7_75t_SL U37618 ( .A1(ic_q[16]), .A2(n22387), .B(n26665), .C(
        n27249), .Y(n26667) );
  NOR2xp33_ASAP7_75t_SL U37619 ( .A(n26664), .B(n31466), .Y(n26665) );
  AOI211xp5_ASAP7_75t_SL U37620 ( .A1(n31004), .A2(dc_q[8]), .B(n29762), .C(
        n29761), .Y(n30482) );
  NOR2xp33_ASAP7_75t_SL U37621 ( .A(n32322), .B(n31470), .Y(n29761) );
  AOI211xp5_ASAP7_75t_SL U37622 ( .A1(dc_q[0]), .A2(n31473), .B(n30476), .C(
        n30475), .Y(n30485) );
  NOR2xp33_ASAP7_75t_SL U37623 ( .A(n32463), .B(n24426), .Y(n30476) );
  AOI211xp5_ASAP7_75t_SL U37624 ( .A1(n31004), .A2(dc_q[11]), .B(n30884), .C(
        n30883), .Y(n30970) );
  NOR2xp33_ASAP7_75t_SL U37625 ( .A(n32333), .B(n31470), .Y(n30883) );
  AOI211xp5_ASAP7_75t_SL U37626 ( .A1(n31473), .A2(dc_q[4]), .B(n31472), .C(
        n31471), .Y(n31489) );
  AOI211xp5_ASAP7_75t_SL U37627 ( .A1(n31004), .A2(dc_q[10]), .B(n31003), .C(
        n31002), .Y(n31046) );
  NOR2xp33_ASAP7_75t_SL U37628 ( .A(n32328), .B(n31470), .Y(n31002) );
  AOI211xp5_ASAP7_75t_SL U37629 ( .A1(dc_q[2]), .A2(n31473), .B(n30998), .C(
        n30997), .Y(n31010) );
  NOR2xp33_ASAP7_75t_SL U37630 ( .A(n32475), .B(n24426), .Y(n30998) );
  AOI211xp5_ASAP7_75t_SL U37631 ( .A1(n28742), .A2(n28615), .B(n27212), .C(
        n27211), .Y(n27213) );
  AOI211xp5_ASAP7_75t_SL U37632 ( .A1(n26278), .A2(n24571), .B(n26155), .C(
        n24475), .Y(n27106) );
  AND2x2_ASAP7_75t_SL U37633 ( .A(n26140), .B(n26139), .Y(n28982) );
  AOI211xp5_ASAP7_75t_SL U37634 ( .A1(n31356), .A2(n28411), .B(n27254), .C(
        n30578), .Y(n3018) );
  AOI211xp5_ASAP7_75t_SL U37635 ( .A1(n30025), .A2(n28411), .B(n26336), .C(
        n30578), .Y(n3015) );
  NOR2xp33_ASAP7_75t_SL U37636 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__21_), .B(n31001), .Y(n26331) );
  NOR2xp33_ASAP7_75t_SL U37637 ( .A(n25417), .B(n30575), .Y(n25418) );
  NOR2xp33_ASAP7_75t_SL U37638 ( .A(n26889), .B(n30575), .Y(n26347) );
  NOR2xp33_ASAP7_75t_SL U37639 ( .A(n23550), .B(n30575), .Y(n26375) );
  NOR2xp33_ASAP7_75t_SL U37640 ( .A(n26224), .B(n30575), .Y(n26225) );
  NOR2xp33_ASAP7_75t_SL U37641 ( .A(n25815), .B(n30575), .Y(n25718) );
  NOR2xp33_ASAP7_75t_SL U37642 ( .A(n26967), .B(n30575), .Y(n26968) );
  NOR2xp33_ASAP7_75t_SL U37643 ( .A(n25050), .B(n30017), .Y(n25051) );
  AOI211xp5_ASAP7_75t_SL U37644 ( .A1(u0_0_leon3x0_p0_divi[52]), .A2(n28782), 
        .B(n27072), .C(n27071), .Y(n27073) );
  NOR2xp33_ASAP7_75t_SL U37645 ( .A(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__17_), .B(n31001), .Y(n27250) );
  NOR2xp33_ASAP7_75t_SL U37646 ( .A(n25067), .B(n25440), .Y(n30015) );
  AOI211xp5_ASAP7_75t_SL U37647 ( .A1(n30130), .A2(n32615), .B(n30129), .C(
        n30128), .Y(n31359) );
  NOR2xp33_ASAP7_75t_SL U37648 ( .A(n31694), .B(n30017), .Y(n25017) );
  NOR2xp33_ASAP7_75t_SL U37649 ( .A(n32730), .B(n30017), .Y(n25049) );
  NOR2xp33_ASAP7_75t_SL U37650 ( .A(n32713), .B(n30017), .Y(n25054) );
  NOR2xp33_ASAP7_75t_SL U37651 ( .A(n32734), .B(n30017), .Y(n25039) );
  AOI211xp5_ASAP7_75t_SL U37652 ( .A1(dc_q[1]), .A2(n31473), .B(n31355), .C(
        n31354), .Y(n31362) );
  OR2x2_ASAP7_75t_SL U37653 ( .A(n25030), .B(n25029), .Y(n24426) );
  NOR2xp33_ASAP7_75t_SL U37654 ( .A(n25584), .B(n32198), .Y(n25027) );
  AOI211xp5_ASAP7_75t_SL U37655 ( .A1(n32883), .A2(sr1_r_MCFG1__IOWIDTH__1_), 
        .B(n32727), .C(n32726), .Y(n1779) );
  NOR2xp33_ASAP7_75t_SL U37656 ( .A(n32721), .B(n32801), .Y(n32724) );
  NOR2xp33_ASAP7_75t_SL U37657 ( .A(n32833), .B(n32875), .Y(n32727) );
  NOR2xp33_ASAP7_75t_SL U37658 ( .A(n28482), .B(n27195), .Y(n30616) );
  NOR2xp33_ASAP7_75t_SL U37659 ( .A(n28734), .B(n25497), .Y(n27195) );
  NOR2xp33_ASAP7_75t_SL U37660 ( .A(n26394), .B(n25820), .Y(n27153) );
  NOR2xp33_ASAP7_75t_SL U37661 ( .A(n28513), .B(n22379), .Y(n28514) );
  AOI211xp5_ASAP7_75t_SL U37662 ( .A1(n32883), .A2(sr1_r_MCFG1__IOWIDTH__0_), 
        .B(n32882), .C(n32881), .Y(n2291) );
  NOR2xp33_ASAP7_75t_SL U37663 ( .A(n32723), .B(n32722), .Y(n32877) );
  NOR2xp33_ASAP7_75t_SL U37664 ( .A(n32876), .B(n32879), .Y(n32878) );
  NOR2xp33_ASAP7_75t_SL U37665 ( .A(n32884), .B(n32875), .Y(n32882) );
  OR2x2_ASAP7_75t_SL U37666 ( .A(n32036), .B(n32002), .Y(n24424) );
  NOR4xp25_ASAP7_75t_SL U37667 ( .A(n31734), .B(n32879), .C(n33029), .D(n33049), .Y(n25259) );
  NOR4xp25_ASAP7_75t_SL U37668 ( .A(n33032), .B(n33039), .C(n33046), .D(n32776), .Y(n25260) );
  AOI211xp5_ASAP7_75t_SL U37669 ( .A1(n30632), .A2(n28497), .B(n28496), .C(
        n28495), .Y(n28501) );
  AOI31xp33_ASAP7_75t_SL U37670 ( .A1(n28489), .A2(n28488), .A3(n28487), .B(
        n24427), .Y(n28496) );
  NAND2xp33_ASAP7_75t_SRAM U37671 ( .A(u0_0_leon3x0_p0_iu_r_W__S__TBA__10_), 
        .B(n28480), .Y(n28484) );
  AOI211xp5_ASAP7_75t_SL U37672 ( .A1(n24578), .A2(n22436), .B(n26155), .C(
        n25791), .Y(n27107) );
  NOR2xp33_ASAP7_75t_SL U37673 ( .A(n27108), .B(n26152), .Y(n25793) );
  AOI211xp5_ASAP7_75t_SL U37674 ( .A1(n28835), .A2(n30240), .B(n26898), .C(
        n26897), .Y(n26899) );
  NOR2xp33_ASAP7_75t_SL U37675 ( .A(n26894), .B(n29594), .Y(n26898) );
  AOI211xp5_ASAP7_75t_SL U37676 ( .A1(n30679), .A2(n29171), .B(n29170), .C(
        n29169), .Y(n29172) );
  NOR2xp33_ASAP7_75t_SL U37677 ( .A(n29168), .B(n29167), .Y(n29169) );
  NOR4xp25_ASAP7_75t_SL U37678 ( .A(u0_0_leon3x0_p0_mulo[10]), .B(
        u0_0_leon3x0_p0_mulo[8]), .C(u0_0_leon3x0_p0_mulo[9]), .D(
        u0_0_leon3x0_p0_mulo[5]), .Y(n29122) );
  NOR4xp25_ASAP7_75t_SL U37679 ( .A(u0_0_leon3x0_p0_mulo[7]), .B(
        u0_0_leon3x0_p0_mulo[6]), .C(u0_0_leon3x0_p0_mulo[3]), .D(
        u0_0_leon3x0_p0_mulo[4]), .Y(n29123) );
  NOR4xp25_ASAP7_75t_SL U37680 ( .A(u0_0_leon3x0_p0_mulo[18]), .B(
        u0_0_leon3x0_p0_mulo[17]), .C(u0_0_leon3x0_p0_mulo[16]), .D(
        u0_0_leon3x0_p0_mulo[2]), .Y(n29124) );
  NOR4xp25_ASAP7_75t_SL U37681 ( .A(u0_0_leon3x0_p0_mulo[12]), .B(
        u0_0_leon3x0_p0_mulo[11]), .C(u0_0_leon3x0_p0_mulo[0]), .D(
        u0_0_leon3x0_p0_mulo[1]), .Y(n29125) );
  NOR4xp25_ASAP7_75t_SL U37682 ( .A(u0_0_leon3x0_p0_mulo[21]), .B(
        u0_0_leon3x0_p0_mulo[20]), .C(u0_0_leon3x0_p0_mulo[19]), .D(
        u0_0_leon3x0_p0_mulo[13]), .Y(n29118) );
  NOR4xp25_ASAP7_75t_SL U37683 ( .A(u0_0_leon3x0_p0_mulo[24]), .B(
        u0_0_leon3x0_p0_mulo[22]), .C(u0_0_leon3x0_p0_mulo[15]), .D(
        u0_0_leon3x0_p0_mulo[14]), .Y(n29119) );
  NOR4xp25_ASAP7_75t_SL U37684 ( .A(u0_0_leon3x0_p0_mulo[27]), .B(
        u0_0_leon3x0_p0_mulo[25]), .C(u0_0_leon3x0_p0_mulo[26]), .D(
        u0_0_leon3x0_p0_mulo[23]), .Y(n29120) );
  NOR4xp25_ASAP7_75t_SL U37685 ( .A(u0_0_leon3x0_p0_mulo[63]), .B(
        u0_0_leon3x0_p0_mulo[30]), .C(u0_0_leon3x0_p0_mulo[28]), .D(
        u0_0_leon3x0_p0_mulo[29]), .Y(n29121) );
  NOR2xp33_ASAP7_75t_SL U37686 ( .A(n28799), .B(n28469), .Y(n28468) );
  OR2x2_ASAP7_75t_SL U37687 ( .A(n24658), .B(n28536), .Y(n28802) );
  AND2x2_ASAP7_75t_SL U37688 ( .A(n22379), .B(n30648), .Y(n28799) );
  NAND2xp33_ASAP7_75t_SRAM U37689 ( .A(n18296), .B(n26278), .Y(n25758) );
  AOI211xp5_ASAP7_75t_SL U37690 ( .A1(n29598), .A2(n29067), .B(n26422), .C(
        n26421), .Y(n26436) );
  AOI211xp5_ASAP7_75t_SL U37691 ( .A1(n29605), .A2(n28497), .B(n28439), .C(
        n28438), .Y(n28442) );
  NOR2xp33_ASAP7_75t_SL U37692 ( .A(n18891), .B(n28941), .Y(n28424) );
  NOR2xp33_ASAP7_75t_SL U37693 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__24_), .B(
        n30007), .Y(n26409) );
  AOI211xp5_ASAP7_75t_SL U37694 ( .A1(n29605), .A2(n28498), .B(n26407), .C(
        n26406), .Y(n26410) );
  AOI211xp5_ASAP7_75t_SL U37695 ( .A1(n29583), .A2(n23002), .B(n26400), .C(
        n26399), .Y(n26401) );
  NAND2xp33_ASAP7_75t_SRAM U37696 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__PC__24_), 
        .B(n28888), .Y(n26398) );
  NOR2xp33_ASAP7_75t_SL U37697 ( .A(n26394), .B(n26674), .Y(n28729) );
  NAND2xp33_ASAP7_75t_SRAM U37698 ( .A(n28742), .B(n28497), .Y(n26403) );
  NOR2xp33_ASAP7_75t_SL U37699 ( .A(n18813), .B(n25782), .Y(n26380) );
  AOI211xp5_ASAP7_75t_SL U37700 ( .A1(n29603), .A2(n18794), .B(n25906), .C(
        n25905), .Y(n25914) );
  AOI211xp5_ASAP7_75t_SL U37701 ( .A1(n29583), .A2(n22968), .B(n25899), .C(
        n25898), .Y(n25903) );
  NOR2xp33_ASAP7_75t_SL U37702 ( .A(n30625), .B(n30225), .Y(n25906) );
  AOI211xp5_ASAP7_75t_SL U37703 ( .A1(n28835), .A2(n30236), .B(n26931), .C(
        n26930), .Y(n26932) );
  NOR2xp33_ASAP7_75t_SL U37704 ( .A(n26927), .B(n29594), .Y(n26931) );
  NAND2xp33_ASAP7_75t_SRAM U37705 ( .A(add_x_735_A_29_), .B(n24578), .Y(n25462) );
  NOR2xp33_ASAP7_75t_SL U37706 ( .A(u0_0_leon3x0_p0_iu_r_E__SHLEFT_), .B(
        n26139), .Y(n24578) );
  NOR2xp33_ASAP7_75t_SL U37707 ( .A(n29160), .B(n29159), .Y(n29161) );
  NOR2xp33_ASAP7_75t_SL U37708 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[27]), .Y(
        n26921) );
  NOR2xp33_ASAP7_75t_SL U37709 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[1]), .Y(
        n28929) );
  NOR2xp33_ASAP7_75t_SL U37710 ( .A(n29561), .B(n28928), .Y(n28930) );
  NOR2xp33_ASAP7_75t_SL U37711 ( .A(n24631), .B(n18909), .Y(n26359) );
  NOR2xp33_ASAP7_75t_SL U37712 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[10]), .Y(
        n28679) );
  NOR2xp33_ASAP7_75t_SL U37713 ( .A(n29148), .B(u0_0_leon3x0_p0_divi[10]), .Y(
        n28678) );
  NOR2xp33_ASAP7_75t_SL U37714 ( .A(u0_0_leon3x0_p0_divi[10]), .B(n29150), .Y(
        n28684) );
  NOR2xp33_ASAP7_75t_SL U37715 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[11]), .Y(
        n28628) );
  NOR2xp33_ASAP7_75t_SL U37716 ( .A(n28621), .B(n28928), .Y(n28629) );
  NOR2xp33_ASAP7_75t_SL U37717 ( .A(n29148), .B(n22721), .Y(n28630) );
  NOR4xp25_ASAP7_75t_SL U37718 ( .A(n30416), .B(n30406), .C(n31416), .D(n30337), .Y(n29162) );
  AOI211xp5_ASAP7_75t_SL U37719 ( .A1(n18406), .A2(n28821), .B(n27200), .C(
        n26682), .Y(n26686) );
  AOI211xp5_ASAP7_75t_SL U37720 ( .A1(n18406), .A2(n29148), .B(n24631), .C(
        u0_0_leon3x0_p0_divi[15]), .Y(n26687) );
  NOR2xp33_ASAP7_75t_SL U37721 ( .A(n28771), .B(n28770), .Y(n28776) );
  NOR2xp33_ASAP7_75t_SL U37722 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[6]), .Y(
        n28778) );
  NOR4xp25_ASAP7_75t_SL U37723 ( .A(n30261), .B(n30349), .C(n30266), .D(n30360), .Y(n29163) );
  AOI211xp5_ASAP7_75t_SL U37724 ( .A1(n29148), .A2(n27196), .B(n24631), .C(
        u0_0_leon3x0_p0_divi[13]), .Y(n27203) );
  AOI211xp5_ASAP7_75t_SL U37725 ( .A1(n29148), .A2(n22418), .B(n24631), .C(
        u0_0_leon3x0_p0_divi[23]), .Y(n26388) );
  AOI211xp5_ASAP7_75t_SL U37726 ( .A1(n28928), .A2(add_x_735_A_9_), .B(n24631), 
        .C(n18904), .Y(n28722) );
  NOR2xp33_ASAP7_75t_SL U37727 ( .A(n29148), .B(n18904), .Y(n28721) );
  AOI211xp5_ASAP7_75t_SL U37728 ( .A1(n28928), .A2(n24571), .B(n24631), .C(
        u0_0_leon3x0_p0_divi[17]), .Y(n25824) );
  NOR2xp33_ASAP7_75t_SL U37729 ( .A(n29148), .B(u0_0_leon3x0_p0_divi[17]), .Y(
        n25823) );
  NOR2xp33_ASAP7_75t_SL U37730 ( .A(n29146), .B(n25822), .Y(n25827) );
  NOR2xp33_ASAP7_75t_SL U37731 ( .A(n29148), .B(u0_0_leon3x0_p0_divi[18]), .Y(
        n25774) );
  NOR2xp33_ASAP7_75t_SL U37732 ( .A(n29146), .B(n25773), .Y(n25778) );
  NOR2xp33_ASAP7_75t_SL U37733 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[2]), .Y(
        n28884) );
  NOR2xp33_ASAP7_75t_SL U37734 ( .A(n23954), .B(n28928), .Y(n28885) );
  NOR2xp33_ASAP7_75t_SL U37735 ( .A(n29148), .B(n22449), .Y(n28886) );
  NOR2xp33_ASAP7_75t_SL U37736 ( .A(n29148), .B(u0_0_leon3x0_p0_divi[3]), .Y(
        n28826) );
  AOI211xp5_ASAP7_75t_SL U37737 ( .A1(n28928), .A2(u0_0_leon3x0_p0_muli[41]), 
        .B(n24631), .C(u0_0_leon3x0_p0_divi[3]), .Y(n28832) );
  NOR2xp33_ASAP7_75t_SL U37738 ( .A(n29148), .B(n22837), .Y(n27140) );
  NOR2xp33_ASAP7_75t_SL U37739 ( .A(n29134), .B(n30246), .Y(n29140) );
  NOR2xp33_ASAP7_75t_SL U37740 ( .A(n29148), .B(u0_0_leon3x0_p0_divi[25]), .Y(
        n25489) );
  AOI211xp5_ASAP7_75t_SL U37741 ( .A1(n28928), .A2(n18606), .B(n24631), .C(
        u0_0_leon3x0_p0_divi[24]), .Y(n28433) );
  NOR2xp33_ASAP7_75t_SL U37742 ( .A(n25488), .B(n24488), .Y(n28928) );
  NOR2xp33_ASAP7_75t_SL U37743 ( .A(n29148), .B(u0_0_leon3x0_p0_divi[24]), .Y(
        n28432) );
  NOR2xp33_ASAP7_75t_SL U37744 ( .A(n29146), .B(n28431), .Y(n28436) );
  AOI31xp33_ASAP7_75t_SL U37745 ( .A1(n24579), .A2(u0_0_leon3x0_p0_divi[0]), 
        .A3(n26742), .B(n26741), .Y(n26745) );
  NOR2xp33_ASAP7_75t_SL U37746 ( .A(n26740), .B(u0_0_leon3x0_p0_divi[0]), .Y(
        n26741) );
  NOR2xp33_ASAP7_75t_SL U37747 ( .A(n32828), .B(n32831), .Y(n32829) );
  NOR2xp33_ASAP7_75t_SL U37748 ( .A(n32823), .B(n32822), .Y(n32825) );
  NAND2xp33_ASAP7_75t_SRAM U37749 ( .A(n24943), .B(n24929), .Y(n24919) );
  NOR2xp33_ASAP7_75t_SL U37750 ( .A(n32489), .B(n25333), .Y(n25332) );
  NOR2xp33_ASAP7_75t_SL U37751 ( .A(n2963), .B(n31697), .Y(n25331) );
  AOI211xp5_ASAP7_75t_SL U37752 ( .A1(rwen[3]), .A2(n32749), .B(n32748), .C(
        n32747), .Y(n1719) );
  AOI211xp5_ASAP7_75t_SL U37753 ( .A1(rwen[0]), .A2(n32749), .B(n32744), .C(
        n32746), .Y(n1722) );
  AOI211xp5_ASAP7_75t_SL U37754 ( .A1(rwen[1]), .A2(n32749), .B(n32744), .C(
        n32747), .Y(n1721) );
  NOR2xp33_ASAP7_75t_SL U37755 ( .A(n1723), .B(n32745), .Y(n32744) );
  AOI211xp5_ASAP7_75t_SL U37756 ( .A1(rwen[2]), .A2(n32749), .B(n32748), .C(
        n32746), .Y(n1720) );
  NOR2xp33_ASAP7_75t_SL U37757 ( .A(address[1]), .B(n32745), .Y(n32748) );
  NOR2xp33_ASAP7_75t_SL U37758 ( .A(u0_0_leon3x0_p0_iu_r_E__SHLEFT_), .B(
        n26139), .Y(n24577) );
  AOI211xp5_ASAP7_75t_SL U37759 ( .A1(n29603), .A2(n29602), .B(n29601), .C(
        n29600), .Y(n29607) );
  AOI211xp5_ASAP7_75t_SL U37760 ( .A1(n30591), .A2(n29598), .B(n29597), .C(
        n29596), .Y(n29599) );
  NAND2xp33_ASAP7_75t_SRAM U37761 ( .A(n30598), .B(n24662), .Y(n30602) );
  NOR2xp33_ASAP7_75t_SL U37762 ( .A(n32719), .B(n22386), .Y(n32991) );
  NOR2xp33_ASAP7_75t_SL U37763 ( .A(n25080), .B(n24989), .Y(n25075) );
  NOR2xp33_ASAP7_75t_SL U37764 ( .A(n26993), .B(n26992), .Y(n29155) );
  NOR2xp33_ASAP7_75t_SL U37765 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[19]), .Y(
        n26990) );
  NOR2xp33_ASAP7_75t_SL U37766 ( .A(n28931), .B(u0_0_leon3x0_p0_divi[19]), .Y(
        n26989) );
  NOR2xp33_ASAP7_75t_SL U37767 ( .A(n29148), .B(u0_0_leon3x0_p0_divi[20]), .Y(
        n27060) );
  NAND2xp33_ASAP7_75t_SRAM U37768 ( .A(n29146), .B(u0_0_leon3x0_p0_divi[20]), 
        .Y(n27062) );
  NOR2xp33_ASAP7_75t_SL U37769 ( .A(u0_0_leon3x0_p0_divi[0]), .B(n18909), .Y(
        n30662) );
  NOR2xp33_ASAP7_75t_SL U37770 ( .A(n18530), .B(u0_0_leon3x0_p0_divi[30]), .Y(
        n30659) );
  AOI211xp5_ASAP7_75t_SL U37771 ( .A1(n29148), .A2(n22493), .B(n24631), .C(
        u0_0_leon3x0_p0_divi[22]), .Y(n26433) );
  AOI211xp5_ASAP7_75t_SL U37772 ( .A1(n24576), .A2(n26377), .B(n25202), .C(
        n25201), .Y(n25203) );
  NOR2xp33_ASAP7_75t_SL U37773 ( .A(n28986), .B(n25463), .Y(n25201) );
  NAND2xp33_ASAP7_75t_SRAM U37774 ( .A(add_x_735_A_10_), .B(n25200), .Y(n25463) );
  NOR2xp33_ASAP7_75t_SL U37775 ( .A(n28977), .B(n28845), .Y(n24576) );
  AOI211xp5_ASAP7_75t_SL U37776 ( .A1(n28894), .A2(n31416), .B(n25186), .C(
        n25185), .Y(n25205) );
  AOI211xp5_ASAP7_75t_SL U37777 ( .A1(n28835), .A2(n31401), .B(n25181), .C(
        n25180), .Y(n25182) );
  NOR2xp33_ASAP7_75t_SL U37778 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .B(
        n25894), .Y(n25173) );
  AOI31xp33_ASAP7_75t_SL U37779 ( .A1(n25901), .A2(n24634), .A3(n26585), .B(
        n26575), .Y(n25183) );
  NOR2xp33_ASAP7_75t_SL U37780 ( .A(n26394), .B(n29910), .Y(n26575) );
  NOR2xp33_ASAP7_75t_SL U37781 ( .A(n26169), .B(n24427), .Y(n27065) );
  AND2x2_ASAP7_75t_SL U37782 ( .A(n24634), .B(n28403), .Y(n29598) );
  AND2x2_ASAP7_75t_SL U37783 ( .A(n24634), .B(n28486), .Y(n29583) );
  AOI211xp5_ASAP7_75t_SL U37784 ( .A1(n24575), .A2(n25910), .B(n25149), .C(
        n25148), .Y(n25150) );
  NOR2xp33_ASAP7_75t_SL U37785 ( .A(n28869), .B(n25907), .Y(n25148) );
  AOI211xp5_ASAP7_75t_SL U37786 ( .A1(n25142), .A2(n23091), .B(n18813), .C(
        n25141), .Y(n25912) );
  NOR2xp33_ASAP7_75t_SL U37787 ( .A(n24572), .B(n25190), .Y(n25141) );
  NOR2xp33_ASAP7_75t_SL U37788 ( .A(n24631), .B(u0_0_leon3x0_p0_divi[30]), .Y(
        n25136) );
  AOI211xp5_ASAP7_75t_SL U37789 ( .A1(n28981), .A2(n26389), .B(n28968), .C(
        n25117), .Y(n25118) );
  NOR2xp33_ASAP7_75t_SL U37790 ( .A(n26298), .B(n25198), .Y(n25142) );
  NOR2xp33_ASAP7_75t_SL U37791 ( .A(u0_0_leon3x0_p0_iu_r_E__SHLEFT_), .B(
        n26139), .Y(n26278) );
  NOR2xp33_ASAP7_75t_SL U37792 ( .A(n22418), .B(n25190), .Y(n25469) );
  NOR2xp33_ASAP7_75t_SL U37793 ( .A(n26140), .B(n26139), .Y(n25200) );
  NOR2xp33_ASAP7_75t_SL U37794 ( .A(n28977), .B(n28845), .Y(n24575) );
  NOR2xp33_ASAP7_75t_SL U37795 ( .A(n31980), .B(n25675), .Y(n25653) );
  NOR2xp33_ASAP7_75t_SL U37796 ( .A(n25323), .B(n22415), .Y(n31700) );
  NOR2xp33_ASAP7_75t_SL U37797 ( .A(n32105), .B(n32104), .Y(n32106) );
  NOR4xp25_ASAP7_75t_SL U37798 ( .A(n26818), .B(n26816), .C(n26817), .D(n26815), .Y(n32103) );
  NOR2xp33_ASAP7_75t_SL U37799 ( .A(n22380), .B(n22378), .Y(n33056) );
  NOR2xp33_ASAP7_75t_SL U37800 ( .A(n32082), .B(n31809), .Y(n25602) );
  NOR2xp33_ASAP7_75t_SL U37801 ( .A(n32085), .B(n25601), .Y(n25603) );
  NOR2xp33_ASAP7_75t_SL U37802 ( .A(n32122), .B(n31934), .Y(n31935) );
  NOR2xp33_ASAP7_75t_SL U37803 ( .A(n31385), .B(n22379), .Y(n31386) );
  NOR2xp33_ASAP7_75t_SL U37804 ( .A(n18842), .B(n31384), .Y(n32049) );
  NAND2xp33_ASAP7_75t_SRAM U37805 ( .A(n24910), .B(n32050), .Y(n31651) );
  NOR2xp33_ASAP7_75t_SL U37806 ( .A(u0_0_leon3x0_p0_iu_r_D__DIVRDY_), .B(
        n32084), .Y(n24910) );
  AOI31xp33_ASAP7_75t_SL U37807 ( .A1(n32123), .A2(n3880), .A3(n32044), .B(
        n32689), .Y(n32045) );
  NOR2xp33_ASAP7_75t_SL U37808 ( .A(n31878), .B(n32123), .Y(n31879) );
  NOR2xp33_ASAP7_75t_SL U37809 ( .A(n31886), .B(n18876), .Y(n31887) );
  NOR2xp33_ASAP7_75t_SL U37810 ( .A(u0_0_leon3x0_p0_ici[29]), .B(n31890), .Y(
        n31888) );
  NOR2xp33_ASAP7_75t_SL U37811 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_UNDERRUN_), 
        .B(n31892), .Y(n31893) );
  NOR2xp33_ASAP7_75t_SL U37812 ( .A(n32713), .B(n31428), .Y(n31430) );
  NOR2xp33_ASAP7_75t_SL U37813 ( .A(n25449), .B(n26352), .Y(n25450) );
  NOR2xp33_ASAP7_75t_SL U37814 ( .A(n24869), .B(n25214), .Y(n24870) );
  NOR2xp33_ASAP7_75t_SL U37815 ( .A(u0_0_leon3x0_p0_iu_r_A__CTRL__ANNUL_), .B(
        n18798), .Y(n30682) );
  AOI31xp33_ASAP7_75t_SL U37816 ( .A1(n31652), .A2(n3725), .A3(n23229), .B(
        n31676), .Y(n28288) );
  NOR2xp33_ASAP7_75t_SL U37817 ( .A(n28285), .B(n31814), .Y(n31652) );
  NOR2xp33_ASAP7_75t_SL U37818 ( .A(u0_0_leon3x0_p0_div0_r_X__31_), .B(n29110), 
        .Y(n28284) );
  NAND2xp33_ASAP7_75t_SRAM U37819 ( .A(n32496), .B(n32662), .Y(n31319) );
  NOR2xp33_ASAP7_75t_SL U37820 ( .A(n32496), .B(n31318), .Y(n32481) );
  NOR2xp33_ASAP7_75t_SL U37821 ( .A(n30206), .B(n31447), .Y(n32199) );
  AND2x2_ASAP7_75t_SL U37822 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_NOMDS_), .B(
        n31574), .Y(n30207) );
  NOR4xp25_ASAP7_75t_SL U37823 ( .A(n22436), .B(add_x_735_A_29_), .C(n22721), 
        .D(add_x_735_A_9_), .Y(n31666) );
  NOR2xp33_ASAP7_75t_SL U37824 ( .A(n4318), .B(n32729), .Y(n32029) );
  NOR2xp33_ASAP7_75t_SL U37825 ( .A(n32664), .B(n32663), .Y(n2936) );
  AOI211xp5_ASAP7_75t_SL U37826 ( .A1(n32668), .A2(n32662), .B(n32674), .C(
        n22405), .Y(n32663) );
  NOR2xp33_ASAP7_75t_SL U37827 ( .A(n32668), .B(n32662), .Y(n32674) );
  NOR2xp33_ASAP7_75t_SL U37828 ( .A(n31594), .B(n31593), .Y(n31595) );
  NOR2xp33_ASAP7_75t_SL U37829 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_RBURST_), 
        .B(n30916), .Y(n31308) );
  NOR2xp33_ASAP7_75t_SL U37830 ( .A(n26658), .B(n26467), .Y(n30790) );
  NOR2xp33_ASAP7_75t_SL U37831 ( .A(n31584), .B(n31572), .Y(n31577) );
  AOI31xp33_ASAP7_75t_SL U37832 ( .A1(n29999), .A2(ahbso_0__HRESP__0_), .A3(
        n25599), .B(n25598), .Y(n32455) );
  NOR2xp33_ASAP7_75t_SL U37833 ( .A(n32037), .B(n31802), .Y(n25598) );
  NOR2xp33_ASAP7_75t_SL U37834 ( .A(n29889), .B(n29888), .Y(n29890) );
  NOR4xp25_ASAP7_75t_SL U37835 ( .A(u0_0_leon3x0_p0_div0_addout_27_), .B(
        u0_0_leon3x0_p0_div0_addout_28_), .C(u0_0_leon3x0_p0_div0_addout_29_), 
        .D(u0_0_leon3x0_p0_div0_addout_30_), .Y(n25932) );
  NOR4xp25_ASAP7_75t_SL U37836 ( .A(u0_0_leon3x0_p0_div0_addout_25_), .B(
        u0_0_leon3x0_p0_div0_addout_26_), .C(u0_0_leon3x0_p0_div0_addout_23_), 
        .D(u0_0_leon3x0_p0_div0_addout_24_), .Y(n25933) );
  NOR4xp25_ASAP7_75t_SL U37837 ( .A(u0_0_leon3x0_p0_div0_addout_19_), .B(
        u0_0_leon3x0_p0_div0_addout_20_), .C(u0_0_leon3x0_p0_div0_addout_21_), 
        .D(u0_0_leon3x0_p0_div0_addout_22_), .Y(n25934) );
  NOR4xp25_ASAP7_75t_SL U37838 ( .A(n25926), .B(u0_0_leon3x0_p0_div0_addout_8_), .C(u0_0_leon3x0_p0_div0_addout_6_), .D(u0_0_leon3x0_p0_div0_addout_7_), .Y(
        n25928) );
  NOR4xp25_ASAP7_75t_SL U37839 ( .A(u0_0_leon3x0_p0_div0_addout_3_), .B(
        u0_0_leon3x0_p0_div0_addout_2_), .C(u0_0_leon3x0_p0_div0_addout_0_), 
        .D(u0_0_leon3x0_p0_div0_addout_1_), .Y(n25924) );
  NOR2xp33_ASAP7_75t_SL U37840 ( .A(u0_0_leon3x0_p0_divi[18]), .B(n24630), .Y(
        n28535) );
  NOR2xp33_ASAP7_75t_SL U37841 ( .A(u0_0_leon3x0_p0_divi[19]), .B(n24630), .Y(
        n28524) );
  NOR2xp33_ASAP7_75t_SL U37842 ( .A(u0_0_leon3x0_p0_divi[21]), .B(n24630), .Y(
        n28517) );
  NOR2xp33_ASAP7_75t_SL U37843 ( .A(u0_0_leon3x0_p0_divi[22]), .B(n24630), .Y(
        n28473) );
  NOR2xp33_ASAP7_75t_SL U37844 ( .A(u0_0_leon3x0_p0_divi[23]), .B(n24630), .Y(
        n28470) );
  NOR2xp33_ASAP7_75t_SL U37845 ( .A(u0_0_leon3x0_p0_divi[24]), .B(n24630), .Y(
        n28460) );
  NOR2xp33_ASAP7_75t_SL U37846 ( .A(u0_0_leon3x0_p0_divi[25]), .B(n24630), .Y(
        n28401) );
  NOR2xp33_ASAP7_75t_SL U37847 ( .A(u0_0_leon3x0_p0_divi[27]), .B(n24630), .Y(
        n28382) );
  NOR4xp25_ASAP7_75t_SL U37848 ( .A(u0_0_leon3x0_p0_div0_addout_11_), .B(
        u0_0_leon3x0_p0_div0_addout_13_), .C(u0_0_leon3x0_p0_div0_addout_14_), 
        .D(u0_0_leon3x0_p0_div0_addout_12_), .Y(n25921) );
  NOR2xp33_ASAP7_75t_SL U37849 ( .A(u0_0_leon3x0_p0_divi[17]), .B(n24630), .Y(
        n28549) );
  NOR2xp33_ASAP7_75t_SL U37850 ( .A(u0_0_leon3x0_p0_divi[3]), .B(n24630), .Y(
        n28867) );
  NOR2xp33_ASAP7_75t_SL U37851 ( .A(u0_0_leon3x0_p0_divi[4]), .B(n24630), .Y(
        n28819) );
  NOR2xp33_ASAP7_75t_SL U37852 ( .A(u0_0_leon3x0_p0_divi[5]), .B(n24630), .Y(
        n28810) );
  NOR2xp33_ASAP7_75t_SL U37853 ( .A(u0_0_leon3x0_p0_divi[6]), .B(n24630), .Y(
        n28804) );
  NOR2xp33_ASAP7_75t_SL U37854 ( .A(n18909), .B(n24630), .Y(n28960) );
  NOR2xp33_ASAP7_75t_SL U37855 ( .A(n22431), .B(u0_0_leon3x0_p0_divi[0]), .Y(
        n29021) );
  NOR2xp33_ASAP7_75t_SL U37856 ( .A(u0_0_leon3x0_p0_divi[1]), .B(n24630), .Y(
        n28959) );
  NOR2xp33_ASAP7_75t_SL U37857 ( .A(u0_0_leon3x0_p0_divi[2]), .B(n24630), .Y(
        n28907) );
  NOR2xp33_ASAP7_75t_SL U37858 ( .A(n18904), .B(n24630), .Y(n28758) );
  NOR2xp33_ASAP7_75t_SL U37859 ( .A(n18890), .B(n24630), .Y(n28717) );
  NOR2xp33_ASAP7_75t_SL U37860 ( .A(u0_0_leon3x0_p0_divi[9]), .B(n24630), .Y(
        n28716) );
  NOR2xp33_ASAP7_75t_SL U37861 ( .A(u0_0_leon3x0_p0_divi[10]), .B(n24630), .Y(
        n28700) );
  NOR2xp33_ASAP7_75t_SL U37862 ( .A(u0_0_leon3x0_p0_divi[11]), .B(n24630), .Y(
        n28657) );
  NOR2xp33_ASAP7_75t_SL U37863 ( .A(u0_0_leon3x0_p0_divi[12]), .B(n24630), .Y(
        n28612) );
  NOR2xp33_ASAP7_75t_SL U37864 ( .A(u0_0_leon3x0_p0_divi[13]), .B(n24630), .Y(
        n28587) );
  NOR2xp33_ASAP7_75t_SL U37865 ( .A(u0_0_leon3x0_p0_divi[14]), .B(n24630), .Y(
        n28582) );
  NOR2xp33_ASAP7_75t_SL U37866 ( .A(u0_0_leon3x0_p0_divi[15]), .B(n24630), .Y(
        n28561) );
  NOR2xp33_ASAP7_75t_SL U37867 ( .A(u0_0_leon3x0_p0_divi[16]), .B(n24630), .Y(
        n28550) );
  AOI31xp33_ASAP7_75t_SL U37868 ( .A1(n31624), .A2(n31623), .A3(n31622), .B(
        n22380), .Y(u0_0_leon3x0_p0_c0mmu_dcache0_v_REQ_) );
  NAND2xp33_ASAP7_75t_SRAM U37869 ( .A(n31460), .B(n32030), .Y(n31622) );
  NOR2xp33_ASAP7_75t_SL U37870 ( .A(n31573), .B(n31572), .Y(n25588) );
  NOR2xp33_ASAP7_75t_SL U37871 ( .A(n32245), .B(n31609), .Y(n32273) );
  NOR2xp33_ASAP7_75t_SL U37872 ( .A(n2963), .B(n31306), .Y(n31608) );
  NOR2xp33_ASAP7_75t_SL U37873 ( .A(n23885), .B(n31601), .Y(n31614) );
  NOR2xp33_ASAP7_75t_SL U37874 ( .A(n31585), .B(n31463), .Y(n31299) );
  NOR2xp33_ASAP7_75t_SL U37875 ( .A(n30172), .B(n30182), .Y(n30173) );
  NOR2xp33_ASAP7_75t_SL U37876 ( .A(n30182), .B(n30175), .Y(n30167) );
  AOI211xp5_ASAP7_75t_SL U37877 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__19_), .A2(n22382), .B(
        n26541), .C(n26540), .Y(n2352) );
  NOR2xp33_ASAP7_75t_SL U37878 ( .A(n26539), .B(n18877), .Y(n26540) );
  AOI211xp5_ASAP7_75t_SL U37879 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__23_), .A2(n22382), .B(
        n26528), .C(n26527), .Y(n4416) );
  NOR2xp33_ASAP7_75t_SL U37880 ( .A(n26526), .B(n31633), .Y(n26527) );
  NOR2xp33_ASAP7_75t_SL U37881 ( .A(n30263), .B(n22376), .Y(n26415) );
  AOI211xp5_ASAP7_75t_SL U37882 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__5_), .A2(n22382), .B(n30028), .C(n30027), .Y(n4744) );
  NOR2xp33_ASAP7_75t_SL U37883 ( .A(n32851), .B(n31633), .Y(n30027) );
  AOI211xp5_ASAP7_75t_SL U37884 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__30_), .A2(n22382), .B(
        n25647), .C(n25646), .Y(n4738) );
  NOR2xp33_ASAP7_75t_SL U37885 ( .A(n32966), .B(n31633), .Y(n25646) );
  NOR2xp33_ASAP7_75t_SL U37886 ( .A(n30213), .B(n22376), .Y(n25643) );
  AOI211xp5_ASAP7_75t_SL U37887 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__22_), .A2(n22382), .B(
        n31636), .C(n31635), .Y(n4575) );
  NOR2xp33_ASAP7_75t_SL U37888 ( .A(n31634), .B(n31633), .Y(n31635) );
  AOI211xp5_ASAP7_75t_SL U37889 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__14_), .A2(n22382), .B(
        n25633), .C(n25632), .Y(n2327) );
  NOR2xp33_ASAP7_75t_SL U37890 ( .A(n25631), .B(n18877), .Y(n25632) );
  NOR2xp33_ASAP7_75t_SL U37891 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__14_), .B(
        n30007), .Y(n25630) );
  NOR2xp33_ASAP7_75t_SL U37892 ( .A(n25624), .B(n25623), .Y(n25628) );
  AOI211xp5_ASAP7_75t_SL U37893 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__17_), .A2(n22382), .B(
        n27289), .C(n27288), .Y(n4034) );
  NOR2xp33_ASAP7_75t_SL U37894 ( .A(n27287), .B(n18877), .Y(n27288) );
  AOI211xp5_ASAP7_75t_SL U37895 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__25_), .A2(n22382), .B(
        n31366), .C(n31365), .Y(n4626) );
  NOR2xp33_ASAP7_75t_SL U37896 ( .A(n32926), .B(n31633), .Y(n31365) );
  AOI211xp5_ASAP7_75t_SL U37897 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__26_), .A2(n22382), .B(
        n26496), .C(n26495), .Y(n4616) );
  NOR2xp33_ASAP7_75t_SL U37898 ( .A(n32934), .B(n31633), .Y(n26495) );
  NOR2xp33_ASAP7_75t_SL U37899 ( .A(n29801), .B(n30007), .Y(n26226) );
  AOI211xp5_ASAP7_75t_SL U37900 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__3_), .A2(n22382), .B(n29508), .C(n29507), .Y(n4692) );
  NOR2xp33_ASAP7_75t_SL U37901 ( .A(n32847), .B(n31633), .Y(n29507) );
  NOR2xp33_ASAP7_75t_SL U37902 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__3_), .B(
        n30007), .Y(n29503) );
  AOI211xp5_ASAP7_75t_SL U37903 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__1_), .A2(n22382), .B(n27492), .C(n27491), .Y(n4534) );
  NOR2xp33_ASAP7_75t_SL U37904 ( .A(n32843), .B(n31633), .Y(n27491) );
  AOI211xp5_ASAP7_75t_SL U37905 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__24_), .A2(n22382), .B(
        n26516), .C(n26515), .Y(n2274) );
  NOR2xp33_ASAP7_75t_SL U37906 ( .A(n32916), .B(n31633), .Y(n26515) );
  AOI211xp5_ASAP7_75t_SL U37907 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__27_), .A2(n22382), .B(
        n30892), .C(n30891), .Y(n4528) );
  NOR2xp33_ASAP7_75t_SL U37908 ( .A(n32942), .B(n31633), .Y(n30891) );
  AOI211xp5_ASAP7_75t_SL U37909 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__21_), .A2(n22382), .B(
        n29293), .C(n29292), .Y(n2328) );
  NOR2xp33_ASAP7_75t_SL U37910 ( .A(n29291), .B(n31633), .Y(n29292) );
  AOI211xp5_ASAP7_75t_SL U37911 ( .A1(n28403), .A2(n28521), .B(n26327), .C(
        n26483), .Y(n26328) );
  AOI211xp5_ASAP7_75t_SL U37912 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__10_), .A2(n22382), .B(
        n26616), .C(n26615), .Y(n4458) );
  NOR2xp33_ASAP7_75t_SL U37913 ( .A(n26614), .B(n18877), .Y(n26615) );
  AOI211xp5_ASAP7_75t_SL U37914 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__12_), .A2(n22382), .B(
        n29850), .C(n29849), .Y(n4755) );
  NOR2xp33_ASAP7_75t_SL U37915 ( .A(n29848), .B(n18877), .Y(n29849) );
  AOI211xp5_ASAP7_75t_SL U37916 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__31_), .A2(n22382), .B(
        n26460), .C(n26459), .Y(n4772) );
  NOR2xp33_ASAP7_75t_SL U37917 ( .A(n32976), .B(n31633), .Y(n26459) );
  AOI211xp5_ASAP7_75t_SL U37918 ( .A1(n28405), .A2(n26585), .B(n26456), .C(
        n26455), .Y(n26458) );
  NOR2xp33_ASAP7_75t_SL U37919 ( .A(n26734), .B(n26522), .Y(n26455) );
  NOR2xp33_ASAP7_75t_SL U37920 ( .A(n25207), .B(n30007), .Y(n26456) );
  AOI211xp5_ASAP7_75t_SL U37921 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__11_), .A2(n22382), .B(
        n28137), .C(n28136), .Y(n4522) );
  NOR2xp33_ASAP7_75t_SL U37922 ( .A(n28135), .B(n18877), .Y(n28136) );
  NOR2xp33_ASAP7_75t_SL U37923 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .B(
        n26169), .Y(n26341) );
  AOI211xp5_ASAP7_75t_SL U37924 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__9_), .A2(n22382), .B(n30133), .C(n30132), .Y(n1805) );
  NOR2xp33_ASAP7_75t_SL U37925 ( .A(n30131), .B(n18877), .Y(n30132) );
  AOI211xp5_ASAP7_75t_SL U37926 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__28_), .A2(n22382), .B(
        n31493), .C(n31492), .Y(n1782) );
  NOR2xp33_ASAP7_75t_SL U37927 ( .A(n32950), .B(n31633), .Y(n31492) );
  NOR2xp33_ASAP7_75t_SL U37928 ( .A(n30235), .B(n22376), .Y(n25429) );
  AOI211xp5_ASAP7_75t_SL U37929 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__13_), .A2(n22382), .B(
        n26603), .C(n26602), .Y(n1767) );
  NOR2xp33_ASAP7_75t_SL U37930 ( .A(n26601), .B(n18877), .Y(n26602) );
  AOI211xp5_ASAP7_75t_SL U37931 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__2_), .A2(n22382), .B(n29567), .C(n29566), .Y(n4672) );
  NOR2xp33_ASAP7_75t_SL U37932 ( .A(n32845), .B(n31633), .Y(n29566) );
  AOI211xp5_ASAP7_75t_SL U37933 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__16_), .A2(n22382), .B(
        n26450), .C(n26449), .Y(n1774) );
  NOR2xp33_ASAP7_75t_SL U37934 ( .A(n26448), .B(n18877), .Y(n26449) );
  AOI211xp5_ASAP7_75t_SL U37935 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__18_), .A2(n22382), .B(
        n25845), .C(n25844), .Y(n4356) );
  NOR2xp33_ASAP7_75t_SL U37936 ( .A(n25843), .B(n18877), .Y(n25844) );
  AOI211xp5_ASAP7_75t_SL U37937 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__20_), .A2(n22382), .B(
        n31524), .C(n31523), .Y(n4499) );
  NOR2xp33_ASAP7_75t_SL U37938 ( .A(n31522), .B(n18877), .Y(n31523) );
  AOI211xp5_ASAP7_75t_SL U37939 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__8_), .A2(n22382), .B(n25524), .C(n25523), .Y(n4686) );
  NOR2xp33_ASAP7_75t_SL U37940 ( .A(n25522), .B(n31633), .Y(n25523) );
  AOI211xp5_ASAP7_75t_SL U37941 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__29_), .A2(n22382), .B(
        n26490), .C(n26489), .Y(n4666) );
  NOR2xp33_ASAP7_75t_SL U37942 ( .A(n32958), .B(n31633), .Y(n26489) );
  NOR2xp33_ASAP7_75t_SL U37943 ( .A(n18381), .B(n22392), .Y(n25893) );
  AOI211xp5_ASAP7_75t_SL U37944 ( .A1(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_WB__DATA2__15_), .A2(n22382), .B(
        n26591), .C(n26590), .Y(n4637) );
  NOR2xp33_ASAP7_75t_SL U37945 ( .A(n26589), .B(n18877), .Y(n26590) );
  NOR2xp33_ASAP7_75t_SL U37946 ( .A(n25901), .B(n25488), .Y(n26574) );
  NOR2xp33_ASAP7_75t_SL U37947 ( .A(n32606), .B(n31632), .Y(n25872) );
  NOR2xp33_ASAP7_75t_SL U37948 ( .A(n29499), .B(n26338), .Y(n25423) );
  NOR2xp33_ASAP7_75t_SL U37949 ( .A(n32612), .B(n31632), .Y(n29936) );
  NOR2xp33_ASAP7_75t_SL U37950 ( .A(n32713), .B(n31632), .Y(n28103) );
  NOR2xp33_ASAP7_75t_SL U37951 ( .A(n30006), .B(n29009), .Y(n28102) );
  NOR2xp33_ASAP7_75t_SL U37952 ( .A(n32610), .B(n31632), .Y(n25858) );
  NOR2xp33_ASAP7_75t_SL U37953 ( .A(n25237), .B(n18891), .Y(n25126) );
  NOR2xp33_ASAP7_75t_SL U37954 ( .A(n26514), .B(n18891), .Y(n26382) );
  NOR2xp33_ASAP7_75t_SL U37955 ( .A(n26562), .B(n18891), .Y(n26564) );
  NOR2xp33_ASAP7_75t_SL U37956 ( .A(n27110), .B(n18891), .Y(n27112) );
  AND2x2_ASAP7_75t_SL U37957 ( .A(n22379), .B(n31824), .Y(n31989) );
  AOI211xp5_ASAP7_75t_SL U37958 ( .A1(n28255), .A2(n24818), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__7_), .C(n32171), .Y(n24824) );
  NOR2xp33_ASAP7_75t_SL U37959 ( .A(n24876), .B(n24741), .Y(n24742) );
  NOR2xp33_ASAP7_75t_SL U37960 ( .A(n26817), .B(n24876), .Y(n24881) );
  NOR2xp33_ASAP7_75t_SL U37961 ( .A(n26192), .B(n26191), .Y(n26193) );
  NAND2xp33_ASAP7_75t_SRAM U37962 ( .A(n24688), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__5_), .Y(n26301) );
  NAND2xp33_ASAP7_75t_SRAM U37963 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__11_), 
        .B(n24688), .Y(n28676) );
  NAND2xp33_ASAP7_75t_SRAM U37964 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__14_), 
        .B(n24688), .Y(n27192) );
  NAND2xp33_ASAP7_75t_SRAM U37965 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__30_), 
        .B(n24688), .Y(n28380) );
  NAND2xp33_ASAP7_75t_SRAM U37966 ( .A(n24688), .B(
        u0_0_leon3x0_p0_iu_r_X__DATA__0__20_), .Y(n26987) );
  NAND2xp33_ASAP7_75t_SRAM U37967 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__22_), 
        .B(n24688), .Y(n28478) );
  OR2x2_ASAP7_75t_SL U37968 ( .A(n24548), .B(n24530), .Y(n24429) );
  AND2x2_ASAP7_75t_SL U37969 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__11_), .B(
        n28769), .Y(n24432) );
  OA21x2_ASAP7_75t_SL U37970 ( .A1(n32333), .A2(n22402), .B(n28518), .Y(n24433) );
  OA21x2_ASAP7_75t_SL U37971 ( .A1(n32322), .A2(n22402), .B(n25573), .Y(n24434) );
  OA21x2_ASAP7_75t_SL U37972 ( .A1(n32328), .A2(n22402), .B(n26969), .Y(n24435) );
  OA21x2_ASAP7_75t_SL U37973 ( .A1(n32354), .A2(n22402), .B(n28383), .Y(n24436) );
  OA21x2_ASAP7_75t_SL U37974 ( .A1(n31032), .A2(n22402), .B(n28412), .Y(n24437) );
  OA21x2_ASAP7_75t_SL U37975 ( .A1(n32410), .A2(n22402), .B(n32061), .Y(n24438) );
  OA21x2_ASAP7_75t_SL U37976 ( .A1(n32419), .A2(n22402), .B(n31942), .Y(n24439) );
  OA21x2_ASAP7_75t_SL U37977 ( .A1(n32361), .A2(n22402), .B(n30919), .Y(n24440) );
  OA21x2_ASAP7_75t_SL U37978 ( .A1(n32399), .A2(n22402), .B(n31332), .Y(n24441) );
  OA21x2_ASAP7_75t_SL U37979 ( .A1(n32430), .A2(n22402), .B(n31957), .Y(n24442) );
  OA21x2_ASAP7_75t_SL U37980 ( .A1(n30876), .A2(n22402), .B(n30875), .Y(n24443) );
  OA21x2_ASAP7_75t_SL U37981 ( .A1(n30557), .A2(n22402), .B(n28461), .Y(n24444) );
  OA21x2_ASAP7_75t_SL U37982 ( .A1(n30155), .A2(n22402), .B(n30154), .Y(n24445) );
  OA21x2_ASAP7_75t_SL U37983 ( .A1(n32371), .A2(n22402), .B(n32009), .Y(n24446) );
  OA21x2_ASAP7_75t_SL U37984 ( .A1(n32380), .A2(n22402), .B(n31856), .Y(n24447) );
  OA21x2_ASAP7_75t_SL U37985 ( .A1(n32384), .A2(n22402), .B(n31979), .Y(n24448) );
  OA21x2_ASAP7_75t_SL U37986 ( .A1(n32377), .A2(n22402), .B(n31536), .Y(n24449) );
  OA21x2_ASAP7_75t_SL U37987 ( .A1(n32382), .A2(n22402), .B(n31650), .Y(n24450) );
  OA21x2_ASAP7_75t_SL U37988 ( .A1(n32367), .A2(n22402), .B(n29574), .Y(n24451) );
  OA21x2_ASAP7_75t_SL U37989 ( .A1(n31509), .A2(n22402), .B(n31508), .Y(n24452) );
  OA21x2_ASAP7_75t_SL U37990 ( .A1(n30904), .A2(n22402), .B(n30903), .Y(n24453) );
  OA21x2_ASAP7_75t_SL U37991 ( .A1(n31378), .A2(n22402), .B(n31377), .Y(n24454) );
  OA21x2_ASAP7_75t_SL U37992 ( .A1(n32315), .A2(n22402), .B(n31253), .Y(n24455) );
  OA21x2_ASAP7_75t_SL U37993 ( .A1(n32391), .A2(n22402), .B(n32047), .Y(n24456) );
  OA21x2_ASAP7_75t_SL U37994 ( .A1(n32311), .A2(n22402), .B(n30113), .Y(n24457) );
  OA21x2_ASAP7_75t_SL U37995 ( .A1(n30808), .A2(n22402), .B(n30807), .Y(n24458) );
  AND2x2_ASAP7_75t_SL U37996 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__14_), .B(
        n28769), .Y(n24459) );
  AND2x2_ASAP7_75t_SL U37997 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__5_), .B(
        n28769), .Y(n24460) );
  AND2x2_ASAP7_75t_SL U37998 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__17_), .B(
        n28769), .Y(n24461) );
  AND2x2_ASAP7_75t_SL U37999 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__10_), .B(
        n28769), .Y(n24462) );
  AND2x2_ASAP7_75t_SL U38000 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__20_), .B(
        n28769), .Y(n24463) );
  AND2x2_ASAP7_75t_SL U38001 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__21_), .B(
        n28769), .Y(n24464) );
  AND2x2_ASAP7_75t_SL U38002 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__23_), .B(
        n28769), .Y(n24465) );
  AND2x2_ASAP7_75t_SL U38003 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__22_), .B(
        n28769), .Y(n24466) );
  AND2x2_ASAP7_75t_SL U38004 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__29_), .B(
        n28769), .Y(n24467) );
  AND2x2_ASAP7_75t_SL U38005 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__30_), .B(
        n28769), .Y(n24468) );
  AO22x1_ASAP7_75t_SL U38006 ( .A1(n26376), .A2(n27098), .B1(n28967), .B2(
        n27091), .Y(n24470) );
  AND3x1_ASAP7_75t_SL U38007 ( .A(n25043), .B(n25042), .C(n25041), .Y(n24471)
         );
  OR2x2_ASAP7_75t_SL U38008 ( .A(n27108), .B(n25908), .Y(n24472) );
  AND2x2_ASAP7_75t_SL U38009 ( .A(add_x_735_A_2_), .B(n22416), .Y(n24473) );
  OR2x2_ASAP7_75t_SL U38010 ( .A(n4391), .B(ahbso_1__HREADY_), .Y(n24474) );
  AND2x2_ASAP7_75t_SL U38011 ( .A(n22449), .B(n22416), .Y(n24475) );
  AND2x2_ASAP7_75t_SL U38012 ( .A(n29899), .B(n22392), .Y(n24476) );
  OR2x2_ASAP7_75t_SL U38013 ( .A(n22902), .B(n24469), .Y(n24477) );
  OR2x2_ASAP7_75t_SL U38014 ( .A(n22902), .B(n22392), .Y(n24478) );
  AND2x2_ASAP7_75t_SL U38015 ( .A(n24579), .B(u0_0_leon3x0_p0_divi[30]), .Y(
        n24480) );
  AND2x2_ASAP7_75t_SL U38016 ( .A(n29680), .B(n22392), .Y(n24481) );
  AO22x1_ASAP7_75t_SL U38017 ( .A1(dc_q[12]), .A2(n31004), .B1(dt_q[8]), .B2(
        n29991), .Y(n24482) );
  AO22x1_ASAP7_75t_SL U38018 ( .A1(dc_q[13]), .A2(n31004), .B1(dt_q[9]), .B2(
        n24573), .Y(n24483) );
  OA21x2_ASAP7_75t_SL U38019 ( .A1(n28824), .A2(n28823), .B(n28822), .Y(n24485) );
  OA21x2_ASAP7_75t_SL U38020 ( .A1(n18296), .A2(n28827), .B(
        u0_0_leon3x0_p0_divi[22]), .Y(n24487) );
  AND2x2_ASAP7_75t_SL U38021 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .B(
        n28824), .Y(n24488) );
  AND2x2_ASAP7_75t_SL U38022 ( .A(n28830), .B(n18904), .Y(n24489) );
  OA211x2_ASAP7_75t_SL U38023 ( .A1(n32306), .A2(n31470), .B(n30880), .C(
        n30879), .Y(n24490) );
  AO21x1_ASAP7_75t_SL U38024 ( .A1(n29148), .A2(n22902), .B(n24631), .Y(n24492) );
  OA21x2_ASAP7_75t_SL U38025 ( .A1(n18876), .A2(n31687), .B(n25885), .Y(n24493) );
  AND3x1_ASAP7_75t_SL U38026 ( .A(n32023), .B(n24896), .C(n25244), .Y(n24494)
         );
  OR2x2_ASAP7_75t_SL U38027 ( .A(n25939), .B(n30580), .Y(n24496) );
  OR2x2_ASAP7_75t_SL U38028 ( .A(n26348), .B(n30580), .Y(n24498) );
  OR2x2_ASAP7_75t_SL U38029 ( .A(n26370), .B(n30580), .Y(n24499) );
  OR2x2_ASAP7_75t_SL U38030 ( .A(n28471), .B(n30580), .Y(n24500) );
  OR2x2_ASAP7_75t_SL U38031 ( .A(n29862), .B(n30580), .Y(n24501) );
  OR2x2_ASAP7_75t_SL U38032 ( .A(n28384), .B(n30580), .Y(n24502) );
  OR2x2_ASAP7_75t_SL U38033 ( .A(n28462), .B(n30580), .Y(n24503) );
  OR2x2_ASAP7_75t_SL U38034 ( .A(n28519), .B(n30580), .Y(n24504) );
  OR2x2_ASAP7_75t_SL U38035 ( .A(n26970), .B(n30580), .Y(n24505) );
  OR2x2_ASAP7_75t_SL U38036 ( .A(n28525), .B(n30580), .Y(n24506) );
  OR2x2_ASAP7_75t_SL U38037 ( .A(u0_0_leon3x0_p0_iu_r_A__CTRL__TT__0_), .B(
        n22378), .Y(n24510) );
  AND2x2_ASAP7_75t_SL U38038 ( .A(ahbso_0__HRDATA__24_), .B(n29999), .Y(n24512) );
  OR2x2_ASAP7_75t_SL U38039 ( .A(u0_0_leon3x0_p0_c0mmu_a0_r_HCACHE_), .B(
        n32451), .Y(n24513) );
  OR2x2_ASAP7_75t_SL U38040 ( .A(n22380), .B(n25402), .Y(n24515) );
  AND2x2_ASAP7_75t_SL U38041 ( .A(u0_0_leon3x0_p0_iu_v_E__RFE1_), .B(n24659), 
        .Y(n24516) );
  AND2x2_ASAP7_75t_SL U38042 ( .A(ahbso_0__HRDATA__12_), .B(n29999), .Y(n24518) );
  OR2x2_ASAP7_75t_SL U38043 ( .A(n22999), .B(add_x_735_A_2_), .Y(n24519) );
  AND2x2_ASAP7_75t_SL U38044 ( .A(uart1_r_THOLD__30__2_), .B(n28018), .Y(
        n24520) );
  AND2x2_ASAP7_75t_SL U38045 ( .A(uart1_r_THOLD__28__5_), .B(n28018), .Y(
        n24522) );
  OR2x2_ASAP7_75t_SL U38046 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__8_), .B(
        n24646), .Y(n24523) );
  OR2x2_ASAP7_75t_SL U38047 ( .A(n22427), .B(n25075), .Y(n24524) );
  OR2x2_ASAP7_75t_SL U38048 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .B(
        n24983), .Y(n24526) );
  AND2x2_ASAP7_75t_SL U38049 ( .A(uart1_r_THOLD__30__3_), .B(n28018), .Y(
        n24529) );
  OR2x2_ASAP7_75t_SL U38050 ( .A(u0_0_leon3x0_p0_dci[2]), .B(n25587), .Y(
        n24530) );
  OR2x2_ASAP7_75t_SL U38051 ( .A(n25534), .B(n27328), .Y(n24531) );
  OR2x2_ASAP7_75t_SL U38052 ( .A(u0_0_leon3x0_p0_div0_r_QMSB_), .B(n31672), 
        .Y(n24532) );
  OA211x2_ASAP7_75t_SL U38053 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__ICS__1_), .A2(u0_0_leon3x0_p0_c0mmu_icache0_r_HIT_), .B(n32482), .C(
        u0_0_leon3x0_p0_c0mmu_a0_r_HCACHE_), .Y(n24533) );
  OR2x2_ASAP7_75t_SL U38054 ( .A(n31276), .B(n31275), .Y(n24534) );
  AND2x2_ASAP7_75t_SL U38055 ( .A(ahbso_0__HRDATA__5_), .B(n29999), .Y(n24535)
         );
  OR2x2_ASAP7_75t_SL U38056 ( .A(n4775), .B(n2851), .Y(n24536) );
  AND2x2_ASAP7_75t_SL U38057 ( .A(ahbso_0__HRDATA__6_), .B(n29999), .Y(n24537)
         );
  OR2x2_ASAP7_75t_SL U38058 ( .A(n25452), .B(n26758), .Y(n24538) );
  OA21x2_ASAP7_75t_SL U38059 ( .A1(n29831), .A2(n31396), .B(n29616), .Y(n24539) );
  AND2x2_ASAP7_75t_SL U38060 ( .A(sr1_r_MCFG1__IOEN_), .B(n32003), .Y(n24540)
         );
  AND3x1_ASAP7_75t_SL U38061 ( .A(n25722), .B(n30685), .C(n30684), .Y(n24542)
         );
  OA21x2_ASAP7_75t_SL U38062 ( .A1(n32290), .A2(n32144), .B(n32143), .Y(n24543) );
  NOR3xp33_ASAP7_75t_SL U38063 ( .A(n31257), .B(n24429), .C(n32198), .Y(n24547) );
  NOR2xp33_ASAP7_75t_SL U38064 ( .A(n24492), .B(u0_0_leon3x0_p0_divi[5]), .Y(
        n26265) );
  HB1xp67_ASAP7_75t_SL U38065 ( .A(ic_address[9]), .Y(it_address[6]) );
  HB1xp67_ASAP7_75t_SL U38066 ( .A(ic_address[8]), .Y(it_address[5]) );
  HB1xp67_ASAP7_75t_SL U38067 ( .A(ic_address[7]), .Y(it_address[4]) );
  HB1xp67_ASAP7_75t_SL U38068 ( .A(ic_address[6]), .Y(it_address[3]) );
  HB1xp67_ASAP7_75t_SL U38069 ( .A(ic_address[5]), .Y(it_address[2]) );
  HB1xp67_ASAP7_75t_SL U38070 ( .A(ic_address[4]), .Y(it_address[1]) );
  HB1xp67_ASAP7_75t_SL U38071 ( .A(clk), .Y(clk_out) );
  HB1xp67_ASAP7_75t_SL U38072 ( .A(ic_address[3]), .Y(it_address[0]) );
  HB1xp67_ASAP7_75t_SL U38073 ( .A(dt_address[6]), .Y(dc_address[9]) );
  HB1xp67_ASAP7_75t_SL U38074 ( .A(dc_address[8]), .Y(dt_address[5]) );
  HB1xp67_ASAP7_75t_SL U38075 ( .A(dc_address[7]), .Y(dt_address[4]) );
  HB1xp67_ASAP7_75t_SL U38076 ( .A(dt_address[0]), .Y(dc_address[3]) );
  HB1xp67_ASAP7_75t_SL U38077 ( .A(dc_address[6]), .Y(dt_address[3]) );
  HB1xp67_ASAP7_75t_SL U38078 ( .A(dc_address[5]), .Y(dt_address[2]) );
  HB1xp67_ASAP7_75t_SL U38079 ( .A(dc_address[4]), .Y(dt_address[1]) );
  TIEHIx1_ASAP7_75t_SL U38080 ( .H(ramoen[4]) );
  NAND2xp33_ASAP7_75t_SRAM U38081 ( .A(n23396), .B(n26278), .Y(n26141) );
  NAND2xp33_ASAP7_75t_SRAM U38082 ( .A(n23396), .B(n22416), .Y(n25461) );
  NOR2xp33_ASAP7_75t_SL U38083 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__31_), .B(
        n18911), .Y(n25236) );
  NOR2xp33_ASAP7_75t_SL U38084 ( .A(n18614), .B(n28928), .Y(n26360) );
  NOR4xp25_ASAP7_75t_SL U38085 ( .A(n18530), .B(n23969), .C(n31668), .D(n31667), .Y(n31670) );
  AOI211xp5_ASAP7_75t_SL U38086 ( .A1(n29583), .A2(n23965), .B(n26708), .C(
        n26707), .Y(n26711) );
  AOI211xp5_ASAP7_75t_SL U38087 ( .A1(n24577), .A2(n23965), .B(n26155), .C(
        n26142), .Y(n26557) );
  AOI211xp5_ASAP7_75t_SL U38088 ( .A1(n22919), .A2(u0_0_leon3x0_p0_muli[8]), 
        .B(n32015), .C(n32014), .Y(n32020) );
  NOR4xp25_ASAP7_75t_SL U38089 ( .A(n32014), .B(u0_0_leon3x0_p0_muli[8]), .C(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_), .D(n32012), .Y(n24971) );
  AOI211xp5_ASAP7_75t_SL U38090 ( .A1(n28928), .A2(n24231), .B(n24631), .C(
        u0_0_leon3x0_p0_divi[18]), .Y(n25775) );
  OR2x2_ASAP7_75t_SL U38091 ( .A(n25177), .B(n25901), .Y(n24579) );
  OR2x2_ASAP7_75t_SL U38092 ( .A(n25177), .B(n25901), .Y(n24580) );
  OR2x2_ASAP7_75t_SL U38093 ( .A(u0_0_leon3x0_p0_iu_r_E__JMPL_), .B(n27067), 
        .Y(n24581) );
  OR2x2_ASAP7_75t_SL U38094 ( .A(u0_0_leon3x0_p0_iu_r_E__JMPL_), .B(n27067), 
        .Y(n24582) );
  NAND3xp33_ASAP7_75t_SL U38095 ( .A(n24599), .B(n24587), .C(n24600), .Y(
        n24586) );
  A2O1A1Ixp33_ASAP7_75t_SL U38096 ( .A1(n24587), .A2(n24600), .B(n24599), .C(
        n24586), .Y(uart1_scaler_10_) );
  NAND3xp33_ASAP7_75t_SL U38097 ( .A(n24607), .B(n24608), .C(n24609), .Y(
        n24588) );
  A2O1A1Ixp33_ASAP7_75t_SL U38098 ( .A1(n24608), .A2(n24609), .B(n24607), .C(
        n24588), .Y(uart1_scaler_2_) );
  NAND3xp33_ASAP7_75t_SL U38099 ( .A(n24606), .B(n24592), .C(n24607), .Y(
        n24589) );
  A2O1A1Ixp33_ASAP7_75t_SL U38100 ( .A1(n24592), .A2(n24607), .B(n24606), .C(
        n24589), .Y(uart1_scaler_3_) );
  NAND3xp33_ASAP7_75t_SL U38101 ( .A(n24605), .B(n24591), .C(n24606), .Y(
        n24590) );
  A2O1A1Ixp33_ASAP7_75t_SL U38102 ( .A1(n24591), .A2(n24606), .B(n24605), .C(
        n24590), .Y(uart1_scaler_4_) );
  NAND3xp33_ASAP7_75t_SL U38103 ( .A(n24600), .B(n24598), .C(n24601), .Y(
        n24597) );
  A2O1A1Ixp33_ASAP7_75t_SL U38104 ( .A1(n24598), .A2(n24601), .B(n24600), .C(
        n24597), .Y(uart1_scaler_9_) );
  NOR2xp33_ASAP7_75t_SL U38105 ( .A(uart1_uarto_SCALER__0_), .B(
        uart1_uarto_SCALER__1_), .Y(n24592) );
  NOR2xp33_ASAP7_75t_SL U38106 ( .A(uart1_uarto_SCALER__4_), .B(n24593), .Y(
        n24595) );
  NOR2xp33_ASAP7_75t_SL U38107 ( .A(uart1_uarto_SCALER__7_), .B(n24596), .Y(
        n24598) );
  NAND3xp33_ASAP7_75t_SL U38108 ( .A(n24626), .B(n24627), .C(n24628), .Y(
        n24610) );
  A2O1A1Ixp33_ASAP7_75t_SL U38109 ( .A1(n24627), .A2(n24628), .B(n24626), .C(
        n24610), .Y(timer0_scaler_2_) );
  NAND3xp33_ASAP7_75t_SL U38110 ( .A(n24625), .B(n24613), .C(n24626), .Y(
        n24611) );
  A2O1A1Ixp33_ASAP7_75t_SL U38111 ( .A1(n24613), .A2(n24626), .B(n24625), .C(
        n24611), .Y(timer0_scaler_3_) );
  NAND3xp33_ASAP7_75t_SL U38112 ( .A(n24624), .B(n24617), .C(n24625), .Y(
        n24612) );
  A2O1A1Ixp33_ASAP7_75t_SL U38113 ( .A1(n24617), .A2(n24625), .B(n24624), .C(
        n24612), .Y(timer0_scaler_4_) );
  NAND3xp33_ASAP7_75t_SL U38114 ( .A(n24623), .B(n24616), .C(n24624), .Y(
        n24615) );
  A2O1A1Ixp33_ASAP7_75t_SL U38115 ( .A1(n24616), .A2(n24624), .B(n24623), .C(
        n24615), .Y(timer0_scaler_5_) );
  NAND3xp33_ASAP7_75t_SL U38116 ( .A(n24622), .B(n24619), .C(n24623), .Y(
        n24618) );
  A2O1A1Ixp33_ASAP7_75t_SL U38117 ( .A1(n24619), .A2(n24623), .B(n24622), .C(
        n24618), .Y(timer0_scaler_6_) );
  NOR3xp33_ASAP7_75t_SL U38118 ( .A(timer0_r_SCALER__1_), .B(
        timer0_r_SCALER__2_), .C(timer0_r_SCALER__0_), .Y(n24617) );
  NOR3xp33_ASAP7_75t_SL U38119 ( .A(n24620), .B(timer0_r_SCALER__5_), .C(
        timer0_r_SCALER__4_), .Y(n24621) );
  NOR2xp33_ASAP7_75t_SL U38120 ( .A(timer0_r_SCALER__0_), .B(
        timer0_r_SCALER__1_), .Y(n24613) );
  NOR2xp33_ASAP7_75t_SL U38121 ( .A(timer0_r_SCALER__3_), .B(n24614), .Y(
        n24616) );
  NOR2xp33_ASAP7_75t_SL U38122 ( .A(timer0_r_SCALER__4_), .B(n24620), .Y(
        n24619) );
  A2O1A1Ixp33_ASAP7_75t_SL U38123 ( .A1(n32140), .A2(n24707), .B(n24678), .C(
        n24706), .Y(n3318) );
  A2O1A1Ixp33_ASAP7_75t_SL U38124 ( .A1(n25689), .A2(
        u0_0_leon3x0_p0_iu_de_icc_2_), .B(u0_0_leon3x0_p0_iu_de_icc_0_), .C(
        n24714), .Y(n24710) );
  NAND3xp33_ASAP7_75t_SL U38125 ( .A(n30677), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__26_), .C(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__25_), .Y(n24708) );
  O2A1O1Ixp5_ASAP7_75t_SL U38126 ( .A1(n24711), .A2(n24714), .B(n24710), .C(
        n24709), .Y(n24717) );
  XOR2xp5_ASAP7_75t_SL U38127 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__25_), 
        .B(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__26_), .Y(n24712) );
  O2A1O1Ixp5_ASAP7_75t_SL U38128 ( .A1(n24873), .A2(n24714), .B(n24713), .C(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__27_), .Y(n24718) );
  NOR3xp33_ASAP7_75t_SL U38129 ( .A(n24718), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__28_), .C(n24717), .Y(n24722) );
  NAND3xp33_ASAP7_75t_SL U38130 ( .A(n24850), .B(n24719), .C(n30952), .Y(
        n24856) );
  NOR3xp33_ASAP7_75t_SL U38131 ( .A(n24856), .B(
        u0_0_leon3x0_p0_iu_r_A__CTRL__ANNUL_), .C(n24720), .Y(n24721) );
  A2O1A1Ixp33_ASAP7_75t_SL U38132 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__28_), .A2(n24723), .B(n24722), .C(
        n24721), .Y(n25882) );
  O2A1O1Ixp5_ASAP7_75t_SL U38133 ( .A1(n25549), .A2(n25537), .B(
        u0_0_leon3x0_p0_iu_de_icc_2_), .C(u0_0_leon3x0_p0_iu_de_icc_0_), .Y(
        n24731) );
  A2O1A1Ixp33_ASAP7_75t_SL U38134 ( .A1(u0_0_leon3x0_p0_iu_de_icc_2_), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__25_), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_), .C(n25553), .Y(n24730) );
  O2A1O1Ixp5_ASAP7_75t_SL U38135 ( .A1(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__27_), .A2(n24873), .B(n24724), .C(n25537), .Y(n24725) );
  A2O1A1Ixp33_ASAP7_75t_SL U38136 ( .A1(n25537), .A2(n24726), .B(n24725), .C(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__26_), .Y(n24729) );
  O2A1O1Ixp5_ASAP7_75t_SL U38137 ( .A1(n24731), .A2(n24730), .B(n24729), .C(
        n24728), .Y(n24732) );
  XNOR2xp5_ASAP7_75t_SL U38138 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__INST__28_), 
        .B(n24732), .Y(n24733) );
  A2O1A1Ixp33_ASAP7_75t_SL U38139 ( .A1(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__29_), .A2(n25217), .B(
        u0_0_leon3x0_p0_iu_r_D__PV_), .C(n30682), .Y(n24737) );
  NAND3xp33_ASAP7_75t_SL U38140 ( .A(n24738), .B(n30503), .C(n24737), .Y(
        n24889) );
  OR2x2_ASAP7_75t_SL U38141 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__30_), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__31_), .Y(n25937) );
  NAND3xp33_ASAP7_75t_SL U38142 ( .A(n32052), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__23_), .C(n24855), .Y(n24739) );
  O2A1O1Ixp5_ASAP7_75t_SL U38143 ( .A1(n32082), .A2(n24743), .B(n32048), .C(
        n24742), .Y(n24770) );
  XNOR2xp5_ASAP7_75t_SL U38144 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__6_), .B(
        n32170), .Y(n24769) );
  A2O1A1Ixp33_ASAP7_75t_SL U38145 ( .A1(n4930), .A2(n3878), .B(n18867), .C(
        u0_0_leon3x0_p0_iu_v_M__CTRL__RD__7_), .Y(n24752) );
  XNOR2xp5_ASAP7_75t_SL U38146 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__0_), .B(
        DP_OP_1196_128_7433_n452), .Y(n24749) );
  XNOR2xp5_ASAP7_75t_SL U38147 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__2_), .B(
        DP_OP_1196_128_7433_n454), .Y(n24757) );
  XNOR2xp5_ASAP7_75t_SL U38148 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__1_), .B(
        DP_OP_1196_128_7433_n453), .Y(n24756) );
  NAND4xp25_ASAP7_75t_SL U38149 ( .A(n24758), .B(n24797), .C(n24757), .D(
        n24756), .Y(n24759) );
  O2A1O1Ixp5_ASAP7_75t_SL U38150 ( .A1(n24762), .A2(n24761), .B(n24760), .C(
        n24759), .Y(n24768) );
  OR2x2_ASAP7_75t_SL U38151 ( .A(n32171), .B(n24765), .Y(n32168) );
  O2A1O1Ixp5_ASAP7_75t_SL U38152 ( .A1(n31857), .A2(n26817), .B(n24772), .C(
        n26818), .Y(n24775) );
  NAND3xp33_ASAP7_75t_SL U38153 ( .A(n24773), .B(
        u0_0_leon3x0_p0_iu_v_A__CWP__0_), .C(n26777), .Y(n24774) );
  XNOR2xp5_ASAP7_75t_SL U38154 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__4_), .B(
        n32183), .Y(n24803) );
  OAI31xp33_ASAP7_75t_SL U38155 ( .A1(n31857), .A2(
        u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__0_), .A3(n26815), .B(n30907), .Y(
        n24791) );
  XNOR2xp5_ASAP7_75t_SL U38156 ( .A(n26829), .B(n30939), .Y(n24793) );
  XNOR2xp5_ASAP7_75t_SL U38157 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__7_), .B(
        n32186), .Y(n24792) );
  XNOR2xp5_ASAP7_75t_SL U38158 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__3_), .B(
        n32179), .Y(n24800) );
  XNOR2xp5_ASAP7_75t_SL U38159 ( .A(u0_0_leon3x0_p0_iu_v_M__CTRL__RD__2_), .B(
        n32178), .Y(n24799) );
  NAND4xp25_ASAP7_75t_SL U38160 ( .A(n24800), .B(n24798), .C(n24799), .D(
        n24797), .Y(n24801) );
  NOR3xp33_ASAP7_75t_SL U38161 ( .A(n24803), .B(n24802), .C(n24801), .Y(n24804) );
  A2O1A1Ixp33_ASAP7_75t_SL U38162 ( .A1(n24806), .A2(n26842), .B(n24805), .C(
        n24804), .Y(n24813) );
  NOR3xp33_ASAP7_75t_SL U38163 ( .A(n24808), .B(n24807), .C(n26778), .Y(n24811) );
  O2A1O1Ixp5_ASAP7_75t_SL U38164 ( .A1(n32173), .A2(n30810), .B(n24815), .C(
        n24814), .Y(n24868) );
  OR2x2_ASAP7_75t_SL U38165 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__1_), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__CNT__0_), .Y(n32084) );
  OAI211xp5_ASAP7_75t_SL U38166 ( .A1(DP_OP_1196_128_7433_n455), .A2(n24818), 
        .B(n24817), .C(n24833), .Y(n24822) );
  XNOR2xp5_ASAP7_75t_SL U38167 ( .A(n24819), .B(DP_OP_1196_128_7433_n454), .Y(
        n24821) );
  XNOR2xp5_ASAP7_75t_SL U38168 ( .A(n26819), .B(DP_OP_1196_128_7433_n452), .Y(
        n24820) );
  NOR3xp33_ASAP7_75t_SL U38169 ( .A(n24822), .B(n24821), .C(n24820), .Y(n24823) );
  A2O1A1Ixp33_ASAP7_75t_SL U38170 ( .A1(n32171), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__7_), .B(n24824), .C(n24823), .Y(
        n24825) );
  O2A1O1Ixp5_ASAP7_75t_SL U38171 ( .A1(n32164), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__4_), .B(n24826), .C(n24825), .Y(
        n24827) );
  A2O1A1Ixp33_ASAP7_75t_SL U38172 ( .A1(n26853), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__5_), .B(n24828), .C(n24827), .Y(
        n24831) );
  XNOR2xp5_ASAP7_75t_SL U38173 ( .A(n24829), .B(n32170), .Y(n24830) );
  XNOR2xp5_ASAP7_75t_SL U38174 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__RD__4_), .B(
        n32183), .Y(n24839) );
  NAND4xp25_ASAP7_75t_SL U38175 ( .A(n24834), .B(n24835), .C(n24836), .D(
        n24833), .Y(n24837) );
  NOR3xp33_ASAP7_75t_SL U38176 ( .A(n24839), .B(n24838), .C(n24837), .Y(n24840) );
  A2O1A1Ixp33_ASAP7_75t_SL U38177 ( .A1(n18870), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__RD__5_), .B(n24841), .C(n24840), .Y(
        n24843) );
  NAND3xp33_ASAP7_75t_SL U38178 ( .A(n26190), .B(n24856), .C(n32102), .Y(
        n25232) );
  NAND3xp33_ASAP7_75t_SL U38179 ( .A(n31858), .B(n18819), .C(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), .Y(n31384) );
  OR2x2_ASAP7_75t_SL U38180 ( .A(n32087), .B(n31384), .Y(n32081) );
  OR2x2_ASAP7_75t_SL U38181 ( .A(n18842), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .Y(n24852) );
  NAND3xp33_ASAP7_75t_SL U38182 ( .A(n24846), .B(n24998), .C(n24852), .Y(
        n29206) );
  O2A1O1Ixp5_ASAP7_75t_SL U38183 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__WY_), 
        .A2(u0_0_leon3x0_p0_iu_v_M__CTRL__WY_), .B(n32050), .C(n24848), .Y(
        n24849) );
  A2O1A1Ixp33_ASAP7_75t_SL U38184 ( .A1(n24851), .A2(n24850), .B(n25232), .C(
        n24849), .Y(n24862) );
  NAND4xp25_ASAP7_75t_SL U38185 ( .A(n32048), .B(n24998), .C(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__20_), .D(n24853), .Y(n32057) );
  NAND4xp25_ASAP7_75t_SL U38186 ( .A(n32055), .B(n25221), .C(n24855), .D(
        n32083), .Y(n24857) );
  O2A1O1Ixp5_ASAP7_75t_SL U38187 ( .A1(n31381), .A2(n32057), .B(n24857), .C(
        n24874), .Y(n24861) );
  NOR3xp33_ASAP7_75t_SL U38188 ( .A(n24862), .B(n24861), .C(n24860), .Y(n24863) );
  A2O1A1Ixp33_ASAP7_75t_SL U38189 ( .A1(n24866), .A2(n24865), .B(n24864), .C(
        n24863), .Y(n24867) );
  OR2x2_ASAP7_75t_SL U38190 ( .A(n24659), .B(n31809), .Y(n32104) );
  NAND3xp33_ASAP7_75t_SL U38191 ( .A(n26190), .B(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_), .C(n30502), .Y(n24894) );
  NAND3xp33_ASAP7_75t_SL U38192 ( .A(n31817), .B(n24911), .C(n24883), .Y(
        n24887) );
  OR2x2_ASAP7_75t_SL U38193 ( .A(n24884), .B(n24900), .Y(n24903) );
  A2O1A1Ixp33_ASAP7_75t_SL U38194 ( .A1(n32102), .A2(n24895), .B(n24894), .C(
        n25219), .Y(n31816) );
  OR2x2_ASAP7_75t_SL U38195 ( .A(n18800), .B(u0_0_leon3x0_p0_c0mmu_a0_r_BO__0_), .Y(n25568) );
  OR2x2_ASAP7_75t_SL U38196 ( .A(n22380), .B(n22422), .Y(n24907) );
  NAND3xp33_ASAP7_75t_SL U38197 ( .A(n25214), .B(n24911), .C(n31651), .Y(
        n24914) );
  OA21x2_ASAP7_75t_SL U38198 ( .A1(n24916), .A2(n31816), .B(n24915), .Y(n4336)
         );
  NAND4xp25_ASAP7_75t_SL U38199 ( .A(n24919), .B(n24918), .C(n24931), .D(
        n24940), .Y(n25077) );
  O2A1O1Ixp5_ASAP7_75t_SL U38200 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__19_), .A2(n25649), .B(n25659), .C(n24939), .Y(n24986) );
  A2O1A1Ixp33_ASAP7_75t_SL U38201 ( .A1(n24943), .A2(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), .B(n25652), .C(n25653), .Y(
        n24946) );
  AO21x1_ASAP7_75t_SL U38202 ( .A1(n24983), .A2(n24987), .B(n25668), .Y(n31945) );
  NAND3xp33_ASAP7_75t_SL U38203 ( .A(n30663), .B(n32016), .C(n22919), .Y(
        n27020) );
  NAND3xp33_ASAP7_75t_SL U38204 ( .A(n24961), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__21_), .C(n25675), .Y(n24962) );
  NAND4xp25_ASAP7_75t_SL U38205 ( .A(n32015), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__20_), .C(n32012), .D(n25172), .Y(
        n24970) );
  A2O1A1Ixp33_ASAP7_75t_SL U38206 ( .A1(n24976), .A2(n24975), .B(n25245), .C(
        n31697), .Y(n31626) );
  OR2x2_ASAP7_75t_SL U38207 ( .A(n18801), .B(n32035), .Y(n10988) );
  OA21x2_ASAP7_75t_SL U38208 ( .A1(n31971), .A2(n32719), .B(n24980), .Y(n32998) );
  OR2x2_ASAP7_75t_SL U38209 ( .A(n24659), .B(n31872), .Y(n25007) );
  A2O1A1Ixp33_ASAP7_75t_SL U38210 ( .A1(n24995), .A2(n24994), .B(n24993), .C(
        n24992), .Y(n31946) );
  A2O1A1Ixp33_ASAP7_75t_SL U38211 ( .A1(n25602), .A2(n25000), .B(n24680), .C(
        n25001), .Y(n3164) );
  A2O1A1Ixp33_ASAP7_75t_SL U38212 ( .A1(u0_0_leon3x0_p0_iu_r_A__JMPL_), .A2(
        n31807), .B(n24680), .C(n25002), .Y(n3162) );
  AND2x2_ASAP7_75t_SL U38213 ( .A(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__29_), 
        .B(n32091), .Y(n25004) );
  AND2x2_ASAP7_75t_SL U38214 ( .A(n22379), .B(n32101), .Y(n26810) );
  OR2x2_ASAP7_75t_SL U38215 ( .A(n25006), .B(n25399), .Y(n13499) );
  OR2x2_ASAP7_75t_SL U38216 ( .A(n25238), .B(n17284), .Y(n17278) );
  A2O1A1Ixp33_ASAP7_75t_SL U38217 ( .A1(u0_0_leon3x0_p0_c0mmu_dcache0_r_READ_), 
        .A2(u0_0_leon3x0_p0_ico_DIAGRDY_), .B(n25008), .C(n31582), .Y(n25016)
         );
  XOR2xp5_ASAP7_75t_SL U38218 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__4_), .B(
        n3133), .Y(n25010) );
  XOR2xp5_ASAP7_75t_SL U38219 ( .A(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__3_), .B(
        n2962), .Y(n25009) );
  NAND3xp33_ASAP7_75t_SL U38220 ( .A(n25010), .B(n25009), .C(n31303), .Y(
        n25012) );
  OR3x1_ASAP7_75t_SL U38221 ( .A(n31303), .B(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_NOMDS_), .C(n32253), .Y(n25011) );
  O2A1O1Ixp5_ASAP7_75t_SL U38222 ( .A1(n2963), .A2(n25012), .B(n25011), .C(
        n3067), .Y(n31450) );
  O2A1O1Ixp5_ASAP7_75t_SL U38223 ( .A1(n25013), .A2(n25012), .B(n25011), .C(
        n32437), .Y(n31449) );
  OR2x2_ASAP7_75t_SL U38224 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__LD_), .B(n30017), .Y(n31474) );
  OR2x2_ASAP7_75t_SL U38225 ( .A(n31259), .B(n31582), .Y(n25044) );
  AND2x2_ASAP7_75t_SL U38226 ( .A(n13499), .B(n25020), .Y(n25026) );
  AOI222xp33_ASAP7_75t_SL U38227 ( .A1(n29999), .A2(ahbso_0__HRDATA__31_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__31_), .C1(n24574), .C2(
        ahb0_r_HRDATAS__31_), .Y(n32430) );
  NAND3xp33_ASAP7_75t_SL U38228 ( .A(n31259), .B(n32602), .C(n32604), .Y(
        n31466) );
  AOI222xp33_ASAP7_75t_SL U38229 ( .A1(n29999), .A2(ahbso_0__HRDATA__15_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__15_), .C1(n30000), .C2(
        ahb0_r_HRDATAS__15_), .Y(n31032) );
  A2O1A1Ixp33_ASAP7_75t_SL U38230 ( .A1(n24471), .A2(n25047), .B(n30207), .C(
        n25046), .Y(n31034) );
  A2O1A1Ixp33_ASAP7_75t_SL U38231 ( .A1(n30017), .A2(
        u0_0_leon3x0_p0_iu_r_X__DCI__SIGNED_), .B(n25051), .C(n25439), .Y(
        n25052) );
  OR2x2_ASAP7_75t_SL U38232 ( .A(n31364), .B(n25052), .Y(n25069) );
  AOI222xp33_ASAP7_75t_SL U38233 ( .A1(n29999), .A2(ahbso_0__HRDATA__7_), .B1(
        n30002), .B2(ahbso_1__HRDATA__7_), .C1(n30000), .C2(ahb0_r_HRDATAS__7_), .Y(n30876) );
  NAND3xp33_ASAP7_75t_SL U38234 ( .A(n25063), .B(n25062), .C(n25061), .Y(
        n29919) );
  NAND3xp33_ASAP7_75t_SL U38235 ( .A(n25067), .B(n25440), .C(n29919), .Y(
        n25064) );
  A2O1A1Ixp33_ASAP7_75t_SL U38236 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__LD_), 
        .A2(n31398), .B(n24524), .C(n25076), .Y(n3314) );
  OR2x2_ASAP7_75t_SL U38237 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL1__2_), .B(
        u0_0_leon3x0_p0_iu_r_A__RSEL1__1_), .Y(n25208) );
  XOR2xp5_ASAP7_75t_SL U38238 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__1_), .B(
        u0_0_leon3x0_p0_iu_r_E__INVOP2_), .Y(n25081) );
  AND2x2_ASAP7_75t_SL U38239 ( .A(n22224), .B(n26351), .Y(n28968) );
  XOR2xp5_ASAP7_75t_SL U38240 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__4_), .B(
        u0_0_leon3x0_p0_iu_r_E__INVOP2_), .Y(n25088) );
  XOR2xp5_ASAP7_75t_SL U38241 ( .A(u0_0_leon3x0_p0_iu_r_X__DATA__0__0_), .B(
        u0_0_leon3x0_p0_iu_r_E__INVOP2_), .Y(n25121) );
  OR2x2_ASAP7_75t_SL U38242 ( .A(n25122), .B(n28992), .Y(n30635) );
  A2O1A1Ixp33_ASAP7_75t_SL U38243 ( .A1(u0_0_leon3x0_p0_iu_r_E__ALUOP__2_), 
        .A2(u0_0_leon3x0_p0_iu_r_E__ALUOP__1_), .B(n25488), .C(n26482), .Y(
        n25127) );
  A2O1A1Ixp33_ASAP7_75t_SL U38244 ( .A1(n25136), .A2(n25135), .B(n24480), .C(
        n25134), .Y(n31416) );
  OR2x2_ASAP7_75t_SL U38245 ( .A(n28968), .B(n29609), .Y(n27208) );
  NAND3xp33_ASAP7_75t_SL U38246 ( .A(n25174), .B(n30664), .C(n25173), .Y(
        n26269) );
  OR2x2_ASAP7_75t_SL U38247 ( .A(u0_0_leon3x0_p0_iu_v_X__CTRL__WY_), .B(n28734), .Y(n28934) );
  OR2x2_ASAP7_75t_SL U38248 ( .A(u0_0_leon3x0_p0_iu_r_E__JMPL_), .B(n27067), 
        .Y(n28888) );
  OAI211xp5_ASAP7_75t_SL U38249 ( .A1(n31678), .A2(n29594), .B(n29591), .C(
        n25179), .Y(n25180) );
  NAND3xp33_ASAP7_75t_SL U38250 ( .A(n25184), .B(n25183), .C(n25182), .Y(
        n25185) );
  OAI211xp5_ASAP7_75t_SL U38251 ( .A1(n29608), .A2(n30635), .B(n25205), .C(
        n25204), .Y(n25206) );
  A2O1A1Ixp33_ASAP7_75t_SL U38252 ( .A1(n31681), .A2(n31398), .B(n25212), .C(
        n22379), .Y(n25213) );
  NAND3xp33_ASAP7_75t_SL U38253 ( .A(n31657), .B(n25220), .C(n32084), .Y(
        n32099) );
  A2O1A1Ixp33_ASAP7_75t_SL U38254 ( .A1(n32099), .A2(n25228), .B(n32083), .C(
        n25227), .Y(n25229) );
  NAND3xp33_ASAP7_75t_SL U38255 ( .A(n25241), .B(n25240), .C(n31949), .Y(
        n30802) );
  OR2x2_ASAP7_75t_SL U38256 ( .A(n17271), .B(n17270), .Y(n25413) );
  A2O1A1Ixp33_ASAP7_75t_SL U38257 ( .A1(n24494), .A2(n25246), .B(n25245), .C(
        n31697), .Y(n31706) );
  NAND3xp33_ASAP7_75t_SL U38258 ( .A(n25260), .B(n25259), .C(n25258), .Y(
        n32002) );
  OA21x2_ASAP7_75t_SL U38259 ( .A1(n31948), .A2(n32719), .B(n25265), .Y(n32992) );
  OA21x2_ASAP7_75t_SL U38260 ( .A1(n30737), .A2(n32719), .B(n25267), .Y(n32996) );
  OA21x2_ASAP7_75t_SL U38261 ( .A1(n31056), .A2(n32719), .B(n25269), .Y(n33000) );
  OA21x2_ASAP7_75t_SL U38262 ( .A1(n30973), .A2(n32719), .B(n25270), .Y(n33002) );
  XNOR2xp5_ASAP7_75t_SL U38263 ( .A(n3133), .B(n25330), .Y(n32986) );
  A2O1A1Ixp33_ASAP7_75t_SL U38264 ( .A1(n31877), .A2(n32496), .B(n31700), .C(
        n25325), .Y(n32988) );
  AO21x1_ASAP7_75t_SL U38265 ( .A1(n2963), .A2(n31697), .B(n25331), .Y(n25328)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U38266 ( .A1(n31877), .A2(n32467), .B(n31700), .C(
        n25333), .Y(n25327) );
  OR2x2_ASAP7_75t_SL U38267 ( .A(n31848), .B(n1637), .Y(n27460) );
  OR2x2_ASAP7_75t_SL U38268 ( .A(n26658), .B(n27460), .Y(n4536) );
  NOR3xp33_ASAP7_75t_SL U38269 ( .A(n31963), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__INST__21_), .C(n31961), .Y(n25339) );
  OR2x2_ASAP7_75t_SL U38270 ( .A(n25339), .B(
        u0_0_leon3x0_p0_iu_ex_jump_address_2_), .Y(n32438) );
  NAND3xp33_ASAP7_75t_SL U38271 ( .A(n25344), .B(n25345), .C(n25346), .Y(
        n25347) );
  NOR3xp33_ASAP7_75t_SL U38272 ( .A(n25347), .B(u0_0_leon3x0_p0_dci[23]), .C(
        u0_0_leon3x0_p0_dci[17]), .Y(n25348) );
  NAND3xp33_ASAP7_75t_SL U38273 ( .A(n25350), .B(n25349), .C(n25348), .Y(
        n25351) );
  A2O1A1Ixp33_ASAP7_75t_SL U38274 ( .A1(n29884), .A2(
        u0_0_leon3x0_p0_iu_de_icc_1_), .B(n25365), .C(n30687), .Y(n25369) );
  NAND3xp33_ASAP7_75t_SL U38275 ( .A(n29708), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__22_), .C(
        u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_), .Y(n29704) );
  A2O1A1Ixp33_ASAP7_75t_SL U38276 ( .A1(irqi_0__IRL__0_), .A2(n30700), .B(
        n25372), .C(n25371), .Y(n25373) );
  O2A1O1Ixp5_ASAP7_75t_SL U38277 ( .A1(n3328), .A2(n25375), .B(n29645), .C(
        n25374), .Y(n25378) );
  OAI211xp5_ASAP7_75t_SL U38278 ( .A1(n3327), .A2(n29882), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__PV_), .C(u0_0_leon3x0_p0_iu_r_W__S__ET_), 
        .Y(n25376) );
  OR2x2_ASAP7_75t_SL U38279 ( .A(u0_0_leon3x0_p0_c0mmu_mmudci[0]), .B(
        u0_0_leon3x0_p0_c0mmu_mmudci[1]), .Y(n29716) );
  A2O1A1Ixp33_ASAP7_75t_SL U38280 ( .A1(n29706), .A2(n25382), .B(n25381), .C(
        n29705), .Y(n25383) );
  A2O1A1Ixp33_ASAP7_75t_SL U38281 ( .A1(n25385), .A2(n25384), .B(n29717), .C(
        n29716), .Y(n25386) );
  OR3x1_ASAP7_75t_SL U38282 ( .A(n25396), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__0_), .C(
        u0_0_leon3x0_p0_iu_v_X__CTRL__CNT__1_), .Y(n29707) );
  O2A1O1Ixp5_ASAP7_75t_SL U38283 ( .A1(n29715), .A2(n25387), .B(n25386), .C(
        n29707), .Y(n29675) );
  OR2x2_ASAP7_75t_SL U38284 ( .A(n3730), .B(n3704), .Y(n32074) );
  OR2x2_ASAP7_75t_SL U38285 ( .A(n31264), .B(n32030), .Y(n25516) );
  AOI222xp33_ASAP7_75t_SL U38286 ( .A1(n29999), .A2(ahbso_0__HRDATA__9_), .B1(
        n30002), .B2(ahbso_1__HRDATA__9_), .C1(n24574), .C2(ahb0_r_HRDATAS__9_), .Y(n30155) );
  AND2x2_ASAP7_75t_SL U38287 ( .A(n4746), .B(n33063), .Y(n33066) );
  AOI222xp33_ASAP7_75t_SL U38288 ( .A1(n29999), .A2(ahbso_0__HRDATA__29_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__29_), .C1(n30000), .C2(
        ahb0_r_HRDATAS__29_), .Y(n32410) );
  NAND3xp33_ASAP7_75t_SL U38289 ( .A(n25416), .B(n25415), .C(n25414), .Y(
        n30024) );
  NAND3xp33_ASAP7_75t_SL U38290 ( .A(n25432), .B(n25426), .C(n25425), .Y(
        n32336) );
  AND2x2_ASAP7_75t_SL U38291 ( .A(n25433), .B(n25432), .Y(n32405) );
  NAND3xp33_ASAP7_75t_SL U38292 ( .A(n25444), .B(n25443), .C(n25442), .Y(
        n31477) );
  NAND4xp25_ASAP7_75t_SL U38293 ( .A(n26755), .B(n29212), .C(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__19_), .D(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__20_), .Y(n25452) );
  OR2x2_ASAP7_75t_SL U38294 ( .A(n22380), .B(n26354), .Y(n25559) );
  A2O1A1Ixp33_ASAP7_75t_SL U38295 ( .A1(n25882), .A2(
        u0_0_leon3x0_p0_iu_r_A__BP_), .B(n22378), .C(n25454), .Y(n3294) );
  NAND3xp33_ASAP7_75t_SL U38296 ( .A(n25458), .B(n25785), .C(n25457), .Y(
        n26555) );
  NAND3xp33_ASAP7_75t_SL U38297 ( .A(n25462), .B(n25785), .C(n25461), .Y(
        n26376) );
  NAND3xp33_ASAP7_75t_SL U38298 ( .A(n25466), .B(n25785), .C(n25465), .Y(
        n26425) );
  NAND3xp33_ASAP7_75t_SL U38299 ( .A(n25479), .B(n25785), .C(n25478), .Y(
        n25790) );
  OAI211xp5_ASAP7_75t_SL U38300 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__26_), 
        .A2(n28637), .B(n25485), .C(n25484), .Y(n25486) );
  A2O1A1Ixp33_ASAP7_75t_SL U38301 ( .A1(u0_0_leon3x0_p0_divi[25]), .A2(n26358), 
        .B(n25489), .C(n22472), .Y(n25490) );
  A2O1A1Ixp33_ASAP7_75t_SL U38302 ( .A1(u0_0_leon3x0_p0_divi[25]), .A2(n28830), 
        .B(n22472), .C(n25490), .Y(n25492) );
  A2O1A1Ixp33_ASAP7_75t_SL U38303 ( .A1(u0_0_leon3x0_p0_divi[25]), .A2(n24580), 
        .B(n25493), .C(n25492), .Y(n30246) );
  AO21x1_ASAP7_75t_SL U38304 ( .A1(n30614), .A2(n30244), .B(n25498), .Y(n25499) );
  NAND4xp25_ASAP7_75t_SL U38305 ( .A(n25503), .B(n25502), .C(n25501), .D(
        n25500), .Y(n25504) );
  OAI211xp5_ASAP7_75t_SL U38306 ( .A1(n27208), .A2(n25915), .B(n25506), .C(
        n25505), .Y(n25507) );
  A2O1A1Ixp33_ASAP7_75t_SL U38307 ( .A1(u0_0_leon3x0_p0_dci[31]), .A2(n22398), 
        .B(n25507), .C(n30007), .Y(n25508) );
  OR2x2_ASAP7_75t_SL U38308 ( .A(n31455), .B(n31306), .Y(n25521) );
  O2A1O1Ixp5_ASAP7_75t_SL U38309 ( .A1(n25512), .A2(n25511), .B(n32198), .C(
        n31605), .Y(n25514) );
  OR2x2_ASAP7_75t_SL U38310 ( .A(n25518), .B(n25517), .Y(n31609) );
  OR2x2_ASAP7_75t_SL U38311 ( .A(ahb0_r_HMASTERD_), .B(n25597), .Y(n32888) );
  NAND3xp33_ASAP7_75t_SL U38312 ( .A(n31252), .B(n2992), .C(n31529), .Y(n25534) );
  NAND3xp33_ASAP7_75t_SL U38313 ( .A(n25527), .B(n25526), .C(n25525), .Y(
        n25532) );
  NAND3xp33_ASAP7_75t_SL U38314 ( .A(n25530), .B(n25529), .C(n25528), .Y(
        n25531) );
  OR2x2_ASAP7_75t_SL U38315 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__26_), .B(
        n26354), .Y(n25556) );
  NOR3xp33_ASAP7_75t_SL U38316 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__28_), 
        .B(u0_0_leon3x0_p0_iu_r_X__CTRL__INST__27_), .C(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__20_), .Y(n25554) );
  NOR3xp33_ASAP7_75t_SL U38317 ( .A(u0_0_dbgo_OPTYPE__0_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__19_), .C(u0_0_dbgo_OPTYPE__1_), 
        .Y(n29178) );
  OR2x2_ASAP7_75t_SL U38318 ( .A(n25555), .B(n26758), .Y(n25557) );
  AOI222xp33_ASAP7_75t_SL U38319 ( .A1(n29999), .A2(ahbso_0__HRDATA__8_), .B1(
        n30002), .B2(ahbso_1__HRDATA__8_), .C1(n30000), .C2(ahb0_r_HRDATAS__8_), .Y(n32322) );
  OR2x2_ASAP7_75t_SL U38320 ( .A(u0_0_leon3x0_p0_dci[41]), .B(n25575), .Y(
        n30195) );
  AO21x1_ASAP7_75t_SL U38321 ( .A1(n30161), .A2(u0_0_leon3x0_p0_dci[37]), .B(
        n25576), .Y(n30194) );
  O2A1O1Ixp5_ASAP7_75t_SL U38322 ( .A1(n25578), .A2(n30194), .B(
        u0_0_leon3x0_p0_dci[38]), .C(n25577), .Y(n25579) );
  NAND3xp33_ASAP7_75t_SL U38323 ( .A(n31575), .B(n31574), .C(
        u0_0_leon3x0_p0_dci[2]), .Y(n31589) );
  NAND3xp33_ASAP7_75t_SL U38324 ( .A(u0_0_leon3x0_p0_c0mmu_dcache0_r_READ_), 
        .B(u0_0_leon3x0_p0_c0mmu_dcache0_r_DSTATE__0_), .C(n25592), .Y(n25589)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U38325 ( .A1(n31613), .A2(n31589), .B(n25590), .C(
        n25589), .Y(n25596) );
  A2O1A1Ixp33_ASAP7_75t_SL U38326 ( .A1(n32272), .A2(n31572), .B(n25593), .C(
        u0_0_leon3x0_p0_c0mmu_mcdi[0]), .Y(n25594) );
  A2O1A1Ixp33_ASAP7_75t_SL U38327 ( .A1(n30418), .A2(n29212), .B(n29214), .C(
        n25609), .Y(n29695) );
  AOI222xp33_ASAP7_75t_SL U38328 ( .A1(n29999), .A2(ahbso_0__HRDATA__14_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__14_), .C1(n24574), .C2(
        ahb0_r_HRDATAS__14_), .Y(n30557) );
  AOI222xp33_ASAP7_75t_SL U38329 ( .A1(n29999), .A2(ahbso_0__HRDATA__30_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__30_), .C1(n30000), .C2(
        ahb0_r_HRDATAS__30_), .Y(n32419) );
  NAND3xp33_ASAP7_75t_SL U38330 ( .A(n25618), .B(n25617), .C(n25616), .Y(
        n25619) );
  OAI211xp5_ASAP7_75t_SL U38331 ( .A1(u0_0_leon3x0_p0_iu_r_E__ALUOP__0_), .A2(
        n28488), .B(n29587), .C(n29504), .Y(n25645) );
  A2O1A1Ixp33_ASAP7_75t_SL U38332 ( .A1(n27215), .A2(n30007), .B(n25630), .C(
        n25629), .Y(n32342) );
  NAND4xp25_ASAP7_75t_SL U38333 ( .A(n31325), .B(n2992), .C(n25952), .D(n25951), .Y(n25638) );
  A2O1A1Ixp33_ASAP7_75t_SL U38334 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_), .A2(n25649), .B(n25705), .C(
        n25648), .Y(n29874) );
  OR2x2_ASAP7_75t_SL U38335 ( .A(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__31_), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__30_), .Y(n25665) );
  NAND4xp25_ASAP7_75t_SL U38336 ( .A(n25653), .B(n25652), .C(n31537), .D(
        n31943), .Y(n25654) );
  NAND3xp33_ASAP7_75t_SL U38337 ( .A(n29874), .B(n29700), .C(n29872), .Y(
        n29223) );
  AO21x1_ASAP7_75t_SL U38338 ( .A1(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__23_), 
        .A2(u0_0_leon3x0_p0_iu_v_E__CTRL__INST__13_), .B(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__24_), .Y(n25660) );
  A2O1A1Ixp33_ASAP7_75t_SL U38339 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__20_), .A2(n25661), .B(n25675), .C(
        n25660), .Y(n25662) );
  OAI211xp5_ASAP7_75t_SL U38340 ( .A1(n25664), .A2(n25676), .B(n25663), .C(
        n25662), .Y(n25674) );
  A2O1A1Ixp33_ASAP7_75t_SL U38341 ( .A1(n25706), .A2(n25705), .B(n25704), .C(
        n29219), .Y(n29230) );
  NAND3xp33_ASAP7_75t_SL U38342 ( .A(n26230), .B(n25713), .C(n25712), .Y(
        n32211) );
  NAND3xp33_ASAP7_75t_SL U38343 ( .A(n25717), .B(n25716), .C(n25715), .Y(
        n31005) );
  NAND3xp33_ASAP7_75t_SL U38344 ( .A(n29737), .B(n24684), .C(n30685), .Y(
        n25723) );
  NOR3xp33_ASAP7_75t_SL U38345 ( .A(n25723), .B(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PV_), .C(n25722), .Y(n25724) );
  OR2x2_ASAP7_75t_SL U38346 ( .A(u0_0_leon3x0_p0_iu_r_X__NPC__1_), .B(
        u0_0_leon3x0_p0_iu_r_X__NPC__0_), .Y(n25732) );
  AND2x2_ASAP7_75t_SL U38347 ( .A(n32077), .B(n32153), .Y(n32162) );
  AND2x2_ASAP7_75t_SL U38348 ( .A(u0_0_leon3x0_p0_iu_r_X__NPC__2_), .B(n33054), 
        .Y(n30724) );
  NAND3xp33_ASAP7_75t_SL U38349 ( .A(n25741), .B(n25740), .C(n25739), .Y(
        rf_di_w[18]) );
  NAND3xp33_ASAP7_75t_SL U38350 ( .A(n25744), .B(n25743), .C(n25742), .Y(
        n30885) );
  NAND3xp33_ASAP7_75t_SL U38351 ( .A(n25756), .B(n25755), .C(n25754), .Y(
        rf_di_w[19]) );
  NAND3xp33_ASAP7_75t_SL U38352 ( .A(n25758), .B(n25785), .C(n25757), .Y(
        n27097) );
  NAND3xp33_ASAP7_75t_SL U38353 ( .A(n25762), .B(n25761), .C(n25760), .Y(
        n26709) );
  OAI211xp5_ASAP7_75t_SL U38354 ( .A1(n25771), .A2(n26675), .B(n25770), .C(
        n25769), .Y(n25781) );
  OA21x2_ASAP7_75t_SL U38355 ( .A1(n28769), .A2(n18327), .B(n25772), .Y(
        u0_0_leon3x0_p0_divi[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38356 ( .A1(u0_0_leon3x0_p0_divi[18]), .A2(n28827), 
        .B(n25774), .C(n23936), .Y(n25777) );
  O2A1O1Ixp5_ASAP7_75t_SL U38357 ( .A1(n23935), .A2(n25778), .B(n25777), .C(
        n25776), .Y(n30304) );
  NAND3xp33_ASAP7_75t_SL U38358 ( .A(n25786), .B(n25785), .C(n25784), .Y(
        n27092) );
  OAI211xp5_ASAP7_75t_SL U38359 ( .A1(n26380), .A2(n28850), .B(n25789), .C(
        n25788), .Y(n26986) );
  AND2x2_ASAP7_75t_SL U38360 ( .A(n30007), .B(n29603), .Y(n28924) );
  A2O1A1Ixp33_ASAP7_75t_SL U38361 ( .A1(n25805), .A2(n25804), .B(n25803), .C(
        n25802), .Y(n30820) );
  OAI211xp5_ASAP7_75t_SL U38362 ( .A1(n31340), .A2(n30821), .B(n25807), .C(
        n25806), .Y(n25808) );
  AO21x1_ASAP7_75t_SL U38363 ( .A1(n31342), .A2(n30820), .B(n25808), .Y(n27035) );
  AO21x1_ASAP7_75t_SL U38364 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__6_), .A2(
        n28480), .B(n25814), .Y(n25818) );
  OA21x2_ASAP7_75t_SL U38365 ( .A1(n28769), .A2(u0_0_leon3x0_p0_muli[26]), .B(
        n25821), .Y(u0_0_leon3x0_p0_divi[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38366 ( .A1(u0_0_leon3x0_p0_divi[17]), .A2(n28827), 
        .B(n25823), .C(n25828), .Y(n25826) );
  O2A1O1Ixp5_ASAP7_75t_SL U38367 ( .A1(n25828), .A2(n25827), .B(n25826), .C(
        n25825), .Y(n30307) );
  OAI211xp5_ASAP7_75t_SL U38368 ( .A1(n30625), .A2(n30307), .B(n25830), .C(
        n25829), .Y(n25831) );
  OAI211xp5_ASAP7_75t_SL U38369 ( .A1(n25836), .A2(n30628), .B(n25835), .C(
        n25834), .Y(n25837) );
  A2O1A1Ixp33_ASAP7_75t_SL U38370 ( .A1(n22375), .A2(n25841), .B(n25839), .C(
        n25838), .Y(n28546) );
  OR2x2_ASAP7_75t_SL U38371 ( .A(n25850), .B(n30134), .Y(n29516) );
  AND2x2_ASAP7_75t_SL U38372 ( .A(n29563), .B(n29584), .Y(n25860) );
  OR2x2_ASAP7_75t_SL U38373 ( .A(n28879), .B(n22375), .Y(n30008) );
  O2A1O1Ixp5_ASAP7_75t_SL U38374 ( .A1(n25860), .A2(n25859), .B(n29937), .C(
        n25858), .Y(n25861) );
  A2O1A1Ixp33_ASAP7_75t_SL U38375 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[10]), .B(n25863), .C(n31638), .Y(n4711) );
  AOI222xp33_ASAP7_75t_SL U38376 ( .A1(n29999), .A2(ahbso_0__HRDATA__4_), .B1(
        n30002), .B2(ahbso_1__HRDATA__4_), .C1(n30000), .C2(ahb0_r_HRDATAS__4_), .Y(n32308) );
  O2A1O1Ixp5_ASAP7_75t_SL U38377 ( .A1(n25874), .A2(n25873), .B(n29937), .C(
        n25872), .Y(n25875) );
  A2O1A1Ixp33_ASAP7_75t_SL U38378 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[8]), .B(n25877), .C(n31638), .Y(n4765) );
  OAI31xp33_ASAP7_75t_SL U38379 ( .A1(n29000), .A2(n28931), .A3(n25894), .B(
        n31812), .Y(n29589) );
  OAI211xp5_ASAP7_75t_SL U38380 ( .A1(n25896), .A2(n29592), .B(n29591), .C(
        n25895), .Y(n25899) );
  A2O1A1Ixp33_ASAP7_75t_SL U38381 ( .A1(n26597), .A2(n25901), .B(n25900), .C(
        n24634), .Y(n25902) );
  NAND3xp33_ASAP7_75t_SL U38382 ( .A(n25904), .B(n25903), .C(n25902), .Y(
        n25905) );
  OAI211xp5_ASAP7_75t_SL U38383 ( .A1(n25915), .A2(n28502), .B(n25914), .C(
        n25913), .Y(n25916) );
  A2O1A1Ixp33_ASAP7_75t_SL U38384 ( .A1(u0_0_leon3x0_p0_dci[34]), .A2(n22398), 
        .B(n25916), .C(n30007), .Y(n25917) );
  NAND3xp33_ASAP7_75t_SL U38385 ( .A(n25919), .B(
        u0_0_leon3x0_p0_iu_r_A__DIVSTART_), .C(n32066), .Y(n28293) );
  NAND3xp33_ASAP7_75t_SL U38386 ( .A(n25922), .B(n25921), .C(n25920), .Y(
        n25931) );
  NOR3xp33_ASAP7_75t_SL U38387 ( .A(u0_0_leon3x0_p0_div0_addout_16_), .B(
        u0_0_leon3x0_p0_div0_addout_9_), .C(u0_0_leon3x0_p0_div0_addout_10_), 
        .Y(n25929) );
  NAND3xp33_ASAP7_75t_SL U38388 ( .A(n25925), .B(n25924), .C(n25923), .Y(
        n25926) );
  NAND3xp33_ASAP7_75t_SL U38389 ( .A(n25929), .B(n25928), .C(n25927), .Y(
        n25930) );
  AO21x1_ASAP7_75t_SL U38390 ( .A1(n23229), .A2(n28377), .B(n25936), .Y(n4313)
         );
  NAND4xp25_ASAP7_75t_SL U38391 ( .A(n26097), .B(n25940), .C(n27476), .D(
        n25952), .Y(n25942) );
  NAND3xp33_ASAP7_75t_SL U38392 ( .A(n31325), .B(n27290), .C(n25952), .Y(
        n25953) );
  AO21x1_ASAP7_75t_SL U38393 ( .A1(n27290), .A2(n30894), .B(n27291), .Y(n25960) );
  OR2x2_ASAP7_75t_SL U38394 ( .A(irqo[1]), .B(n3325), .Y(n29329) );
  A2O1A1Ixp33_ASAP7_75t_SL U38395 ( .A1(n25960), .A2(irqctrl0_r_IFORCE__0__11_), .B(n25959), .C(n25958), .Y(n4526) );
  A2O1A1Ixp33_ASAP7_75t_SL U38396 ( .A1(apbi[11]), .A2(n29745), .B(n25968), 
        .C(n25967), .Y(n4525) );
  AND2x2_ASAP7_75t_SL U38397 ( .A(n29985), .B(n31057), .Y(n28192) );
  OR2x2_ASAP7_75t_SL U38398 ( .A(uart1_r_RWADDR__0_), .B(uart1_r_RWADDR__1_), 
        .Y(n26021) );
  A2O1A1Ixp33_ASAP7_75t_SL U38399 ( .A1(uart1_r_RWADDR__1_), .A2(n28192), .B(
        n28191), .C(n25973), .Y(n2454) );
  INVx1_ASAP7_75t_SL U38400 ( .A(uart1_r_RWADDR__2_), .Y(n26023) );
  OR2x2_ASAP7_75t_SL U38401 ( .A(n26023), .B(n26001), .Y(n25975) );
  O2A1O1Ixp5_ASAP7_75t_SL U38402 ( .A1(n2456), .A2(n25975), .B(n28191), .C(
        n28192), .Y(n25977) );
  O2A1O1Ixp5_ASAP7_75t_SL U38403 ( .A1(n25976), .A2(n25975), .B(n2456), .C(
        n25977), .Y(uart1_v_RWADDR__3_) );
  INVx1_ASAP7_75t_SL U38404 ( .A(uart1_r_RWADDR__4_), .Y(n26003) );
  INVx1_ASAP7_75t_SL U38405 ( .A(n2456), .Y(n26004) );
  OAI21xp5_ASAP7_75t_SL U38406 ( .A1(n29369), .A2(n25980), .B(n26012), .Y(
        n26051) );
  OR2x2_ASAP7_75t_SL U38407 ( .A(n26065), .B(n26051), .Y(n31061) );
  OR2x2_ASAP7_75t_SL U38408 ( .A(n28108), .B(n31057), .Y(n26069) );
  OR2x2_ASAP7_75t_SL U38409 ( .A(uart1_r_RCNT__5_), .B(uart1_r_RCNT__4_), .Y(
        n29746) );
  NAND3xp33_ASAP7_75t_SL U38410 ( .A(n25983), .B(n30898), .C(n31503), .Y(
        n27510) );
  NAND3xp33_ASAP7_75t_SL U38411 ( .A(n25985), .B(n25984), .C(n2992), .Y(n25987) );
  OR3x1_ASAP7_75t_SL U38412 ( .A(n1637), .B(n25987), .C(n25986), .Y(n25989) );
  O2A1O1Ixp5_ASAP7_75t_SL U38413 ( .A1(n2389), .A2(n25994), .B(n2388), .C(
        n25993), .Y(n17458) );
  OR2x2_ASAP7_75t_SL U38414 ( .A(n2387), .B(n25995), .Y(n25996) );
  OR2x2_ASAP7_75t_SL U38415 ( .A(n2387), .B(n2388), .Y(n27449) );
  OAI21xp5_ASAP7_75t_SL U38416 ( .A1(n29369), .A2(n25998), .B(n26012), .Y(
        n26041) );
  OR2x2_ASAP7_75t_SL U38417 ( .A(n26065), .B(n26041), .Y(n31065) );
  OR2x2_ASAP7_75t_SL U38418 ( .A(n26031), .B(n26041), .Y(n31069) );
  OAI21xp5_ASAP7_75t_SL U38419 ( .A1(n29369), .A2(n26005), .B(n26012), .Y(
        n26064) );
  OR2x2_ASAP7_75t_SL U38420 ( .A(n26052), .B(n26064), .Y(n31073) );
  OR2x2_ASAP7_75t_SL U38421 ( .A(n26038), .B(n26041), .Y(n31077) );
  OR2x2_ASAP7_75t_SL U38422 ( .A(n26042), .B(n26064), .Y(n31081) );
  OR2x2_ASAP7_75t_SL U38423 ( .A(n26038), .B(n26064), .Y(n31085) );
  OAI21xp5_ASAP7_75t_SL U38424 ( .A1(n29369), .A2(n26013), .B(n26012), .Y(
        n26058) );
  OR2x2_ASAP7_75t_SL U38425 ( .A(n26048), .B(n26058), .Y(n31089) );
  OR2x2_ASAP7_75t_SL U38426 ( .A(n26031), .B(n26058), .Y(n31093) );
  OR2x2_ASAP7_75t_SL U38427 ( .A(n26042), .B(n26058), .Y(n31097) );
  OR2x2_ASAP7_75t_SL U38428 ( .A(n26048), .B(n26041), .Y(n31101) );
  OR2x2_ASAP7_75t_SL U38429 ( .A(n26031), .B(n26051), .Y(n31105) );
  OR2x2_ASAP7_75t_SL U38430 ( .A(n26035), .B(n26041), .Y(n31109) );
  OR2x2_ASAP7_75t_SL U38431 ( .A(n26059), .B(n26051), .Y(n31113) );
  OR2x2_ASAP7_75t_SL U38432 ( .A(n26038), .B(n26058), .Y(n31117) );
  OR2x2_ASAP7_75t_SL U38433 ( .A(n26035), .B(n26058), .Y(n31121) );
  OR2x2_ASAP7_75t_SL U38434 ( .A(n26052), .B(n26041), .Y(n31125) );
  OR2x2_ASAP7_75t_SL U38435 ( .A(n26048), .B(n26064), .Y(n31129) );
  OR2x2_ASAP7_75t_SL U38436 ( .A(n26042), .B(n26051), .Y(n31133) );
  OR2x2_ASAP7_75t_SL U38437 ( .A(n26059), .B(n26041), .Y(n31137) );
  OR2x2_ASAP7_75t_SL U38438 ( .A(n26035), .B(n26064), .Y(n31141) );
  OR2x2_ASAP7_75t_SL U38439 ( .A(n26031), .B(n26064), .Y(n31145) );
  OR2x2_ASAP7_75t_SL U38440 ( .A(n26052), .B(n26058), .Y(n31149) );
  OR2x2_ASAP7_75t_SL U38441 ( .A(n26035), .B(n26051), .Y(n31153) );
  OR2x2_ASAP7_75t_SL U38442 ( .A(n26038), .B(n26051), .Y(n31157) );
  OR2x2_ASAP7_75t_SL U38443 ( .A(n26042), .B(n26041), .Y(n31161) );
  OR2x2_ASAP7_75t_SL U38444 ( .A(n26059), .B(n26064), .Y(n31165) );
  OR2x2_ASAP7_75t_SL U38445 ( .A(n26048), .B(n26051), .Y(n31169) );
  OR2x2_ASAP7_75t_SL U38446 ( .A(n26052), .B(n26051), .Y(n31173) );
  OR2x2_ASAP7_75t_SL U38447 ( .A(n26065), .B(n26058), .Y(n31177) );
  OR2x2_ASAP7_75t_SL U38448 ( .A(n26059), .B(n26058), .Y(n31181) );
  OR2x2_ASAP7_75t_SL U38449 ( .A(n26065), .B(n26064), .Y(n31187) );
  AND2x2_ASAP7_75t_SL U38450 ( .A(n31372), .B(n27309), .Y(n29356) );
  AND2x2_ASAP7_75t_SL U38451 ( .A(n4518), .B(n4517), .Y(n27540) );
  NAND3xp33_ASAP7_75t_SL U38452 ( .A(n26075), .B(uart1_r_FLOW_), .C(
        uart1_r_LOOPB_), .Y(n26076) );
  XNOR2xp5_ASAP7_75t_SL U38453 ( .A(uart1_r_TICK_), .B(n26082), .Y(n26083) );
  NAND3xp33_ASAP7_75t_SL U38454 ( .A(n33065), .B(uart1_uarto_RXEN_), .C(
        uart1_r_RXDB__1_), .Y(n27537) );
  NAND3xp33_ASAP7_75t_SL U38455 ( .A(n27534), .B(n26091), .C(n27525), .Y(
        n26092) );
  OR2x2_ASAP7_75t_SL U38456 ( .A(n27537), .B(n28189), .Y(n30774) );
  OR2x2_ASAP7_75t_SL U38457 ( .A(n27493), .B(n31057), .Y(n26127) );
  OR2x2_ASAP7_75t_SL U38458 ( .A(n26129), .B(n28036), .Y(n27581) );
  AND2x2_ASAP7_75t_SL U38459 ( .A(n30007), .B(n29605), .Y(n28855) );
  OAI211xp5_ASAP7_75t_SL U38460 ( .A1(n23974), .A2(n26147), .B(n26146), .C(
        n26145), .Y(n27101) );
  OA21x2_ASAP7_75t_SL U38461 ( .A1(n28769), .A2(u0_0_leon3x0_p0_muli[23]), .B(
        n26161), .Y(u0_0_leon3x0_p0_divi[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38462 ( .A1(n26168), .A2(n26167), .B(n26166), .C(
        n26165), .Y(n30369) );
  AO21x1_ASAP7_75t_SL U38463 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__TBA__1_), .A2(
        n28480), .B(n26170), .Y(n26173) );
  A2O1A1Ixp33_ASAP7_75t_SL U38464 ( .A1(n26341), .A2(n27064), .B(n26177), .C(
        n24634), .Y(n26178) );
  NAND3xp33_ASAP7_75t_SL U38465 ( .A(n26180), .B(n26179), .C(n26178), .Y(
        n26183) );
  A2O1A1Ixp33_ASAP7_75t_SL U38466 ( .A1(u0_0_leon3x0_p0_dci[18]), .A2(n22398), 
        .B(n26183), .C(n26182), .Y(n26184) );
  OR2x2_ASAP7_75t_SL U38467 ( .A(u0_0_leon3x0_p0_divo[31]), .B(n29110), .Y(
        n26186) );
  OR2x2_ASAP7_75t_SL U38468 ( .A(n24658), .B(n28292), .Y(n31677) );
  O2A1O1Ixp5_ASAP7_75t_SL U38469 ( .A1(n29177), .A2(n26194), .B(n26193), .C(
        n18876), .Y(n26202) );
  OR2x2_ASAP7_75t_SL U38470 ( .A(n31884), .B(n18876), .Y(n26199) );
  NAND3xp33_ASAP7_75t_SL U38471 ( .A(n28489), .B(n27489), .C(n28506), .Y(
        n26218) );
  NAND3xp33_ASAP7_75t_SL U38472 ( .A(n26223), .B(n26222), .C(n26221), .Y(
        n30563) );
  AOI222xp33_ASAP7_75t_SL U38473 ( .A1(n29999), .A2(ahbso_0__HRDATA__26_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__26_), .C1(n24574), .C2(
        ahb0_r_HRDATAS__26_), .Y(n32399) );
  NAND3xp33_ASAP7_75t_SL U38474 ( .A(n26229), .B(n26228), .C(n26227), .Y(
        n26231) );
  NAND3xp33_ASAP7_75t_SL U38475 ( .A(n26235), .B(n26234), .C(n26233), .Y(
        n31044) );
  AND2x2_ASAP7_75t_SL U38476 ( .A(n3725), .B(n31676), .Y(n29925) );
  AO21x1_ASAP7_75t_SL U38477 ( .A1(n31830), .A2(u0_0_leon3x0_p0_iu_N5470), .B(
        n26238), .Y(n26239) );
  NAND3xp33_ASAP7_75t_SL U38478 ( .A(n26257), .B(n26256), .C(n26255), .Y(
        n28763) );
  OA21x2_ASAP7_75t_SL U38479 ( .A1(n28769), .A2(u0_0_leon3x0_p0_muli[17]), .B(
        n26261), .Y(u0_0_leon3x0_p0_divi[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38480 ( .A1(n26265), .A2(n26264), .B(n24486), .C(
        n26263), .Y(n30416) );
  OAI211xp5_ASAP7_75t_SL U38481 ( .A1(n30412), .A2(n29595), .B(n26267), .C(
        n26266), .Y(n26274) );
  OR2x2_ASAP7_75t_SL U38482 ( .A(n26270), .B(n26269), .Y(n26308) );
  OAI211xp5_ASAP7_75t_SL U38483 ( .A1(n29594), .A2(n30413), .B(n26272), .C(
        n26271), .Y(n26273) );
  AO21x1_ASAP7_75t_SL U38484 ( .A1(n28845), .A2(n27101), .B(n26277), .Y(n28873) );
  A2O1A1Ixp33_ASAP7_75t_SL U38485 ( .A1(n26284), .A2(n26283), .B(n26282), .C(
        n26281), .Y(n31016) );
  OAI222xp33_ASAP7_75t_SL U38486 ( .A1(n22373), .A2(n26285), .B1(n32610), .B2(
        n18806), .C1(n28352), .C2(n22374), .Y(n28806) );
  AO21x1_ASAP7_75t_SL U38487 ( .A1(n29150), .A2(n26307), .B(n18381), .Y(n26304) );
  NAND3xp33_ASAP7_75t_SL U38488 ( .A(n26304), .B(n24632), .C(n26307), .Y(
        n26306) );
  AND2x2_ASAP7_75t_SL U38489 ( .A(n28821), .B(u0_0_leon3x0_p0_divi[4]), .Y(
        n26309) );
  A2O1A1Ixp33_ASAP7_75t_SL U38490 ( .A1(n29148), .A2(n26307), .B(n26309), .C(
        n18381), .Y(n26303) );
  O2A1O1Ixp5_ASAP7_75t_SL U38491 ( .A1(n28771), .A2(n26307), .B(n26306), .C(
        n26305), .Y(n30425) );
  AO21x1_ASAP7_75t_SL U38492 ( .A1(u0_0_leon3x0_p0_iu_r_W__S__WIM__5_), .A2(
        n30611), .B(n26309), .Y(n26310) );
  A2O1A1Ixp33_ASAP7_75t_SL U38493 ( .A1(n27064), .A2(n28879), .B(n26310), .C(
        n24634), .Y(n26314) );
  NAND4xp25_ASAP7_75t_SL U38494 ( .A(n26314), .B(n26313), .C(n26312), .D(
        n26311), .Y(n26315) );
  A2O1A1Ixp33_ASAP7_75t_SL U38495 ( .A1(u0_0_leon3x0_p0_dci[10]), .A2(n22398), 
        .B(n26320), .C(n26319), .Y(n26321) );
  NAND3xp33_ASAP7_75t_SL U38496 ( .A(n26340), .B(n26339), .C(n26887), .Y(
        n26342) );
  NAND3xp33_ASAP7_75t_SL U38497 ( .A(n26346), .B(n26345), .C(n26344), .Y(
        n30968) );
  NOR3xp33_ASAP7_75t_SL U38498 ( .A(u0_0_leon3x0_p0_iu_r_X__CTRL__WY_), .B(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__25_), .C(
        u0_0_leon3x0_p0_iu_r_X__CTRL__INST__29_), .Y(n26357) );
  A2O1A1Ixp33_ASAP7_75t_SL U38499 ( .A1(n18614), .A2(n28931), .B(n26360), .C(
        n26359), .Y(n26361) );
  A2O1A1Ixp33_ASAP7_75t_SL U38500 ( .A1(n26364), .A2(n26363), .B(n26362), .C(
        n26361), .Y(n30626) );
  OAI211xp5_ASAP7_75t_SL U38501 ( .A1(n26380), .A2(n28986), .B(n26379), .C(
        n26378), .Y(n28498) );
  A2O1A1Ixp33_ASAP7_75t_SL U38502 ( .A1(n26388), .A2(n26387), .B(n26384), .C(
        n26386), .Y(n30261) );
  OAI211xp5_ASAP7_75t_SL U38503 ( .A1(n29592), .A2(n26397), .B(n26396), .C(
        n26395), .Y(n26400) );
  OAI211xp5_ASAP7_75t_SL U38504 ( .A1(n30258), .A2(n29594), .B(n29591), .C(
        n26398), .Y(n26399) );
  NAND4xp25_ASAP7_75t_SL U38505 ( .A(n26404), .B(n26403), .C(n26402), .D(
        n26401), .Y(n26407) );
  NAND3xp33_ASAP7_75t_SL U38506 ( .A(n28736), .B(n28405), .C(n24634), .Y(
        n26408) );
  A2O1A1Ixp33_ASAP7_75t_SL U38507 ( .A1(n26411), .A2(n26410), .B(n26409), .C(
        n26408), .Y(n29767) );
  AO21x1_ASAP7_75t_SL U38508 ( .A1(n31342), .A2(n29767), .B(n26414), .Y(n29791) );
  OAI211xp5_ASAP7_75t_SL U38509 ( .A1(n30265), .A2(n29594), .B(n26420), .C(
        n26419), .Y(n26421) );
  NAND3xp33_ASAP7_75t_SL U38510 ( .A(n26428), .B(n26427), .C(n26426), .Y(
        n28499) );
  A2O1A1Ixp33_ASAP7_75t_SL U38511 ( .A1(n26433), .A2(n26432), .B(n24487), .C(
        n26431), .Y(n30266) );
  NAND4xp25_ASAP7_75t_SL U38512 ( .A(n26437), .B(n26436), .C(n26435), .D(
        n26434), .Y(n26439) );
  A2O1A1Ixp33_ASAP7_75t_SL U38513 ( .A1(u0_0_leon3x0_p0_dci[28]), .A2(n22398), 
        .B(n26439), .C(n26438), .Y(n26440) );
  OR2x2_ASAP7_75t_SL U38514 ( .A(n31396), .B(n26523), .Y(n29072) );
  A2O1A1Ixp33_ASAP7_75t_SL U38515 ( .A1(n29073), .A2(n29072), .B(n31343), .C(
        n26442), .Y(n26443) );
  NAND3xp33_ASAP7_75t_SL U38516 ( .A(n26447), .B(n26446), .C(n26445), .Y(
        n32209) );
  NAND3xp33_ASAP7_75t_SL U38517 ( .A(n26588), .B(n26458), .C(n26457), .Y(
        n32233) );
  NAND3xp33_ASAP7_75t_SL U38518 ( .A(n26600), .B(n26487), .C(n26486), .Y(
        n32228) );
  OR2x2_ASAP7_75t_SL U38519 ( .A(n31954), .B(n1637), .Y(n31323) );
  NAND3xp33_ASAP7_75t_SL U38520 ( .A(n26513), .B(n26512), .C(n26511), .Y(
        n30479) );
  AO21x1_ASAP7_75t_SL U38521 ( .A1(n22375), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__19_), .B(n30006), .Y(n26533) );
  NAND3xp33_ASAP7_75t_SL U38522 ( .A(n26537), .B(n26536), .C(n26535), .Y(
        n32212) );
  A2O1A1Ixp33_ASAP7_75t_SL U38523 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[23]), .B(n26542), .C(n31638), .Y(n2351) );
  A2O1A1Ixp33_ASAP7_75t_SL U38524 ( .A1(n26570), .A2(n26569), .B(n26566), .C(
        n26568), .Y(n30349) );
  NAND4xp25_ASAP7_75t_SL U38525 ( .A(n26579), .B(n26578), .C(n26577), .D(
        n26576), .Y(n26581) );
  A2O1A1Ixp33_ASAP7_75t_SL U38526 ( .A1(u0_0_leon3x0_p0_dci[20]), .A2(n22398), 
        .B(n26581), .C(n26580), .Y(n26582) );
  NAND3xp33_ASAP7_75t_SL U38527 ( .A(n26588), .B(n26587), .C(n26586), .Y(
        n32343) );
  NAND3xp33_ASAP7_75t_SL U38528 ( .A(n26600), .B(n26599), .C(n26598), .Y(
        n32339) );
  AO21x1_ASAP7_75t_SL U38529 ( .A1(n28132), .A2(n27155), .B(n26611), .Y(n26613) );
  AOI222xp33_ASAP7_75t_SL U38530 ( .A1(n29999), .A2(ahbso_0__HRDATA__16_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__16_), .C1(n30000), .C2(
        ahb0_r_HRDATAS__16_), .Y(n32354) );
  NAND3xp33_ASAP7_75t_SL U38531 ( .A(n26668), .B(n26667), .C(n26666), .Y(
        n26669) );
  OAI211xp5_ASAP7_75t_SL U38532 ( .A1(n29594), .A2(n30334), .B(n26677), .C(
        n26676), .Y(n26678) );
  A2O1A1Ixp33_ASAP7_75t_SL U38533 ( .A1(n26688), .A2(n26687), .B(n26686), .C(
        n26685), .Y(n30337) );
  NAND3xp33_ASAP7_75t_SL U38534 ( .A(n26691), .B(n26690), .C(n26689), .Y(
        n26694) );
  A2O1A1Ixp33_ASAP7_75t_SL U38535 ( .A1(u0_0_leon3x0_p0_dci[21]), .A2(n22398), 
        .B(n26694), .C(n26693), .Y(n26695) );
  NAND3xp33_ASAP7_75t_SL U38536 ( .A(n27240), .B(n31542), .C(n27242), .Y(
        n26720) );
  OAI211xp5_ASAP7_75t_SL U38537 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__17_), 
        .A2(n28637), .B(n26701), .C(n26700), .Y(n26708) );
  NAND3xp33_ASAP7_75t_SL U38538 ( .A(n26706), .B(n26705), .C(n26704), .Y(
        n26707) );
  OAI211xp5_ASAP7_75t_SL U38539 ( .A1(n27209), .A2(n28502), .B(n26711), .C(
        n26710), .Y(n26713) );
  A2O1A1Ixp33_ASAP7_75t_SL U38540 ( .A1(u0_0_leon3x0_p0_dci[22]), .A2(n22398), 
        .B(n26713), .C(n26712), .Y(n26714) );
  OAI211xp5_ASAP7_75t_SL U38541 ( .A1(n31340), .A2(n27267), .B(n26717), .C(
        n26716), .Y(n26718) );
  OAI211xp5_ASAP7_75t_SL U38542 ( .A1(n24681), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__16_), .B(n26720), .C(n26719), .Y(n3986)
         );
  NAND3xp33_ASAP7_75t_SL U38543 ( .A(n26728), .B(n26727), .C(n26726), .Y(
        rf_di_w[31]) );
  OR2x2_ASAP7_75t_SL U38544 ( .A(u0_0_leon3x0_p0_iu_r_A__RSEL2__2_), .B(
        u0_0_leon3x0_p0_iu_r_A__RSEL2__1_), .Y(n26731) );
  OR2x2_ASAP7_75t_SL U38545 ( .A(u0_0_leon3x0_p0_iu_r_W__S__CWP__0_), .B(
        u0_0_leon3x0_p0_iu_r_W__S__CWP__1_), .Y(n26787) );
  A2O1A1Ixp33_ASAP7_75t_SL U38546 ( .A1(n26788), .A2(n26760), .B(n32158), .C(
        n26800), .Y(n26768) );
  NAND3xp33_ASAP7_75t_SL U38547 ( .A(n26789), .B(
        u0_0_leon3x0_p0_iu_r_W__S__CWP__0_), .C(n32158), .Y(n26763) );
  A2O1A1Ixp33_ASAP7_75t_SL U38548 ( .A1(n26796), .A2(n26769), .B(n26765), .C(
        n29179), .Y(n26766) );
  O2A1O1Ixp5_ASAP7_75t_SL U38549 ( .A1(n26800), .A2(n26769), .B(n26768), .C(
        n26767), .Y(n26776) );
  NAND3xp33_ASAP7_75t_SL U38550 ( .A(n26770), .B(n26800), .C(n32157), .Y(
        n26771) );
  A2O1A1Ixp33_ASAP7_75t_SL U38551 ( .A1(n26772), .A2(n26800), .B(n32157), .C(
        n26771), .Y(n26773) );
  XOR2xp5_ASAP7_75t_SL U38552 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__1_), .B(
        u0_0_leon3x0_p0_iu_v_A__CWP__0_), .Y(n26781) );
  OR2x2_ASAP7_75t_SL U38553 ( .A(u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(
        u0_0_leon3x0_p0_iu_v_A__CWP__1_), .Y(n26804) );
  XNOR2xp5_ASAP7_75t_SL U38554 ( .A(n32159), .B(n26790), .Y(n26793) );
  A2O1A1Ixp33_ASAP7_75t_SL U38555 ( .A1(n26796), .A2(n26801), .B(n26795), .C(
        n29179), .Y(n26797) );
  O2A1O1Ixp5_ASAP7_75t_SL U38556 ( .A1(n26801), .A2(n26800), .B(n26799), .C(
        n26798), .Y(n26802) );
  AOI222xp33_ASAP7_75t_SL U38557 ( .A1(n29999), .A2(ahbso_0__HRDATA__1_), .B1(
        n30002), .B2(ahbso_1__HRDATA__1_), .C1(n30000), .C2(ahb0_r_HRDATAS__1_), .Y(n32301) );
  NAND3xp33_ASAP7_75t_SL U38558 ( .A(n26847), .B(n26846), .C(n26845), .Y(
        n26848) );
  OR2x2_ASAP7_75t_SL U38559 ( .A(n28257), .B(n18825), .Y(n30811) );
  AO21x1_ASAP7_75t_SL U38560 ( .A1(u0_0_leon3x0_p0_iu_v_X__CTRL__RD__4_), .A2(
        n26855), .B(n30925), .Y(n26856) );
  NAND3xp33_ASAP7_75t_SL U38561 ( .A(n26867), .B(n26866), .C(n26865), .Y(
        n30809) );
  NAND3xp33_ASAP7_75t_SL U38562 ( .A(n32055), .B(n32083), .C(n32078), .Y(
        n26871) );
  NAND3xp33_ASAP7_75t_SL U38563 ( .A(n26871), .B(n26870), .C(n32090), .Y(
        n30812) );
  A2O1A1Ixp33_ASAP7_75t_SL U38564 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_27_), .A2(
        n31833), .B(n26878), .C(n26877), .Y(n4394) );
  OA21x2_ASAP7_75t_SL U38565 ( .A1(n28769), .A2(u0_0_leon3x0_p0_muli[34]), .B(
        n26890), .Y(u0_0_leon3x0_p0_divi[26]) );
  OAI211xp5_ASAP7_75t_SL U38566 ( .A1(n30241), .A2(n30625), .B(n26900), .C(
        n26899), .Y(n26901) );
  OAI211xp5_ASAP7_75t_SL U38567 ( .A1(n28443), .A2(n28502), .B(n26905), .C(
        n26904), .Y(n26907) );
  A2O1A1Ixp33_ASAP7_75t_SL U38568 ( .A1(u0_0_leon3x0_p0_dci[32]), .A2(n22398), 
        .B(n26907), .C(n26906), .Y(n26908) );
  OAI211xp5_ASAP7_75t_SL U38569 ( .A1(n26924), .A2(n29146), .B(
        u0_0_leon3x0_p0_divi[27]), .C(n24579), .Y(n26926) );
  A2O1A1Ixp33_ASAP7_75t_SL U38570 ( .A1(add_x_735_A_29_), .A2(n29150), .B(
        n26922), .C(n26921), .Y(n26925) );
  OAI211xp5_ASAP7_75t_SL U38571 ( .A1(n26929), .A2(n29592), .B(n29591), .C(
        n26928), .Y(n26930) );
  OAI211xp5_ASAP7_75t_SL U38572 ( .A1(n30237), .A2(n30625), .B(n26933), .C(
        n26932), .Y(n26934) );
  NAND4xp25_ASAP7_75t_SL U38573 ( .A(n26939), .B(n26941), .C(n26940), .D(
        n26942), .Y(n26943) );
  A2O1A1Ixp33_ASAP7_75t_SL U38574 ( .A1(u0_0_leon3x0_p0_dci[33]), .A2(n22398), 
        .B(n26943), .C(n30007), .Y(n26944) );
  OAI211xp5_ASAP7_75t_SL U38575 ( .A1(n31340), .A2(n26953), .B(n26952), .C(
        n26951), .Y(n26954) );
  O2A1O1Ixp5_ASAP7_75t_SL U38576 ( .A1(n22375), .A2(n28825), .B(n27002), .C(
        n26962), .Y(n32376) );
  NAND3xp33_ASAP7_75t_SL U38577 ( .A(n26966), .B(n26965), .C(n26964), .Y(
        n31480) );
  AOI222xp33_ASAP7_75t_SL U38578 ( .A1(n29999), .A2(ahbso_0__HRDATA__10_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__10_), .C1(n24574), .C2(
        ahb0_r_HRDATAS__10_), .Y(n32328) );
  AO21x1_ASAP7_75t_SL U38579 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5484), .B(
        n26973), .Y(n26974) );
  NAND3xp33_ASAP7_75t_SL U38580 ( .A(n26985), .B(n26984), .C(n26983), .Y(
        rf_di_w[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38581 ( .A1(u0_0_leon3x0_p0_divi[19]), .A2(n28821), 
        .B(n26989), .C(n22952), .Y(n29137) );
  OAI211xp5_ASAP7_75t_SL U38582 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__20_), 
        .A2(n28637), .B(n26995), .C(n26994), .Y(n26996) );
  NAND4xp25_ASAP7_75t_SL U38583 ( .A(n27001), .B(n27000), .C(n26999), .D(
        n26998), .Y(n27003) );
  A2O1A1Ixp33_ASAP7_75t_SL U38584 ( .A1(n28894), .A2(n30295), .B(n27003), .C(
        n27002), .Y(n27004) );
  NAND3xp33_ASAP7_75t_SL U38585 ( .A(n27006), .B(n27005), .C(n27004), .Y(
        n27007) );
  AO21x1_ASAP7_75t_SL U38586 ( .A1(n28902), .A2(u0_0_leon3x0_p0_dci[25]), .B(
        n27007), .Y(n27032) );
  AO21x1_ASAP7_75t_SL U38587 ( .A1(u0_0_leon3x0_p0_iu_de_icc_0_), .A2(n30652), 
        .B(n24647), .Y(n27019) );
  OR2x2_ASAP7_75t_SL U38588 ( .A(n30946), .B(n24679), .Y(n30679) );
  OR2x2_ASAP7_75t_SL U38589 ( .A(u0_0_leon3x0_p0_iu_r_E__CTRL__WICC_), .B(
        u0_0_leon3x0_p0_iu_r_M__CTRL__WICC_), .Y(n30667) );
  OR2x2_ASAP7_75t_SL U38590 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUSEL__1_), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_), .Y(n29870) );
  XNOR2xp5_ASAP7_75t_SL U38591 ( .A(u0_0_leon3x0_p0_iu_r_E__ALUADD_), .B(
        n27021), .Y(n27022) );
  OAI211xp5_ASAP7_75t_SL U38592 ( .A1(n22420), .A2(n27036), .B(n27023), .C(
        n31422), .Y(n27024) );
  OAI211xp5_ASAP7_75t_SL U38593 ( .A1(n31340), .A2(n27030), .B(n27029), .C(
        n27028), .Y(n27031) );
  A2O1A1Ixp33_ASAP7_75t_SL U38594 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_21_), .A2(
        n31833), .B(n27044), .C(n27043), .Y(n3240) );
  NAND3xp33_ASAP7_75t_SL U38595 ( .A(n27055), .B(n27054), .C(n27053), .Y(
        rf_di_w[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38596 ( .A1(u0_0_leon3x0_p0_divi[20]), .A2(n28827), 
        .B(n27060), .C(n23061), .Y(n27061) );
  A2O1A1Ixp33_ASAP7_75t_SL U38597 ( .A1(n27063), .A2(n27062), .B(n23061), .C(
        n27061), .Y(n29154) );
  OAI211xp5_ASAP7_75t_SL U38598 ( .A1(n23061), .A2(n27075), .B(n27074), .C(
        n27073), .Y(n27076) );
  NAND4xp25_ASAP7_75t_SL U38599 ( .A(n27082), .B(n27081), .C(n27080), .D(
        n27079), .Y(n27083) );
  A2O1A1Ixp33_ASAP7_75t_SL U38600 ( .A1(u0_0_leon3x0_p0_dci[26]), .A2(n22398), 
        .B(n27083), .C(n30007), .Y(n27084) );
  NAND3xp33_ASAP7_75t_SL U38601 ( .A(n27095), .B(n27094), .C(n27093), .Y(
        n28669) );
  AO21x1_ASAP7_75t_SL U38602 ( .A1(n29588), .A2(n18890), .B(n28887), .Y(n27114) );
  OAI211xp5_ASAP7_75t_SL U38603 ( .A1(n30389), .A2(n30625), .B(n27118), .C(
        n28426), .Y(n27119) );
  OAI211xp5_ASAP7_75t_SL U38604 ( .A1(n28666), .A2(n28790), .B(n27121), .C(
        n27120), .Y(n27123) );
  A2O1A1Ixp33_ASAP7_75t_SL U38605 ( .A1(u0_0_leon3x0_p0_dci[14]), .A2(n22398), 
        .B(n27123), .C(n27122), .Y(n27124) );
  A2O1A1Ixp33_ASAP7_75t_SL U38606 ( .A1(n27135), .A2(n28802), .B(n27134), .C(
        n27133), .Y(n2310) );
  OAI211xp5_ASAP7_75t_SL U38607 ( .A1(n27144), .A2(n29146), .B(
        u0_0_leon3x0_p0_divi[9]), .C(n24580), .Y(n27146) );
  A2O1A1Ixp33_ASAP7_75t_SL U38608 ( .A1(n29150), .A2(n22837), .B(n27140), .C(
        n27139), .Y(n27145) );
  NAND3xp33_ASAP7_75t_SL U38609 ( .A(n27151), .B(n27150), .C(n27149), .Y(
        n27152) );
  A2O1A1Ixp33_ASAP7_75t_SL U38610 ( .A1(n27155), .A2(n28737), .B(n27154), .C(
        n24634), .Y(n27156) );
  OAI211xp5_ASAP7_75t_SL U38611 ( .A1(n30386), .A2(n30625), .B(n27157), .C(
        n27156), .Y(n27158) );
  OAI211xp5_ASAP7_75t_SL U38612 ( .A1(n27161), .A2(n27208), .B(n27160), .C(
        n27159), .Y(n27162) );
  A2O1A1Ixp33_ASAP7_75t_SL U38613 ( .A1(u0_0_leon3x0_p0_dci[15]), .A2(n22398), 
        .B(n27162), .C(n30007), .Y(n27163) );
  AO21x1_ASAP7_75t_SL U38614 ( .A1(n31342), .A2(n31055), .B(n27167), .Y(n31050) );
  OAI211xp5_ASAP7_75t_SL U38615 ( .A1(n31340), .A2(n27172), .B(n27171), .C(
        n27170), .Y(n27173) );
  NAND3xp33_ASAP7_75t_SL U38616 ( .A(n27187), .B(n27186), .C(n27185), .Y(
        rf_di_w[14]) );
  OAI222xp33_ASAP7_75t_SL U38617 ( .A1(n22374), .A2(n28336), .B1(n32624), .B2(
        n18806), .C1(n27191), .C2(n22373), .Y(n28601) );
  A2O1A1Ixp33_ASAP7_75t_SL U38618 ( .A1(n27203), .A2(n27202), .B(n27198), .C(
        n27201), .Y(n30360) );
  OAI211xp5_ASAP7_75t_SL U38619 ( .A1(n29594), .A2(n30357), .B(n27205), .C(
        n27204), .Y(n27206) );
  A2O1A1Ixp33_ASAP7_75t_SL U38620 ( .A1(n27215), .A2(n27214), .B(n24427), .C(
        n27213), .Y(n27216) );
  A2O1A1Ixp33_ASAP7_75t_SL U38621 ( .A1(u0_0_leon3x0_p0_dci[19]), .A2(n22398), 
        .B(n27216), .C(n30007), .Y(n27217) );
  OAI211xp5_ASAP7_75t_SL U38622 ( .A1(n31340), .A2(n30496), .B(n27220), .C(
        n27219), .Y(n27221) );
  AO21x1_ASAP7_75t_SL U38623 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5480), .B(
        n27227), .Y(n27228) );
  NAND3xp33_ASAP7_75t_SL U38624 ( .A(n27239), .B(n27238), .C(n27237), .Y(
        rf_di_w[16]) );
  AOI222xp33_ASAP7_75t_SL U38625 ( .A1(n29999), .A2(ahbso_0__HRDATA__17_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__17_), .C1(n30000), .C2(
        ahb0_r_HRDATAS__17_), .Y(n32361) );
  AO21x1_ASAP7_75t_SL U38626 ( .A1(n22375), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__17_), .B(n30006), .Y(n27244) );
  NAND3xp33_ASAP7_75t_SL U38627 ( .A(n27247), .B(n27246), .C(n27245), .Y(
        n32210) );
  A2O1A1Ixp33_ASAP7_75t_SL U38628 ( .A1(n24647), .A2(n27255), .B(n28759), .C(
        n28701), .Y(n27256) );
  AO21x1_ASAP7_75t_SL U38629 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5481), .B(
        n27269), .Y(n27270) );
  NAND3xp33_ASAP7_75t_SL U38630 ( .A(n27278), .B(n27277), .C(n27276), .Y(
        rf_di_w[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38631 ( .A1(irqctrl0_r_IFORCE__0__1_), .A2(n27296), 
        .B(n27295), .C(n27297), .Y(n2700) );
  AND2x2_ASAP7_75t_SL U38632 ( .A(uart1_r_TRADDR__0_), .B(uart1_r_TRADDR__1_), 
        .Y(n27895) );
  INVx1_ASAP7_75t_SL U38633 ( .A(uart1_r_TWADDR__0_), .Y(n27357) );
  NAND3xp33_ASAP7_75t_SL U38634 ( .A(n27306), .B(n24694), .C(n27307), .Y(n2268) );
  XNOR2xp5_ASAP7_75t_SL U38635 ( .A(n27394), .B(n27895), .Y(n27312) );
  XNOR2xp5_ASAP7_75t_SL U38636 ( .A(uart1_r_TRADDR__4_), .B(n27318), .Y(n27319) );
  NAND3xp33_ASAP7_75t_SL U38637 ( .A(n31325), .B(n2267), .C(n27327), .Y(n27329) );
  NAND3xp33_ASAP7_75t_SL U38638 ( .A(n27343), .B(uart1_r_TWADDR__0_), .C(
        uart1_r_TWADDR__2_), .Y(n27353) );
  NAND3xp33_ASAP7_75t_SL U38639 ( .A(n27343), .B(n27355), .C(
        uart1_r_TWADDR__0_), .Y(n27351) );
  NAND3xp33_ASAP7_75t_SL U38640 ( .A(n27355), .B(n27357), .C(
        uart1_r_TWADDR__1_), .Y(n27369) );
  NAND3xp33_ASAP7_75t_SL U38641 ( .A(n27357), .B(uart1_r_TWADDR__1_), .C(
        uart1_r_TWADDR__2_), .Y(n27364) );
  OR2x2_ASAP7_75t_SL U38642 ( .A(uart1_r_TWADDR__2_), .B(n27373), .Y(n27385)
         );
  OR2x2_ASAP7_75t_SL U38643 ( .A(n27391), .B(n27390), .Y(n27405) );
  NAND3xp33_ASAP7_75t_SL U38644 ( .A(n27393), .B(uart1_r_TRADDR__4_), .C(
        uart1_r_TRADDR__2_), .Y(n27407) );
  NAND4xp25_ASAP7_75t_SL U38645 ( .A(n27399), .B(n27398), .C(n27397), .D(
        n27396), .Y(n27400) );
  NAND4xp25_ASAP7_75t_SL U38646 ( .A(n27404), .B(n27403), .C(n27402), .D(
        n27401), .Y(n27423) );
  AO21x1_ASAP7_75t_SL U38647 ( .A1(uart1_r_THOLD__24__1_), .A2(n28017), .B(
        uart1_r_TRADDR__1_), .Y(n27406) );
  NAND4xp25_ASAP7_75t_SL U38648 ( .A(n27415), .B(n27414), .C(n27413), .D(
        n27412), .Y(n27422) );
  AO21x1_ASAP7_75t_SL U38649 ( .A1(uart1_r_THOLD__18__1_), .A2(n28010), .B(
        n28016), .Y(n27416) );
  NAND4xp25_ASAP7_75t_SL U38650 ( .A(n27420), .B(n27419), .C(n27418), .D(
        n27417), .Y(n27421) );
  A2O1A1Ixp33_ASAP7_75t_SL U38651 ( .A1(uart1_r_TRADDR__0_), .A2(n27423), .B(
        n27422), .C(n27421), .Y(n27424) );
  NAND3xp33_ASAP7_75t_SL U38652 ( .A(n27428), .B(n2389), .C(n2386), .Y(n27448)
         );
  NAND3xp33_ASAP7_75t_SL U38653 ( .A(n27428), .B(n27445), .C(n2389), .Y(n27471) );
  OR2x2_ASAP7_75t_SL U38654 ( .A(n2386), .B(n27444), .Y(n27447) );
  NAND4xp25_ASAP7_75t_SL U38655 ( .A(n27433), .B(n27436), .C(n27435), .D(
        n27434), .Y(n27458) );
  NAND4xp25_ASAP7_75t_SL U38656 ( .A(n27443), .B(n27442), .C(n27441), .D(
        n27440), .Y(n27457) );
  OR2x2_ASAP7_75t_SL U38657 ( .A(n27445), .B(n27444), .Y(n27470) );
  NAND4xp25_ASAP7_75t_SL U38658 ( .A(n27455), .B(n27454), .C(n27453), .D(
        n27452), .Y(n27456) );
  OAI31xp33_ASAP7_75t_SL U38659 ( .A1(n27458), .A2(n27457), .A3(n27456), .B(
        n30870), .Y(n27468) );
  AND2x2_ASAP7_75t_SL U38660 ( .A(n27461), .B(n27463), .Y(n31245) );
  NAND4xp25_ASAP7_75t_SL U38661 ( .A(n27468), .B(n27467), .C(n27466), .D(
        n27465), .Y(n27488) );
  OR2x2_ASAP7_75t_SL U38662 ( .A(n27469), .B(n31238), .Y(n27472) );
  NAND3xp33_ASAP7_75t_SL U38663 ( .A(n27486), .B(n27485), .C(n27484), .Y(
        n27487) );
  A2O1A1Ixp33_ASAP7_75t_SL U38664 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[5]), .B(n27494), .C(n31638), .Y(n4533) );
  O2A1O1Ixp5_ASAP7_75t_SL U38665 ( .A1(uart1_r_RCNT__2_), .A2(n27506), .B(
        n27505), .C(n27504), .Y(n27512) );
  NAND3xp33_ASAP7_75t_SL U38666 ( .A(n27521), .B(uart1_r_RCNT__5_), .C(n31940), 
        .Y(n27514) );
  XOR2xp5_ASAP7_75t_SL U38667 ( .A(uart1_r_DPAR_), .B(uart1_v_RXDB__1_), .Y(
        n27527) );
  A2O1A1Ixp33_ASAP7_75t_SL U38668 ( .A1(n29961), .A2(n27529), .B(n27528), .C(
        n27527), .Y(n27530) );
  O2A1O1Ixp5_ASAP7_75t_SL U38669 ( .A1(n29950), .A2(n27531), .B(n27530), .C(
        n27533), .Y(n27532) );
  AND2x2_ASAP7_75t_SL U38670 ( .A(n2867), .B(n24694), .Y(n29336) );
  OR2x2_ASAP7_75t_SL U38671 ( .A(n28187), .B(n27535), .Y(n29973) );
  OR2x2_ASAP7_75t_SL U38672 ( .A(n29951), .B(n28036), .Y(n29948) );
  OAI211xp5_ASAP7_75t_SL U38673 ( .A1(n27985), .A2(n27626), .B(n27625), .C(
        n27624), .Y(n27634) );
  NAND4xp25_ASAP7_75t_SL U38674 ( .A(n27632), .B(n27631), .C(n27630), .D(
        n27629), .Y(n27633) );
  O2A1O1Ixp5_ASAP7_75t_SL U38675 ( .A1(n27635), .A2(n27634), .B(
        uart1_r_TRADDR__0_), .C(n27633), .Y(n27649) );
  NAND4xp25_ASAP7_75t_SL U38676 ( .A(n27639), .B(n27638), .C(n27637), .D(
        n27636), .Y(n27647) );
  NAND3xp33_ASAP7_75t_SL U38677 ( .A(n27644), .B(n27643), .C(n27642), .Y(
        n27645) );
  AOI222xp33_ASAP7_75t_SL U38678 ( .A1(n29954), .A2(uart1_r_TSHIFT__7_), .B1(
        n29951), .B2(uart1_r_TSHIFT__8_), .C1(n28030), .C2(n31239), .Y(n4707)
         );
  NAND4xp25_ASAP7_75t_SL U38679 ( .A(n27693), .B(n27692), .C(n27691), .D(
        n27690), .Y(n27713) );
  NAND4xp25_ASAP7_75t_SL U38680 ( .A(n27697), .B(n27696), .C(n27695), .D(
        n27694), .Y(n27712) );
  NAND4xp25_ASAP7_75t_SL U38681 ( .A(n27701), .B(n27700), .C(n27699), .D(
        n27698), .Y(n27702) );
  AO21x1_ASAP7_75t_SL U38682 ( .A1(uart1_r_THOLD__26__5_), .A2(n28017), .B(
        n28016), .Y(n27705) );
  NAND4xp25_ASAP7_75t_SL U38683 ( .A(n27710), .B(n27709), .C(n27708), .D(
        n27707), .Y(n27711) );
  A2O1A1Ixp33_ASAP7_75t_SL U38684 ( .A1(uart1_r_TRADDR__0_), .A2(n27713), .B(
        n27712), .C(n27711), .Y(n30077) );
  OAI211xp5_ASAP7_75t_SL U38685 ( .A1(n27771), .A2(n27756), .B(n27755), .C(
        n27754), .Y(n27767) );
  NAND4xp25_ASAP7_75t_SL U38686 ( .A(n27764), .B(n27763), .C(n27762), .D(
        n27761), .Y(n27765) );
  O2A1O1Ixp5_ASAP7_75t_SL U38687 ( .A1(n27767), .A2(n27766), .B(
        uart1_r_TRADDR__0_), .C(n27765), .Y(n27785) );
  OAI211xp5_ASAP7_75t_SL U38688 ( .A1(n27771), .A2(n27770), .B(n27769), .C(
        n27768), .Y(n27783) );
  NAND4xp25_ASAP7_75t_SL U38689 ( .A(n27780), .B(n27779), .C(n27778), .D(
        n27777), .Y(n27781) );
  O2A1O1Ixp5_ASAP7_75t_SL U38690 ( .A1(n27783), .A2(n27782), .B(
        uart1_r_TRADDR__0_), .C(n27781), .Y(n27784) );
  AOI222xp33_ASAP7_75t_SL U38691 ( .A1(n29954), .A2(uart1_r_TSHIFT__5_), .B1(
        n29951), .B2(uart1_r_TSHIFT__6_), .C1(n28030), .C2(n30782), .Y(n4705)
         );
  NAND4xp25_ASAP7_75t_SL U38692 ( .A(n27829), .B(n27828), .C(n27827), .D(
        n27826), .Y(n27849) );
  NAND4xp25_ASAP7_75t_SL U38693 ( .A(n27833), .B(n27832), .C(n27831), .D(
        n27830), .Y(n27848) );
  NAND4xp25_ASAP7_75t_SL U38694 ( .A(n27837), .B(n27836), .C(n27835), .D(
        n27834), .Y(n27838) );
  AO21x1_ASAP7_75t_SL U38695 ( .A1(uart1_r_THOLD__24__3_), .A2(n28017), .B(
        uart1_r_TRADDR__1_), .Y(n27841) );
  NAND4xp25_ASAP7_75t_SL U38696 ( .A(n27846), .B(n27845), .C(n27844), .D(
        n27843), .Y(n27847) );
  NAND4xp25_ASAP7_75t_SL U38697 ( .A(n27893), .B(n27892), .C(n27891), .D(
        n27890), .Y(n27894) );
  NAND4xp25_ASAP7_75t_SL U38698 ( .A(n27899), .B(n27898), .C(n27897), .D(
        n27896), .Y(n27912) );
  NAND4xp25_ASAP7_75t_SL U38699 ( .A(n27905), .B(n27904), .C(n27903), .D(
        n27902), .Y(n27911) );
  NAND4xp25_ASAP7_75t_SL U38700 ( .A(n27909), .B(n27908), .C(n27907), .D(
        n27906), .Y(n27910) );
  A2O1A1Ixp33_ASAP7_75t_SL U38701 ( .A1(uart1_r_TRADDR__0_), .A2(n27912), .B(
        n27911), .C(n27910), .Y(n27913) );
  AOI222xp33_ASAP7_75t_SL U38702 ( .A1(n29559), .A2(n28030), .B1(
        uart1_r_TSHIFT__4_), .B2(n29951), .C1(n29954), .C2(uart1_r_TSHIFT__3_), 
        .Y(n4703) );
  OAI211xp5_ASAP7_75t_SL U38703 ( .A1(n27985), .A2(n27984), .B(n27983), .C(
        n27982), .Y(n27994) );
  NAND4xp25_ASAP7_75t_SL U38704 ( .A(n27992), .B(n27991), .C(n27990), .D(
        n27989), .Y(n27993) );
  NAND4xp25_ASAP7_75t_SL U38705 ( .A(n28007), .B(n28006), .C(n28005), .D(
        n28004), .Y(n28024) );
  NAND3xp33_ASAP7_75t_SL U38706 ( .A(n28021), .B(n28020), .C(n28019), .Y(
        n28022) );
  AO21x1_ASAP7_75t_SL U38707 ( .A1(n28030), .A2(n28084), .B(n28029), .Y(n17443) );
  AO21x1_ASAP7_75t_SL U38708 ( .A1(n28034), .A2(n28033), .B(n4519), .Y(n28035)
         );
  OAI211xp5_ASAP7_75t_SL U38709 ( .A1(n29351), .A2(n28043), .B(n28049), .C(
        n24694), .Y(n4515) );
  O2A1O1Ixp5_ASAP7_75t_SL U38710 ( .A1(uart1_r_TCNT__2_), .A2(n28048), .B(
        uart1_r_TCNT__3_), .C(n28051), .Y(n28050) );
  AO21x1_ASAP7_75t_SL U38711 ( .A1(n28050), .A2(n28049), .B(n28055), .Y(n5592)
         );
  XNOR2xp5_ASAP7_75t_SL U38712 ( .A(uart1_r_TCNT__4_), .B(n28052), .Y(n28054)
         );
  NAND3xp33_ASAP7_75t_SL U38713 ( .A(n28063), .B(n28062), .C(n28061), .Y(
        n28069) );
  NAND4xp25_ASAP7_75t_SL U38714 ( .A(n28067), .B(n28066), .C(n28065), .D(
        n28064), .Y(n28068) );
  NAND4xp25_ASAP7_75t_SL U38715 ( .A(n28073), .B(n28072), .C(n28071), .D(
        n28070), .Y(n28079) );
  NAND4xp25_ASAP7_75t_SL U38716 ( .A(n28077), .B(n28076), .C(n28075), .D(
        n28074), .Y(n28078) );
  OR2x2_ASAP7_75t_SL U38717 ( .A(n4536), .B(n28085), .Y(n31236) );
  NAND3xp33_ASAP7_75t_SL U38718 ( .A(n28087), .B(n28086), .C(n31236), .Y(
        n28088) );
  NAND3xp33_ASAP7_75t_SL U38719 ( .A(n28092), .B(n28091), .C(n28090), .Y(
        n28099) );
  O2A1O1Ixp5_ASAP7_75t_SL U38720 ( .A1(n28099), .A2(n28098), .B(n31954), .C(
        n28097), .Y(n4368) );
  AND2x2_ASAP7_75t_SL U38721 ( .A(u0_0_leon3x0_p0_iu_r_E__OP1__0_), .B(n22375), 
        .Y(n29009) );
  AND2x2_ASAP7_75t_SL U38722 ( .A(n29563), .B(n29003), .Y(n28105) );
  O2A1O1Ixp5_ASAP7_75t_SL U38723 ( .A1(n28105), .A2(n28104), .B(n29937), .C(
        n28103), .Y(n28106) );
  A2O1A1Ixp33_ASAP7_75t_SL U38724 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[4]), .B(n28109), .C(n31638), .Y(n4365) );
  NAND3xp33_ASAP7_75t_SL U38725 ( .A(n18882), .B(n4770), .C(n28115), .Y(n28112) );
  A2O1A1Ixp33_ASAP7_75t_SL U38726 ( .A1(timer0_vtimers_1__ENABLE_), .A2(n28112), .B(n28111), .C(n30030), .Y(n28113) );
  A2O1A1Ixp33_ASAP7_75t_SL U38727 ( .A1(apbi[0]), .A2(n30738), .B(n28114), .C(
        n24694), .Y(n4364) );
  A2O1A1Ixp33_ASAP7_75t_SL U38728 ( .A1(n28128), .A2(n28127), .B(
        apb0_r_CFGSEL_), .C(n28126), .Y(n28129) );
  AOI222xp33_ASAP7_75t_SL U38729 ( .A1(n29999), .A2(ahbso_0__HRDATA__11_), 
        .B1(n30002), .B2(ahbso_1__HRDATA__11_), .C1(n30000), .C2(
        ahb0_r_HRDATAS__11_), .Y(n32333) );
  A2O1A1Ixp33_ASAP7_75t_SL U38730 ( .A1(n28140), .A2(n28172), .B(n28139), .C(
        n28138), .Y(uart1_v_SCALER__11_) );
  A2O1A1Ixp33_ASAP7_75t_SL U38731 ( .A1(uart1_scaler_10_), .A2(n28174), .B(
        n28146), .C(n28145), .Y(n2874) );
  A2O1A1Ixp33_ASAP7_75t_SL U38732 ( .A1(uart1_scaler_9_), .A2(n28174), .B(
        n28150), .C(n28149), .Y(n1799) );
  A2O1A1Ixp33_ASAP7_75t_SL U38733 ( .A1(uart1_scaler_4_), .A2(n28174), .B(
        n28158), .C(n28157), .Y(n2878) );
  A2O1A1Ixp33_ASAP7_75t_SL U38734 ( .A1(uart1_scaler_3_), .A2(n28174), .B(
        n28162), .C(n28161), .Y(n2877) );
  A2O1A1Ixp33_ASAP7_75t_SL U38735 ( .A1(uart1_scaler_2_), .A2(n28174), .B(
        n28166), .C(n28165), .Y(n2876) );
  A2O1A1Ixp33_ASAP7_75t_SL U38736 ( .A1(uart1_scaler_1_), .A2(n28174), .B(
        n28171), .C(n28170), .Y(n2875) );
  OR2x2_ASAP7_75t_SL U38737 ( .A(uart1_r_EXTCLKEN_), .B(n28179), .Y(n4683) );
  XNOR2xp5_ASAP7_75t_SL U38738 ( .A(n28184), .B(n28185), .Y(n28183) );
  NAND3xp33_ASAP7_75t_SL U38739 ( .A(n29961), .B(uart1_r_PAREN_), .C(n29956), 
        .Y(n29964) );
  A2O1A1Ixp33_ASAP7_75t_SL U38740 ( .A1(uart1_r_RXTICK_), .A2(n28189), .B(
        n28186), .C(n24694), .Y(n29974) );
  OR2x2_ASAP7_75t_SL U38741 ( .A(n29510), .B(n31057), .Y(n28225) );
  NAND4xp25_ASAP7_75t_SL U38742 ( .A(n28230), .B(n28229), .C(n28228), .D(
        n28227), .Y(n31192) );
  A2O1A1Ixp33_ASAP7_75t_SL U38743 ( .A1(irqctrl0_r_IFORCE__0__3_), .A2(n28240), 
        .B(n28239), .C(n28238), .Y(n2349) );
  A2O1A1Ixp33_ASAP7_75t_SL U38744 ( .A1(n29510), .A2(n29325), .B(n28245), .C(
        n28244), .Y(n2348) );
  AO21x1_ASAP7_75t_SL U38745 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5492), .B(
        n28260), .Y(n28261) );
  NAND3xp33_ASAP7_75t_SL U38746 ( .A(n28270), .B(n28269), .C(n28268), .Y(
        rf_di_w[28]) );
  OAI222xp33_ASAP7_75t_SL U38747 ( .A1(n22374), .A2(n28302), .B1(n32656), .B2(
        n18805), .C1(n29023), .C2(n22373), .Y(n29866) );
  A2O1A1Ixp33_ASAP7_75t_SL U38748 ( .A1(u0_0_leon3x0_p0_div0_addout_32_), .A2(
        n29110), .B(n28284), .C(n22431), .Y(n28290) );
  A2O1A1Ixp33_ASAP7_75t_SL U38749 ( .A1(n28290), .A2(n28289), .B(n28288), .C(
        n28287), .Y(n18168) );
  OAI211xp5_ASAP7_75t_SL U38750 ( .A1(n2307), .A2(n31660), .B(n28297), .C(
        n28296), .Y(u0_0_leon3x0_p0_div0_vaddin1[32]) );
  OAI211xp5_ASAP7_75t_SL U38751 ( .A1(n31675), .A2(n31660), .B(n28300), .C(
        n28299), .Y(u0_0_leon3x0_p0_div0_vaddin1[31]) );
  OAI211xp5_ASAP7_75t_SL U38752 ( .A1(n22420), .A2(n29792), .B(n28307), .C(
        n31422), .Y(n28308) );
  OAI211xp5_ASAP7_75t_SL U38753 ( .A1(n22420), .A2(n28312), .B(n28311), .C(
        n31422), .Y(n28313) );
  OAI211xp5_ASAP7_75t_SL U38754 ( .A1(n28316), .A2(n31660), .B(n28315), .C(
        n28314), .Y(u0_0_leon3x0_p0_div0_vaddin1[23]) );
  OAI211xp5_ASAP7_75t_SL U38755 ( .A1(n28319), .A2(n31660), .B(n28318), .C(
        n28317), .Y(u0_0_leon3x0_p0_div0_vaddin1[21]) );
  OAI211xp5_ASAP7_75t_SL U38756 ( .A1(n28327), .A2(n31660), .B(n28326), .C(
        n28325), .Y(u0_0_leon3x0_p0_div0_vaddin1[17]) );
  OAI211xp5_ASAP7_75t_SL U38757 ( .A1(n28333), .A2(n31660), .B(n28332), .C(
        n28331), .Y(u0_0_leon3x0_p0_div0_vaddin1[15]) );
  OAI211xp5_ASAP7_75t_SL U38758 ( .A1(n28648), .A2(n31660), .B(n28339), .C(
        n28338), .Y(u0_0_leon3x0_p0_div0_vaddin1[12]) );
  OAI211xp5_ASAP7_75t_SL U38759 ( .A1(n28697), .A2(n31660), .B(n28341), .C(
        n28340), .Y(u0_0_leon3x0_p0_div0_vaddin1[11]) );
  OAI211xp5_ASAP7_75t_SL U38760 ( .A1(n28344), .A2(n31660), .B(n28343), .C(
        n28342), .Y(u0_0_leon3x0_p0_div0_vaddin1[10]) );
  OAI211xp5_ASAP7_75t_SL U38761 ( .A1(n28347), .A2(n31660), .B(n28346), .C(
        n28345), .Y(u0_0_leon3x0_p0_div0_vaddin1[9]) );
  OAI211xp5_ASAP7_75t_SL U38762 ( .A1(n28749), .A2(n31660), .B(n28349), .C(
        n28348), .Y(u0_0_leon3x0_p0_div0_vaddin1[8]) );
  OAI211xp5_ASAP7_75t_SL U38763 ( .A1(n28794), .A2(n31660), .B(n28351), .C(
        n28350), .Y(u0_0_leon3x0_p0_div0_vaddin1[7]) );
  OAI211xp5_ASAP7_75t_SL U38764 ( .A1(n28356), .A2(n31660), .B(n28355), .C(
        n28354), .Y(u0_0_leon3x0_p0_div0_vaddin1[5]) );
  OAI211xp5_ASAP7_75t_SL U38765 ( .A1(n28860), .A2(n31660), .B(n28359), .C(
        n28358), .Y(u0_0_leon3x0_p0_div0_vaddin1[4]) );
  OAI211xp5_ASAP7_75t_SL U38766 ( .A1(n28903), .A2(n31660), .B(n28361), .C(
        n28360), .Y(u0_0_leon3x0_p0_div0_vaddin1[3]) );
  OAI211xp5_ASAP7_75t_SL U38767 ( .A1(n28364), .A2(n31660), .B(n28363), .C(
        n28362), .Y(u0_0_leon3x0_p0_div0_vaddin1[2]) );
  AO21x1_ASAP7_75t_SL U38768 ( .A1(n30453), .A2(n30609), .B(n24647), .Y(n28366) );
  OAI211xp5_ASAP7_75t_SL U38769 ( .A1(n28370), .A2(n31660), .B(n28369), .C(
        n28368), .Y(u0_0_leon3x0_p0_div0_vaddin1[1]) );
  NAND3xp33_ASAP7_75t_SL U38770 ( .A(n28376), .B(n28375), .C(n28374), .Y(
        u0_0_leon3x0_p0_div0_vaddin1[0]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38771 ( .A1(u0_0_leon3x0_p0_divi[27]), .A2(n22410), 
        .B(n28382), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[28]) );
  AO21x1_ASAP7_75t_SL U38772 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5490), .B(
        n28387), .Y(n28388) );
  NAND3xp33_ASAP7_75t_SL U38773 ( .A(n28399), .B(n28398), .C(n28397), .Y(
        rf_di_w[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38774 ( .A1(u0_0_leon3x0_p0_divi[25]), .A2(n22410), 
        .B(n28401), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[26]) );
  NAND3xp33_ASAP7_75t_SL U38775 ( .A(n28410), .B(n28409), .C(n28408), .Y(
        n31357) );
  AO21x1_ASAP7_75t_SL U38776 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5489), .B(
        n28415), .Y(n28416) );
  OAI211xp5_ASAP7_75t_SL U38777 ( .A1(n28422), .A2(n29592), .B(n28421), .C(
        n29591), .Y(n28423) );
  NAND4xp25_ASAP7_75t_SL U38778 ( .A(n28429), .B(n28428), .C(n28427), .D(
        n28426), .Y(n28439) );
  OA21x2_ASAP7_75t_SL U38779 ( .A1(n28769), .A2(u0_0_leon3x0_p0_muli[33]), .B(
        n28430), .Y(u0_0_leon3x0_p0_divi[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38780 ( .A1(u0_0_leon3x0_p0_divi[24]), .A2(n28827), 
        .B(n28432), .C(n24691), .Y(n28435) );
  OAI211xp5_ASAP7_75t_SL U38781 ( .A1(n28790), .A2(n28443), .B(n28442), .C(
        n28441), .Y(n28445) );
  A2O1A1Ixp33_ASAP7_75t_SL U38782 ( .A1(u0_0_leon3x0_p0_dci[30]), .A2(n22398), 
        .B(n28445), .C(n28444), .Y(n28446) );
  AO21x1_ASAP7_75t_SL U38783 ( .A1(n23229), .A2(n29789), .B(n28449), .Y(n4123)
         );
  OAI222xp33_ASAP7_75t_SL U38784 ( .A1(n22374), .A2(n28452), .B1(n32648), .B2(
        n18805), .C1(n28451), .C2(n22373), .Y(n29787) );
  NAND3xp33_ASAP7_75t_SL U38785 ( .A(n28459), .B(n28458), .C(n28457), .Y(
        rf_di_w[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38786 ( .A1(u0_0_leon3x0_p0_divi[24]), .A2(n22410), 
        .B(n28460), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38787 ( .A1(n28469), .A2(n28802), .B(n28468), .C(
        n28467), .Y(n2490) );
  A2O1A1Ixp33_ASAP7_75t_SL U38788 ( .A1(u0_0_leon3x0_p0_divi[23]), .A2(n22410), 
        .B(n28470), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38789 ( .A1(u0_0_leon3x0_p0_divi[22]), .A2(n22410), 
        .B(n28473), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[23]) );
  AO21x1_ASAP7_75t_SL U38790 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5486), .B(
        n28476), .Y(n28477) );
  OAI211xp5_ASAP7_75t_SL U38791 ( .A1(n28827), .A2(n28491), .B(n28484), .C(
        n28483), .Y(n28485) );
  OAI211xp5_ASAP7_75t_SL U38792 ( .A1(n28503), .A2(n28502), .B(n28501), .C(
        n28500), .Y(n28504) );
  A2O1A1Ixp33_ASAP7_75t_SL U38793 ( .A1(u0_0_leon3x0_p0_dci[27]), .A2(n22398), 
        .B(n28504), .C(n30007), .Y(n28505) );
  A2O1A1Ixp33_ASAP7_75t_SL U38794 ( .A1(u0_0_leon3x0_p0_divi[21]), .A2(n22410), 
        .B(n28517), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[22]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38795 ( .A1(u0_0_leon3x0_p0_divi[19]), .A2(n22410), 
        .B(n28524), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38796 ( .A1(n28534), .A2(n28802), .B(n28533), .C(
        n28532), .Y(n2540) );
  A2O1A1Ixp33_ASAP7_75t_SL U38797 ( .A1(u0_0_leon3x0_p0_divi[18]), .A2(n22410), 
        .B(n28535), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[19]) );
  OA21x2_ASAP7_75t_SL U38798 ( .A1(n30645), .A2(n31823), .B(n28541), .Y(n28544) );
  A2O1A1Ixp33_ASAP7_75t_SL U38799 ( .A1(n31821), .A2(n28543), .B(n28542), .C(
        n28544), .Y(n28548) );
  A2O1A1Ixp33_ASAP7_75t_SL U38800 ( .A1(n28546), .A2(n22432), .B(n28545), .C(
        n28799), .Y(n28547) );
  OAI211xp5_ASAP7_75t_SL U38801 ( .A1(n24681), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP2__18_), .B(n28548), .C(n28547), .Y(n4002)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U38802 ( .A1(u0_0_leon3x0_p0_divi[17]), .A2(n22410), 
        .B(n28549), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38803 ( .A1(u0_0_leon3x0_p0_divi[16]), .A2(n22410), 
        .B(n28550), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38804 ( .A1(n28560), .A2(n28802), .B(n28559), .C(
        n28558), .Y(n2612) );
  A2O1A1Ixp33_ASAP7_75t_SL U38805 ( .A1(u0_0_leon3x0_p0_divi[15]), .A2(n22410), 
        .B(n28561), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[16]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38806 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_15_), .A2(
        n31833), .B(n28570), .C(n28569), .Y(n3228) );
  A2O1A1Ixp33_ASAP7_75t_SL U38807 ( .A1(n28581), .A2(n28802), .B(n28580), .C(
        n28579), .Y(n3982) );
  A2O1A1Ixp33_ASAP7_75t_SL U38808 ( .A1(u0_0_leon3x0_p0_divi[14]), .A2(n22410), 
        .B(n28582), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38809 ( .A1(u0_0_leon3x0_p0_divi[13]), .A2(n22410), 
        .B(n28587), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[14]) );
  AO21x1_ASAP7_75t_SL U38810 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5477), .B(
        n28591), .Y(n28592) );
  NAND3xp33_ASAP7_75t_SL U38811 ( .A(n28600), .B(n28599), .C(n28598), .Y(
        rf_di_w[13]) );
  NAND4xp25_ASAP7_75t_SL U38812 ( .A(n28606), .B(n28605), .C(n28604), .D(
        n28603), .Y(n28607) );
  A2O1A1Ixp33_ASAP7_75t_SL U38813 ( .A1(n28611), .A2(n28802), .B(n28610), .C(
        n28609), .Y(n2636) );
  A2O1A1Ixp33_ASAP7_75t_SL U38814 ( .A1(u0_0_leon3x0_p0_divi[12]), .A2(n22410), 
        .B(n28612), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[13]) );
  OAI211xp5_ASAP7_75t_SL U38815 ( .A1(n28667), .A2(n28618), .B(n28617), .C(
        n28616), .Y(n28647) );
  OA21x2_ASAP7_75t_SL U38816 ( .A1(n28769), .A2(n18316), .B(n28624), .Y(
        u0_0_leon3x0_p0_divi[11]) );
  O2A1O1Ixp5_ASAP7_75t_SL U38817 ( .A1(n28630), .A2(n28629), .B(n28628), .C(
        n28627), .Y(n30380) );
  AO21x1_ASAP7_75t_SL U38818 ( .A1(u0_0_leon3x0_p0_iu_r_E__JMPL_), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__12_), .B(n22375), .Y(n28634) );
  OAI211xp5_ASAP7_75t_SL U38819 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__12_), 
        .A2(n28637), .B(n28636), .C(n28635), .Y(n28638) );
  A2O1A1Ixp33_ASAP7_75t_SL U38820 ( .A1(n28642), .A2(n28641), .B(n24427), .C(
        n28640), .Y(n28644) );
  A2O1A1Ixp33_ASAP7_75t_SL U38821 ( .A1(u0_0_leon3x0_p0_dci[17]), .A2(n22398), 
        .B(n28644), .C(n28643), .Y(n28645) );
  OAI222xp33_ASAP7_75t_SL U38822 ( .A1(n22373), .A2(n29098), .B1(n32622), .B2(
        n18805), .C1(n28648), .C2(n22374), .Y(n29846) );
  OAI211xp5_ASAP7_75t_SL U38823 ( .A1(n29865), .A2(n29831), .B(n28650), .C(
        n28649), .Y(n28651) );
  A2O1A1Ixp33_ASAP7_75t_SL U38824 ( .A1(n28809), .A2(n28656), .B(n28655), .C(
        n28654), .Y(n2660) );
  A2O1A1Ixp33_ASAP7_75t_SL U38825 ( .A1(u0_0_leon3x0_p0_divi[11]), .A2(n22410), 
        .B(n28657), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[12]) );
  AO21x1_ASAP7_75t_SL U38826 ( .A1(n31830), .A2(u0_0_leon3x0_p0_iu_N5475), .B(
        n28660), .Y(n28661) );
  NAND3xp33_ASAP7_75t_SL U38827 ( .A(n28665), .B(n28664), .C(n28663), .Y(
        rf_di_w[11]) );
  O2A1O1Ixp5_ASAP7_75t_SL U38828 ( .A1(n28684), .A2(n28683), .B(n28682), .C(
        n28681), .Y(n30384) );
  NAND4xp25_ASAP7_75t_SL U38829 ( .A(n28688), .B(n28687), .C(n28686), .D(
        n28685), .Y(n28689) );
  A2O1A1Ixp33_ASAP7_75t_SL U38830 ( .A1(u0_0_leon3x0_p0_dci[16]), .A2(n22398), 
        .B(n28694), .C(n28693), .Y(n28695) );
  A2O1A1Ixp33_ASAP7_75t_SL U38831 ( .A1(u0_0_leon3x0_p0_divi[10]), .A2(n22410), 
        .B(n28700), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[11]) );
  OAI222xp33_ASAP7_75t_SL U38832 ( .A1(n24495), .A2(DP_OP_1196_128_7433_n452), 
        .B1(n28701), .B2(u0_0_leon3x0_p0_iu_v_A__CTRL__INST__10_), .C1(
        u0_0_leon3x0_p0_iu_r_A__IMM__10_), .C2(n23229), .Y(n3472) );
  NAND3xp33_ASAP7_75t_SL U38833 ( .A(n28712), .B(n28711), .C(n28710), .Y(
        rf_di_w[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38834 ( .A1(u0_0_leon3x0_p0_divi[9]), .A2(n22410), 
        .B(n28716), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38835 ( .A1(n18890), .A2(n22410), .B(n28717), .C(
        n24629), .Y(u0_0_leon3x0_p0_div0_b[9]) );
  OAI211xp5_ASAP7_75t_SL U38836 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__8_), .A2(
        n30813), .B(n28760), .C(n24523), .Y(n3660) );
  A2O1A1Ixp33_ASAP7_75t_SL U38837 ( .A1(n18904), .A2(n28827), .B(n28721), .C(
        n28725), .Y(n28724) );
  OAI211xp5_ASAP7_75t_SL U38838 ( .A1(n28734), .A2(n30393), .B(n28733), .C(
        n28732), .Y(n28735) );
  A2O1A1Ixp33_ASAP7_75t_SL U38839 ( .A1(n28737), .A2(n28736), .B(n28735), .C(
        n24634), .Y(n28738) );
  OAI211xp5_ASAP7_75t_SL U38840 ( .A1(n30396), .A2(n30625), .B(n28739), .C(
        n28738), .Y(n28740) );
  OAI211xp5_ASAP7_75t_SL U38841 ( .A1(n28745), .A2(n28790), .B(n28744), .C(
        n28743), .Y(n28746) );
  A2O1A1Ixp33_ASAP7_75t_SL U38842 ( .A1(n18887), .A2(n22398), .B(n28746), .C(
        n30007), .Y(n28747) );
  A2O1A1Ixp33_ASAP7_75t_SL U38843 ( .A1(n28757), .A2(n28802), .B(n28756), .C(
        n28755), .Y(n2319) );
  A2O1A1Ixp33_ASAP7_75t_SL U38844 ( .A1(n18904), .A2(n22410), .B(n28758), .C(
        n24629), .Y(u0_0_leon3x0_p0_div0_b[8]) );
  OAI211xp5_ASAP7_75t_SL U38845 ( .A1(u0_0_leon3x0_p0_iu_r_A__IMM__7_), .A2(
        n30813), .B(n28760), .C(n30877), .Y(n3669) );
  A2O1A1Ixp33_ASAP7_75t_SL U38846 ( .A1(n28778), .A2(n28777), .B(n28776), .C(
        n28775), .Y(n30406) );
  OAI211xp5_ASAP7_75t_SL U38847 ( .A1(n29595), .A2(n30402), .B(n28781), .C(
        n28780), .Y(n28787) );
  OAI211xp5_ASAP7_75t_SL U38848 ( .A1(n29910), .A2(n28785), .B(n28784), .C(
        n28783), .Y(n28786) );
  A2O1A1Ixp33_ASAP7_75t_SL U38849 ( .A1(u0_0_leon3x0_p0_dci[12]), .A2(n22398), 
        .B(n28792), .C(n28791), .Y(n28793) );
  A2O1A1Ixp33_ASAP7_75t_SL U38850 ( .A1(n28803), .A2(n28802), .B(n28801), .C(
        n28800), .Y(n3926) );
  A2O1A1Ixp33_ASAP7_75t_SL U38851 ( .A1(u0_0_leon3x0_p0_divi[6]), .A2(n22410), 
        .B(n28804), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38852 ( .A1(u0_0_leon3x0_p0_divi[5]), .A2(n22410), 
        .B(n28810), .C(n29018), .Y(u0_0_leon3x0_p0_div0_b[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38853 ( .A1(u0_0_leon3x0_p0_divi[4]), .A2(n22410), 
        .B(n28819), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38854 ( .A1(u0_0_leon3x0_p0_divi[3]), .A2(n28827), 
        .B(n28826), .C(n28829), .Y(n28828) );
  A2O1A1Ixp33_ASAP7_75t_SL U38855 ( .A1(n28830), .A2(u0_0_leon3x0_p0_divi[3]), 
        .B(n28829), .C(n28828), .Y(n28831) );
  A2O1A1Ixp33_ASAP7_75t_SL U38856 ( .A1(n24579), .A2(u0_0_leon3x0_p0_divi[3]), 
        .B(n28832), .C(n28831), .Y(n30438) );
  OAI211xp5_ASAP7_75t_SL U38857 ( .A1(n29594), .A2(n30441), .B(n28837), .C(
        n28836), .Y(n28838) );
  A2O1A1Ixp33_ASAP7_75t_SL U38858 ( .A1(n24485), .A2(n28840), .B(n24427), .C(
        n28839), .Y(n28842) );
  OAI211xp5_ASAP7_75t_SL U38859 ( .A1(n28858), .A2(n28914), .B(n28857), .C(
        n28856), .Y(n28859) );
  OAI222xp33_ASAP7_75t_SL U38860 ( .A1(n29104), .A2(n22373), .B1(n32606), .B2(
        n18805), .C1(n28860), .C2(n22374), .Y(n29623) );
  OAI211xp5_ASAP7_75t_SL U38861 ( .A1(n29865), .A2(n29499), .B(n28862), .C(
        n28861), .Y(n28863) );
  AO21x1_ASAP7_75t_SL U38862 ( .A1(n31868), .A2(n29623), .B(n28863), .Y(n28864) );
  A2O1A1Ixp33_ASAP7_75t_SL U38863 ( .A1(u0_0_leon3x0_p0_divi[3]), .A2(n22410), 
        .B(n28867), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38864 ( .A1(n28992), .A2(n30631), .B(n28874), .C(
        n28968), .Y(n28900) );
  A2O1A1Ixp33_ASAP7_75t_SL U38865 ( .A1(n28992), .A2(n28876), .B(n28875), .C(
        n28987), .Y(n28899) );
  OR2x2_ASAP7_75t_SL U38866 ( .A(n22256), .B(n28880), .Y(
        u0_0_leon3x0_p0_divi[2]) );
  O2A1O1Ixp5_ASAP7_75t_SL U38867 ( .A1(n28886), .A2(n28885), .B(n28884), .C(
        n28883), .Y(n30449) );
  A2O1A1Ixp33_ASAP7_75t_SL U38868 ( .A1(n28900), .A2(n28899), .B(n28898), .C(
        n28897), .Y(n28901) );
  OAI222xp33_ASAP7_75t_SL U38869 ( .A1(n29105), .A2(n22373), .B1(n32604), .B2(
        n18805), .C1(n28903), .C2(n22374), .Y(n29887) );
  A2O1A1Ixp33_ASAP7_75t_SL U38870 ( .A1(u0_0_leon3x0_p0_divi[2]), .A2(n22410), 
        .B(n28907), .C(n29018), .Y(u0_0_leon3x0_p0_div0_b[3]) );
  NAND4xp25_ASAP7_75t_SL U38871 ( .A(n32667), .B(n24681), .C(n32666), .D(
        n32665), .Y(n28909) );
  NAND3xp33_ASAP7_75t_SL U38872 ( .A(n28912), .B(n28911), .C(n28910), .Y(
        rf_di_w[2]) );
  OR2x2_ASAP7_75t_SL U38873 ( .A(n28926), .B(n30604), .Y(
        u0_0_leon3x0_p0_divi[1]) );
  NAND3xp33_ASAP7_75t_SL U38874 ( .A(n28927), .B(n24579), .C(
        u0_0_leon3x0_p0_divi[1]), .Y(n28933) );
  A2O1A1Ixp33_ASAP7_75t_SL U38875 ( .A1(n29561), .A2(n28931), .B(n28930), .C(
        n28929), .Y(n28932) );
  NAND3xp33_ASAP7_75t_SL U38876 ( .A(n28938), .B(n28937), .C(n28936), .Y(
        n28939) );
  A2O1A1Ixp33_ASAP7_75t_SL U38877 ( .A1(n30620), .A2(n29564), .B(n28939), .C(
        n24634), .Y(n28945) );
  AO21x1_ASAP7_75t_SL U38878 ( .A1(u0_0_leon3x0_p0_iu_r_E__JMPL_), .A2(
        u0_0_leon3x0_p0_iu_v_M__CTRL__PC__2_), .B(n22375), .Y(n28942) );
  OAI211xp5_ASAP7_75t_SL U38879 ( .A1(n30451), .A2(n30625), .B(n28945), .C(
        n28944), .Y(n28948) );
  A2O1A1Ixp33_ASAP7_75t_SL U38880 ( .A1(n32438), .A2(n22398), .B(n28948), .C(
        n28947), .Y(n28949) );
  A2O1A1Ixp33_ASAP7_75t_SL U38881 ( .A1(u0_0_leon3x0_p0_divi[1]), .A2(n22410), 
        .B(n28959), .C(n24629), .Y(u0_0_leon3x0_p0_div0_b[2]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38882 ( .A1(n18908), .A2(n22410), .B(n28960), .C(
        n24629), .Y(u0_0_leon3x0_p0_div0_b[1]) );
  OAI211xp5_ASAP7_75t_SL U38883 ( .A1(n22216), .A2(n28970), .B(n28969), .C(
        n28968), .Y(n28973) );
  A2O1A1Ixp33_ASAP7_75t_SL U38884 ( .A1(n28975), .A2(n28974), .B(n28973), .C(
        n28972), .Y(n30634) );
  OAI211xp5_ASAP7_75t_SL U38885 ( .A1(n28986), .A2(n28985), .B(n28984), .C(
        n28983), .Y(n28989) );
  A2O1A1Ixp33_ASAP7_75t_SL U38886 ( .A1(n30634), .A2(n28992), .B(n28991), .C(
        u0_0_leon3x0_p0_iu_r_E__ALUSEL__0_), .Y(n28993) );
  NAND4xp25_ASAP7_75t_SL U38887 ( .A(n28999), .B(n28998), .C(n28997), .D(
        n28996), .Y(n29002) );
  A2O1A1Ixp33_ASAP7_75t_SL U38888 ( .A1(n30620), .A2(n29003), .B(n29002), .C(
        n29001), .Y(n29005) );
  O2A1O1Ixp5_ASAP7_75t_SL U38889 ( .A1(n29007), .A2(n29006), .B(n29005), .C(
        n29004), .Y(n29008) );
  OAI222xp33_ASAP7_75t_SL U38890 ( .A1(n29011), .A2(n22374), .B1(n32713), .B2(
        n18806), .C1(n22373), .C2(n29107), .Y(n31424) );
  A2O1A1Ixp33_ASAP7_75t_SL U38891 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_29_), .A2(
        n31833), .B(n29030), .C(n29029), .Y(n3292) );
  AO21x1_ASAP7_75t_SL U38892 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5487), .B(
        n29064), .Y(n29065) );
  NAND3xp33_ASAP7_75t_SL U38893 ( .A(n29070), .B(n29069), .C(n29068), .Y(
        rf_di_w[23]) );
  OAI211xp5_ASAP7_75t_SL U38894 ( .A1(n31340), .A2(n29081), .B(n29076), .C(
        n29075), .Y(n29077) );
  NAND3xp33_ASAP7_75t_SL U38895 ( .A(n29113), .B(n31676), .C(n31653), .Y(
        n29117) );
  NAND4xp25_ASAP7_75t_SL U38896 ( .A(n29121), .B(n29120), .C(n29119), .D(
        n29118), .Y(n29127) );
  NAND4xp25_ASAP7_75t_SL U38897 ( .A(n29125), .B(n29124), .C(n29123), .D(
        n29122), .Y(n29126) );
  NOR3xp33_ASAP7_75t_SL U38898 ( .A(n22373), .B(n29127), .C(n29126), .Y(n29129) );
  A2O1A1Ixp33_ASAP7_75t_SL U38899 ( .A1(u0_0_leon3x0_p0_divo[32]), .A2(n24491), 
        .B(n29129), .C(u0_0_leon3x0_p0_iu_v_X__CTRL__INST__23_), .Y(n29130) );
  NAND4xp25_ASAP7_75t_SL U38900 ( .A(n29137), .B(
        u0_0_leon3x0_p0_iu_r_E__ALUSEL__1_), .C(n29136), .D(n29135), .Y(n29138) );
  NOR3xp33_ASAP7_75t_SL U38901 ( .A(n30438), .B(n30449), .C(n29138), .Y(n29139) );
  NAND4xp25_ASAP7_75t_SL U38902 ( .A(n29140), .B(n30241), .C(n30386), .D(
        n29139), .Y(n29142) );
  NAND4xp25_ASAP7_75t_SL U38903 ( .A(n30304), .B(n30307), .C(n30396), .D(
        n30389), .Y(n29141) );
  NOR3xp33_ASAP7_75t_SL U38904 ( .A(n29142), .B(n30369), .C(n29141), .Y(n29164) );
  NAND4xp25_ASAP7_75t_SL U38905 ( .A(n30425), .B(n29153), .C(n30384), .D(
        n30214), .Y(n29160) );
  NAND3xp33_ASAP7_75t_SL U38906 ( .A(n30626), .B(n30451), .C(n29155), .Y(
        n29156) );
  NOR3xp33_ASAP7_75t_SL U38907 ( .A(n29157), .B(n29156), .C(n30276), .Y(n29158) );
  NAND3xp33_ASAP7_75t_SL U38908 ( .A(n29158), .B(n30225), .C(n30237), .Y(
        n29159) );
  NAND4xp25_ASAP7_75t_SL U38909 ( .A(n29164), .B(n29163), .C(n29162), .D(
        n29161), .Y(n29868) );
  A2O1A1Ixp33_ASAP7_75t_SL U38910 ( .A1(n29176), .A2(n30666), .B(n29175), .C(
        n29174), .Y(n4579) );
  OR2x2_ASAP7_75t_SL U38911 ( .A(n29195), .B(n29202), .Y(n29199) );
  A2O1A1Ixp33_ASAP7_75t_SL U38912 ( .A1(n29624), .A2(n29195), .B(n29194), .C(
        n29202), .Y(n29201) );
  NAND3xp33_ASAP7_75t_SL U38913 ( .A(n32153), .B(n24681), .C(
        u0_0_leon3x0_p0_iu_r_W__S__PS_), .Y(n29208) );
  NAND3xp33_ASAP7_75t_SL U38914 ( .A(n29218), .B(n32075), .C(n29694), .Y(
        n29221) );
  AO21x1_ASAP7_75t_SL U38915 ( .A1(n29230), .A2(n29229), .B(n29228), .Y(n3342)
         );
  OR2x2_ASAP7_75t_SL U38916 ( .A(irqo[0]), .B(n29239), .Y(n29653) );
  A2O1A1Ixp33_ASAP7_75t_SL U38917 ( .A1(irqctrl0_r_IFORCE__0__12_), .A2(n29242), .B(n29241), .C(n29240), .Y(n1778) );
  A2O1A1Ixp33_ASAP7_75t_SL U38918 ( .A1(apbi[12]), .A2(n29745), .B(n29247), 
        .C(n29246), .Y(n1777) );
  A2O1A1Ixp33_ASAP7_75t_SL U38919 ( .A1(irqctrl0_r_IFORCE__0__9_), .A2(n29253), 
        .B(n29252), .C(n29254), .Y(n1798) );
  NOR3xp33_ASAP7_75t_SL U38920 ( .A(n29376), .B(n24695), .C(n30139), .Y(n29257) );
  A2O1A1Ixp33_ASAP7_75t_SL U38921 ( .A1(n29258), .A2(n29325), .B(n29257), .C(
        n29256), .Y(n1797) );
  A2O1A1Ixp33_ASAP7_75t_SL U38922 ( .A1(irqctrl0_r_IFORCE__0__10_), .A2(n29264), .B(n29263), .C(n29262), .Y(n2385) );
  A2O1A1Ixp33_ASAP7_75t_SL U38923 ( .A1(n30978), .A2(n29325), .B(n29269), .C(
        n29268), .Y(n2384) );
  A2O1A1Ixp33_ASAP7_75t_SL U38924 ( .A1(n29278), .A2(n29277), .B(n29276), .C(
        n29742), .Y(n1745) );
  A2O1A1Ixp33_ASAP7_75t_SL U38925 ( .A1(irqctrl0_r_IFORCE__0__7_), .A2(n29281), 
        .B(n29280), .C(n29282), .Y(n2698) );
  A2O1A1Ixp33_ASAP7_75t_SL U38926 ( .A1(n30833), .A2(n29325), .B(n29286), .C(
        n29285), .Y(n2695) );
  A2O1A1Ixp33_ASAP7_75t_SL U38927 ( .A1(irqctrl0_r_IFORCE__0__5_), .A2(n29297), 
        .B(n29296), .C(n29295), .Y(n2699) );
  A2O1A1Ixp33_ASAP7_75t_SL U38928 ( .A1(n30073), .A2(n29325), .B(n29302), .C(
        n29301), .Y(n2696) );
  A2O1A1Ixp33_ASAP7_75t_SL U38929 ( .A1(n29310), .A2(n31641), .B(n29309), .C(
        n29308), .Y(n1733) );
  A2O1A1Ixp33_ASAP7_75t_SL U38930 ( .A1(n31197), .A2(n29325), .B(n29315), .C(
        n29314), .Y(n1732) );
  A2O1A1Ixp33_ASAP7_75t_SL U38931 ( .A1(irqctrl0_r_IFORCE__0__4_), .A2(n29319), 
        .B(n29318), .C(n29317), .Y(n2693) );
  A2O1A1Ixp33_ASAP7_75t_SL U38932 ( .A1(n30780), .A2(n29325), .B(n29324), .C(
        n29323), .Y(n2692) );
  A2O1A1Ixp33_ASAP7_75t_SL U38933 ( .A1(irqctrl0_r_IFORCE__0__2_), .A2(n29332), 
        .B(n29331), .C(n29330), .Y(n2694) );
  NAND3xp33_ASAP7_75t_SL U38934 ( .A(n29338), .B(uart1_r_IRQCNT__1_), .C(
        uart1_r_IRQCNT__2_), .Y(n29341) );
  A2O1A1Ixp33_ASAP7_75t_SL U38935 ( .A1(uart1_r_IRQCNT__1_), .A2(n29338), .B(
        uart1_r_IRQCNT__2_), .C(n29341), .Y(n29339) );
  OR2x2_ASAP7_75t_SL U38936 ( .A(n29339), .B(n29342), .Y(n1762) );
  AND2x2_ASAP7_75t_SL U38937 ( .A(uart1_r_IRQCNT__5_), .B(uart1_r_IRQCNT__4_), 
        .Y(n29359) );
  A2O1A1Ixp33_ASAP7_75t_SL U38938 ( .A1(uart1_r_IRQCNT__4_), .A2(n29344), .B(
        uart1_r_IRQCNT__5_), .C(n29343), .Y(n1759) );
  NAND3xp33_ASAP7_75t_SL U38939 ( .A(n29746), .B(uart1_r_RFIFOIRQEN_), .C(
        uart1_uarto_RXEN_), .Y(n29362) );
  A2O1A1Ixp33_ASAP7_75t_SL U38940 ( .A1(n29350), .A2(n29349), .B(n29348), .C(
        n29362), .Y(n1758) );
  NOR3xp33_ASAP7_75t_SL U38941 ( .A(n29357), .B(n29356), .C(n29355), .Y(n29373) );
  NAND3xp33_ASAP7_75t_SL U38942 ( .A(n29358), .B(uart1_r_RIRQEN_), .C(n33068), 
        .Y(n29371) );
  NAND3xp33_ASAP7_75t_SL U38943 ( .A(n29364), .B(n29363), .C(n29362), .Y(
        n29365) );
  A2O1A1Ixp33_ASAP7_75t_SL U38944 ( .A1(n29371), .A2(n29370), .B(n29369), .C(
        n29368), .Y(n29372) );
  A2O1A1Ixp33_ASAP7_75t_SL U38945 ( .A1(n29382), .A2(n29381), .B(
        apbo_1__PIRQ__2_), .C(n29380), .Y(n1756) );
  A2O1A1Ixp33_ASAP7_75t_SL U38946 ( .A1(irqctrl0_r_IFORCE__0__15_), .A2(n29393), .B(n29392), .C(n29394), .Y(n2691) );
  A2O1A1Ixp33_ASAP7_75t_SL U38947 ( .A1(apbi[15]), .A2(n29657), .B(n29398), 
        .C(n29397), .Y(n2690) );
  OA21x2_ASAP7_75t_SL U38948 ( .A1(irqctrl0_r_IPEND__1_), .A2(
        irqctrl0_r_IFORCE__0__1_), .B(irqctrl0_r_IMASK__0__1_), .Y(n29443) );
  OR2x2_ASAP7_75t_SL U38949 ( .A(irqctrl0_r_IPEND__2_), .B(
        irqctrl0_r_IFORCE__0__2_), .Y(n29417) );
  OR2x2_ASAP7_75t_SL U38950 ( .A(n29407), .B(n29414), .Y(n29659) );
  OR2x2_ASAP7_75t_SL U38951 ( .A(irqctrl0_r_IPEND__8_), .B(
        irqctrl0_r_IFORCE__0__8_), .Y(n29431) );
  NAND3xp33_ASAP7_75t_SL U38952 ( .A(n29423), .B(n29448), .C(n29445), .Y(
        n29450) );
  O2A1O1Ixp5_ASAP7_75t_SL U38953 ( .A1(n29441), .A2(n29440), .B(n29442), .C(
        n29439), .Y(n29666) );
  NAND3xp33_ASAP7_75t_SL U38954 ( .A(n29666), .B(n29634), .C(n29442), .Y(
        n29627) );
  A2O1A1Ixp33_ASAP7_75t_SL U38955 ( .A1(n29455), .A2(n29454), .B(n29453), .C(
        n29877), .Y(n29466) );
  A2O1A1Ixp33_ASAP7_75t_SL U38956 ( .A1(n29466), .A2(n29465), .B(n29633), .C(
        n29464), .Y(n29628) );
  OAI211xp5_ASAP7_75t_SL U38957 ( .A1(n24585), .A2(n29481), .B(n29478), .C(
        n29477), .Y(n29479) );
  AO21x1_ASAP7_75t_SL U38958 ( .A1(n23229), .A2(n32692), .B(n29480), .Y(n4731)
         );
  NAND3xp33_ASAP7_75t_SL U38959 ( .A(n29485), .B(n29484), .C(n29483), .Y(
        rf_di_w[4]) );
  NAND3xp33_ASAP7_75t_SL U38960 ( .A(n29493), .B(n29492), .C(n29491), .Y(
        rf_di_w[3]) );
  A2O1A1Ixp33_ASAP7_75t_SL U38961 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[7]), .B(n29509), .C(n31638), .Y(n4691) );
  OR2x2_ASAP7_75t_SL U38962 ( .A(n29568), .B(n31057), .Y(n29556) );
  A2O1A1Ixp33_ASAP7_75t_SL U38963 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[6]), .B(n29569), .C(n31638), .Y(n4671) );
  NAND3xp33_ASAP7_75t_SL U38964 ( .A(n29582), .B(n29581), .C(n29580), .Y(
        rf_di_w[29]) );
  OAI211xp5_ASAP7_75t_SL U38965 ( .A1(n29593), .A2(n29592), .B(n29591), .C(
        n29590), .Y(n29597) );
  OAI211xp5_ASAP7_75t_SL U38966 ( .A1(n29609), .A2(n29608), .B(n29607), .C(
        n29606), .Y(n29610) );
  A2O1A1Ixp33_ASAP7_75t_SL U38967 ( .A1(u0_0_leon3x0_p0_dci[35]), .A2(n22398), 
        .B(n29610), .C(n30007), .Y(n29611) );
  OR2x2_ASAP7_75t_SL U38968 ( .A(n31396), .B(n29613), .Y(n30599) );
  NAND3xp33_ASAP7_75t_SL U38969 ( .A(n29618), .B(n31054), .C(n29617), .Y(
        n29621) );
  OAI211xp5_ASAP7_75t_SL U38970 ( .A1(n29622), .A2(n29843), .B(n29621), .C(
        n29620), .Y(n3969) );
  O2A1O1Ixp5_ASAP7_75t_SL U38971 ( .A1(n29662), .A2(n29661), .B(n29664), .C(
        n29633), .Y(n29878) );
  OAI321xp33_ASAP7_75t_SL U38972 ( .A1(n29637), .A2(n29879), .A3(n29636), .B1(
        n29635), .B2(n29634), .C(n29878), .Y(irqctrl0_v_IRL__0__2_) );
  O2A1O1Ixp5_ASAP7_75t_SL U38973 ( .A1(n29673), .A2(n31443), .B(n29672), .C(
        n29671), .Y(n3358) );
  AO21x1_ASAP7_75t_SL U38974 ( .A1(n31830), .A2(u0_0_leon3x0_p0_iu_N5469), .B(
        n29678), .Y(n29679) );
  NAND3xp33_ASAP7_75t_SL U38975 ( .A(n29683), .B(n29682), .C(n29681), .Y(
        rf_di_w[5]) );
  NAND3xp33_ASAP7_75t_SL U38976 ( .A(n29686), .B(n31054), .C(n29685), .Y(
        n29690) );
  NAND3xp33_ASAP7_75t_SL U38977 ( .A(n29688), .B(n31542), .C(n29687), .Y(
        n29689) );
  OAI211xp5_ASAP7_75t_SL U38978 ( .A1(n24681), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__4_), .B(n29690), .C(n29689), .Y(n2731) );
  A2O1A1Ixp33_ASAP7_75t_SL U38979 ( .A1(n29725), .A2(n29724), .B(n29723), .C(
        n29722), .Y(n30703) );
  NAND3xp33_ASAP7_75t_SL U38980 ( .A(n30708), .B(u0_0_leon3x0_p0_iu_r_M__DIVZ_), .C(n24491), .Y(n29885) );
  A2O1A1Ixp33_ASAP7_75t_SL U38981 ( .A1(n29755), .A2(n29754), .B(
        apb0_r_CFGSEL_), .C(n29753), .Y(n29756) );
  AO21x1_ASAP7_75t_SL U38982 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5488), .B(
        n29771), .Y(n29772) );
  NAND3xp33_ASAP7_75t_SL U38983 ( .A(n29781), .B(n29780), .C(n29779), .Y(
        rf_di_w[24]) );
  O2A1O1Ixp5_ASAP7_75t_SL U38984 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), 
        .A2(n29812), .B(n29811), .C(n30667), .Y(n29813) );
  A2O1A1Ixp33_ASAP7_75t_SL U38985 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_12_), .A2(
        n31833), .B(n29824), .C(n29823), .Y(n2677) );
  NAND3xp33_ASAP7_75t_SL U38986 ( .A(n29835), .B(n29834), .C(n29833), .Y(
        rf_di_w[12]) );
  OAI211xp5_ASAP7_75t_SL U38987 ( .A1(n31340), .A2(n30381), .B(n29839), .C(
        n29838), .Y(n29840) );
  A2O1A1Ixp33_ASAP7_75t_SL U38988 ( .A1(n29856), .A2(n29855), .B(
        apb0_r_CFGSEL_), .C(n29854), .Y(n29857) );
  OAI211xp5_ASAP7_75t_SL U38989 ( .A1(n29870), .A2(n29869), .B(n24681), .C(
        n29868), .Y(n29871) );
  NAND4xp25_ASAP7_75t_SL U38990 ( .A(n29874), .B(u0_0_leon3x0_p0_iu_r_A__TICC_), .C(n29873), .D(n29872), .Y(n29876) );
  OAI211xp5_ASAP7_75t_SL U38991 ( .A1(n29880), .A2(n29879), .B(n29878), .C(
        n29877), .Y(irqctrl0_v_IRL__0__3_) );
  NAND3xp33_ASAP7_75t_SL U38992 ( .A(n29897), .B(n29896), .C(n29895), .Y(
        rf_di_w[7]) );
  OAI211xp5_ASAP7_75t_SL U38993 ( .A1(n31340), .A2(n29907), .B(n29901), .C(
        n29900), .Y(n29902) );
  AO21x1_ASAP7_75t_SL U38994 ( .A1(n30016), .A2(n29912), .B(n31364), .Y(n29923) );
  O2A1O1Ixp5_ASAP7_75t_SL U38995 ( .A1(u0_0_leon3x0_p0_iu_r_X__DATA__0__7_), 
        .A2(n30575), .B(n29923), .C(n29922), .Y(n3033) );
  OR2x2_ASAP7_75t_SL U38996 ( .A(n31340), .B(n29932), .Y(n30731) );
  NAND3xp33_ASAP7_75t_SL U38997 ( .A(n30732), .B(n31054), .C(n30731), .Y(
        n29933) );
  O2A1O1Ixp5_ASAP7_75t_SL U38998 ( .A1(n29939), .A2(n29938), .B(n29937), .C(
        n29936), .Y(n29940) );
  A2O1A1Ixp33_ASAP7_75t_SL U38999 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[11]), .B(n29942), .C(n31638), .Y(n4776) );
  NAND3xp33_ASAP7_75t_SL U39000 ( .A(n29961), .B(n24694), .C(
        uart1_r_RSHIFT__0_), .Y(n29962) );
  A2O1A1Ixp33_ASAP7_75t_SL U39001 ( .A1(n29987), .A2(n29986), .B(n29985), .C(
        n29984), .Y(n2458) );
  NAND3xp33_ASAP7_75t_SL U39002 ( .A(n30020), .B(
        u0_0_leon3x0_p0_iu_v_X__CTRL__LD_), .C(n31694), .Y(n30019) );
  A2O1A1Ixp33_ASAP7_75t_SL U39003 ( .A1(n22397), .A2(
        u0_0_leon3x0_p0_c0mmu_mcdi[9]), .B(n30029), .C(n31638), .Y(n4743) );
  OR2x2_ASAP7_75t_SL U39004 ( .A(n30073), .B(n31057), .Y(n30063) );
  A2O1A1Ixp33_ASAP7_75t_SL U39005 ( .A1(n30071), .A2(n30070), .B(n30069), .C(
        n30068), .Y(n1748) );
  OAI211xp5_ASAP7_75t_SL U39006 ( .A1(n30872), .A2(n30077), .B(n30076), .C(
        n30075), .Y(n30112) );
  NAND3xp33_ASAP7_75t_SL U39007 ( .A(n30080), .B(n30079), .C(n30078), .Y(
        n30104) );
  NAND3xp33_ASAP7_75t_SL U39008 ( .A(n30083), .B(n30082), .C(n30081), .Y(
        n30089) );
  NAND4xp25_ASAP7_75t_SL U39009 ( .A(n30087), .B(n30086), .C(n30085), .D(
        n30084), .Y(n30088) );
  NAND4xp25_ASAP7_75t_SL U39010 ( .A(n30093), .B(n30092), .C(n30091), .D(
        n30090), .Y(n30099) );
  NAND4xp25_ASAP7_75t_SL U39011 ( .A(n30097), .B(n30096), .C(n30095), .D(
        n30094), .Y(n30098) );
  A2O1A1Ixp33_ASAP7_75t_SL U39012 ( .A1(n30102), .A2(n30101), .B(n31238), .C(
        n30100), .Y(n30103) );
  A2O1A1Ixp33_ASAP7_75t_SL U39013 ( .A1(n30123), .A2(n23229), .B(n30122), .C(
        n30121), .Y(n3364) );
  A2O1A1Ixp33_ASAP7_75t_SL U39014 ( .A1(apbi[9]), .A2(n30136), .B(n30135), .C(
        n24694), .Y(n1794) );
  NAND3xp33_ASAP7_75t_SL U39015 ( .A(n30144), .B(n30143), .C(n30142), .Y(
        n30149) );
  OAI211xp5_ASAP7_75t_SL U39016 ( .A1(n31236), .A2(n30147), .B(n30146), .C(
        n30145), .Y(n30148) );
  OR2x2_ASAP7_75t_SL U39017 ( .A(n3055), .B(n22380), .Y(n30180) );
  A2O1A1Ixp33_ASAP7_75t_SL U39018 ( .A1(n30163), .A2(n30165), .B(n23882), .C(
        n30177), .Y(n3051) );
  O2A1O1Ixp5_ASAP7_75t_SL U39019 ( .A1(n30170), .A2(n30169), .B(n30168), .C(
        n30167), .Y(n30171) );
  O2A1O1Ixp5_ASAP7_75t_SL U39020 ( .A1(n30175), .A2(n30180), .B(n30174), .C(
        n30173), .Y(n30176) );
  XOR2xp5_ASAP7_75t_SL U39021 ( .A(n30179), .B(
        u0_0_leon3x0_p0_c0mmu_dcache0_r_FADDR__5_), .Y(n30178) );
  OR2x2_ASAP7_75t_SL U39022 ( .A(n22380), .B(n18851), .Y(n30191) );
  NAND3xp33_ASAP7_75t_SL U39023 ( .A(n30189), .B(n30186), .C(n30185), .Y(
        n30187) );
  OR2x2_ASAP7_75t_SL U39024 ( .A(n30196), .B(n30195), .Y(n32194) );
  OR2x2_ASAP7_75t_SL U39025 ( .A(n32455), .B(n31306), .Y(n30206) );
  A2O1A1Ixp33_ASAP7_75t_SL U39026 ( .A1(n30223), .A2(n31415), .B(n30222), .C(
        n30221), .Y(n2760) );
  NAND3xp33_ASAP7_75t_SL U39027 ( .A(n30229), .B(n30228), .C(n30227), .Y(
        n30232) );
  A2O1A1Ixp33_ASAP7_75t_SL U39028 ( .A1(n30233), .A2(n31415), .B(n30232), .C(
        n30231), .Y(n1786) );
  OAI211xp5_ASAP7_75t_SL U39029 ( .A1(n24638), .A2(n30255), .B(n30254), .C(
        n30253), .Y(n30256) );
  AO21x1_ASAP7_75t_SL U39030 ( .A1(n30453), .A2(n30257), .B(n30256), .Y(n30260) );
  A2O1A1Ixp33_ASAP7_75t_SL U39031 ( .A1(n30261), .A2(n31415), .B(n30260), .C(
        n30259), .Y(n2488) );
  OAI211xp5_ASAP7_75t_SL U39032 ( .A1(n30270), .A2(n24514), .B(n30269), .C(
        n30268), .Y(n30271) );
  AO21x1_ASAP7_75t_SL U39033 ( .A1(n30453), .A2(n30272), .B(n30271), .Y(n30275) );
  A2O1A1Ixp33_ASAP7_75t_SL U39034 ( .A1(n30276), .A2(n31415), .B(n30275), .C(
        n30274), .Y(n2515) );
  A2O1A1Ixp33_ASAP7_75t_SL U39035 ( .A1(n30672), .A2(n31415), .B(n30284), .C(
        n30283), .Y(n4344) );
  A2O1A1Ixp33_ASAP7_75t_SL U39036 ( .A1(n30295), .A2(n31415), .B(n30294), .C(
        n30293), .Y(n4047) );
  OAI211xp5_ASAP7_75t_SL U39037 ( .A1(n24638), .A2(n30300), .B(n30299), .C(
        n30298), .Y(n30301) );
  A2O1A1Ixp33_ASAP7_75t_SL U39038 ( .A1(n30316), .A2(n31415), .B(n30315), .C(
        n30314), .Y(n3995) );
  OAI211xp5_ASAP7_75t_SL U39039 ( .A1(n30320), .A2(n24514), .B(n30319), .C(
        n30318), .Y(n30321) );
  AO21x1_ASAP7_75t_SL U39040 ( .A1(n30453), .A2(n30322), .B(n30321), .Y(n30325) );
  A2O1A1Ixp33_ASAP7_75t_SL U39041 ( .A1(n30326), .A2(n31415), .B(n30325), .C(
        n30324), .Y(n3993) );
  OAI211xp5_ASAP7_75t_SL U39042 ( .A1(n24638), .A2(n30331), .B(n30330), .C(
        n30329), .Y(n30332) );
  AO21x1_ASAP7_75t_SL U39043 ( .A1(n30453), .A2(n30333), .B(n30332), .Y(n30336) );
  A2O1A1Ixp33_ASAP7_75t_SL U39044 ( .A1(n30337), .A2(n31415), .B(n30336), .C(
        n30335), .Y(n3991) );
  A2O1A1Ixp33_ASAP7_75t_SL U39045 ( .A1(n30349), .A2(n31415), .B(n30348), .C(
        n30347), .Y(n3980) );
  OAI211xp5_ASAP7_75t_SL U39046 ( .A1(n24638), .A2(n30354), .B(n30353), .C(
        n30352), .Y(n30355) );
  AO21x1_ASAP7_75t_SL U39047 ( .A1(n30453), .A2(n30356), .B(n30355), .Y(n30359) );
  A2O1A1Ixp33_ASAP7_75t_SL U39048 ( .A1(n30360), .A2(n31415), .B(n30359), .C(
        n30358), .Y(n3978) );
  A2O1A1Ixp33_ASAP7_75t_SL U39049 ( .A1(n30369), .A2(n31415), .B(n30368), .C(
        n30367), .Y(n3976) );
  A2O1A1Ixp33_ASAP7_75t_SL U39050 ( .A1(n30380), .A2(n31415), .B(n30379), .C(
        n30378), .Y(n3974) );
  A2O1A1Ixp33_ASAP7_75t_SL U39051 ( .A1(n30406), .A2(n31415), .B(n30405), .C(
        n30404), .Y(n3924) );
  A2O1A1Ixp33_ASAP7_75t_SL U39052 ( .A1(n30416), .A2(n31415), .B(n30415), .C(
        n30414), .Y(n3922) );
  OAI211xp5_ASAP7_75t_SL U39053 ( .A1(n24638), .A2(n30421), .B(n30420), .C(
        n30419), .Y(n30422) );
  OAI211xp5_ASAP7_75t_SL U39054 ( .A1(n24638), .A2(n30433), .B(n30432), .C(
        n30431), .Y(n30434) );
  AO21x1_ASAP7_75t_SL U39055 ( .A1(n30453), .A2(n30435), .B(n30434), .Y(n30437) );
  A2O1A1Ixp33_ASAP7_75t_SL U39056 ( .A1(n30438), .A2(n31415), .B(n30437), .C(
        n30436), .Y(n2751) );
  A2O1A1Ixp33_ASAP7_75t_SL U39057 ( .A1(n30449), .A2(n31415), .B(n30448), .C(
        n30447), .Y(n2747) );
  OAI211xp5_ASAP7_75t_SL U39058 ( .A1(n24514), .A2(n30458), .B(n30457), .C(
        n30456), .Y(n30461) );
  A2O1A1Ixp33_ASAP7_75t_SL U39059 ( .A1(n30462), .A2(n31415), .B(n30461), .C(
        n30460), .Y(n3949) );
  AO21x1_ASAP7_75t_SL U39060 ( .A1(n30471), .A2(n31345), .B(n30470), .Y(n3955)
         );
  OAI211xp5_ASAP7_75t_SL U39061 ( .A1(n30482), .A2(n31483), .B(n30481), .C(
        n30480), .Y(n30483) );
  A2O1A1Ixp33_ASAP7_75t_SL U39062 ( .A1(n22413), .A2(n30485), .B(n31488), .C(
        n30484), .Y(n30486) );
  NAND3xp33_ASAP7_75t_SL U39063 ( .A(n30492), .B(n31054), .C(n30491), .Y(
        n30493) );
  OAI211xp5_ASAP7_75t_SL U39064 ( .A1(n24681), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__14_), .B(n30494), .C(n30493), .Y(n4425)
         );
  AO21x1_ASAP7_75t_SL U39065 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5478), .B(
        n30500), .Y(n30501) );
  NAND3xp33_ASAP7_75t_SL U39066 ( .A(n30503), .B(n32253), .C(n30502), .Y(
        n30505) );
  NAND3xp33_ASAP7_75t_SL U39067 ( .A(n30508), .B(n31570), .C(n31447), .Y(
        n30510) );
  OAI211xp5_ASAP7_75t_SL U39068 ( .A1(n30552), .A2(n30983), .B(n30551), .C(
        n30550), .Y(n30553) );
  OR3x1_ASAP7_75t_SL U39069 ( .A(n31027), .B(n1637), .C(n2925), .Y(n31199) );
  AO21x1_ASAP7_75t_SL U39070 ( .A1(ic_q[6]), .A2(n22387), .B(n30559), .Y(
        n30560) );
  OAI211xp5_ASAP7_75t_SL U39071 ( .A1(n30566), .A2(n31483), .B(n30565), .C(
        n30564), .Y(n30567) );
  A2O1A1Ixp33_ASAP7_75t_SL U39072 ( .A1(n30570), .A2(n30569), .B(n31488), .C(
        n30568), .Y(n30571) );
  NAND3xp33_ASAP7_75t_SL U39073 ( .A(n30589), .B(n30588), .C(n30587), .Y(
        rf_di_w[30]) );
  NAND3xp33_ASAP7_75t_SL U39074 ( .A(n30600), .B(n31542), .C(n30599), .Y(
        n30601) );
  A2O1A1Ixp33_ASAP7_75t_SL U39075 ( .A1(n32110), .A2(n30602), .B(n30949), .C(
        n30601), .Y(n4463) );
  NAND3xp33_ASAP7_75t_SL U39076 ( .A(n30617), .B(n30616), .C(n30615), .Y(
        n30618) );
  A2O1A1Ixp33_ASAP7_75t_SL U39077 ( .A1(n30620), .A2(n30619), .B(n30618), .C(
        n24634), .Y(n30624) );
  OAI211xp5_ASAP7_75t_SL U39078 ( .A1(n30626), .A2(n30625), .B(n30624), .C(
        n30623), .Y(n30630) );
  A2O1A1Ixp33_ASAP7_75t_SL U39079 ( .A1(u0_0_leon3x0_p0_dci[7]), .A2(n22398), 
        .B(n30636), .C(n30007), .Y(n30638) );
  O2A1O1Ixp5_ASAP7_75t_SL U39080 ( .A1(n30651), .A2(n31874), .B(n30650), .C(
        n30649), .Y(n4469) );
  NAND3xp33_ASAP7_75t_SL U39081 ( .A(n30665), .B(n30664), .C(n30663), .Y(
        n30675) );
  O2A1O1Ixp5_ASAP7_75t_SL U39082 ( .A1(u0_0_leon3x0_p0_iu_r_X__CTRL__WICC_), 
        .A2(n30669), .B(n30668), .C(n30667), .Y(n30670) );
  A2O1A1Ixp33_ASAP7_75t_SL U39083 ( .A1(n30676), .A2(n30675), .B(n30674), .C(
        n30673), .Y(n30945) );
  NAND3xp33_ASAP7_75t_SL U39084 ( .A(n30689), .B(n30688), .C(n30687), .Y(
        n30691) );
  NAND3xp33_ASAP7_75t_SL U39085 ( .A(n30729), .B(n30728), .C(n30727), .Y(
        rf_di_w[8]) );
  NAND3xp33_ASAP7_75t_SL U39086 ( .A(n30732), .B(n31542), .C(n30731), .Y(
        n30735) );
  OAI211xp5_ASAP7_75t_SL U39087 ( .A1(n24681), .A2(
        u0_0_leon3x0_p0_iu_r_E__OP1__8_), .B(n30735), .C(n30734), .Y(n4438) );
  OR2x2_ASAP7_75t_SL U39088 ( .A(n30780), .B(n31057), .Y(n30772) );
  A2O1A1Ixp33_ASAP7_75t_SL U39089 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_19_), .A2(
        n31833), .B(n30827), .C(n30826), .Y(n2556) );
  OR2x2_ASAP7_75t_SL U39090 ( .A(n30833), .B(n31057), .Y(n30866) );
  AO21x1_ASAP7_75t_SL U39091 ( .A1(ic_q[11]), .A2(n22387), .B(n30882), .Y(
        n30884) );
  OAI211xp5_ASAP7_75t_SL U39092 ( .A1(n30970), .A2(n31483), .B(n30887), .C(
        n30886), .Y(n30888) );
  A2O1A1Ixp33_ASAP7_75t_SL U39093 ( .A1(n22413), .A2(n24490), .B(n31488), .C(
        n30889), .Y(n30890) );
  AO21x1_ASAP7_75t_SL U39094 ( .A1(n31833), .A2(u0_0_leon3x0_p0_iu_fe_npc_3_), 
        .B(n30911), .Y(n32679) );
  XNOR2xp5_ASAP7_75t_SL U39095 ( .A(n31607), .B(n31608), .Y(n30918) );
  NAND3xp33_ASAP7_75t_SL U39096 ( .A(n30915), .B(u0_0_leon3x0_p0_dci[2]), .C(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DCS__1_), .Y(n31298) );
  NOR3xp33_ASAP7_75t_SL U39097 ( .A(n30926), .B(n30925), .C(n30924), .Y(n30930) );
  NAND4xp25_ASAP7_75t_SL U39098 ( .A(n30931), .B(n30930), .C(n30929), .D(
        n30928), .Y(n30932) );
  XNOR2xp5_ASAP7_75t_SL U39099 ( .A(n30948), .B(n30947), .Y(n30951) );
  AO21x1_ASAP7_75t_SL U39100 ( .A1(n31054), .A2(n30951), .B(n30950), .Y(n4488)
         );
  NOR3xp33_ASAP7_75t_SL U39101 ( .A(n30957), .B(n30956), .C(n30955), .Y(n30960) );
  A2O1A1Ixp33_ASAP7_75t_SL U39102 ( .A1(
        u0_0_leon3x0_p0_iu_v_E__CTRL__INST__22_), .A2(n30963), .B(n30962), .C(
        n30961), .Y(n30964) );
  A2O1A1Ixp33_ASAP7_75t_SL U39103 ( .A1(n30990), .A2(n30989), .B(
        apb0_r_CFGSEL_), .C(n30988), .Y(n30991) );
  OAI211xp5_ASAP7_75t_SL U39104 ( .A1(n31046), .A2(n31483), .B(n31007), .C(
        n31006), .Y(n31008) );
  A2O1A1Ixp33_ASAP7_75t_SL U39105 ( .A1(n22413), .A2(n31010), .B(n31488), .C(
        n31009), .Y(n31011) );
  AO21x1_ASAP7_75t_SL U39106 ( .A1(n31054), .A2(n31053), .B(n31052), .Y(n4459)
         );
  OR2x2_ASAP7_75t_SL U39107 ( .A(n31197), .B(n31057), .Y(n31184) );
  NAND4xp25_ASAP7_75t_SL U39108 ( .A(n31270), .B(n31269), .C(n31268), .D(
        n31267), .Y(n31276) );
  NAND4xp25_ASAP7_75t_SL U39109 ( .A(n31274), .B(n31273), .C(n31272), .D(
        n31271), .Y(n31275) );
  A2O1A1Ixp33_ASAP7_75t_SL U39110 ( .A1(n31309), .A2(n32245), .B(n31308), .C(
        n32437), .Y(n31310) );
  OAI211xp5_ASAP7_75t_SL U39111 ( .A1(n32735), .A2(n32602), .B(n31311), .C(
        n31310), .Y(u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__2_) );
  NAND3xp33_ASAP7_75t_SL U39112 ( .A(n31608), .B(n3133), .C(n31607), .Y(n31316) );
  A2O1A1Ixp33_ASAP7_75t_SL U39113 ( .A1(n31317), .A2(n31316), .B(n24645), .C(
        n31315), .Y(u0_0_leon3x0_p0_c0mmu_dcache0_v_WB__ADDR__4_) );
  A2O1A1Ixp33_ASAP7_75t_SL U39114 ( .A1(n31318), .A2(n32496), .B(n32481), .C(
        n31892), .Y(n31320) );
  A2O1A1Ixp33_ASAP7_75t_SL U39115 ( .A1(n31320), .A2(n31319), .B(n22405), .C(
        n32683), .Y(u0_0_leon3x0_p0_c0mmu_icache0_v_WADDRESS__4_) );
  OAI211xp5_ASAP7_75t_SL U39116 ( .A1(n31340), .A2(n31339), .B(n31338), .C(
        n31337), .Y(n31341) );
  AO21x1_ASAP7_75t_SL U39117 ( .A1(n31342), .A2(n31350), .B(n31341), .Y(n32109) );
  AO21x1_ASAP7_75t_SL U39118 ( .A1(n31346), .A2(n31345), .B(n31344), .Y(n4471)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U39119 ( .A1(n22413), .A2(n31362), .B(n31488), .C(
        n31361), .Y(n31363) );
  OAI211xp5_ASAP7_75t_SL U39120 ( .A1(n31396), .A2(n31395), .B(n31394), .C(
        n31393), .Y(n31397) );
  A2O1A1Ixp33_ASAP7_75t_SL U39121 ( .A1(n31416), .A2(n31415), .B(n31414), .C(
        n31413), .Y(n2816) );
  A2O1A1Ixp33_ASAP7_75t_SL U39122 ( .A1(n18793), .A2(
        u0_0_leon3x0_p0_iu_v_A__CWP__0_), .B(n31434), .C(n31433), .Y(n31436)
         );
  NAND3xp33_ASAP7_75t_SL U39123 ( .A(n31452), .B(u0_0_leon3x0_p0_dci[3]), .C(
        n31451), .Y(n31453) );
  AO21x1_ASAP7_75t_SL U39124 ( .A1(ic_q[4]), .A2(n22387), .B(n31468), .Y(
        n31472) );
  OAI211xp5_ASAP7_75t_SL U39125 ( .A1(n31484), .A2(n31483), .B(n31482), .C(
        n31481), .Y(n31485) );
  A2O1A1Ixp33_ASAP7_75t_SL U39126 ( .A1(n22413), .A2(n31489), .B(n31488), .C(
        n31487), .Y(n31490) );
  OAI211xp5_ASAP7_75t_SL U39127 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__0_), .A2(n32583), .B(n32545), 
        .C(n32566), .Y(n3057) );
  XNOR2xp5_ASAP7_75t_SL U39128 ( .A(u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__1_), 
        .B(n32566), .Y(n31550) );
  A2O1A1Ixp33_ASAP7_75t_SL U39129 ( .A1(n32545), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__3_), .B(n31554), .C(n31553), 
        .Y(n3060) );
  A2O1A1Ixp33_ASAP7_75t_SL U39130 ( .A1(n32545), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__4_), .B(n31555), .C(n31556), 
        .Y(n3061) );
  A2O1A1Ixp33_ASAP7_75t_SL U39131 ( .A1(n32545), .A2(
        u0_0_leon3x0_p0_c0mmu_icache0_r_FADDR__5_), .B(n31557), .C(n31560), 
        .Y(n3062) );
  OR2x2_ASAP7_75t_SL U39132 ( .A(n31569), .B(n31568), .Y(n31587) );
  A2O1A1Ixp33_ASAP7_75t_SL U39133 ( .A1(n32250), .A2(n31598), .B(n31590), .C(
        n31596), .Y(n31581) );
  NOR3xp33_ASAP7_75t_SL U39134 ( .A(n31579), .B(n32198), .C(n31578), .Y(n31580) );
  OAI211xp5_ASAP7_75t_SL U39135 ( .A1(n3071), .A2(n31593), .B(n31581), .C(
        n31588), .Y(n18100) );
  AO21x1_ASAP7_75t_SL U39136 ( .A1(n31592), .A2(n31591), .B(n31590), .Y(n31597) );
  OAI31xp33_ASAP7_75t_SL U39137 ( .A1(n24549), .A2(n31617), .A3(n31600), .B(
        n31599), .Y(n31616) );
  OAI211xp5_ASAP7_75t_SL U39138 ( .A1(n3046), .A2(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__DCS__1_), .B(n31605), .C(
        u0_0_leon3x0_p0_c0mmu_mcdi[1]), .Y(n31606) );
  A2O1A1Ixp33_ASAP7_75t_SL U39139 ( .A1(n31614), .A2(n31613), .B(n31612), .C(
        n31611), .Y(n31615) );
  A2O1A1Ixp33_ASAP7_75t_SL U39140 ( .A1(n31616), .A2(n31618), .B(n31615), .C(
        n24684), .Y(n4083) );
  A2O1A1Ixp33_ASAP7_75t_SL U39141 ( .A1(n31620), .A2(n31619), .B(n32272), .C(
        n31618), .Y(n31624) );
  AO21x1_ASAP7_75t_SL U39142 ( .A1(n31897), .A2(n31626), .B(n31625), .Y(n4079)
         );
  OR2x2_ASAP7_75t_SL U39143 ( .A(n31877), .B(n31630), .Y(n31695) );
  OAI211xp5_ASAP7_75t_SL U39144 ( .A1(apbi[32]), .A2(n22408), .B(n31837), .C(
        n24694), .Y(n4072) );
  A2O1A1Ixp33_ASAP7_75t_SL U39145 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_31_), .A2(
        n31833), .B(n31686), .C(n31685), .Y(n4334) );
  AND2x2_ASAP7_75t_SL U39146 ( .A(n32875), .B(n32723), .Y(n32883) );
  OR2x2_ASAP7_75t_SL U39147 ( .A(sr1_r_WS__3_), .B(sr1_r_WS__2_), .Y(n31712)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U39148 ( .A1(n24583), .A2(n31701), .B(n31700), .C(
        n31699), .Y(n31702) );
  NAND3xp33_ASAP7_75t_SL U39149 ( .A(n32879), .B(sr1_r_MCFG2__RAMWIDTH__1_), 
        .C(sr1_r_MCFG2__RMW_), .Y(n31704) );
  A2O1A1Ixp33_ASAP7_75t_SL U39150 ( .A1(sr1_r_READY_), .A2(n31732), .B(n32832), 
        .C(n31719), .Y(n31721) );
  NAND3xp33_ASAP7_75t_SL U39151 ( .A(n31750), .B(n32716), .C(n2357), .Y(n32696) );
  OR2x2_ASAP7_75t_SL U39152 ( .A(n32786), .B(n11260), .Y(n32787) );
  AND2x2_ASAP7_75t_SL U39153 ( .A(u0_0_leon3x0_p0_ici[86]), .B(n22405), .Y(
        n32554) );
  AND2x2_ASAP7_75t_SL U39154 ( .A(u0_0_leon3x0_p0_ici[80]), .B(n22405), .Y(
        n32537) );
  AND2x2_ASAP7_75t_SL U39155 ( .A(u0_0_leon3x0_p0_ici[82]), .B(n22405), .Y(
        n32544) );
  NAND4xp25_ASAP7_75t_SL U39156 ( .A(n33032), .B(n33020), .C(n33046), .D(
        n33008), .Y(n31797) );
  NAND4xp25_ASAP7_75t_SL U39157 ( .A(n31794), .B(n31793), .C(n32879), .D(
        n33023), .Y(n31796) );
  NAND4xp25_ASAP7_75t_SL U39158 ( .A(n33011), .B(n33017), .C(n33029), .D(
        n33049), .Y(n31795) );
  NOR3xp33_ASAP7_75t_SL U39159 ( .A(n31797), .B(n31796), .C(n31795), .Y(n31801) );
  NAND3xp33_ASAP7_75t_SL U39160 ( .A(n31801), .B(n31800), .C(n31799), .Y(
        n32039) );
  A2O1A1Ixp33_ASAP7_75t_SL U39161 ( .A1(n31892), .A2(n31806), .B(n18900), .C(
        n31805), .Y(n3702) );
  AO21x1_ASAP7_75t_SL U39162 ( .A1(n31828), .A2(u0_0_leon3x0_p0_dci[23]), .B(
        n31827), .Y(n31829) );
  AO21x1_ASAP7_75t_SL U39163 ( .A1(n31830), .A2(u0_0_leon3x0_p0_iu_N5482), .B(
        n31829), .Y(n31832) );
  A2O1A1Ixp33_ASAP7_75t_SL U39164 ( .A1(u0_0_leon3x0_p0_iu_fe_npc_18_), .A2(
        n31833), .B(n31832), .C(n31831), .Y(n2584) );
  AO21x1_ASAP7_75t_SL U39165 ( .A1(n31838), .A2(n31837), .B(n24695), .Y(n4716)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U39166 ( .A1(
        u0_0_leon3x0_p0_iu_v_A__CTRL__INST__19_), .A2(n31858), .B(n32087), .C(
        n23898), .Y(n31861) );
  A2O1A1Ixp33_ASAP7_75t_SL U39167 ( .A1(n18844), .A2(n31861), .B(n31860), .C(
        n22379), .Y(n31863) );
  A2O1A1Ixp33_ASAP7_75t_SL U39168 ( .A1(n32114), .A2(n31870), .B(n31869), .C(
        n22379), .Y(n31871) );
  NAND3xp33_ASAP7_75t_SL U39169 ( .A(n31877), .B(u0_0_leon3x0_p0_c0mmu_mcii[0]), .C(n31897), .Y(n31880) );
  OAI211xp5_ASAP7_75t_SL U39170 ( .A1(n32511), .A2(n32662), .B(
        u0_0_leon3x0_p0_dco_ICDIAG__CCTRL__BURST_), .C(
        u0_0_leon3x0_p0_c0mmu_icache0_r_BURST_), .Y(n31881) );
  NAND3xp33_ASAP7_75t_SL U39171 ( .A(n31884), .B(n3730), .C(n32153), .Y(n31886) );
  A2O1A1Ixp33_ASAP7_75t_SL U39172 ( .A1(n31890), .A2(n31889), .B(n31888), .C(
        n31887), .Y(n31896) );
  O2A1O1Ixp5_ASAP7_75t_SL U39173 ( .A1(u0_0_leon3x0_p0_ici[62]), .A2(n31906), 
        .B(n31905), .C(n32459), .Y(n31933) );
  OR2x2_ASAP7_75t_SL U39174 ( .A(n31916), .B(n31915), .Y(n31932) );
  AO21x1_ASAP7_75t_SL U39175 ( .A1(n31938), .A2(n31937), .B(n22380), .Y(n3906)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U39176 ( .A1(timer0_vtimers_1__RELOAD__31_), .A2(
        n31956), .B(n31955), .C(n31954), .Y(n4070) );
  A2O1A1Ixp33_ASAP7_75t_SL U39177 ( .A1(n31968), .A2(n31967), .B(n31966), .C(
        n31965), .Y(n31969) );
  AO21x1_ASAP7_75t_SL U39178 ( .A1(n31994), .A2(u0_0_leon3x0_p0_iu_N5494), .B(
        n31993), .Y(n31995) );
  A2O1A1Ixp33_ASAP7_75t_SL U39179 ( .A1(n18903), .A2(n32029), .B(n32028), .C(
        n32027), .Y(n32031) );
  A2O1A1Ixp33_ASAP7_75t_SL U39180 ( .A1(n32034), .A2(n32033), .B(n32032), .C(
        n32031), .Y(n4074) );
  A2O1A1Ixp33_ASAP7_75t_SL U39181 ( .A1(
        u0_0_leon3x0_p0_c0mmu_icache0_r_OVERRUN_), .A2(n24684), .B(n32129), 
        .C(n32046), .Y(n3894) );
  AO21x1_ASAP7_75t_SL U39182 ( .A1(n32052), .A2(n32051), .B(n32050), .Y(n32053) );
  A2O1A1Ixp33_ASAP7_75t_SL U39183 ( .A1(n32075), .A2(n32074), .B(n22380), .C(
        n32073), .Y(n18276) );
  A2O1A1Ixp33_ASAP7_75t_SL U39184 ( .A1(n32099), .A2(n32098), .B(n32097), .C(
        n32096), .Y(n32100) );
  OAI31xp33_ASAP7_75t_SL U39185 ( .A1(n32103), .A2(n32102), .A3(n32101), .B(
        n32100), .Y(n32105) );
  OAI222xp33_ASAP7_75t_SL U39186 ( .A1(n32213), .A2(n32218), .B1(n32232), .B2(
        n32376), .C1(n32217), .C2(n32638), .Y(dt_data[16]) );
  OAI222xp33_ASAP7_75t_SL U39187 ( .A1(n32216), .A2(n32218), .B1(n32232), .B2(
        n32383), .C1(n32642), .C2(n32217), .Y(dt_data[18]) );
  OAI222xp33_ASAP7_75t_SL U39188 ( .A1(n32219), .A2(n32218), .B1(n32232), .B2(
        n32387), .C1(n32217), .C2(n32644), .Y(dt_data[19]) );
  OAI211xp5_ASAP7_75t_SL U39189 ( .A1(n32235), .A2(n32656), .B(n32230), .C(
        n32229), .Y(dt_data[25]) );
  OAI211xp5_ASAP7_75t_SL U39190 ( .A1(n4318), .A2(n32255), .B(n32253), .C(
        n32256), .Y(n32248) );
  AO21x1_ASAP7_75t_SL U39191 ( .A1(n32446), .A2(u0_0_leon3x0_p0_c0mmu_mcdi[38]), .B(n33067), .Y(n32257) );
  A2O1A1Ixp33_ASAP7_75t_SL U39192 ( .A1(n32263), .A2(n32262), .B(n33067), .C(
        n32261), .Y(dc_address[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U39193 ( .A1(n32266), .A2(n32265), .B(n33067), .C(
        n32264), .Y(dc_address[5]) );
  AO21x1_ASAP7_75t_SL U39194 ( .A1(n32446), .A2(u0_0_leon3x0_p0_c0mmu_mcdi[44]), .B(n33067), .Y(n32267) );
  AO21x1_ASAP7_75t_SL U39195 ( .A1(n32270), .A2(n32284), .B(n32271), .Y(n3044)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U39196 ( .A1(n32278), .A2(n32277), .B(n32276), .C(
        n32275), .Y(n32279) );
  A2O1A1Ixp33_ASAP7_75t_SL U39197 ( .A1(n32286), .A2(n32390), .B(n32285), .C(
        n24543), .Y(n32348) );
  OAI211xp5_ASAP7_75t_SL U39198 ( .A1(n32394), .A2(n32348), .B(n32324), .C(
        n32323), .Y(dc_data[8]) );
  OAI211xp5_ASAP7_75t_SL U39199 ( .A1(n32397), .A2(n32348), .B(n32327), .C(
        n32326), .Y(dc_data[9]) );
  OAI211xp5_ASAP7_75t_SL U39200 ( .A1(n32341), .A2(n32398), .B(n32331), .C(
        n32330), .Y(dc_data[10]) );
  OAI211xp5_ASAP7_75t_SL U39201 ( .A1(n32404), .A2(n32348), .B(n32335), .C(
        n32334), .Y(dc_data[11]) );
  OAI211xp5_ASAP7_75t_SL U39202 ( .A1(n32407), .A2(n32348), .B(n32338), .C(
        n32337), .Y(dc_data[12]) );
  OAI211xp5_ASAP7_75t_SL U39203 ( .A1(n32436), .A2(n32348), .B(n32347), .C(
        n32346), .Y(dc_data[15]) );
  OAI211xp5_ASAP7_75t_SL U39204 ( .A1(n32360), .A2(n32431), .B(n32359), .C(
        n32358), .Y(dc_data[16]) );
  OAI211xp5_ASAP7_75t_SL U39205 ( .A1(n32365), .A2(n32431), .B(n32364), .C(
        n32363), .Y(dc_data[17]) );
  OAI211xp5_ASAP7_75t_SL U39206 ( .A1(n32375), .A2(n32431), .B(n32374), .C(
        n32373), .Y(dc_data[19]) );
  OR2x2_ASAP7_75t_SL U39207 ( .A(n32388), .B(n32435), .Y(n32425) );
  OAI211xp5_ASAP7_75t_SL U39208 ( .A1(n32417), .A2(n32431), .B(n32416), .C(
        n32415), .Y(dc_data[29]) );
  AO21x1_ASAP7_75t_SL U39209 ( .A1(dc_q[30]), .A2(n33069), .B(n32420), .Y(
        n32421) );
  A2O1A1Ixp33_ASAP7_75t_SL U39210 ( .A1(u0_0_leon3x0_p0_c0mmu_mcdi[62]), .A2(
        n2972), .B(u0_0_leon3x0_p0_c0mmu_mcdi[63]), .C(n32451), .Y(n32453) );
  A2O1A1Ixp33_ASAP7_75t_SL U39211 ( .A1(n24513), .A2(n32453), .B(n32452), .C(
        n24684), .Y(n2290) );
  OAI211xp5_ASAP7_75t_SL U39212 ( .A1(n32457), .A2(n24643), .B(n3065), .C(
        n32597), .Y(it_wren) );
  OR2x2_ASAP7_75t_SL U39213 ( .A(n32511), .B(n32503), .Y(n32508) );
  OR2x2_ASAP7_75t_SL U39214 ( .A(n32511), .B(n32510), .Y(n32521) );
  OAI31xp33_ASAP7_75t_SL U39215 ( .A1(n32598), .A2(n14803), .A3(n24643), .B(
        n32597), .Y(ic_wren) );
  NAND3xp33_ASAP7_75t_SL U39216 ( .A(n18858), .B(n32666), .C(n32665), .Y(
        n32671) );
  A2O1A1Ixp33_ASAP7_75t_SL U39217 ( .A1(n32686), .A2(n32671), .B(n32670), .C(
        n14803), .Y(n32672) );
  AO21x1_ASAP7_75t_SL U39218 ( .A1(u0_0_leon3x0_p0_dco_ICDIAG__ADDR__4_), .A2(
        n32694), .B(n32693), .Y(ic_address[2]) );
  NOR3xp33_ASAP7_75t_SL U39219 ( .A(n32706), .B(n32705), .C(sr1_r_IOSN__1_), 
        .Y(n32708) );
  AND2x2_ASAP7_75t_SL U39220 ( .A(n32708), .B(n32707), .Y(n2304) );
  OR2x2_ASAP7_75t_SL U39221 ( .A(n32883), .B(n2304), .Y(n2302) );
  AND2x2_ASAP7_75t_SL U39222 ( .A(n32712), .B(n22381), .Y(n32739) );
  A2O1A1Ixp33_ASAP7_75t_SL U39223 ( .A1(n32801), .A2(sr1_r_MCFG1__ROMWIDTH__1_), .B(n32724), .C(n32877), .Y(n32725) );
  OR4x1_ASAP7_75t_SL U39224 ( .A(n32749), .B(sr1_sdi_HSIZE__1_), .C(n32742), 
        .D(n32833), .Y(n32745) );
  OAI31xp33_ASAP7_75t_SL U39225 ( .A1(sr1_sdi_HSIZE__0_), .A2(n1724), .A3(
        n32745), .B(n32743), .Y(n32746) );
  OAI31xp33_ASAP7_75t_SL U39226 ( .A1(sr1_sdi_HSIZE__0_), .A2(address[0]), 
        .A3(n32745), .B(n32743), .Y(n32747) );
  A2O1A1Ixp33_ASAP7_75t_SL U39227 ( .A1(n2924), .A2(n33033), .B(n32750), .C(
        n32774), .Y(n32760) );
  A2O1A1Ixp33_ASAP7_75t_SL U39228 ( .A1(n32756), .A2(n32774), .B(n32755), .C(
        n32754), .Y(n32757) );
  A2O1A1Ixp33_ASAP7_75t_SL U39229 ( .A1(n32760), .A2(n32759), .B(n32758), .C(
        n32757), .Y(n32785) );
  OAI211xp5_ASAP7_75t_SL U39230 ( .A1(n32780), .A2(n32767), .B(n32766), .C(
        n32765), .Y(n32768) );
  O2A1O1Ixp5_ASAP7_75t_SL U39231 ( .A1(n32774), .A2(n32782), .B(n32768), .C(
        sr1_r_MCFG2__RAMBANKSZ__0_), .Y(n32769) );
  OAI211xp5_ASAP7_75t_SL U39232 ( .A1(n32780), .A2(n32779), .B(n32778), .C(
        n32777), .Y(n32781) );
  O2A1O1Ixp5_ASAP7_75t_SL U39233 ( .A1(sr1_r_MCFG2__RAMBANKSZ__1_), .A2(n32782), .B(n32781), .C(n32784), .Y(n32783) );
  NAND3xp33_ASAP7_75t_SL U39234 ( .A(n32817), .B(n32815), .C(n32808), .Y(
        n32799) );
  NOR3xp33_ASAP7_75t_SL U39235 ( .A(n32802), .B(n32801), .C(n22393), .Y(n32803) );
  NAND3xp33_ASAP7_75t_SL U39236 ( .A(n32817), .B(n32816), .C(n32815), .Y(
        n32818) );
  NAND3xp33_ASAP7_75t_SL U39237 ( .A(n32886), .B(n32835), .C(n32834), .Y(
        n32887) );
  OR2x2_ASAP7_75t_SL U39238 ( .A(n1724), .B(n1723), .Y(n32908) );
  A2O1A1Ixp33_ASAP7_75t_SL U39239 ( .A1(sr1_r_MCFG2__RAMWIDTH__0_), .A2(n32879), .B(n32878), .C(n32877), .Y(n32880) );
  OR2x2_ASAP7_75t_SL U39240 ( .A(sr1_r_BUSW__1_), .B(sr1_r_BUSW__0_), .Y(
        n32918) );
  OR2x2_ASAP7_75t_SL U39241 ( .A(n32910), .B(n32912), .Y(n32977) );
  OAI211xp5_ASAP7_75t_SL U39242 ( .A1(n32977), .A2(n32916), .B(n32915), .C(
        n32914), .Y(n32921) );
  OAI211xp5_ASAP7_75t_SL U39243 ( .A1(n32977), .A2(n32926), .B(n32925), .C(
        n32924), .Y(n32929) );
  A2O1A1Ixp33_ASAP7_75t_SL U39244 ( .A1(dataout[26]), .A2(n22433), .B(n32972), 
        .C(n32931), .Y(n32933) );
  OAI211xp5_ASAP7_75t_SL U39245 ( .A1(n32934), .A2(n32977), .B(n32933), .C(
        n32932), .Y(n32937) );
  OAI211xp5_ASAP7_75t_SL U39246 ( .A1(n32977), .A2(n32942), .B(n32941), .C(
        n32940), .Y(n32945) );
  OAI211xp5_ASAP7_75t_SL U39247 ( .A1(n32977), .A2(n32950), .B(n32949), .C(
        n32948), .Y(n32953) );
  OAI211xp5_ASAP7_75t_SL U39248 ( .A1(n32977), .A2(n32958), .B(n32957), .C(
        n32956), .Y(n32961) );
  OAI211xp5_ASAP7_75t_SL U39249 ( .A1(n32977), .A2(n32966), .B(n32965), .C(
        n32964), .Y(n32969) );
  OAI211xp5_ASAP7_75t_SL U39250 ( .A1(n32977), .A2(n32976), .B(n32975), .C(
        n32974), .Y(n32981) );
  AO21x1_ASAP7_75t_SL U39251 ( .A1(n33055), .A2(n33054), .B(n33057), .Y(
        u0_0_leon3x0_p0_iu_vp_ERROR_) );
endmodule

