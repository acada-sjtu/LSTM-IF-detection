
module or1200_top ( clk_i, rst_i, pic_ints_i, clmode_i, iwb_clk_i, iwb_rst_i, 
        iwb_ack_i, iwb_err_i, iwb_rty_i, iwb_dat_i, iwb_cyc_o, iwb_adr_o, 
        iwb_stb_o, iwb_we_o, iwb_sel_o, iwb_dat_o, iwb_cti_o, iwb_bte_o, 
        dwb_clk_i, dwb_rst_i, dwb_ack_i, dwb_err_i, dwb_rty_i, dwb_dat_i, 
        dwb_cyc_o, dwb_adr_o, dwb_stb_o, dwb_we_o, dwb_sel_o, dwb_dat_o, 
        dwb_cti_o, dwb_bte_o, dbg_stall_i, dbg_ewt_i, dbg_lss_o, dbg_is_o, 
        dbg_wp_o, dbg_bp_o, dbg_stb_i, dbg_we_i, dbg_adr_i, dbg_dat_i, 
        dbg_dat_o, dbg_ack_o, pm_cpustall_i, pm_clksd_o, pm_dc_gate_o, 
        pm_ic_gate_o, pm_dmmu_gate_o, pm_immu_gate_o, pm_tt_gate_o, 
        pm_cpu_gate_o, pm_wakeup_o, pm_lvolt_o, sig_tick, finish );
  input [19:0] pic_ints_i;
  input [1:0] clmode_i;
  input [31:0] iwb_dat_i;
  output [31:0] iwb_adr_o;
  output [3:0] iwb_sel_o;
  output [31:0] iwb_dat_o;
  output [2:0] iwb_cti_o;
  output [1:0] iwb_bte_o;
  input [31:0] dwb_dat_i;
  output [31:0] dwb_adr_o;
  output [3:0] dwb_sel_o;
  output [31:0] dwb_dat_o;
  output [2:0] dwb_cti_o;
  output [1:0] dwb_bte_o;
  output [3:0] dbg_lss_o;
  output [1:0] dbg_is_o;
  output [10:0] dbg_wp_o;
  input [31:0] dbg_adr_i;
  input [31:0] dbg_dat_i;
  output [31:0] dbg_dat_o;
  output [3:0] pm_clksd_o;
  input clk_i, rst_i, iwb_clk_i, iwb_rst_i, iwb_ack_i, iwb_err_i, iwb_rty_i,
         dwb_clk_i, dwb_rst_i, dwb_ack_i, dwb_err_i, dwb_rty_i, dbg_stall_i,
         dbg_ewt_i, dbg_stb_i, dbg_we_i, pm_cpustall_i;
  output iwb_cyc_o, iwb_stb_o, iwb_we_o, dwb_cyc_o, dwb_stb_o, dwb_we_o,
         dbg_bp_o, dbg_ack_o, pm_dc_gate_o, pm_ic_gate_o, pm_dmmu_gate_o,
         pm_immu_gate_o, pm_tt_gate_o, pm_cpu_gate_o, pm_wakeup_o, pm_lvolt_o,
         sig_tick, finish;
  wire   ic_en, supv, id_insn_22_, dc_en, or1200_immu_top_N34,
         or1200_immu_top_N33, or1200_immu_top_N30, or1200_immu_top_N29,
         or1200_immu_top_N27, or1200_immu_top_N26, or1200_immu_top_N25,
         or1200_immu_top_N24, or1200_immu_top_N21, or1200_immu_top_N20,
         or1200_immu_top_N15, or1200_immu_top_N14, or1200_immu_top_N13,
         or1200_immu_top_N12, or1200_immu_top_N10, or1200_immu_top_N9,
         or1200_immu_top_N8, or1200_immu_top_N7, or1200_immu_top_N6,
         or1200_immu_top_N5, or1200_immu_top_N3,
         or1200_immu_top_icpu_adr_default_8_, or1200_ic_top_icram_we_3_,
         or1200_ic_top_tag_v, or1200_ic_top_ictag_v, or1200_ic_top_ictag_en,
         or1200_ic_top_ictag_we, or1200_cpu_rf_dataa_0_, or1200_cpu_alu_op_2_,
         or1200_cpu_rf_rdb, or1200_cpu_epcr_1_, or1200_cpu_epcr_31_,
         or1200_cpu_except_type_1_, or1200_cpu_sr_15_, or1200_dc_top_dirty,
         or1200_dc_top_tag_v, or1200_dc_top_tag_0_, or1200_dc_top_tag_1_,
         or1200_dc_top_tag_2_, or1200_dc_top_tag_3_, or1200_dc_top_tag_4_,
         or1200_dc_top_tag_5_, or1200_dc_top_tag_6_, or1200_dc_top_tag_7_,
         or1200_dc_top_tag_8_, or1200_dc_top_tag_9_, or1200_dc_top_tag_10_,
         or1200_dc_top_tag_11_, or1200_dc_top_tag_12_, or1200_dc_top_tag_13_,
         or1200_dc_top_tag_14_, or1200_dc_top_tag_15_, or1200_dc_top_tag_16_,
         or1200_dc_top_tag_17_, or1200_dc_top_tag_18_, or1200_dc_top_tag_19_,
         or1200_dc_top_from_dcram_0_, or1200_dc_top_from_dcram_1_,
         or1200_dc_top_from_dcram_2_, or1200_dc_top_from_dcram_3_,
         or1200_dc_top_from_dcram_4_, or1200_dc_top_from_dcram_5_,
         or1200_dc_top_from_dcram_6_, or1200_dc_top_from_dcram_7_,
         or1200_dc_top_from_dcram_8_, or1200_dc_top_from_dcram_9_,
         or1200_dc_top_from_dcram_10_, or1200_dc_top_from_dcram_11_,
         or1200_dc_top_from_dcram_12_, or1200_dc_top_from_dcram_13_,
         or1200_dc_top_from_dcram_14_, or1200_dc_top_from_dcram_15_,
         or1200_dc_top_from_dcram_16_, or1200_dc_top_from_dcram_17_,
         or1200_dc_top_from_dcram_18_, or1200_dc_top_from_dcram_19_,
         or1200_dc_top_from_dcram_20_, or1200_dc_top_from_dcram_21_,
         or1200_dc_top_from_dcram_22_, or1200_dc_top_from_dcram_23_,
         or1200_dc_top_from_dcram_24_, or1200_dc_top_from_dcram_25_,
         or1200_dc_top_from_dcram_26_, or1200_dc_top_from_dcram_27_,
         or1200_dc_top_from_dcram_28_, or1200_dc_top_from_dcram_29_,
         or1200_dc_top_from_dcram_30_, or1200_dc_top_from_dcram_31_,
         or1200_dc_top_dctag_v, or1200_dc_top_dctag_en, or1200_dc_top_dctag_we,
         or1200_dc_top_dcfsm_tag_we, or1200_du_N108, or1200_du_N107,
         or1200_du_N106, or1200_du_N105, or1200_du_N104, or1200_du_N103,
         or1200_du_N98, or1200_du_N97, or1200_du_N96, or1200_du_N95,
         or1200_du_N76, or1200_du_dbg_ack, or1200_pic_N66, or1200_pic_N65,
         or1200_pic_N64, or1200_pic_N63, or1200_pic_N62, or1200_pic_N61,
         or1200_pic_N60, or1200_pic_N59, or1200_pic_N58, or1200_pic_N57,
         or1200_pic_N56, or1200_pic_N55, or1200_pic_N54, or1200_pic_N53,
         or1200_pic_N52, or1200_pic_N51, or1200_pic_N50, or1200_pic_N49,
         or1200_pic_N48, or1200_pic_N47, or1200_pic_picmr_19_, iwb_biu_N62,
         iwb_biu_N36, dwb_biu_N62, dwb_biu_N36, or1200_cpu_or1200_if_if_bypass,
         or1200_cpu_or1200_fpu_fpu_op_valid_re_r,
         or1200_cpu_or1200_fpu_b_is_zero, or1200_cpu_or1200_fpu_a_is_zero,
         or1200_cpu_or1200_fpu_a_b_sign_xor, or1200_cpu_or1200_fpu_b_is_inf,
         or1200_cpu_or1200_fpu_a_is_inf, or1200_cpu_or1200_fpu_b_is_qnan,
         or1200_cpu_or1200_fpu_a_is_qnan, or1200_cpu_or1200_fpu_b_is_snan,
         or1200_cpu_or1200_fpu_a_is_snan, or1200_cpu_or1200_fpu_dbz,
         or1200_cpu_or1200_fpu_inf, or1200_cpu_or1200_fpu_ine_conv,
         or1200_cpu_or1200_fpu_ine, or1200_cpu_or1200_fpu_zero_conv,
         or1200_cpu_or1200_fpu_zero, or1200_cpu_or1200_fpu_qnan,
         or1200_cpu_or1200_fpu_snan, or1200_cpu_or1200_fpu_underflow,
         or1200_cpu_or1200_fpu_overflow, or1200_cpu_or1200_fpu_snan_conv,
         or1200_cpu_or1200_fpu_fpu_arith_done,
         or1200_cpu_or1200_fpu_fpu_op_r_0_, or1200_cpu_or1200_fpu_fpu_op_r_1_,
         or1200_cpu_or1200_fpu_fpu_op_r_2_, or1200_cpu_or1200_fpu_fpu_op_r_3_,
         or1200_cpu_or1200_fpu_fpu_op_r_4_, or1200_cpu_or1200_fpu_fpu_op_r_5_,
         or1200_cpu_or1200_fpu_fpu_op_r_6_,
         or1200_cpu_or1200_fpu_fpu_arith_N114,
         or1200_cpu_or1200_fpu_fpu_arith_N105,
         or1200_cpu_or1200_fpu_fpu_arith_N104,
         or1200_cpu_or1200_fpu_fpu_arith_N103,
         or1200_cpu_or1200_fpu_fpu_arith_N102,
         or1200_cpu_or1200_fpu_fpu_arith_N101,
         or1200_cpu_or1200_fpu_fpu_arith_N100,
         or1200_cpu_or1200_fpu_fpu_arith_N99,
         or1200_cpu_or1200_fpu_fpu_arith_N98,
         or1200_cpu_or1200_fpu_fpu_arith_N97,
         or1200_cpu_or1200_fpu_fpu_arith_N96,
         or1200_cpu_or1200_fpu_fpu_arith_N95,
         or1200_cpu_or1200_fpu_fpu_arith_N94,
         or1200_cpu_or1200_fpu_fpu_arith_N93,
         or1200_cpu_or1200_fpu_fpu_arith_N92,
         or1200_cpu_or1200_fpu_fpu_arith_N91,
         or1200_cpu_or1200_fpu_fpu_arith_N90,
         or1200_cpu_or1200_fpu_fpu_arith_N89,
         or1200_cpu_or1200_fpu_fpu_arith_N88,
         or1200_cpu_or1200_fpu_fpu_arith_N87,
         or1200_cpu_or1200_fpu_fpu_arith_N86,
         or1200_cpu_or1200_fpu_fpu_arith_N85,
         or1200_cpu_or1200_fpu_fpu_arith_N84,
         or1200_cpu_or1200_fpu_fpu_arith_N83,
         or1200_cpu_or1200_fpu_fpu_arith_s_output1_23_,
         or1200_cpu_or1200_fpu_fpu_arith_s_state,
         or1200_cpu_or1200_fpu_fpu_arith_s_count_0_,
         or1200_cpu_or1200_fpu_fpu_arith_s_count_1_,
         or1200_cpu_or1200_fpu_fpu_arith_s_count_2_,
         or1200_cpu_or1200_fpu_fpu_arith_s_count_3_,
         or1200_cpu_or1200_fpu_fpu_arith_s_count_4_,
         or1200_cpu_or1200_fpu_fpu_arith_s_count_5_,
         or1200_cpu_or1200_fpu_fpu_arith_s_ine_o,
         or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_ine,
         or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_ine,
         or1200_cpu_or1200_fpu_fpu_arith_serial_mul_sign,
         or1200_cpu_or1200_fpu_fpu_arith_s_start_i,
         or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_ine_o,
         or1200_cpu_or1200_fpu_fpu_arith_addsub_sign_o,
         or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_,
         or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_,
         or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_,
         or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_,
         or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_27_,
         or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_,
         or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_29_,
         or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_30_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_sign,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_0_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_2_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_3_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_4_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_5_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_6_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_7_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_8_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_9_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_10_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_11_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_12_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_13_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_14_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_15_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_16_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_17_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_18_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_19_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_20_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_21_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_nan,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_qnan_d,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_inf_d,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_0_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_0_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_2_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_0_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_0_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_3_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_4_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_5_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_6_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_7_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_8_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_9_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_10_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_11_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_12_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_13_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_14_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_15_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_16_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_17_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_18_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_19_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_20_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_21_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_22_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_30_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_31_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_27_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_25_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_26_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_27_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_N190,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_s_exp_10_o_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_26_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_27_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_28_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_29_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_30_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_31_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_32_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_33_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_34_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_35_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_36_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_37_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_38_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_39_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_40_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_41_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_42_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_43_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_44_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_45_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_46_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_47_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_48_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_49_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_N586,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_N139,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_25_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_v_shl_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_output_o_31_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_25_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_26_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_25_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_26_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_27_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_28_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_29_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_30_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_snan_r_a,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_r_a,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_infa_f_r,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_expa_ff, n235, n527, n529,
         n531, n533, n535, n537, n539, n541, n543, n545, n547, n549, n551,
         n553, n555, n557, n559, n561, n563, n565, n572, n579, n589, n596,
         n603, n610, n617, n626, n631, n636, n643, n648, n653, n658, n663,
         n668, n673, n678, n683, n688, n693, n698, n703, n708, n713, n720,
         n727, n748, n749, n751, n753, n755, n757, n759, n761, n763, n765,
         n767, n769, n771, n773, n775, n777, n779, n781, n783, n785, n787,
         n789, n791, n793, n795, n797, n799, n801, n803, n805, n807, n809,
         n811, n813, n815, n817, n819, n821, n823, n825, n826, n829, n831,
         n833, n835, n837, n839, n840, n843, n845, n847, n849, n850, n852,
         n854, n856, n858, n860, n861, n863, n865, n867, n869, n870, n872,
         n874, n876, n878, n879, n881, n883, n885, n887, n888, n890, n892,
         n894, n896, n897, n899, n901, n903, n905, n906, n908, n910, n912,
         n914, n915, n917, n919, n921, n923, n924, n926, n928, n930, n932,
         n933, n935, n937, n939, n941, n942, n944, n946, n948, n950, n951,
         n953, n955, n957, n959, n960, n962, n964, n966, n968, n971, n973,
         n975, n977, n978, n980, n982, n984, n986, n989, n991, n993, n995,
         n998, n1000, n1002, n1004, n1007, n1009, n1011, n1013, n1014, n1016,
         n1018, n1020, n1022, n1023, n1025, n1027, n1028, n1031, n1033, n1035,
         n1036, n1038, n1039, n1042, n1044, n1046, n1047, n1049, n1050, n1053,
         n1055, n1057, n1058, n1060, n1061, n1064, n1066, n1068, n1069, n1071,
         n1073, n1075, n1076, n1079, n1080, n1082, n1084, n1086, n1088, n1090,
         n1091, n1093, n1095, n1097, n1099, n1101, n1102, n1104, n1106, n1108,
         n1110, n1112, n1113, n1115, n1117, n1119, n1121, n1123, n1125, n1127,
         n1129, n1131, n1133, n1135, n1137, n1139, n1141, n1143, n1145, n1147,
         n1149, n1151, n1153, n1155, n1157, n1159, n1161, n1163, n1165, n1167,
         n1169, n1171, n1173, n1175, n1177, n1179, n1181, n1183, n1185, n1187,
         n1188, n1190, n1192, n1193, n1195, n1197, n1200, n1202, n1205, n1207,
         n1210, n1212, n1215, n1217, n1220, n1222, n1223, n1225, n1227, n1230,
         n1232, n1235, n1237, n1238, n1240, n1242, n1245, n1247, n1250, n1252,
         n1253, n1255, n1257, n1260, n1262, n1263, n1265, n1267, n1270, n1272,
         n1275, n1277, n1278, n1280, n1282, n1285, n1287, n1288, n1290, n1292,
         n1293, n1295, n1297, n1298, n1300, n1302, n1303, n1305, n1307, n1308,
         n1310, n1312, n1313, n1315, n1317, n1318, n1320, n1322, n1323, n1325,
         n1327, n1328, n1330, n1332, n1333, n1335, n1337, n1339, n1341, n1343,
         n1345, n1347, n1349, n1350, n1352, n1353, n1356, n1358, n1360, n1362,
         n1364, n1366, n1368, n1370, n1372, n1374, n1376, n1378, n1380, n1382,
         n1384, n1386, n1388, n1390, n1392, n1394, n1396, n1398, n1400, n1402,
         n1404, n1406, n1408, n1410, n1412, n1414, n1416, n1418, n1420, n1422,
         n1424, n1426, n1428, n1430, n1432, n1434, n1436, n1438, n1440, n1442,
         n1444, n1446, n1448, n1450, n1452, n1454, n1456, n1458, n1460, n1462,
         n1464, n1466, n1468, n1470, n1472, n1474, n1476, n1478, n1480, n1482,
         n1484, n1486, n1487, n1489, n1492, n1494, n1496, n1497, n1499, n1501,
         n1502, n1504, n1505, n1506, n1508, n1510, n1511, n1512, n1514, n1516,
         n1517, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1531, n1533, n1534, n1536, n1537, n1539, n1540, n1543, n1546,
         n1547, n1550, n1551, n1552, n1553, n1556, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1566, n1567, n1568, n1571, n1573, n1574, n1576,
         n1577, n1580, n1581, n1582, n1584, n1588, n1590, n1591, n1593, n1594,
         n1597, n1598, n1599, n1600, n1602, n1603, n1606, n1608, n1609, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1621, n1622, n1623,
         n1626, n1628, n1629, n1631, n1632, n1633, n1634, n1636, n1637, n1638,
         n1640, n1642, n1643, n1645, n1646, n1647, n1648, n1651, n1652, n1653,
         n1656, n1658, n1659, n1661, n1662, n1663, n1664, n1667, n1668, n1669,
         n1672, n1674, n1677, n1678, n1679, n1680, n1683, n1684, n1686, n1687,
         n1690, n1692, n1693, n1695, n1696, n1697, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1717, n1719, n1721, n1722, n1725, n1727, n1728,
         n1729, n1733, n1735, n1737, n1739, n1740, n1743, n1746, n1749, n1753,
         n1755, n1757, n1758, n1761, n1762, n1763, n1764, n1766, n1768, n1770,
         n1771, n1774, n1776, n1777, n1779, n1780, n1782, n1785, n1787, n1788,
         n1790, n1791, n1792, n1793, n1796, n1798, n1799, n1802, n1804, n1805,
         n1807, n1808, n1809, n1810, n1813, n1815, n1816, n1819, n1821, n1822,
         n1824, n1826, n1828, n1830, n1832, n1833, n1836, n1837, n1838, n1839,
         n1842, n1844, n1847, n1849, n1851, n1853, n1854, n1857, n1859, n1862,
         n1865, n1868, n1871, n1874, n1876, n1877, n1879, n1880, n1882, n1883,
         n1885, n1886, n1888, n1889, n1891, n1892, n1894, n1895, n1897, n1898,
         n1900, n1901, n1903, n1904, n1906, n1907, n1909, n1910, n1912, n1913,
         n1915, n1916, n1918, n1919, n1921, n1922, n1924, n1925, n1926, n1929,
         n1931, n1934, n1936, n1938, n1939, n1941, n1943, n1945, n1946, n1949,
         n1951, n1952, n1953, n1956, n1958, n1959, n1961, n1963, n1964, n1967,
         n1968, n1969, n1971, n1973, n1974, n1976, n1978, n1979, n1981, n1983,
         n1985, n1986, n1989, n1990, n1991, n1992, n1995, n1996, n1997, n1998,
         n2001, n2002, n2003, n2006, n2007, n2008, n2009, n2011, n2012, n2013,
         n2016, n2017, n2018, n2021, n2023, n2024, n2026, n2028, n2029, n2031,
         n2033, n2035, n2037, n2039, n2040, n2042, n2043, n2045, n2047, n2048,
         n2050, n2052, n2054, n2056, n2057, n2059, n2060, n2062, n2064, n2065,
         n2067, n2069, n2071, n2073, n2074, n2076, n2077, n2079, n2080, n2083,
         n2086, n2087, n2090, n2091, n2093, n2095, n2096, n2098, n2100, n2101,
         n2103, n2105, n2107, n2108, n2110, n2112, n2113, n2115, n2117, n2119,
         n2120, n2122, n2124, n2125, n2127, n2129, n2131, n2132, n2134, n2136,
         n2137, n2139, n2141, n2142, n2145, n2146, n2148, n2150, n2151, n2153,
         n2154, n2157, n2158, n2160, n2162, n2163, n2165, n2166, n2169, n2170,
         n2172, n2179, n2181, n2182, n2184, n2186, n2188, n2189, n2191, n2193,
         n2194, n2196, n2197, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2210, n2216, n2218, n2220, n2226, n2228, n2230,
         n2232, n2234, n2236, n2238, n2240, n2242, n2244, n2246, n2248, n2250,
         n2254, n2258, n2260, n2262, n2263, n2265, n2267, n2269, n2271, n2273,
         n2275, n2277, n2279, n2281, n2283, n2285, n2287, n2289, n2291, n2293,
         n2295, n2297, n2299, n2301, n2303, n2305, n2307, n2309, n2311, n2313,
         n2316, n2317, n2318, n2320, n2322, n2323, n2324, n2326, n2327, n2328,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2338, n2339, n2340,
         n2342, n2343, n2344, n2345, n2346, n2348, n2349, n2350, n2352, n2353,
         n2354, n2356, n2358, n2360, n2362, n2363, n2364, n2366, n2368, n2369,
         n2370, n2372, n2373, n2374, n2376, n2377, n2378, n2379, n2380, n2382,
         n2383, n2384, n2386, n2388, n2389, n2390, n2392, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2402, n2404, n2405, n2406, n2408, n2409,
         n2410, n2411, n2412, n2414, n2417, n2418, n2419, n2421, n2422, n2423,
         n2424, n2425, n2427, n2428, n2429, n2431, n2432, n2433, n2435, n2436,
         n2437, n2439, n2440, n2441, n2442, n2443, n2445, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2461,
         n2462, n2464, n2466, n2467, n2469, n2470, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2487,
         n2488, n2489, n2490, n2491, n2493, n2496, n2497, n2499, n2501, n2503,
         n2504, n2506, n2508, n2511, n2514, n2515, n2517, n2519, n2521, n2522,
         n2524, n2526, n2527, n2529, n2532, n2533, n2536, n2539, n2540, n2542,
         n2544, n2545, n2547, n2549, n2550, n2552, n2555, n2556, n2558, n2559,
         n2561, n2562, n2564, n2565, n2567, n2569, n2572, n2573, n2575, n2577,
         n2579, n2581, n2583, n2585, n2587, n2589, n2591, n2592, n2594, n2596,
         n2598, n2600, n2601, n2604, n2607, n2609, n2611, n2612, n2614, n2616,
         n2618, n2619, n2621, n2623, n2625, n2626, n2628, n2630, n2632, n2633,
         n2635, n2637, n2639, n2640, n2642, n2644, n2646, n2647, n2649, n2651,
         n2654, n2657, n2659, n2660, n2662, n2664, n2666, n2667, n2669, n2671,
         n2673, n2674, n2676, n2678, n2680, n2681, n2683, n2685, n2687, n2688,
         n2691, n2693, n2694, n2696, n2698, n2700, n2703, n2705, n2707, n2709,
         n2711, n2713, n2715, n2717, n2719, n2721, n2723, n2725, n2727, n2729,
         n2731, n2733, n2735, n2737, n2739, n2741, n2743, n2745, n2747, n2749,
         n2751, n2753, n2755, n2757, n2759, n2761, n2763, n2765, n2767, n2769,
         n2770, n2773, n2775, n2777, n2779, n2781, n2783, n2785, n2786, n2789,
         n2791, n2792, n2794, n2796, n2798, n2799, n2802, n2804, n2805, n2807,
         n2808, n2811, n2814, n2816, n2817, n2819, n2821, n2822, n2824, n2826,
         n2827, n2830, n2832, n2835, n2837, n2838, n2841, n2843, n2844, n2845,
         n2848, n2850, n2852, n2853, n2854, n2856, n2858, n2859, n2860, n2862,
         n2864, n2865, n2867, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2902, n2934, n2935, n2936, n2939,
         n2941, n2942, n2944, n2945, n2946, n2949, n2950, n2951, n2952, n2953,
         n2956, n2958, n2959, n2961, n2963, n2964, n2966, n2967, n2970, n2972,
         n2974, n2976, n2977, n2979, n2980, n2982, n2983, n2985, n2986, n2988,
         n2989, n2991, n2992, n2994, n2995, n2997, n2998, n3000, n3001, n3003,
         n3004, n3006, n3007, n3009, n3010, n3012, n3013, n3015, n3016, n3018,
         n3019, n3021, n3022, n3024, n3025, n3027, n3028, n3030, n3031, n3033,
         n3034, n3036, n3037, n3039, n3040, n3042, n3043, n3045, n3046, n3048,
         n3049, n3051, n3052, n3054, n3055, n3057, n3058, n3060, n3061, n3063,
         n3064, n3066, n3068, n3069, n3071, n3072, n3074, n3076, n3078, n3080,
         n3082, n3084, n3086, n3088, n3090, n3092, n3095, n3097, n3100, n3103,
         n3105, n3107, n3109, n3111, n3112, n3115, n3117, n3119, n3121, n3123,
         n3124, n3127, n3128, n3130, n3132, n3134, n3136, n3138, n3141, n3142,
         n3143, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3174, n3176, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3254, n3256, n3257, n3258,
         n3259, n3260, n3262, n3265, n3266, n3271, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3313, n3321, n3327, n3331, n3337, n3338, n3339,
         n3340, n3341, n3351, n3374, n3375, n3376, n3390, n3392, n3417, n3418,
         n3419, n3423, n3426, n3645, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3920, n3921, n3922, n3923, n4041, n4042, n4045, n4046, n4049, n4050,
         n4053, n4054, n4057, n4058, n4061, n4062, n4066, n4067, n4070, n4071,
         n4089, n4090, n4091, n4092, n4093, n4095, n4097, n4099, n4101, n4103,
         n4106, n4108, n4110, n4112, n4114, n4116, n4118, n4120, n4122, n4124,
         n4126, n4128, n4130, n4132, n4133, n4134, n4135, n4136, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4152, n4183,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4320,
         n4743, n4747, n5349, n5503, n5505, n5506, n5507, n5508, n5509, n5510,
         n5513, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n6731, n6739, n7192, n7615, n7616,
         n7617, n7620, n7621, n7622, n7625, n7626, n7627, n7630, n7631, n7632,
         n7635, n7636, n7637, n8750, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9206,
         n9208, n9209, n9210, n9212, n9213, n9214, n9215, n9216, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9235, n9236, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9380, n9381, n9382, n9383,
         n9384, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9427, n9429, n9430, n9431, n9433, n9434, n9435, n9436, n9437, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9479, n9480, n9481, n9482,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9559, n9560, n9562, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, or1200_cpu_or1200_rf_n145,
         or1200_cpu_or1200_rf_n144, or1200_cpu_or1200_rf_n142,
         or1200_cpu_or1200_rf_n141, or1200_cpu_or1200_rf_n140,
         or1200_cpu_or1200_rf_n139, or1200_cpu_or1200_rf_n138,
         or1200_cpu_or1200_rf_n137, or1200_cpu_or1200_rf_n136,
         or1200_cpu_or1200_rf_n135, or1200_cpu_or1200_rf_n134,
         or1200_cpu_or1200_rf_n133, or1200_cpu_or1200_rf_n132,
         or1200_cpu_or1200_rf_n131, or1200_cpu_or1200_rf_n130,
         or1200_cpu_or1200_rf_n129, or1200_cpu_or1200_rf_n128,
         or1200_cpu_or1200_rf_n125, or1200_cpu_or1200_rf_n124,
         or1200_cpu_or1200_rf_n123, or1200_cpu_or1200_rf_n122,
         or1200_cpu_or1200_rf_n121, or1200_cpu_or1200_rf_n120,
         or1200_cpu_or1200_rf_n119, or1200_cpu_or1200_rf_n118,
         or1200_cpu_or1200_rf_n117, or1200_cpu_or1200_rf_n116,
         or1200_cpu_or1200_rf_n113, or1200_cpu_or1200_rf_n112,
         or1200_cpu_or1200_rf_n111, or1200_cpu_or1200_rf_n110,
         or1200_cpu_or1200_rf_n109, or1200_cpu_or1200_rf_n108,
         or1200_cpu_or1200_rf_n107, or1200_cpu_or1200_rf_n106,
         or1200_cpu_or1200_rf_n105, or1200_cpu_or1200_rf_n104,
         or1200_cpu_or1200_rf_n103, or1200_cpu_or1200_rf_n102,
         or1200_cpu_or1200_rf_n101, or1200_cpu_or1200_rf_n100,
         or1200_cpu_or1200_rf_n99, or1200_cpu_or1200_rf_n98,
         or1200_cpu_or1200_rf_n97, or1200_cpu_or1200_rf_n96,
         or1200_cpu_or1200_rf_n95, or1200_cpu_or1200_rf_n94,
         or1200_cpu_or1200_rf_n93, or1200_cpu_or1200_rf_n92,
         or1200_cpu_or1200_rf_n91, or1200_cpu_or1200_rf_n90,
         or1200_cpu_or1200_rf_n89, or1200_cpu_or1200_rf_n88,
         or1200_cpu_or1200_rf_n87, or1200_cpu_or1200_rf_n86,
         or1200_cpu_or1200_rf_n85, or1200_cpu_or1200_rf_n84,
         or1200_cpu_or1200_rf_n83, or1200_cpu_or1200_rf_n82,
         or1200_cpu_or1200_rf_n81, or1200_cpu_or1200_rf_n80,
         or1200_cpu_or1200_rf_n79, or1200_cpu_or1200_rf_n78,
         or1200_cpu_or1200_rf_n77, or1200_cpu_or1200_rf_n76,
         or1200_cpu_or1200_rf_n75, or1200_cpu_or1200_rf_n74,
         or1200_cpu_or1200_rf_n73, or1200_cpu_or1200_rf_n72,
         or1200_cpu_or1200_rf_n71, or1200_cpu_or1200_rf_n70,
         or1200_cpu_or1200_rf_n69, or1200_cpu_or1200_rf_n68,
         or1200_cpu_or1200_rf_n67, or1200_cpu_or1200_rf_n66,
         or1200_cpu_or1200_rf_n65, or1200_cpu_or1200_rf_n64,
         or1200_cpu_or1200_rf_n63, or1200_cpu_or1200_rf_n62,
         or1200_cpu_or1200_rf_n61, or1200_cpu_or1200_rf_n60,
         or1200_cpu_or1200_rf_n59, or1200_cpu_or1200_rf_n58,
         or1200_cpu_or1200_rf_n57, or1200_cpu_or1200_rf_n56,
         or1200_cpu_or1200_rf_n55, or1200_cpu_or1200_rf_n54,
         or1200_cpu_or1200_rf_n53, or1200_cpu_or1200_rf_n52,
         or1200_cpu_or1200_rf_n44, or1200_cpu_or1200_rf_n12,
         or1200_cpu_or1200_rf_n11, or1200_cpu_or1200_rf_n10,
         or1200_cpu_or1200_rf_n9, or1200_cpu_or1200_rf_n8,
         or1200_cpu_or1200_rf_n7, or1200_cpu_or1200_rf_N36,
         or1200_cpu_or1200_rf_N31, or1200_cpu_or1200_rf_rf_enb,
         or1200_cpu_or1200_rf_rf_we, or1200_cpu_or1200_rf_rf_we_allow,
         or1200_cpu_or1200_rf_spr_du_cs, or1200_cpu_or1200_rf_addra_last_0_,
         or1200_cpu_or1200_rf_addra_last_1_,
         or1200_cpu_or1200_rf_addra_last_2_,
         or1200_cpu_or1200_rf_addra_last_3_,
         or1200_cpu_or1200_rf_addra_last_4_, or1200_cpu_or1200_rf_rf_ena,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N1,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N3,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N5,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N6,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N9,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N10,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N11,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N13,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N14,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N15,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N17,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N19,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N22,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N34,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n66,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n68,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n70,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n72,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n74,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n76,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n78,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n80,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n82,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n84,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n86,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n88,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n90,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n92,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n94,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n96,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n98,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n100,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n102,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n104,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n106,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n108,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n110,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n112,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n114,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n116,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n118,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n120,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n122,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n124,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n126,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n128,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n130,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n132,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n134,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n136,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n138,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n140,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n142,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n144,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n146,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n148,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n150,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n152,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n154,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n156,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n158,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n160,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n162,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n164,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n166,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n168,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n170,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n172,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n174,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n176,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n178,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n180,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n182,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n184,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n186,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n188,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n190,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n192,
         or1200_cpu_or1200_mult_mac_n1625, or1200_cpu_or1200_mult_mac_n1624,
         or1200_cpu_or1200_mult_mac_n1623, or1200_cpu_or1200_mult_mac_n1622,
         or1200_cpu_or1200_mult_mac_n1621, or1200_cpu_or1200_mult_mac_n1620,
         or1200_cpu_or1200_mult_mac_n1619, or1200_cpu_or1200_mult_mac_n1618,
         or1200_cpu_or1200_mult_mac_n1617, or1200_cpu_or1200_mult_mac_n1616,
         or1200_cpu_or1200_mult_mac_n1615, or1200_cpu_or1200_mult_mac_n1614,
         or1200_cpu_or1200_mult_mac_n1613, or1200_cpu_or1200_mult_mac_n1612,
         or1200_cpu_or1200_mult_mac_n1611, or1200_cpu_or1200_mult_mac_n1610,
         or1200_cpu_or1200_mult_mac_n1609, or1200_cpu_or1200_mult_mac_n1608,
         or1200_cpu_or1200_mult_mac_n1607, or1200_cpu_or1200_mult_mac_n1606,
         or1200_cpu_or1200_mult_mac_n1605, or1200_cpu_or1200_mult_mac_n1604,
         or1200_cpu_or1200_mult_mac_n1603, or1200_cpu_or1200_mult_mac_n1602,
         or1200_cpu_or1200_mult_mac_n1601, or1200_cpu_or1200_mult_mac_n1600,
         or1200_cpu_or1200_mult_mac_n1599, or1200_cpu_or1200_mult_mac_n1598,
         or1200_cpu_or1200_mult_mac_n1597, or1200_cpu_or1200_mult_mac_n1596,
         or1200_cpu_or1200_mult_mac_n1595, or1200_cpu_or1200_mult_mac_n1594,
         or1200_cpu_or1200_mult_mac_n1593, or1200_cpu_or1200_mult_mac_n1592,
         or1200_cpu_or1200_mult_mac_n1591, or1200_cpu_or1200_mult_mac_n1590,
         or1200_cpu_or1200_mult_mac_n1589, or1200_cpu_or1200_mult_mac_n1588,
         or1200_cpu_or1200_mult_mac_n1587, or1200_cpu_or1200_mult_mac_n1586,
         or1200_cpu_or1200_mult_mac_n1585, or1200_cpu_or1200_mult_mac_n1584,
         or1200_cpu_or1200_mult_mac_n1583, or1200_cpu_or1200_mult_mac_n1582,
         or1200_cpu_or1200_mult_mac_n1581, or1200_cpu_or1200_mult_mac_n1580,
         or1200_cpu_or1200_mult_mac_n1579, or1200_cpu_or1200_mult_mac_n1578,
         or1200_cpu_or1200_mult_mac_n1577, or1200_cpu_or1200_mult_mac_n1576,
         or1200_cpu_or1200_mult_mac_n1575, or1200_cpu_or1200_mult_mac_n1574,
         or1200_cpu_or1200_mult_mac_n1573, or1200_cpu_or1200_mult_mac_n1572,
         or1200_cpu_or1200_mult_mac_n1571, or1200_cpu_or1200_mult_mac_n1570,
         or1200_cpu_or1200_mult_mac_n1569, or1200_cpu_or1200_mult_mac_n1568,
         or1200_cpu_or1200_mult_mac_n1567, or1200_cpu_or1200_mult_mac_n1566,
         or1200_cpu_or1200_mult_mac_n1565, or1200_cpu_or1200_mult_mac_n1564,
         or1200_cpu_or1200_mult_mac_n1563, or1200_cpu_or1200_mult_mac_n1562,
         or1200_cpu_or1200_mult_mac_n1560, or1200_cpu_or1200_mult_mac_n1559,
         or1200_cpu_or1200_mult_mac_n1558, or1200_cpu_or1200_mult_mac_n1557,
         or1200_cpu_or1200_mult_mac_n1556, or1200_cpu_or1200_mult_mac_n1555,
         or1200_cpu_or1200_mult_mac_n1554, or1200_cpu_or1200_mult_mac_n1553,
         or1200_cpu_or1200_mult_mac_n1552, or1200_cpu_or1200_mult_mac_n1551,
         or1200_cpu_or1200_mult_mac_n1550, or1200_cpu_or1200_mult_mac_n1549,
         or1200_cpu_or1200_mult_mac_n1548, or1200_cpu_or1200_mult_mac_n1544,
         or1200_cpu_or1200_mult_mac_n1542, or1200_cpu_or1200_mult_mac_n1541,
         or1200_cpu_or1200_mult_mac_n1539, or1200_cpu_or1200_mult_mac_n1537,
         or1200_cpu_or1200_mult_mac_n1535, or1200_cpu_or1200_mult_mac_n1534,
         or1200_cpu_or1200_mult_mac_n1531, or1200_cpu_or1200_mult_mac_n1530,
         or1200_cpu_or1200_mult_mac_n1529, or1200_cpu_or1200_mult_mac_n1528,
         or1200_cpu_or1200_mult_mac_n1527, or1200_cpu_or1200_mult_mac_n1526,
         or1200_cpu_or1200_mult_mac_n1525, or1200_cpu_or1200_mult_mac_n1524,
         or1200_cpu_or1200_mult_mac_n1523, or1200_cpu_or1200_mult_mac_n1522,
         or1200_cpu_or1200_mult_mac_n1521, or1200_cpu_or1200_mult_mac_n1520,
         or1200_cpu_or1200_mult_mac_n1519, or1200_cpu_or1200_mult_mac_n1518,
         or1200_cpu_or1200_mult_mac_n1517, or1200_cpu_or1200_mult_mac_n1516,
         or1200_cpu_or1200_mult_mac_n1515, or1200_cpu_or1200_mult_mac_n1514,
         or1200_cpu_or1200_mult_mac_n1513, or1200_cpu_or1200_mult_mac_n1512,
         or1200_cpu_or1200_mult_mac_n1511, or1200_cpu_or1200_mult_mac_n1510,
         or1200_cpu_or1200_mult_mac_n1509, or1200_cpu_or1200_mult_mac_n1508,
         or1200_cpu_or1200_mult_mac_n1507, or1200_cpu_or1200_mult_mac_n1506,
         or1200_cpu_or1200_mult_mac_n1505, or1200_cpu_or1200_mult_mac_n1504,
         or1200_cpu_or1200_mult_mac_n1503, or1200_cpu_or1200_mult_mac_n1502,
         or1200_cpu_or1200_mult_mac_n1501, or1200_cpu_or1200_mult_mac_n1500,
         or1200_cpu_or1200_mult_mac_n1499, or1200_cpu_or1200_mult_mac_n1498,
         or1200_cpu_or1200_mult_mac_n1497, or1200_cpu_or1200_mult_mac_n1496,
         or1200_cpu_or1200_mult_mac_n1107, or1200_cpu_or1200_mult_mac_n1106,
         or1200_cpu_or1200_mult_mac_n1105, or1200_cpu_or1200_mult_mac_n1104,
         or1200_cpu_or1200_mult_mac_n1103, or1200_cpu_or1200_mult_mac_n413,
         or1200_cpu_or1200_mult_mac_n411, or1200_cpu_or1200_mult_mac_n409,
         or1200_cpu_or1200_mult_mac_n407, or1200_cpu_or1200_mult_mac_n405,
         or1200_cpu_or1200_mult_mac_n403, or1200_cpu_or1200_mult_mac_n401,
         or1200_cpu_or1200_mult_mac_n399, or1200_cpu_or1200_mult_mac_n397,
         or1200_cpu_or1200_mult_mac_n395, or1200_cpu_or1200_mult_mac_n393,
         or1200_cpu_or1200_mult_mac_n391, or1200_cpu_or1200_mult_mac_n389,
         or1200_cpu_or1200_mult_mac_n387, or1200_cpu_or1200_mult_mac_n385,
         or1200_cpu_or1200_mult_mac_n383, or1200_cpu_or1200_mult_mac_n381,
         or1200_cpu_or1200_mult_mac_n379, or1200_cpu_or1200_mult_mac_n377,
         or1200_cpu_or1200_mult_mac_n375, or1200_cpu_or1200_mult_mac_n373,
         or1200_cpu_or1200_mult_mac_n371, or1200_cpu_or1200_mult_mac_n369,
         or1200_cpu_or1200_mult_mac_n367, or1200_cpu_or1200_mult_mac_n365,
         or1200_cpu_or1200_mult_mac_n363, or1200_cpu_or1200_mult_mac_n361,
         or1200_cpu_or1200_mult_mac_n359, or1200_cpu_or1200_mult_mac_n357,
         or1200_cpu_or1200_mult_mac_n355, or1200_cpu_or1200_mult_mac_n353,
         or1200_cpu_or1200_mult_mac_n351, or1200_cpu_or1200_mult_mac_n349,
         or1200_cpu_or1200_mult_mac_n347, or1200_cpu_or1200_mult_mac_n345,
         or1200_cpu_or1200_mult_mac_n343, or1200_cpu_or1200_mult_mac_n341,
         or1200_cpu_or1200_mult_mac_n339, or1200_cpu_or1200_mult_mac_n337,
         or1200_cpu_or1200_mult_mac_n335, or1200_cpu_or1200_mult_mac_n333,
         or1200_cpu_or1200_mult_mac_n331, or1200_cpu_or1200_mult_mac_n329,
         or1200_cpu_or1200_mult_mac_n327, or1200_cpu_or1200_mult_mac_n325,
         or1200_cpu_or1200_mult_mac_n323, or1200_cpu_or1200_mult_mac_n321,
         or1200_cpu_or1200_mult_mac_n319, or1200_cpu_or1200_mult_mac_n317,
         or1200_cpu_or1200_mult_mac_n315, or1200_cpu_or1200_mult_mac_n313,
         or1200_cpu_or1200_mult_mac_n311, or1200_cpu_or1200_mult_mac_n309,
         or1200_cpu_or1200_mult_mac_n307, or1200_cpu_or1200_mult_mac_n305,
         or1200_cpu_or1200_mult_mac_n303, or1200_cpu_or1200_mult_mac_n301,
         or1200_cpu_or1200_mult_mac_n299, or1200_cpu_or1200_mult_mac_n297,
         or1200_cpu_or1200_mult_mac_n295, or1200_cpu_or1200_mult_mac_n293,
         or1200_cpu_or1200_mult_mac_n291, or1200_cpu_or1200_mult_mac_n289,
         or1200_cpu_or1200_mult_mac_n287, or1200_cpu_or1200_mult_mac_n285,
         or1200_cpu_or1200_mult_mac_n282, or1200_cpu_or1200_mult_mac_n280,
         or1200_cpu_or1200_mult_mac_n278, or1200_cpu_or1200_mult_mac_n273,
         or1200_cpu_or1200_mult_mac_n271, or1200_cpu_or1200_mult_mac_n269,
         or1200_cpu_or1200_mult_mac_n267, or1200_cpu_or1200_mult_mac_n265,
         or1200_cpu_or1200_mult_mac_n263, or1200_cpu_or1200_mult_mac_n261,
         or1200_cpu_or1200_mult_mac_n259, or1200_cpu_or1200_mult_mac_n257,
         or1200_cpu_or1200_mult_mac_n255, or1200_cpu_or1200_mult_mac_n253,
         or1200_cpu_or1200_mult_mac_n251, or1200_cpu_or1200_mult_mac_n249,
         or1200_cpu_or1200_mult_mac_n247, or1200_cpu_or1200_mult_mac_n245,
         or1200_cpu_or1200_mult_mac_n243, or1200_cpu_or1200_mult_mac_n241,
         or1200_cpu_or1200_mult_mac_n239, or1200_cpu_or1200_mult_mac_n237,
         or1200_cpu_or1200_mult_mac_n235, or1200_cpu_or1200_mult_mac_n233,
         or1200_cpu_or1200_mult_mac_n231, or1200_cpu_or1200_mult_mac_n229,
         or1200_cpu_or1200_mult_mac_n227, or1200_cpu_or1200_mult_mac_n225,
         or1200_cpu_or1200_mult_mac_n223, or1200_cpu_or1200_mult_mac_n221,
         or1200_cpu_or1200_mult_mac_n219, or1200_cpu_or1200_mult_mac_n217,
         or1200_cpu_or1200_mult_mac_n215, or1200_cpu_or1200_mult_mac_n213,
         or1200_cpu_or1200_mult_mac_n211, or1200_cpu_or1200_mult_mac_n209,
         or1200_cpu_or1200_mult_mac_n207, or1200_cpu_or1200_mult_mac_n205,
         or1200_cpu_or1200_mult_mac_n203, or1200_cpu_or1200_mult_mac_n201,
         or1200_cpu_or1200_mult_mac_n199, or1200_cpu_or1200_mult_mac_n197,
         or1200_cpu_or1200_mult_mac_n195, or1200_cpu_or1200_mult_mac_n193,
         or1200_cpu_or1200_mult_mac_n191, or1200_cpu_or1200_mult_mac_n189,
         or1200_cpu_or1200_mult_mac_n187, or1200_cpu_or1200_mult_mac_n185,
         or1200_cpu_or1200_mult_mac_n183, or1200_cpu_or1200_mult_mac_n181,
         or1200_cpu_or1200_mult_mac_n179, or1200_cpu_or1200_mult_mac_n177,
         or1200_cpu_or1200_mult_mac_n175, or1200_cpu_or1200_mult_mac_n173,
         or1200_cpu_or1200_mult_mac_n171, or1200_cpu_or1200_mult_mac_n169,
         or1200_cpu_or1200_mult_mac_n167, or1200_cpu_or1200_mult_mac_n165,
         or1200_cpu_or1200_mult_mac_n163, or1200_cpu_or1200_mult_mac_n161,
         or1200_cpu_or1200_mult_mac_n159, or1200_cpu_or1200_mult_mac_n157,
         or1200_cpu_or1200_mult_mac_n155, or1200_cpu_or1200_mult_mac_n153,
         or1200_cpu_or1200_mult_mac_n151, or1200_cpu_or1200_mult_mac_n149,
         or1200_cpu_or1200_mult_mac_n147, or1200_cpu_or1200_mult_mac_n145,
         or1200_cpu_or1200_mult_mac_n143, or1200_cpu_or1200_mult_mac_n141,
         or1200_cpu_or1200_mult_mac_n139, or1200_cpu_or1200_mult_mac_n136,
         or1200_cpu_or1200_mult_mac_n135, or1200_cpu_or1200_mult_mac_n128,
         or1200_cpu_or1200_mult_mac_n126, or1200_cpu_or1200_mult_mac_n124,
         or1200_cpu_or1200_mult_mac_n122, or1200_cpu_or1200_mult_mac_n120,
         or1200_cpu_or1200_mult_mac_n118, or1200_cpu_or1200_mult_mac_n116,
         or1200_cpu_or1200_mult_mac_n114, or1200_cpu_or1200_mult_mac_n112,
         or1200_cpu_or1200_mult_mac_n110, or1200_cpu_or1200_mult_mac_n108,
         or1200_cpu_or1200_mult_mac_n106, or1200_cpu_or1200_mult_mac_n104,
         or1200_cpu_or1200_mult_mac_n102, or1200_cpu_or1200_mult_mac_n100,
         or1200_cpu_or1200_mult_mac_n98, or1200_cpu_or1200_mult_mac_n96,
         or1200_cpu_or1200_mult_mac_n94, or1200_cpu_or1200_mult_mac_n92,
         or1200_cpu_or1200_mult_mac_n90, or1200_cpu_or1200_mult_mac_n88,
         or1200_cpu_or1200_mult_mac_n86, or1200_cpu_or1200_mult_mac_n84,
         or1200_cpu_or1200_mult_mac_n82, or1200_cpu_or1200_mult_mac_n80,
         or1200_cpu_or1200_mult_mac_n78, or1200_cpu_or1200_mult_mac_n76,
         or1200_cpu_or1200_mult_mac_n74, or1200_cpu_or1200_mult_mac_n72,
         or1200_cpu_or1200_mult_mac_n70, or1200_cpu_or1200_mult_mac_n68,
         or1200_cpu_or1200_mult_mac_n66, or1200_cpu_or1200_mult_mac_n64,
         or1200_cpu_or1200_mult_mac_n62, or1200_cpu_or1200_mult_mac_n60,
         or1200_cpu_or1200_mult_mac_n58, or1200_cpu_or1200_mult_mac_n56,
         or1200_cpu_or1200_mult_mac_n54, or1200_cpu_or1200_mult_mac_n52,
         or1200_cpu_or1200_mult_mac_n50, or1200_cpu_or1200_mult_mac_n48,
         or1200_cpu_or1200_mult_mac_n46, or1200_cpu_or1200_mult_mac_n44,
         or1200_cpu_or1200_mult_mac_n42, or1200_cpu_or1200_mult_mac_n40,
         or1200_cpu_or1200_mult_mac_n38, or1200_cpu_or1200_mult_mac_n36,
         or1200_cpu_or1200_mult_mac_n34, or1200_cpu_or1200_mult_mac_n32,
         or1200_cpu_or1200_mult_mac_n30, or1200_cpu_or1200_mult_mac_n28,
         or1200_cpu_or1200_mult_mac_n26, or1200_cpu_or1200_mult_mac_n24,
         or1200_cpu_or1200_mult_mac_n22, or1200_cpu_or1200_mult_mac_n20,
         or1200_cpu_or1200_mult_mac_n18, or1200_cpu_or1200_mult_mac_n16,
         or1200_cpu_or1200_mult_mac_n14, or1200_cpu_or1200_mult_mac_n12,
         or1200_cpu_or1200_mult_mac_n10, or1200_cpu_or1200_mult_mac_n8,
         or1200_cpu_or1200_mult_mac_n6, or1200_cpu_or1200_mult_mac_n4,
         or1200_cpu_or1200_mult_mac_n2, or1200_cpu_or1200_mult_mac_div_free,
         or1200_cpu_or1200_mult_mac_div_cntr_0_,
         or1200_cpu_or1200_mult_mac_div_cntr_1_,
         or1200_cpu_or1200_mult_mac_div_cntr_2_,
         or1200_cpu_or1200_mult_mac_div_cntr_3_,
         or1200_cpu_or1200_mult_mac_div_cntr_4_,
         or1200_cpu_or1200_mult_mac_N503,
         or1200_cpu_or1200_mult_mac_mac_op_r2_0_,
         or1200_cpu_or1200_mult_mac_mac_op_r2_1_,
         or1200_cpu_or1200_mult_mac_mac_op_r2_2_,
         or1200_cpu_or1200_mult_mac_N294, or1200_cpu_or1200_mult_mac_N293,
         or1200_cpu_or1200_mult_mac_N292, or1200_cpu_or1200_mult_mac_N290,
         or1200_cpu_or1200_mult_mac_mul_stall_count_1_,
         or1200_cpu_or1200_mult_mac_ex_freeze_r, DP_OP_742J1_130_9702_n59,
         DP_OP_741J1_129_6992_n46,
         or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_mult_x_1_n211, n12827,
         n12855, n12856, n12861, n12863, n12864, n12871, n12873, n12874,
         n12875, n12876, n12970, n12980, n12981, n12986, n14249, n14251,
         n14253, n14494, n17027, n17028, n17031, n17032, n17033, n17034,
         n17035, n17036, n18256, n18405, n21879, n22057,
         or1200_cpu_or1200_except_n1831, or1200_cpu_or1200_except_n1830,
         or1200_cpu_or1200_except_n1827, or1200_cpu_or1200_except_n1826,
         or1200_cpu_or1200_except_n1825, or1200_cpu_or1200_except_n1824,
         or1200_cpu_or1200_except_n1821, or1200_cpu_or1200_except_n1820,
         or1200_cpu_or1200_except_n1819, or1200_cpu_or1200_except_n1818,
         or1200_cpu_or1200_except_n1817, or1200_cpu_or1200_except_n1816,
         or1200_cpu_or1200_except_n1815, or1200_cpu_or1200_except_n1814,
         or1200_cpu_or1200_except_n1813, or1200_cpu_or1200_except_n1812,
         or1200_cpu_or1200_except_n1811, or1200_cpu_or1200_except_n1810,
         or1200_cpu_or1200_except_n1809, or1200_cpu_or1200_except_n1808,
         or1200_cpu_or1200_except_n1807, or1200_cpu_or1200_except_n1806,
         or1200_cpu_or1200_except_n1805, or1200_cpu_or1200_except_n1804,
         or1200_cpu_or1200_except_n1803, or1200_cpu_or1200_except_n1802,
         or1200_cpu_or1200_except_n1801, or1200_cpu_or1200_except_n1800,
         or1200_cpu_or1200_except_n1799, or1200_cpu_or1200_except_n1798,
         or1200_cpu_or1200_except_n1797, or1200_cpu_or1200_except_n1796,
         or1200_cpu_or1200_except_n1795, or1200_cpu_or1200_except_n1794,
         or1200_cpu_or1200_except_n1793, or1200_cpu_or1200_except_n1792,
         or1200_cpu_or1200_except_n1791, or1200_cpu_or1200_except_n1788,
         or1200_cpu_or1200_except_n1787, or1200_cpu_or1200_except_n1786,
         or1200_cpu_or1200_except_n1785, or1200_cpu_or1200_except_n1784,
         or1200_cpu_or1200_except_n1783, or1200_cpu_or1200_except_n1782,
         or1200_cpu_or1200_except_n1781, or1200_cpu_or1200_except_n1780,
         or1200_cpu_or1200_except_n1779, or1200_cpu_or1200_except_n1778,
         or1200_cpu_or1200_except_n1777, or1200_cpu_or1200_except_n1776,
         or1200_cpu_or1200_except_n1775, or1200_cpu_or1200_except_n1774,
         or1200_cpu_or1200_except_n1773, or1200_cpu_or1200_except_n1772,
         or1200_cpu_or1200_except_n1771, or1200_cpu_or1200_except_n1770,
         or1200_cpu_or1200_except_n1769, or1200_cpu_or1200_except_n1768,
         or1200_cpu_or1200_except_n1767, or1200_cpu_or1200_except_n1766,
         or1200_cpu_or1200_except_n1765, or1200_cpu_or1200_except_n1764,
         or1200_cpu_or1200_except_n1763, or1200_cpu_or1200_except_n1762,
         or1200_cpu_or1200_except_n1761, or1200_cpu_or1200_except_n1760,
         or1200_cpu_or1200_except_n1759, or1200_cpu_or1200_except_n1758,
         or1200_cpu_or1200_except_n1757, or1200_cpu_or1200_except_n1756,
         or1200_cpu_or1200_except_n1755, or1200_cpu_or1200_except_n1754,
         or1200_cpu_or1200_except_n1753, or1200_cpu_or1200_except_n1751,
         or1200_cpu_or1200_except_n1750, or1200_cpu_or1200_except_n1749,
         or1200_cpu_or1200_except_n1748, or1200_cpu_or1200_except_n1747,
         or1200_cpu_or1200_except_n1746, or1200_cpu_or1200_except_n1745,
         or1200_cpu_or1200_except_n1744, or1200_cpu_or1200_except_n1743,
         or1200_cpu_or1200_except_n1742, or1200_cpu_or1200_except_n1741,
         or1200_cpu_or1200_except_n1740, or1200_cpu_or1200_except_n1739,
         or1200_cpu_or1200_except_n1738, or1200_cpu_or1200_except_n1736,
         or1200_cpu_or1200_except_n1735, or1200_cpu_or1200_except_n1734,
         or1200_cpu_or1200_except_n1733, or1200_cpu_or1200_except_n1732,
         or1200_cpu_or1200_except_n1731, or1200_cpu_or1200_except_n1730,
         or1200_cpu_or1200_except_n1729, or1200_cpu_or1200_except_n1728,
         or1200_cpu_or1200_except_n1727, or1200_cpu_or1200_except_n1726,
         or1200_cpu_or1200_except_n1725, or1200_cpu_or1200_except_n1724,
         or1200_cpu_or1200_except_n1723, or1200_cpu_or1200_except_n1722,
         or1200_cpu_or1200_except_n1721, or1200_cpu_or1200_except_n1720,
         or1200_cpu_or1200_except_n1719, or1200_cpu_or1200_except_n1718,
         or1200_cpu_or1200_except_n1717, or1200_cpu_or1200_except_n1716,
         or1200_cpu_or1200_except_n1715, or1200_cpu_or1200_except_n1714,
         or1200_cpu_or1200_except_n1713, or1200_cpu_or1200_except_n1712,
         or1200_cpu_or1200_except_n1711, or1200_cpu_or1200_except_n1710,
         or1200_cpu_or1200_except_n1709, or1200_cpu_or1200_except_n1708,
         or1200_cpu_or1200_except_n1707, or1200_cpu_or1200_except_n1706,
         or1200_cpu_or1200_except_n1705, or1200_cpu_or1200_except_n1704,
         or1200_cpu_or1200_except_n1703, or1200_cpu_or1200_except_n1702,
         or1200_cpu_or1200_except_n1701, or1200_cpu_or1200_except_n1700,
         or1200_cpu_or1200_except_n1699, or1200_cpu_or1200_except_n1697,
         or1200_cpu_or1200_except_n1696, or1200_cpu_or1200_except_n1694,
         or1200_cpu_or1200_except_n691, or1200_cpu_or1200_except_n690,
         or1200_cpu_or1200_except_n687, or1200_cpu_or1200_except_n685,
         or1200_cpu_or1200_except_n684, or1200_cpu_or1200_except_n682,
         or1200_cpu_or1200_except_n681, or1200_cpu_or1200_except_n679,
         or1200_cpu_or1200_except_n677, or1200_cpu_or1200_except_n671,
         or1200_cpu_or1200_except_n670, or1200_cpu_or1200_except_n668,
         or1200_cpu_or1200_except_n667, or1200_cpu_or1200_except_n665,
         or1200_cpu_or1200_except_n664, or1200_cpu_or1200_except_n662,
         or1200_cpu_or1200_except_n661, or1200_cpu_or1200_except_n659,
         or1200_cpu_or1200_except_n658, or1200_cpu_or1200_except_n656,
         or1200_cpu_or1200_except_n655, or1200_cpu_or1200_except_n653,
         or1200_cpu_or1200_except_n652, or1200_cpu_or1200_except_n650,
         or1200_cpu_or1200_except_n649, or1200_cpu_or1200_except_n647,
         or1200_cpu_or1200_except_n646, or1200_cpu_or1200_except_n644,
         or1200_cpu_or1200_except_n643, or1200_cpu_or1200_except_n641,
         or1200_cpu_or1200_except_n640, or1200_cpu_or1200_except_n638,
         or1200_cpu_or1200_except_n637, or1200_cpu_or1200_except_n635,
         or1200_cpu_or1200_except_n634, or1200_cpu_or1200_except_n632,
         or1200_cpu_or1200_except_n631, or1200_cpu_or1200_except_n629,
         or1200_cpu_or1200_except_n628, or1200_cpu_or1200_except_n626,
         or1200_cpu_or1200_except_n625, or1200_cpu_or1200_except_n623,
         or1200_cpu_or1200_except_n622, or1200_cpu_or1200_except_n620,
         or1200_cpu_or1200_except_n619, or1200_cpu_or1200_except_n617,
         or1200_cpu_or1200_except_n616, or1200_cpu_or1200_except_n614,
         or1200_cpu_or1200_except_n613, or1200_cpu_or1200_except_n611,
         or1200_cpu_or1200_except_n610, or1200_cpu_or1200_except_n608,
         or1200_cpu_or1200_except_n607, or1200_cpu_or1200_except_n605,
         or1200_cpu_or1200_except_n604, or1200_cpu_or1200_except_n602,
         or1200_cpu_or1200_except_n601, or1200_cpu_or1200_except_n599,
         or1200_cpu_or1200_except_n598, or1200_cpu_or1200_except_n596,
         or1200_cpu_or1200_except_n595, or1200_cpu_or1200_except_n593,
         or1200_cpu_or1200_except_n592, or1200_cpu_or1200_except_n590,
         or1200_cpu_or1200_except_n589, or1200_cpu_or1200_except_n587,
         or1200_cpu_or1200_except_n586, or1200_cpu_or1200_except_n584,
         or1200_cpu_or1200_except_n583, or1200_cpu_or1200_except_n575,
         or1200_cpu_or1200_except_n571, or1200_cpu_or1200_except_n567,
         or1200_cpu_or1200_except_n565, or1200_cpu_or1200_except_n563,
         or1200_cpu_or1200_except_n561, or1200_cpu_or1200_except_n555,
         or1200_cpu_or1200_except_n553, or1200_cpu_or1200_except_n552,
         or1200_cpu_or1200_except_n550, or1200_cpu_or1200_except_n548,
         or1200_cpu_or1200_except_n546, or1200_cpu_or1200_except_n544,
         or1200_cpu_or1200_except_n542, or1200_cpu_or1200_except_n540,
         or1200_cpu_or1200_except_n538, or1200_cpu_or1200_except_n536,
         or1200_cpu_or1200_except_n534, or1200_cpu_or1200_except_n532,
         or1200_cpu_or1200_except_n530, or1200_cpu_or1200_except_n528,
         or1200_cpu_or1200_except_n526, or1200_cpu_or1200_except_n524,
         or1200_cpu_or1200_except_n522, or1200_cpu_or1200_except_n520,
         or1200_cpu_or1200_except_n518, or1200_cpu_or1200_except_n516,
         or1200_cpu_or1200_except_n514, or1200_cpu_or1200_except_n512,
         or1200_cpu_or1200_except_n510, or1200_cpu_or1200_except_n508,
         or1200_cpu_or1200_except_n506, or1200_cpu_or1200_except_n504,
         or1200_cpu_or1200_except_n502, or1200_cpu_or1200_except_n500,
         or1200_cpu_or1200_except_n498, or1200_cpu_or1200_except_n496,
         or1200_cpu_or1200_except_n494, or1200_cpu_or1200_except_n492,
         or1200_cpu_or1200_except_n486, or1200_cpu_or1200_except_n483,
         or1200_cpu_or1200_except_n482, or1200_cpu_or1200_except_n480,
         or1200_cpu_or1200_except_n477, or1200_cpu_or1200_except_n476,
         or1200_cpu_or1200_except_n474, or1200_cpu_or1200_except_n471,
         or1200_cpu_or1200_except_n468, or1200_cpu_or1200_except_n467,
         or1200_cpu_or1200_except_n465, or1200_cpu_or1200_except_n462,
         or1200_cpu_or1200_except_n461, or1200_cpu_or1200_except_n459,
         or1200_cpu_or1200_except_n456, or1200_cpu_or1200_except_n453,
         or1200_cpu_or1200_except_n450, or1200_cpu_or1200_except_n447,
         or1200_cpu_or1200_except_n446, or1200_cpu_or1200_except_n444,
         or1200_cpu_or1200_except_n441, or1200_cpu_or1200_except_n440,
         or1200_cpu_or1200_except_n438, or1200_cpu_or1200_except_n437,
         or1200_cpu_or1200_except_n435, or1200_cpu_or1200_except_n434,
         or1200_cpu_or1200_except_n432, or1200_cpu_or1200_except_n431,
         or1200_cpu_or1200_except_n429, or1200_cpu_or1200_except_n428,
         or1200_cpu_or1200_except_n426, or1200_cpu_or1200_except_n425,
         or1200_cpu_or1200_except_n423, or1200_cpu_or1200_except_n422,
         or1200_cpu_or1200_except_n420, or1200_cpu_or1200_except_n419,
         or1200_cpu_or1200_except_n417, or1200_cpu_or1200_except_n416,
         or1200_cpu_or1200_except_n414, or1200_cpu_or1200_except_n413,
         or1200_cpu_or1200_except_n411, or1200_cpu_or1200_except_n410,
         or1200_cpu_or1200_except_n408, or1200_cpu_or1200_except_n407,
         or1200_cpu_or1200_except_n405, or1200_cpu_or1200_except_n404,
         or1200_cpu_or1200_except_n402, or1200_cpu_or1200_except_n401,
         or1200_cpu_or1200_except_n399, or1200_cpu_or1200_except_n398,
         or1200_cpu_or1200_except_n390, or1200_cpu_or1200_except_n389,
         or1200_cpu_or1200_except_n387, or1200_cpu_or1200_except_n386,
         or1200_cpu_or1200_except_n384, or1200_cpu_or1200_except_n383,
         or1200_cpu_or1200_except_n381, or1200_cpu_or1200_except_n380,
         or1200_cpu_or1200_except_n378, or1200_cpu_or1200_except_n377,
         or1200_cpu_or1200_except_n375, or1200_cpu_or1200_except_n374,
         or1200_cpu_or1200_except_n372, or1200_cpu_or1200_except_n371,
         or1200_cpu_or1200_except_n369, or1200_cpu_or1200_except_n368,
         or1200_cpu_or1200_except_n366, or1200_cpu_or1200_except_n365,
         or1200_cpu_or1200_except_n363, or1200_cpu_or1200_except_n362,
         or1200_cpu_or1200_except_n360, or1200_cpu_or1200_except_n359,
         or1200_cpu_or1200_except_n357, or1200_cpu_or1200_except_n356,
         or1200_cpu_or1200_except_n354, or1200_cpu_or1200_except_n353,
         or1200_cpu_or1200_except_n351, or1200_cpu_or1200_except_n350,
         or1200_cpu_or1200_except_n348, or1200_cpu_or1200_except_n347,
         or1200_cpu_or1200_except_n345, or1200_cpu_or1200_except_n344,
         or1200_cpu_or1200_except_n342, or1200_cpu_or1200_except_n341,
         or1200_cpu_or1200_except_n339, or1200_cpu_or1200_except_n338,
         or1200_cpu_or1200_except_n336, or1200_cpu_or1200_except_n335,
         or1200_cpu_or1200_except_n333, or1200_cpu_or1200_except_n332,
         or1200_cpu_or1200_except_n330, or1200_cpu_or1200_except_n329,
         or1200_cpu_or1200_except_n327, or1200_cpu_or1200_except_n326,
         or1200_cpu_or1200_except_n324, or1200_cpu_or1200_except_n323,
         or1200_cpu_or1200_except_n321, or1200_cpu_or1200_except_n320,
         or1200_cpu_or1200_except_n318, or1200_cpu_or1200_except_n317,
         or1200_cpu_or1200_except_n315, or1200_cpu_or1200_except_n314,
         or1200_cpu_or1200_except_n312, or1200_cpu_or1200_except_n311,
         or1200_cpu_or1200_except_n309, or1200_cpu_or1200_except_n308,
         or1200_cpu_or1200_except_n306, or1200_cpu_or1200_except_n305,
         or1200_cpu_or1200_except_n303, or1200_cpu_or1200_except_n302,
         or1200_cpu_or1200_except_n294, or1200_cpu_or1200_except_n292,
         or1200_cpu_or1200_except_n290, or1200_cpu_or1200_except_n288,
         or1200_cpu_or1200_except_n286, or1200_cpu_or1200_except_n283,
         or1200_cpu_or1200_except_n282, or1200_cpu_or1200_except_n280,
         or1200_cpu_or1200_except_n278, or1200_cpu_or1200_except_n276,
         or1200_cpu_or1200_except_n274, or1200_cpu_or1200_except_n272,
         or1200_cpu_or1200_except_n270, or1200_cpu_or1200_except_n268,
         or1200_cpu_or1200_except_n266, or1200_cpu_or1200_except_n264,
         or1200_cpu_or1200_except_n262, or1200_cpu_or1200_except_n260,
         or1200_cpu_or1200_except_n258, or1200_cpu_or1200_except_n256,
         or1200_cpu_or1200_except_n253, or1200_cpu_or1200_except_n252,
         or1200_cpu_or1200_except_n248, or1200_cpu_or1200_except_n246,
         or1200_cpu_or1200_except_n244, or1200_cpu_or1200_except_n242,
         or1200_cpu_or1200_except_n240, or1200_cpu_or1200_except_n238,
         or1200_cpu_or1200_except_n236, or1200_cpu_or1200_except_n234,
         or1200_cpu_or1200_except_n232, or1200_cpu_or1200_except_n230,
         or1200_cpu_or1200_except_n228, or1200_cpu_or1200_except_n226,
         or1200_cpu_or1200_except_n224, or1200_cpu_or1200_except_n222,
         or1200_cpu_or1200_except_n220, or1200_cpu_or1200_except_n218,
         or1200_cpu_or1200_except_n216, or1200_cpu_or1200_except_n214,
         or1200_cpu_or1200_except_n212, or1200_cpu_or1200_except_n210,
         or1200_cpu_or1200_except_n208, or1200_cpu_or1200_except_n206,
         or1200_cpu_or1200_except_n204, or1200_cpu_or1200_except_n202,
         or1200_cpu_or1200_except_n200, or1200_cpu_or1200_except_n198,
         or1200_cpu_or1200_except_n196, or1200_cpu_or1200_except_n194,
         or1200_cpu_or1200_except_n192, or1200_cpu_or1200_except_n188,
         or1200_cpu_or1200_except_n186, or1200_cpu_or1200_except_n184,
         or1200_cpu_or1200_except_n182, or1200_cpu_or1200_except_n180,
         or1200_cpu_or1200_except_n178, or1200_cpu_or1200_except_n176,
         or1200_cpu_or1200_except_n174, or1200_cpu_or1200_except_n172,
         or1200_cpu_or1200_except_n170, or1200_cpu_or1200_except_n168,
         or1200_cpu_or1200_except_n166, or1200_cpu_or1200_except_n164,
         or1200_cpu_or1200_except_n162, or1200_cpu_or1200_except_n160,
         or1200_cpu_or1200_except_n158, or1200_cpu_or1200_except_n156,
         or1200_cpu_or1200_except_n154, or1200_cpu_or1200_except_n152,
         or1200_cpu_or1200_except_n150, or1200_cpu_or1200_except_n148,
         or1200_cpu_or1200_except_n146, or1200_cpu_or1200_except_n144,
         or1200_cpu_or1200_except_n142, or1200_cpu_or1200_except_n140,
         or1200_cpu_or1200_except_n138, or1200_cpu_or1200_except_n136,
         or1200_cpu_or1200_except_n134, or1200_cpu_or1200_except_n132,
         or1200_cpu_or1200_except_n130, or1200_cpu_or1200_except_n128,
         or1200_cpu_or1200_except_n126, or1200_cpu_or1200_except_n124,
         or1200_cpu_or1200_except_n122, or1200_cpu_or1200_except_n120,
         or1200_cpu_or1200_except_n116,
         or1200_cpu_or1200_except_ex_freeze_prev,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n137,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n136,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n135,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n134,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n133,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n132,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n131,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n130,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n129,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n128,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n127,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n126,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n125,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n124,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n123,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n122,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n121,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n120,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n119,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n118,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n117,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n116,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n115,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n114,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n113,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n112,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n111,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n110,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n109,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n108,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n106,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n105,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n103,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n102,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n101,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n100,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n99,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n98,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n97,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n96,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n95,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n94,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n93,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n92,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n91,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n90,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n89,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n88,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n87,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n86,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n85,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n84,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n83,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n82,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n81,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n80,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n79,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n78,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n77,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n76,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n75,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n74,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n73,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n72,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n71,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n70,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n69,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n68,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n67,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n66,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n65,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n64,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n63,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n62,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n61,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n60,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n59,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n58,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n57,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n56,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n55,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n54,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n53,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n52,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n51,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n50,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n49,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n48,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n47,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n46,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n45,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n44,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n43,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n42,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n41,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n40,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n39,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n38,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n37,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n36,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n35,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n34,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n33,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n32,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n31,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n30,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n29,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n27,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n26,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n25,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n23,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n22,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n21,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n19,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n18,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n17,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n15,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n14,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n13,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n11,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n10,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n9,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n7,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n6,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n5,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n4,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n3,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n2,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n1,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_N2648,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_25_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_26_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_27_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_28_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_29_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_30_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_31_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_32_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_33_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_34_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_35_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_36_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_37_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_38_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_39_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_40_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_41_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_42_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_43_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_44_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_45_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_47_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_N2435,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_output_o_31_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_25_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_32_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_33_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_35_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_36_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_37_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n254,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n253,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n252,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n251,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n250,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n249,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n248,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n244,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n241,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n238,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n235,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n232,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n229,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n226,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n223,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n220,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n217,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n214,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n211,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n208,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n205,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n202,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n199,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n196,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n193,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n190,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n187,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n184,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n181,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n178,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n175,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n172,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n169,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n166,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n163,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n160,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n157,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n154,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n151,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n148,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n145,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n142,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n139,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n136,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n133,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n130,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n127,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n124,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n121,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n118,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n115,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n112,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n109,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n106,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n103,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_state,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_0_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_1_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_2_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_3_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_4_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_5_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_6_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_7_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_8_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_9_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_10_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_11_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_12_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_13_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_14_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_15_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_16_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_17_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_18_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_19_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_20_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_21_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_22_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_23_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_24_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_25_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_26_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_27_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_28_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_29_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_30_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_31_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_32_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_33_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_34_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_35_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_36_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_37_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_38_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_39_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_40_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_41_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_42_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_43_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_44_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_45_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_46_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_47_,
         or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_start_i,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n63,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n62,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n61,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n60,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n59,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n58,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n57,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n56,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n55,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n54,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n53,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n52,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n51,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n50,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n49,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n48,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n47,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n46,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n45,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n44,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n43,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n42,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n41,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n40,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n39,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n38,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n37,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n36,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n35,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n34,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n33,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n32,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n31,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n30,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n29,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n28,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n27,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n26,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n25,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n24,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n23,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n22,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n21,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n20,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n19,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n18,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n17,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n16,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n15,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n14,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n13,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n12,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n11,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n10,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n9,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n8,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n7,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n6,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n5,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n4,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n3,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n2,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n1,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_N398,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_0_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_2_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_3_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_4_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_5_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_6_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_7_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_8_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_9_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_10_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_11_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_12_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_13_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_14_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_15_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_16_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_17_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_18_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_19_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_20_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_21_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_22_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_23_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_24_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_in_00,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_0_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_2_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_3_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_4_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_5_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_6_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_7_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_8_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_9_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_10_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_11_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_12_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_13_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_14_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_15_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_16_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_17_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_18_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_19_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_20_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_21_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_22_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_0_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_2_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_3_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_4_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_5_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_6_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_7_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_1_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_2_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_3_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_4_,
         or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_5_, n27027, n27028,
         n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036,
         n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
         n27045, n27046, n27047, n27066, n27067, n27068, n27069, n27070,
         n27071, n27072, n27073, n27074, n27075, n27100, n27324, n27420,
         n27421, n27433, n27447, n27448, n27456, n27472, n27477, n27495,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27531, n27532, n27533, n27534, n27535,
         n27536, n27627, n27713, n27721, n27728, n27729, n27731, n27733,
         n27735, n27738, n27977, n27978, n27979, n27980, n27981, n27982,
         n28105, n28158, n28160, n28161, n28162, n28163, n28164, n28165,
         n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173,
         n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181,
         n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189,
         n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197,
         n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205,
         n28206, n28207, n28208, n28210, n28213, n28256, n51945, n51946,
         n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954,
         n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962,
         n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970,
         n51971, n51972, n51973, n51974, n51975, n51976, n51978, n51979,
         n51980, n51981, n51982, n51985, n51986, n51987, n51988, n51990,
         n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998,
         n51999, n52000, n52001, n52003, n52004, n52005, n52006, n52007,
         n52008, n52009, n52010, n52011, n52012, n52013, n52014, n52047,
         n52048, n52049, n52050, n52051, n52052, n52053, n52054, n52055,
         n52056, n52057, n52058, n52059, n52060, n52061, n52469, n52470,
         n52471, n52472, n52473, n52474, n52475, n52484, n52485, n52486,
         n52489, n52490, n52491, n52492, n52493, n52494, n52496, n52497,
         n52498, n52499, n52500, n52501, n52502, n52503, n52504, n52505,
         n52506, n52507, n52508, n52509, n52517, n52518, n52519, n52520,
         n52521, n52522, n52523, n52524, n52526, n52545, n52546, n52547,
         n52549, n53175, n53176, n53189, n53190, n53191, n53192, n53193,
         n53194, n53195, n53196, n53197, n53198, n53199, n53200, n53201,
         n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209,
         n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217,
         n53218, n53219, n53220, n53221, n53222, n53223, n53224, n53225,
         n53226, n53227, n53228, n53229, n53230, n53231, n53232, n53233,
         n53234, n53235, n53236, n53237, n53238, n53239, n53240, n53241,
         n53242, n53243, n53244, n53245, n53246, n53247, n53248, n53249,
         n53250, n53251, n53252, n53253, n53254, n53255, n53256, n53257,
         n53258, n53259, n53260, n53261, n53262, n53263, n53264, n53265,
         n53266, n53267, n53268, n53269, n53270, n53271, n53272, n53273,
         n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281,
         n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289,
         n53290, n53291, n53292, n53293, n53294, n53295, n53296, n53297,
         n53298, n53299, n53300, n53301, n53302, n53303, n53304, n53305,
         n53306, n53307, n53308, n53309, n53310, n53311, n53312, n53313,
         n53314, n53315, n53316, n53317, n53318, n53319, n53320, n53321,
         n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329,
         n53330, n53331, n53332, n53333, n53334, n53335, n53336, n53337,
         n53338, n53339, n53340, n53341, n53342, n53343, n53344, n53345,
         n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353,
         n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361,
         n53362, n53363, n53364, n53365, n53366, n53367, n53368, n53369,
         n53370, n53371, n53372, n53373, n53374, n53375, n53376, n53377,
         n53378, n53379, n53380, n53381, n53382, n53383, n53384, n53385,
         n53386, n53387, n53388, n53389, n53390, n53391, n53392, n53393,
         n53394, n53395, n53396, n53397, n53398, n53399, n53400, n53401,
         n53402, n53403, n53404, n53405, n53406, n53407, n53408, n53409,
         n53410, n53411, n53412, n53413, n53414, n53415, n53416, n53417,
         n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425,
         n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433,
         n53434, n53435, n53436, n53437, n53438, n53439, n53440, n53441,
         n53442, n53443, n53444, n53445, n53446, n53447, n53448, n53449,
         n53450, n53451, n53452, n53453, n53454, n53455, n53456, n53457,
         n53458, n53459, n53460, n53461, n53462, n53463, n53464, n53465,
         n53466, n53467, n53468, n53469, n53470, n53471, n53472, n53473,
         n53474, n53475, n53476, n53477, n53478, n53479, n53480, n53481,
         n53482, n53483, n53484, n53485, n53486, n53487, n53488, n53489,
         n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497,
         n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505,
         n53506, n53507, n53508, n53509, n53510, n53511, n53512, n53513,
         n53514, n53515, n53516, n53517, n53518, n53519, n53520, n53521,
         n53522, n53523, n53524, n53525, n53526, n53527, n53528, n53529,
         n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537,
         n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545,
         n53546, n53547, n53548, n53549, n53550, n53551, n53552, n53553,
         n53554, n53555, n53556, n53557, n53558, n53559, n53560, n53561,
         n53562, n53563, n53564, n53565, n53566, n53567, n53568, n53569,
         n53570, n53571, n53572, n53573, n53574, n53575, n53576, n53577,
         n53578, n53579, n53580, n53581, n53582, n53583, n53584, n53585,
         n53586, n53587, n53588, n53589, n53590, n53591, n53592, n53593,
         n53594, n53595, n53596, n53597, n53598, n53599, n53600, n53601,
         n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609,
         n53610, n53611, n53612, n53613, n53614, n53615, n53616, n53617,
         n53618, n53619, n53620, n53621, n53622, n53623, n53624, n53625,
         n53626, n53627, n53628, n53629, n53630, n53631, n53632, n53633,
         n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641,
         n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649,
         n53650, n53651, n53652, n53653, n53654, n53655, n53656, n53657,
         n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665,
         n53666, n53667, n53668, n53669, n53670, n53671, n53672, n53673,
         n53674, n53675, n53676, n53677, n53678, n53679, n53680, n53681,
         n53682, n53683, n53684, n53685, n53686, n53687, n53688, n53689,
         n53690, n53691, n53692, n53693, n53694, n53695, n53696, n53697,
         n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705,
         n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713,
         n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721,
         n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729,
         n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737,
         n53738, n53739, n53740, n53741, n53742, n53743, n53744, n53745,
         n53746, n53747, n53748, n53749, n53750, n53751, n53752, n53753,
         n53754, n53755, n53756, n53757, n53758, n53759, n53760, n53761,
         n53762, n53763, n53764, n53765, n53766, n53767, n53768, n53769,
         n53770, n53771, n53772, n53773, n53774, n53775, n53776, n53777,
         n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785,
         n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793,
         n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801,
         n53802, n53803, n53804, n53805, n53806, n53807, n53808, n53809,
         n53810, n53811, n53812, n53813, n53814, n53815, n53816, n53817,
         n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825,
         n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833,
         n53834, n53835, n53836, n53837, n53838, n53839, n53840, n53841,
         n53842, n53843, n53844, n53845, n53846, n53847, n53848, n53849,
         n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857,
         n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865,
         n53866, n53867, n53868, n53869, n53870, n53871, n53872, n53873,
         n53874, n53875, n53876, n53877, n53878, n53879, n53880, n53881,
         n53882, n53883, n53884, n53885, n53886, n53887, n53888, n53889,
         n53890, n53891, n53892, n53893, n53894, n53895, n53896, n53897,
         n53898, n53899, n53900, n53901, n53902, n53903, n53904, n53905,
         n53906, n53907, n53908, n53909, n53910, n53911, n53912, n53913,
         n53914, n53915, n53916, n53917, n53918, n53919, n53920, n53921,
         n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929,
         n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937,
         n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945,
         n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953,
         n53954, n53955, n53956, n53957, n53958, n53959, n53960, n53961,
         n53962, n53963, n53964, n53965, n53966, n53967, n53968, n53969,
         n53970, n53971, n53972, n53973, n53974, n53975, n53976, n53977,
         n53978, n53979, n53980, n53981, n53982, n53983, n53984, n53985,
         n53986, n53987, n53988, n53989, n53990, n53991, n53992, n53993,
         n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001,
         n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009,
         n54010, n54011, n54012, n54013, n54014, n54015, n54016, n54017,
         n54018, n54019, n54020, n54021, n54022, n54023, n54024, n54025,
         n54026, n54027, n54028, n54029, n54030, n54031, n54032, n54033,
         n54034, n54035, n54036, n54037, n54038, n54039, n54040, n54041,
         n54042, n54043, n54044, n54045, n54046, n54047, n54048, n54049,
         n54050, n54051, n54052, n54053, n54054, n54055, n54056, n54057,
         n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065,
         n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073,
         n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081,
         n54082, n54083, n54084, n54085, n54086, n54087, n54088, n54089,
         n54090, n54091, n54092, n54093, n54094, n54095, n54096, n54097,
         n54098, n54099, n54100, n54101, n54102, n54103, n54104, n54105,
         n54106, n54107, n54108, n54109, n54110, n54111, n54112, n54113,
         n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121,
         n54122, n54123, n54124, n54125, n54126, n54127, n54128, n54129,
         n54130, n54131, n54132, n54133, n54134, n54135, n54136, n54137,
         n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145,
         n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153,
         n54154, n54155, n54156, n54157, n54158, n54159, n54160, n54161,
         n54162, n54163, n54164, n54165, n54166, n54167, n54168, n54169,
         n54170, n54171, n54172, n54173, n54174, n54175, n54176, n54177,
         n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185,
         n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193,
         n54194, n54195, n54196, n54197, n54198, n54199, n54200, n54201,
         n54202, n54203, n54204, n54205, n54206, n54207, n54208, n54209,
         n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217,
         n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225,
         n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233,
         n54234, n54235, n54236, n54237, n54238, n54239, n54240, n54241,
         n54242, n54243, n54244, n54245, n54246, n54247, n54248, n54249,
         n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257,
         n54258, n54259, n54260, n54261, n54262, n54263, n54264, n54265,
         n54266, n54267, n54268, n54269, n54270, n54271, n54272, n54273,
         n54274, n54275, n54276, n54277, n54278, n54279, n54280, n54281,
         n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289,
         n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297,
         n54298, n54299, n54300, n54301, n54302, n54303, n54304, n54305,
         n54306, n54307, n54308, n54309, n54310, n54311, n54312, n54313,
         n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321,
         n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329,
         n54330, n54331, n54332, n54333, n54334, n54335, n54336, n54337,
         n54338, n54339, n54340, n54341, n54342, n54343, n54344, n54345,
         n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353,
         n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361,
         n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369,
         n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377,
         n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385,
         n54386, n54387, n54388, n54389, n54390, n54391, n54392, n54393,
         n54394, n54395, n54396, n54397, n54398, n54399, n54400, n54401,
         n54402, n54403, n54404, n54405, n54406, n54407, n54408, n54409,
         n54410, n54411, n54412, n54413, n54414, n54415, n54416, n54417,
         n54418, n54419, n54420, n54421, n54422, n54423, n54424, n54425,
         n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433,
         n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441,
         n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449,
         n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457,
         n54458, n54459, n54460, n54461, n54462, n54463, n54464, n54465,
         n54466, n54467, n54468, n54469, n54470, n54471, n54472, n54473,
         n54474, n54475, n54476, n54477, n54478, n54479, n54480, n54481,
         n54482, n54483, n54484, n54485, n54486, n54487, n54488, n54489,
         n54490, n54491, n54492, n54493, n54494, n54495, n54496, n54497,
         n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505,
         n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513,
         n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521,
         n54522, n54523, n54524, n54525, n54526, n54527, n54528, n54529,
         n54530, n54531, n54532, n54533, n54534, n54535, n54536, n54537,
         n54538, n54539, n54540, n54541, n54542, n54543, n54544, n54545,
         n54546, n54547, n54548, n54549, n54550, n54551, n54552, n54553,
         n54554, n54555, n54556, n54557, n54558, n54559, n54560, n54561,
         n54562, n54563, n54564, n54565, n54566, n54567, n54568, n54569,
         n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577,
         n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585,
         n54586, n54587, n54588, n54589, n54590, n54591, n54592, n54593,
         n54594, n54595, n54596, n54597, n54598, n54599, n54600, n54601,
         n54602, n54603, n54604, n54605, n54606, n54607, n54608, n54609,
         n54610, n54611, n54612, n54613, n54614, n54615, n54616, n54617,
         n54618, n54619, n54620, n54621, n54622, n54623, n54624, n54625,
         n54626, n54627, n54628, n54629, n54630, n54631, n54632, n54633,
         n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641,
         n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649,
         n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657,
         n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665,
         n54666, n54667, n54668, n54669, n54670, n54671, n54672, n54673,
         n54674, n54675, n54676, n54677, n54678, n54679, n54680, n54681,
         n54682, n54683, n54684, n54685, n54686, n54687, n54688, n54689,
         n54690, n54691, n54692, n54693, n54694, n54695, n54696, n54697,
         n54698, n54699, n54700, n54701, n54702, n54703, n54704, n54705,
         n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713,
         n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721,
         n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729,
         n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737,
         n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745,
         n54746, n54747, n54748, n54749, n54750, n54751, n54752, n54753,
         n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761,
         n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769,
         n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777,
         n54778, n54779, n54780, n54781, n54782, n54783, n54784, n54785,
         n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793,
         n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801,
         n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809,
         n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817,
         n54818, n54819, n54820, n54821, n54822, n54823, n54824, n54825,
         n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833,
         n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841,
         n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849,
         n54850, n54851, n54852, n54853, n54854, n54855, n54856, n54857,
         n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865,
         n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873,
         n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881,
         n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889,
         n54890, n54891, n54892, n54893, n54894, n54895, n54896, n54897,
         n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905,
         n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913,
         n54914, n54915, n54916, n54917, n54918, n54919, n54920, n54921,
         n54922, n54923, n54924, n54925, n54926, n54927, n54928, n54929,
         n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937,
         n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945,
         n54946, n54947, n54948, n54949, n54950, n54951, n54952, n54953,
         n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961,
         n54962, n54963, n54964, n54965, n54966, n54967, n54968, n54969,
         n54970, n54971, n54972, n54973, n54974, n54975, n54976, n54977,
         n54978, n54979, n54980, n54981, n54982, n54983, n54984, n54985,
         n54986, n54987, n54988, n54989, n54990, n54991, n54992, n54993,
         n54994, n54995, n54996, n54997, n54998, n54999, n55000, n55001,
         n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009,
         n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017,
         n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025,
         n55026, n55027, n55028, n55029, n55030, n55031, n55032, n55033,
         n55034, n55035, n55036, n55037, n55038, n55039, n55040, n55041,
         n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049,
         n55050, n55051, n55052, n55053, n55054, n55055, n55056, n55057,
         n55058, n55059, n55060, n55061, n55062, n55063, n55064, n55065,
         n55066, n55067, n55068, n55069, n55070, n55071, n55072, n55073,
         n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081,
         n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089,
         n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097,
         n55098, n55099, n55100, n55101, n55102, n55103, n55104, n55105,
         n55106, n55107, n55108, n55109, n55110, n55111, n55112, n55113,
         n55114, n55115, n55116, n55117, n55118, n55119, n55120, n55121,
         n55122, n55123, n55124, n55125, n55126, n55127, n55128, n55129,
         n55130, n55131, n55132, n55133, n55134, n55135, n55136, n55137,
         n55138, n55139, n55140, n55141, n55142, n55143, n55144, n55145,
         n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153,
         n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161,
         n55162, n55163, n55164, n55165, n55166, n55167, n55168, n55169,
         n55170, n55171, n55172, n55173, n55174, n55175, n55176, n55177,
         n55178, n55179, n55180, n55181, n55182, n55183, n55184, n55185,
         n55186, n55187, n55188, n55189, n55190, n55191, n55192, n55193,
         n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201,
         n55202, n55203, n55204, n55205, n55206, n55207, n55208, n55209,
         n55210, n55211, n55212, n55213, n55214, n55215, n55216, n55217,
         n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225,
         n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233,
         n55234, n55235, n55236, n55237, n55238, n55239, n55240, n55241,
         n55242, n55243, n55244, n55245, n55246, n55247, n55248, n55249,
         n55250, n55251, n55252, n55253, n55254, n55255, n55256, n55257,
         n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265,
         n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273,
         n55274, n55275, n55276, n55277, n55278, n55279, n55280, n55281,
         n55282, n55283, n55284, n55285, n55286, n55287, n55288, n55289,
         n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297,
         n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305,
         n55306, n55307, n55308, n55309, n55310, n55311, n55312, n55313,
         n55314, n55315, n55316, n55317, n55318, n55319, n55320, n55321,
         n55322, n55323, n55324, n55325, n55326, n55327, n55328, n55329,
         n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337,
         n55338, n55339, n55340, n55341, n55342, n55343, n55344, n55345,
         n55346, n55347, n55348, n55349, n55350, n55351, n55352, n55353,
         n55354, n55355, n55356, n55357, n55358, n55359, n55360, n55361,
         n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369,
         n55370, n55371, n55372, n55373, n55374, n55375, n55376, n55377,
         n55378, n55379, n55380, n55381, n55382, n55383, n55384, n55385,
         n55386, n55387, n55388, n55389, n55390, n55391, n55392, n55393,
         n55394, n55395, n55396, n55397, n55398, n55399, n55400, n55401,
         n55402, n55403, n55404, n55405, n55406, n55407, n55408, n55409,
         n55410, n55411, n55412, n55413, n55414, n55415, n55416, n55417,
         n55418, n55419, n55420, n55421, n55422, n55423, n55424, n55425,
         n55426, n55427, n55428, n55429, n55430, n55431, n55432, n55433,
         n55434, n55435, n55436, n55437, n55438, n55439, n55440, n55441,
         n55442, n55443, n55444, n55445, n55446, n55447, n55448, n55449,
         n55450, n55451, n55452, n55453, n55454, n55455, n55456, n55457,
         n55458, n55459, n55460, n55461, n55462, n55463, n55464, n55465,
         n55466, n55467, n55468, n55469, n55470, n55471, n55472, n55473,
         n55474, n55475, n55476, n55477, n55478, n55479, n55480, n55481,
         n55482, n55483, n55484, n55485, n55486, n55487, n55488, n55489,
         n55490, n55491, n55492, n55493, n55494, n55495, n55496, n55497,
         n55498, n55499, n55500, n55501, n55502, n55503, n55504, n55505,
         n55506, n55507, n55508, n55509, n55510, n55511, n55512, n55513,
         n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521,
         n55522, n55523, n55524, n55525, n55526, n55527, n55528, n55529,
         n55530, n55531, n55532, n55533, n55534, n55535, n55536, n55537,
         n55538, n55539, n55540, n55541, n55542, n55543, n55544, n55545,
         n55546, n55547, n55548, n55549, n55550, n55551, n55552, n55553,
         n55554, n55555, n55556, n55557, n55558, n55559, n55560, n55561,
         n55562, n55563, n55564, n55565, n55566, n55567, n55568, n55569,
         n55570, n55571, n55572, n55573, n55574, n55575, n55576, n55577,
         n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585,
         n55586, n55587, n55588, n55589, n55590, n55591, n55592, n55593,
         n55594, n55595, n55596, n55597, n55598, n55599, n55600, n55601,
         n55602, n55603, n55604, n55605, n55606, n55607, n55608, n55609,
         n55610, n55611, n55612, n55613, n55614, n55615, n55616, n55617,
         n55618, n55619, n55620, n55621, n55622, n55623, n55624, n55625,
         n55626, n55627, n55628, n55629, n55630, n55631, n55632, n55633,
         n55634, n55635, n55636, n55637, n55638, n55639, n55640, n55641,
         n55642, n55643, n55644, n55645, n55646, n55647, n55648, n55649,
         n55650, n55651, n55652, n55653, n55654, n55655, n55656, n55657,
         n55658, n55659, n55660, n55661, n55662, n55663, n55664, n55665,
         n55666, n55667, n55668, n55669, n55670, n55671, n55672, n55673,
         n55674, n55675, n55676, n55677, n55678, n55679, n55680, n55681,
         n55682, n55683, n55684, n55685, n55686, n55687, n55688, n55689,
         n55690, n55691, n55692, n55693, n55694, n55695, n55696, n55697,
         n55698, n55699, n55700, n55701, n55702, n55703, n55704, n55705,
         n55706, n55707, n55708, n55709, n55710, n55711, n55712, n55713,
         n55714, n55715, n55716, n55717, n55718, n55719, n55720, n55721,
         n55722, n55723, n55724, n55725, n55726, n55727, n55728, n55729,
         n55730, n55731, n55732, n55733, n55734, n55735, n55736, n55737,
         n55738, n55739, n55740, n55741, n55742, n55743, n55744, n55745,
         n55746, n55747, n55748, n55749, n55750, n55751, n55752, n55753,
         n55754, n55755, n55756, n55757, n55758, n55759, n55760, n55761,
         n55762, n55763, n55764, n55765, n55766, n55767, n55768, n55769,
         n55770, n55771, n55772, n55773, n55774, n55775, n55776, n55777,
         n55778, n55779, n55780, n55781, n55782, n55783, n55784, n55785,
         n55786, n55787, n55788, n55789, n55790, n55791, n55792, n55793,
         n55794, n55795, n55796, n55797, n55798, n55799, n55800, n55801,
         n55802, n55803, n55804, n55805, n55806, n55807, n55808, n55809,
         n55810, n55811, n55812, n55813, n55814, n55815, n55816, n55817,
         n55818, n55819, n55820, n55821, n55822, n55823, n55824, n55825,
         n55826, n55827, n55828, n55829, n55830, n55831, n55832, n55833,
         n55834, n55835, n55836, n55837, n55838, n55839, n55840, n55841,
         n55842, n55843, n55844, n55845, n55846, n55847, n55848, n55849,
         n55850, n55851, n55852, n55853, n55854, n55855, n55856, n55857,
         n55858, n55859, n55860, n55861, n55862, n55863, n55864, n55865,
         n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873,
         n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881,
         n55882, n55883, n55884, n55885, n55886, n55887, n55888, n55889,
         n55890, n55891, n55892, n55893, n55894, n55895, n55896, n55897,
         n55898, n55899, n55900, n55901, n55902, n55903, n55904, n55905,
         n55906, n55907, n55908, n55909, n55910, n55911, n55912, n55913,
         n55914, n55915, n55916, n55917, n55918, n55919, n55920, n55921,
         n55922, n55923, n55924, n55925, n55926, n55927, n55928, n55929,
         n55930, n55931, n55932, n55933, n55934, n55935, n55936, n55937,
         n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945,
         n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953,
         n55954, n55955, n55956, n55957, n55958, n55959, n55960, n55961,
         n55962, n55963, n55964, n55965, n55966, n55967, n55968, n55969,
         n55970, n55971, n55972, n55973, n55974, n55975, n55976, n55977,
         n55978, n55979, n55980, n55981, n55982, n55983, n55984, n55985,
         n55986, n55987, n55988, n55989, n55990, n55991, n55992, n55993,
         n55994, n55995, n55996, n55997, n55998, n55999, n56000, n56001,
         n56002, n56003, n56004, n56005, n56006, n56007, n56008, n56009,
         n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017,
         n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025,
         n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033,
         n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041,
         n56042, n56043, n56044, n56045, n56046, n56047, n56048, n56049,
         n56050, n56051, n56052, n56053, n56054, n56055, n56056, n56057,
         n56058, n56059, n56060, n56061, n56062, n56063, n56064, n56065,
         n56066, n56067, n56068, n56069, n56070, n56071, n56072, n56073,
         n56074, n56075, n56076, n56077, n56078, n56079, n56080, n56081,
         n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089,
         n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097,
         n56098, n56099, n56100, n56101, n56102, n56103, n56104, n56105,
         n56106, n56107, n56108, n56109, n56110, n56111, n56112, n56113,
         n56114, n56115, n56116, n56117, n56118, n56119, n56120, n56121,
         n56122, n56123, n56124, n56125, n56126, n56127, n56128, n56129,
         n56130, n56131, n56132, n56133, n56134, n56135, n56136, n56137,
         n56138, n56139, n56140, n56141, n56142, n56143, n56144, n56145,
         n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153,
         n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161,
         n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169,
         n56170, n56171, n56172, n56173, n56174, n56175, n56176, n56177,
         n56178, n56179, n56180, n56181, n56182, n56183, n56184, n56185,
         n56186, n56187, n56188, n56189, n56190, n56191, n56192, n56193,
         n56194, n56195, n56196, n56197, n56198, n56199, n56200, n56201,
         n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209,
         n56210, n56211, n56212, n56213, n56214, n56215, n56216, n56217,
         n56218, n56219, n56220, n56221, n56222, n56223, n56224, n56225,
         n56226, n56227, n56228, n56229, n56230, n56231, n56232, n56233,
         n56234, n56235, n56236, n56237, n56238, n56239, n56240, n56241,
         n56242, n56243, n56244, n56245, n56246, n56247, n56248, n56249,
         n56250, n56251, n56252, n56253, n56254, n56255, n56256, n56257,
         n56258, n56259, n56260, n56261, n56262, n56263, n56264, n56265,
         n56266, n56267, n56268, n56269, n56270, n56271, n56272, n56273,
         n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281,
         n56282, n56283, n56284, n56285, n56286, n56287, n56288, n56289,
         n56290, n56291, n56292, n56293, n56294, n56295, n56296, n56297,
         n56298, n56299, n56300, n56301, n56302, n56303, n56304, n56305,
         n56306, n56307, n56308, n56309, n56310, n56311, n56312, n56313,
         n56314, n56315, n56316, n56317, n56318, n56319, n56320, n56321,
         n56322, n56323, n56324, n56325, n56326, n56327, n56328, n56329,
         n56330, n56331, n56332, n56333, n56334, n56335, n56336, n56337,
         n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345,
         n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353,
         n56354, n56355, n56356, n56357, n56358, n56359, n56360, n56361,
         n56362, n56363, n56364, n56365, n56366, n56367, n56368, n56369,
         n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377,
         n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385,
         n56386, n56387, n56388, n56389, n56390, n56391, n56392, n56393,
         n56394, n56395, n56396, n56397, n56398, n56399, n56400, n56401,
         n56402, n56403, n56404, n56405, n56406, n56407, n56408, n56409,
         n56410, n56411, n56412, n56413, n56414, n56415, n56416, n56417,
         n56418, n56419, n56420, n56421, n56422, n56423, n56424, n56425,
         n56426, n56427, n56428, n56429, n56430, n56431, n56432, n56433,
         n56434, n56435, n56436, n56437, n56438, n56439, n56440, n56441,
         n56442, n56443, n56444, n56445, n56446, n56447, n56448, n56449,
         n56450, n56451, n56452, n56453, n56454, n56455, n56456, n56457,
         n56458, n56459, n56460, n56461, n56462, n56463, n56464, n56465,
         n56466, n56467, n56468, n56469, n56470, n56471, n56472, n56473,
         n56474, n56475, n56476, n56477, n56478, n56479, n56480, n56481,
         n56482, n56483, n56484, n56485, n56486, n56487, n56488, n56489,
         n56490, n56491, n56492, n56493, n56494, n56495, n56496, n56497,
         n56498, n56499, n56500, n56501, n56502, n56503, n56504, n56505,
         n56506, n56507, n56508, n56509, n56510, n56511, n56512, n56513,
         n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521,
         n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529,
         n56530, n56531, n56532, n56533, n56534, n56535, n56536, n56537,
         n56538, n56539, n56540, n56541, n56542, n56543, n56544, n56545,
         n56546, n56547, n56548, n56549, n56550, n56551, n56552, n56553,
         n56554, n56555, n56556, n56557, n56558, n56559, n56560, n56561,
         n56562, n56563, n56564, n56565, n56566, n56567, n56568, n56569,
         n56570, n56571, n56572, n56573, n56574, n56575, n56576, n56577,
         n56578, n56579, n56580, n56581, n56582, n56583, n56584, n56585,
         n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593,
         n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601,
         n56602, n56603, n56604, n56605, n56606, n56607, n56608, n56609,
         n56610, n56611, n56612, n56613, n56614, n56615, n56616, n56617,
         n56618, n56619, n56620, n56621, n56622, n56623, n56624, n56625,
         n56626, n56627, n56628, n56629, n56630, n56631, n56632, n56633,
         n56634, n56635, n56636, n56637, n56638, n56639, n56640, n56641,
         n56642, n56643, n56644, n56645, n56646, n56647, n56648, n56649,
         n56650, n56651, n56652, n56653, n56654, n56655, n56656, n56657,
         n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665,
         n56666, n56667, n56668, n56669, n56670, n56671, n56672, n56673,
         n56674, n56675, n56676, n56677, n56678, n56679, n56680, n56681,
         n56682, n56683, n56684, n56685, n56686, n56687, n56688, n56689,
         n56690, n56691, n56692, n56693, n56694, n56695, n56696, n56697,
         n56698, n56699, n56700, n56701, n56702, n56703, n56704, n56705,
         n56706, n56707, n56708, n56709, n56710, n56711, n56712, n56713,
         n56714, n56715, n56716, n56717, n56718, n56719, n56720, n56721,
         n56722, n56723, n56724, n56725, n56726, n56727, n56728, n56729,
         n56730, n56731, n56732, n56733, n56734, n56735, n56736, n56737,
         n56738, n56739, n56740, n56741, n56742, n56743, n56744, n56745,
         n56746, n56747, n56748, n56749, n56750, n56751, n56752, n56753,
         n56754, n56755, n56756, n56757, n56758, n56759, n56760, n56761,
         n56762, n56763, n56764, n56765, n56766, n56767, n56768, n56769,
         n56770, n56771, n56772, n56773, n56774, n56775, n56776, n56777,
         n56778, n56779, n56780, n56781, n56782, n56783, n56784, n56785,
         n56786, n56787, n56788, n56789, n56790, n56791, n56792, n56793,
         n56794, n56795, n56796, n56797, n56798, n56799, n56800, n56801,
         n56802, n56803, n56804, n56805, n56806, n56807, n56808, n56809,
         n56810, n56811, n56812, n56813, n56814, n56815, n56816, n56817,
         n56818, n56819, n56820, n56821, n56822, n56823, n56824, n56825,
         n56826, n56827, n56828, n56829, n56830, n56831, n56832, n56833,
         n56834, n56835, n56836, n56837, n56838, n56839, n56840, n56841,
         n56842, n56843, n56844, n56845, n56846, n56847, n56848, n56849,
         n56850, n56851, n56852, n56853, n56854, n56855, n56856, n56857,
         n56858, n56859, n56860, n56861, n56862, n56863, n56864, n56941,
         n56942, n56943, n56944, n56945, n56946, n56947, n56948, n56949,
         n56950, n56951, n56952, n56953, n56954, n56955, n56956, n56957,
         n56958, n56959, n56960, n56961, n56962, n56963, n56964, n56965,
         n56966, n56967, n56968, n56969, n56970, n56971, n56972, n56973,
         n56974, n56975, n56976, n56977, n56978, n56979, n56980, n56981,
         n56982, n56983, n56984, n56985, n56986, n56987, n56988, n56989,
         n56990, n56991, n56992, n56993, n56994, n56995, n56996, n56997,
         n56998, n56999, n57000, n57001, n57002, n57003, n57004, n57005,
         n57006, n57007, n57008, n57009, n57010, n57011, n57012, n57013,
         n57014, n57015, n57016, n57017, n57018, n57019, n57020, n57021,
         n57022, n57023, n57024, n57025, n57026, n57027, n57028, n57029,
         n57030, n57031, n57032, n57033, n57034, n57035, n57036, n57037,
         n57038, n57039, n57040, n57041, n57042, n57043, n57044, n57045,
         n57046, n57047, n57048, n57049, n57050, n57051, n57052, n57053,
         n57054, n57055, n57056, n57057, n57058, n57059, n57060, n57061,
         n57062, n57063, n57064, n57065, n57066, n57067, n57068, n57069,
         n57070, n57071, n57072, n57073, n57074, n57075, n57076, n57077,
         n57078, n57079, n57080, n57081, n57082, n57083, n57084, n57085,
         n57086, n57087, n57088, n57089, n57090, n57091, n57092, n57093,
         n57094, n57095, n57096, n57097, n57098, n57099, n57100, n57101,
         n57102, n57103, n57104, n57105, n57106, n57107, n57108, n57109,
         n57110, n57111, n57112, n57113, n57114, n57115, n57116, n57117,
         n57118, n57119, n57120, n57121, n57122, n57123, n57124, n57125,
         n57126, n57127, n57128, n57129, n57130, n57131, n57132, n57133,
         n57134, n57135, n57136, n57137, n57138, n57139, n57140, n57141,
         n57142, n57143, n57144, n57145, n57146, n57147, n57148, n57149,
         n57150, n57151, n57152, n57153, n57154, n57155, n57156, n57157,
         n57158, n57159, n57160, n57161, n57162, n57163, n57164, n57165,
         n57166, n57167, n57168, n57169, n57170, n57171, n57172, n57173,
         n57174, n57175, n57176, n57177, n57178, n57179, n57180, n57181,
         n57182, n57183, n57184, n57185, n57186, n57187, n57188, n57189,
         n57190, n57191, n57192, n57193, n57194, n57195, n57196, n57197,
         n57198, n57199, n57200, n57201, n57202, n57203, n57204, n57205,
         n57206, n57207, n57208, n57209, n57210, n57211, n57212, n57213,
         n57214, n57215, n57216, n57217, n57218, n57219, n57220, n57221,
         n57222, n57223, n57224, n57225, n57226, n57227, n57228, n57229,
         n57230, n57231, n57232, n57233, n57234, n57235, n57236, n57237,
         n57238, n57239, n57240, n57241, n57242, n57243, n57244, n57245,
         n57246, n57247, n57248, n57249, n57250, n57251, n57252, n57253,
         n57254, n57255, n57256, n57257, n57258, n57259, n57260, n57261,
         n57262, n57263, n57264, n57265, n57266, n57267, n57268, n57269,
         n57270, n57271, n57272, n57273, n57274, n57275, n57276, n57277,
         n57278, n57279, n57280, n57281, n57282, n57283, n57284, n57285,
         n57286, n57287, n57288, n57289, n57290, n57291, n57292, n57293,
         n57294, n57295, n57296, n57297, n57298, n57299, n57300, n57301,
         n57302, n57303, n57304, n57305, n57306, n57307, n57308, n57309,
         n57310, n57311, n57312, n57313, n57314, n57315, n57316, n57317,
         n57318, n57319, n57320, n57321, n57322, n57323, n57324, n57325,
         n57326, n57327, n57328, n57329, n57330, n57331, n57332, n57333,
         n57334, n57335, n57336, n57337, n57338, n57339, n57340, n57341,
         n57342, n57343, n57344, n57345, n57346, n57347, n57348, n57349,
         n57350, n57351, n57352, n57353, n57354, n57355, n57356, n57357,
         n57358, n57359, n57360, n57361, n57362, n57363, n57364, n57365,
         n57366, n57367, n57368, n57369, n57370, n57371, n57372, n57373,
         n57374, n57375, n57376, n57377, n57378, n57379, n57380, n57381,
         n57382, n57383, n57384, n57385, n57386, n57387, n57388, n57389,
         n57390, n57391, n57392, n57393, n57394, n57395, n57396, n57397,
         n57398, n57399, n57400, n57401, n57402, n57403, n57404, n57405,
         n57406, n57407, n57408, n57409, n57410, n57411, n57412, n57413,
         n57414, n57415, n57416, n57417, n57418, n57419, n57420, n57421,
         n57422, n57423, n57424, n57425, n57426, n57427, n57428, n57429,
         n57430, n57431, n57432, n57433, n57434, n57435, n57436, n57437,
         n57438, n57439, n57440, n57441, n57442, n57443, n57444, n57445,
         n57446, n57447, n57448, n57449, n57450, n57451, n57452, n57453,
         n57454, n57455, n57456, n57457, n57458, n57459, n57460, n57461,
         n57462, n57463, n57464, n57465, n57466, n57467, n57468, n57469,
         n57470, n57471, n57472, n57473, n57474, n57475, n57476, n57477,
         n57478, n57479, n57480, n57481, n57482, n57483, n57484, n57485,
         n57486, n57487, n57488, n57489, n57490, n57491, n57492, n57493,
         n57494, n57495, n57496, n57497, n57498, n57499, n57500, n57501,
         n57502, n57503, n57504, n57505, n57506, n57507, n57508, n57509,
         n57510, n57511, n57512, n57513, n57514, n57515, n57516, n57517,
         n57518, n57519, n57520, n57521, n57522, n57523, n57524, n57525,
         n57526, n57527, n57528, n57529, n57530, n57531, n57532, n57533,
         n57534, n57535, n57536, n57537, n57538, n57539, n57540, n57541,
         n57542, n57543, n57544, n57545, n57546, n57547, n57548, n57549,
         n57550, n57551, n57552, n57553, n57554, n57555, n57556, n57557,
         n57558, n57559, n57560, n57561, n57562, n57563, n57564, n57565,
         n57566, n57567, n57568, n57569, n57570, n57571, n57572, n57573,
         n57574, n57575, n57576, n57577, n57578, n57579, n57580, n57581,
         n57582, n57583, n57584, n57585, n57586, n57587, n57588, n57589,
         n57590, n57591, n57592, n57593, n57594, n57595, n57596, n57597,
         n57598, n57599, n57600, n57601, n57602, n57603, n57604, n57605,
         n57606, n57607, n57608, n57609, n57610, n57611, n57612, n57613,
         n57614, n57615, n57616, n57617, n57618, n57619, n57620, n57621,
         n57622, n57623, n57624, n57625, n57626, n57627, n57628, n57629,
         n57630, n57631, n57632, n57633, n57634, n57635, n57636, n57637,
         n57638, n57639, n57640, n57641, n57642, n57643, n57644, n57645,
         n57646, n57647, n57648, n57649, n57650, n57651, n57652, n57653,
         n57654, n57655, n57656, n57657, n57658, n57659, n57660, n57661,
         n57662, n57663, n57664, n57665, n57666, n57667, n57668, n57669,
         n57670, n57671, n57672, n57673, n57674, n57675, n57676, n57677,
         n57678, n57679, n57680, n57681, n57682, n57683, n57684, n57685,
         n57686, n57687, n57688, n57689, n57690, n57691, n57692, n57693,
         n57694, n57695, n57696, n57697, n57698, n57699, n57700, n57701,
         n57702, n57703, n57704, n57705, n57706, n57707, n57708, n57709,
         n57710, n57711, n57712, n57713, n57714, n57715, n57716, n57717,
         n57718, n57719, n57720, n57721, n57722, n57723, n57724, n57725,
         n57726, n57727, n57728, n57729, n57730, n57731, n57732, n57733,
         n57734, n57735, n57736, n57737, n57738, n57739, n57740, n57741,
         n57742, n57743, n57744, n57745, n57746, n57747, n57748, n57749,
         n57750, n57751, n57752, n57753, n57754, n57755, n57756, n57757,
         n57758, n57759, n57760, n57761, n57762, n57763, n57764, n57765,
         n57766, n57767, n57768, n57769, n57770, n57771, n57772, n57773,
         n57774, n57775, n57776, n57777, n57778, n57779, n57780, n57781,
         n57782, n57783, n57784, n57785, n57786, n57787, n57788, n57789,
         n57790, n57791, n57792, n57793, n57794, n57795, n57796, n57797,
         n57798, n57799, n57800, n57801, n57802, n57803, n57804, n57805,
         n57806, n57807, n57808, n57809, n57810, n57811, n57812, n57813,
         n57814, n57815, n57816, n57817, n57818, n57819, n57820, n57821,
         n57822, n57823, n57824, n57825, n57826, n57827, n57828, n57829,
         n57830, n57831, n57832, n57833, n57834, n57835, n57836, n57837,
         n57838, n57839, n57840, n57841, n57842, n57843, n57844, n57845,
         n57846, n57847, n57848, n57849, n57850, n57851, n57852, n57853,
         n57854, n57855, n57856, n57857, n57858, n57859, n57860, n57861,
         n57862, n57863, n57864, n57865, n57866, n57867, n57868, n57869,
         n57870, n57871, n57872, n57873, n57874, n57875, n57876, n57877,
         n57878, n57879, n57880, n57881, n57882, n57883, n57884, n57885,
         n57886, n57887, n57888, n57889, n57890, n57891, n57892, n57893,
         n57894, n57895, n57896, n57897, n57898, n57899, n57900, n57901,
         n57902, n57903, n57904, n57905, n57906, n57907, n57908, n57909,
         n57910, n57911, n57912, n57913, n57914, n57915, n57916, n57917,
         n57918, n57919, n57920, n57921, n57922, n57923, n57924, n57925,
         n57926, n57927, n57928, n57929, n57930, n57931, n57932, n57933,
         n57934, n57935, n57936, n57937, n57938, n57939, n57940, n57941,
         n57942, n57943, n57944, n57945, n57946, n57947, n57948, n57949,
         n57950, n57951, n57952, n57953, n57954, n57955, n57956, n57957,
         n57958, n57959, n57960, n57961, n57962, n57963, n57964, n57965,
         n57966, n57967, n57968, n57969, n57970, n57971, n57972, n57973,
         n57974, n57975, n57976, n57977, n57978, n57979, n57980, n57981,
         n57982, n57983, n57984, n57985, n57986, n57987, n57988, n57989,
         n57990, n57991, n57992, n57993, n57994, n57995, n57996, n57997,
         n57998, n57999, n58000, n58001, n58002, n58003, n58004, n58005,
         n58006, n58007, n58008, n58009, n58010, n58011, n58012, n58013,
         n58014, n58015, n58016, n58017, n58018, n58019, n58020, n58021,
         n58022, n58023, n58024, n58025, n58026, n58027, n58028, n58029,
         n58030, n58031, n58032, n58033, n58034, n58035, n58036, n58037,
         n58038, n58039, n58040, n58041, n58042, n58043, n58044, n58045,
         n58046, n58047, n58048, n58049, n58050, n58051, n58052, n58053,
         n58054, n58055, n58056, n58057, n58058, n58059, n58060, n58061,
         n58062, n58063, n58064, n58065, n58066, n58067, n58068, n58069,
         n58070, n58071, n58072, n58073, n58074, n58075, n58076, n58077,
         n58078, n58079, n58080, n58081, n58082, n58083, n58084, n58085,
         n58086, n58087, n58088, n58089, n58090, n58091, n58092, n58093,
         n58094, n58095, n58096, n58097, n58098, n58099, n58100, n58101,
         n58102, n58103, n58104, n58105, n58106, n58107, n58108, n58109,
         n58110, n58111, n58112, n58113, n58114, n58115, n58116, n58117,
         n58118, n58119, n58120, n58121, n58122, n58123, n58124, n58125,
         n58126, n58127, n58128, n58129, n58130, n58131, n58132, n58133,
         n58134, n58135, n58136, n58137, n58138, n58139, n58140, n58141,
         n58142, n58143, n58144, n58145, n58146, n58147, n58148, n58149,
         n58150, n58151, n58152, n58153, n58154, n58155, n58156, n58157,
         n58158, n58159, n58160, n58161, n58162, n58163, n58164, n58165,
         n58166, n58167, n58168, n58169, n58170, n58171, n58172, n58173,
         n58174, n58175, n58176, n58177, n58178, n58179, n58180, n58181,
         n58182, n58183, n58184, n58185, n58186, n58187, n58188, n58189,
         n58190, n58191, n58192, n58193, n58194, n58195, n58196, n58197,
         n58198, n58199, n58200, n58201, n58202, n58203, n58204, n58205,
         n58206, n58207, n58208, n58209, n58210, n58211, n58212, n58213,
         n58214, n58215, n58216, n58217, n58218, n58219, n58220, n58221,
         n58222, n58223, n58224, n58225, n58226, n58227, n58228, n58229,
         n58230, n58231, n58232, n58233, n58234, n58235, n58236, n58237,
         n58238, n58239, n58240, n58241, n58242, n58243, n58244, n58245,
         n58246, n58247, n58248, n58249, n58250, n58251, n58252, n58253,
         n58254, n58255, n58256, n58257, n58258, n58259, n58260, n58261,
         n58262, n58263, n58264, n58265, n58266, n58267, n58268, n58269,
         n58270, n58271, n58272, n58273, n58274, n58275, n58276, n58277,
         n58278, n58279, n58280, n58281, n58282, n58283, n58284, n58285,
         n58286, n58287, n58288, n58289, n58290, n58291, n58292, n58293,
         n58294, n58295, n58296, n58297, n58298, n58299, n58300, n58301,
         n58302, n58303, n58304, n58305, n58306, n58307, n58308, n58309,
         n58310, n58311, n58312, n58313, n58314, n58315, n58316, n58317,
         n58318, n58319, n58320, n58321, n58322, n58323, n58324, n58325,
         n58326, n58327, n58328, n58329, n58330, n58331, n58332, n58333,
         n58334, n58335, n58336, n58337, n58338, n58339, n58340, n58341,
         n58342, n58343, n58344, n58345, n58346, n58347, n58348, n58349,
         n58350, n58351, n58352, n58353, n58354, n58355, n58356, n58357,
         n58358, n58359, n58360, n58361, n58362, n58363, n58364, n58365,
         n58366, n58367, n58368, n58369, n58370, n58371, n58372, n58373,
         n58374, n58375, n58376, n58377, n58378, n58379, n58380, n58381,
         n58382, n58383, n58384, n58385, n58386, n58387, n58388, n58389,
         n58390, n58391, n58392, n58393, n58394, n58395, n58396, n58397,
         n58398, n58399, n58400, n58401, n58402, n58403, n58404, n58405,
         n58406, n58407, n58408, n58409, n58410, n58411, n58412, n58413,
         n58414, n58415, n58416, n58417, n58418, n58419, n58420, n58421,
         n58422, n58423, n58424, n58425, n58426, n58427, n58428, n58429,
         n58430, n58431, n58432, n58433, n58434, n58435, n58436, n58437,
         n58438, n58439, n58440, n58441, n58442, n58443, n58444, n58445,
         n58446, n58447, n58448, n58449, n58450, n58451, n58452, n58453,
         n58454, n58455, n58456, n58457, n58458, n58459, n58460, n58461,
         n58462, n58463, n58464, n58465, n58466, n58467, n58468, n58469,
         n58470, n58471, n58472, n58473, n58474, n58475, n58476, n58477,
         n58478, n58479, n58480, n58481, n58482, n58483, n58484, n58485,
         n58486, n58487, n58488, n58489, n58490, n58491, n58492, n58493,
         n58494, n58495, n58496, n58497, n58498, n58499, n58500, n58501,
         n58502, n58503, n58504, n58505, n58506, n58507, n58508, n58509,
         n58510, n58511, n58512, n58513, n58514, n58515, n58516, n58517,
         n58518, n58519, n58520, n58521, n58522, n58523, n58524, n58525,
         n58526, n58527, n58528, n58529, n58530, n58531, n58532, n58533,
         n58534, n58535, n58536, n58537, n58538, n58539, n58540, n58541,
         n58542, n58543, n58544, n58545, n58546, n58547, n58548, n58549,
         n58550, n58551, n58552, n58553, n58554, n58555, n58556, n58557,
         n58558, n58559, n58560, n58561, n58562, n58563, n58564, n58565,
         n58566, n58567, n58568, n58569, n58570, n58571, n58572, n58573,
         n58574, n58575, n58576, n58577, n58578, n58579, n58580, n58581,
         n58582, n58583, n58584, n58585, n58586, n58587, n58588, n58589,
         n58590, n58591, n58592, n58593, n58594, n58595, n58596, n58597,
         n58598, n58599, n58600, n58601, n58602, n58603, n58604, n58605,
         n58606, n58607, n58608, n58609, n58610, n58611, n58612, n58613,
         n58614, n58615, n58616, n58617, n58618, n58619, n58620, n58621,
         n58622, n58623, n58624, n58625, n58626, n58627, n58628, n58629,
         n58630, n58631, n58632, n58633, n58634, n58635, n58636, n58637,
         n58638, n58639, n58640, n58641, n58642, n58643, n58644, n58645,
         n58646, n58647, n58648, n58649, n58650, n58651, n58652, n58653,
         n58654, n58655, n58656, n58657, n58658, n58659, n58660, n58661,
         n58662, n58663, n58664, n58665, n58666, n58667, n58668, n58669,
         n58670, n58671, n58672, n58673, n58674, n58675, n58676, n58677,
         n58678, n58679, n58680, n58681, n58682, n58683, n58684, n58685,
         n58686, n58687, n58688, n58689, n58690, n58691, n58692, n58693,
         n58694, n58695, n58696, n58697, n58698, n58699, n58700, n58701,
         n58702, n58703, n58704, n58705, n58706, n58707, n58708, n58709,
         n58710, n58711, n58712, n58713, n58714, n58715, n58716, n58717,
         n58718, n58719, n58720, n58721, n58722, n58723, n58724, n58725,
         n58726, n58727, n58728, n58729, n58730, n58731, n58732, n58733,
         n58734, n58735, n58736, n58737, n58738, n58739, n58740, n58741,
         n58742, n58743, n58744, n58745, n58746, n58747, n58748, n58749,
         n58750, n58751, n58752, n58753, n58754, n58755, n58756, n58757,
         n58758, n58759, n58760, n58761, n58762, n58763, n58764, n58765,
         n58766, n58767, n58768, n58769, n58770, n58771, n58772, n58773,
         n58774, n58775, n58776, n58777, n58778, n58779, n58780, n58781,
         n58782, n58783, n58784, n58785, n58786, n58787, n58788, n58789,
         n58790, n58791, n58792, n58793, n58794, n58795, n58796, n58797,
         n58798, n58799, n58800, n58801, n58802, n58803, n58804, n58805,
         n58806, n58807, n58808, n58809, n58810, n58811, n58812, n58813,
         n58814, n58815, n58816, n58817, n58818, n58819, n58820, n58821,
         n58822, n58823, n58824, n58825, n58826, n58827, n58828, n58829,
         n58830, n58831, n58832, n58833, n58834, n58835, n58836, n58837,
         n58838, n58839, n58840, n58841, n58842, n58843, n58844, n58845,
         n58846, n58847, n58848, n58849, n58850, n58851, n58852, n58853,
         n58854, n58855, n58856, n58857, n58858, n58859, n58860, n58861,
         n58862, n58863, n58864, n58865, n58866, n58867, n58868, n58869,
         n58870, n58871, n58872, n58873, n58874, n58875, n58876, n58877,
         n58878, n58879, n58880, n58881, n58882, n58883, n58884, n58885,
         n58886, n58887, n58888, n58889, n58890, n58891, n58892, n58893,
         n58894, n58895, n58896, n58897, n58898, n58899, n58900, n58901,
         n58902, n58903, n58904, n58905, n58906, n58907, n58908, n58909,
         n58910, n58911, n58912, n58913, n58914, n58915, n58916, n58917,
         n58918, n58919, n58920, n58921, n58922, n58923, n58924, n58925,
         n58926, n58927, n58928, n58929, n58930, n58931, n58932, n58933,
         n58934, n58935, n58936, n58937, n58938, n58939, n58940, n58941,
         n58942, n58943, n58944, n58945, n58946, n58947, n58948, n58949,
         n58950, n58951, n58952, n58953, n58954, n58955, n58956, n58957,
         n58958, n58959, n58960, n58961, n58962, n58963, n58964, n58965,
         n58966, n58967, n58968, n58969, n58970, n58971, n58972, n58973,
         n58974, n58975, n58976, n58977, n58978, n58979, n58980, n58981,
         n58982, n58983, n58984, n58985, n58986, n58987, n58988, n58989,
         n58990, n58991, n58992, n58993, n58994, n58995, n58996, n58997,
         n58998, n58999, n59000, n59001, n59002, n59003, n59004, n59005,
         n59006, n59007, n59008, n59009, n59010, n59011, n59012, n59013,
         n59014, n59015, n59016, n59017, n59018, n59019, n59020, n59021,
         n59022, n59023, n59024, n59025, n59026, n59027, n59028, n59029,
         n59030, n59031, n59032, n59033, n59034, n59035, n59036, n59037,
         n59038, n59039, n59040, n59041, n59042, n59043, n59044, n59045,
         n59046, n59047, n59048, n59049, n59050, n59051, n59052, n59053,
         n59054, n59055, n59056, n59057, n59058, n59059, n59060, n59061,
         n59062, n59063, n59064, n59065, n59066, n59067, n59068, n59069,
         n59070, n59071, n59072, n59073, n59074, n59075, n59076, n59077,
         n59078, n59079, n59080, n59081, n59082, n59083, n59084, n59085,
         n59086, n59087, n59088, n59089, n59090, n59091, n59092, n59093,
         n59094, n59095, n59096, n59097, n59098, n59099, n59100, n59101,
         n59102, n59103, n59104, n59105, n59106, n59107, n59108, n59109,
         n59110, n59111, n59112, n59113, n59114, n59115, n59116, n59117,
         n59118, n59119, n59120, n59121, n59122, n59123, n59124, n59125,
         n59126, n59127, n59128, n59129, n59130, n59131, n59132, n59133,
         n59134, n59135, n59136, n59137, n59138, n59139, n59140, n59141,
         n59142, n59143, n59144, n59145, n59146, n59147, n59148, n59149,
         n59150, n59151, n59152, n59153, n59154, n59155, n59156, n59157,
         n59158, n59159, n59160, n59161, n59162, n59163, n59164, n59165,
         n59166, n59167, n59168, n59169, n59170, n59171, n59172, n59173,
         n59174, n59175, n59176, n59177, n59178, n59179, n59180, n59181,
         n59182, n59183, n59184, n59185, n59186, n59187, n59188, n59189,
         n59190, n59191, n59192, n59193, n59194, n59195, n59196, n59197,
         n59198, n59199, n59200, n59201, n59202, n59203, n59204, n59205,
         n59206, n59207, n59208, n59209, n59210, n59211, n59212, n59213,
         n59214, n59215, n59216, n59217, n59218, n59219, n59220, n59221,
         n59222, n59223, n59224, n59225, n59226, n59227, n59228, n59229,
         n59230, n59231, n59232, n59233, n59234, n59235, n59236, n59237,
         n59238, n59239, n59240, n59241, n59242, n59243, n59244, n59245,
         n59246, n59247, n59248, n59249, n59250, n59251, n59252, n59253,
         n59254, n59255, n59256, n59257, n59258, n59259, n59260, n59261,
         n59262, n59263, n59264, n59265, n59266, n59267, n59268, n59269,
         n59270, n59271, n59272, n59273, n59274, n59275, n59276, n59277,
         n59278, n59279, n59280, n59281, n59282, n59283, n59284, n59285,
         n59286, n59287, n59288, n59289, n59290, n59291, n59292, n59293,
         n59294, n59295, n59296, n59297, n59298, n59299, n59300, n59301,
         n59302, n59303, n59304, n59305, n59306, n59307, n59308, n59309,
         n59310, n59311, n59312, n59313, n59314, n59315, n59316, n59317,
         n59318, n59319, n59320, n59321, n59322, n59323, n59324, n59325,
         n59326, n59327, n59328, n59329, n59330, n59331, n59332, n59333,
         n59334, n59335, n59336, n59337, n59338, n59339, n59340, n59341,
         n59342, n59343, n59344, n59345, n59346, n59347, n59348, n59349,
         n59350, n59351, n59352, n59353, n59354, n59355, n59356, n59357,
         n59358, n59359, n59360, n59361, n59362, n59363, n59364, n59365,
         n59366, n59367, n59368, n59369, n59370, n59371, n59372, n59373,
         n59374, n59375, n59376, n59377, n59378, n59379, n59380, n59381,
         n59382, n59383, n59384, n59385, n59386, n59387, n59388, n59389,
         n59390, n59391, n59392, n59393, n59394, n59395, n59396, n59397,
         n59398, n59399, n59400, n59401, n59402, n59403, n59404, n59405,
         n59406, n59407, n59408, n59409, n59410, n59411, n59412, n59413,
         n59414, n59415, n59416, n59417, n59418, n59419, n59420, n59421,
         n59422, n59423, n59424, n59425, n59426, n59427, n59428, n59429,
         n59430, n59431, n59433, n59434, n59435, n59436, n59437, n59438,
         n59439, n59440, n59441, n59442, n59443, n59444, n59445, n59446,
         n59447, n59448, n59449, n59450, n59451, n59452, n59453, n59454,
         n59455, n59456, n59457, n59458, n59459, n59460, n59461, n59462,
         n59463, n59464, n59465, n59466, n59467, n59468, n59469, n59470,
         n59471, n59472, n59473, n59474, n59475, n59476, n59477, n59478,
         n59479, n59480, n59481, n59482, n59483, n59484, n59485, n59486,
         n59487, n59488, n59489, n59490, n59491, n59492, n59493, n59494,
         n59495, n59496, n59497, n59498, n59499, n59500, n59501, n59502,
         n59503, n59504, n59505, n59506, n59507, n59508, n59509, n59510,
         n59511, n59512, n59513, n59514, n59515, n59516, n59517, n59518,
         n59519, n59520, n59521, n59522, n59523, n59524, n59525, n59526,
         n59527, n59528, n59529, n59530, n59531, n59532, n59533, n59534,
         n59535, n59536, n59537, n59538, n59539, n59540, n59541, n59542,
         n59543, n59544, n59545, n59546, n59547, n59548, n59549, n59550,
         n59551, n59552, n59553, n59554, n59555, n59556, n59557, n59558,
         n59559, n59560, n59561, n59562, n59563, n59564, n59565, n59566,
         n59567, n59568, n59569, n59570, n59571, n59572, n59573, n59574,
         n59575, n59576, n59577, n59578, n59579, n59580, n59581, n59582,
         n59583, n59584, n59585, n59586, n59587, n59588, n59589, n59590,
         n59591, n59592, n59593, n59594, n59595, n59596, n59597, n59598,
         n59599, n59600, n59601, n59602, n59603, n59604, n59605, n59606,
         n59607, n59608, n59609, n59610, n59611, n59612, n59613, n59614,
         n59615, n59616, n59617, n59618, n59619, n59620, n59621, n59622,
         n59623, n59624, n59625, n59626, n59627, n59628, n59629, n59630,
         n59631, n59632, n59633, n59634, n59635, n59636, n59637, n59638,
         n59639, n59640, n59641, n59642, n59643, n59644, n59645, n59646,
         n59647, n59648, n59649, n59650, n59651, n59652, n59653, n59654,
         n59655, n59656, n59657, n59658, n59659, n59660, n59661, n59662,
         n59663, n59664, n59665, n59666, n59667, n59668, n59669, n59670,
         n59671, n59672, n59673, n59674, n59675, n59676, n59677, n59678,
         n59679, n59680, n59681, n59682, n59683, n59684, n59685, n59686,
         n59687, n59688, n59689, n59690, n59691, n59692, n59693, n59694,
         n59695, n59696, n59697, n59698, n59699, n59700, n59701, n59702,
         n59703, n59704, n59705, n59706, n59707, n59708, n59709, n59710,
         n59711, n59712, n59713, n59714, n59715, n59716, n59717, n59718,
         n59719, n59720, n59721, n59722, n59723, n59724, n59725, n59726,
         n59727, n59728, n59729, n59730, n59731, n59732, n59733, n59734,
         n59735, n59736, n59737, n59738, n59739, n59740, n59741, n59742,
         n59743, n59744, n59745, n59746, n59747, n59748, n59749, n59750,
         n59751, n59752, n59753, n59754, n59755, n59756, n59757, n59758,
         n59759, n59760, n59761, n59762, n59763, n59764, n59765, n59766,
         n59767, n59768, n59769, n59770, n59771, n59772, n59773, n59774,
         n59775, n59776, n59777, n59778, n59779, n59780, n59781, n59782,
         n59783, n59784, n59785, n59786, n59787, n59788, n59789, n59790,
         n59791, n59792, n59793, n59794, n59795, n59796, n59797, n59798,
         n59799, n59800, n59801, n59802, n59803, n59804, n59805, n59806,
         n59807, n59808, n59809, n59810, n59811, n59812, n59813, n59814,
         n59815, n59816, n59817, n59818, n59819, n59820, n59821, n59822,
         n59823, n59824, n59825, n59826, n59827, n59828, n59829, n59830,
         n59831, n59832, n59833, n59834, n59835, n59836, n59837, n59838,
         n59839, n59840, n59841, n59842, n59843, n59844, n59845, n59846,
         n59847, n59848, n59849, n59850, n59851, n59852, n59853, n59854,
         n59855, n59856, n59857, n59858, n59859, n59860, n59861, n59862,
         n59863, n59864, n59865, n59866, n59867, n59868, n59869, n59870,
         n59871, n59872, n59873, n59874, n59875, n59876, n59877, n59878,
         n59879, n59880, n59881, n59882, n59883, n59884, n59885, n59886,
         n59887, n59888, n59889, n59890, n59891, n59892, n59893, n59894,
         n59895, n59896, n59897, n59898, n59899, n59900, n59901, n59902,
         n59903, n59904, n59905, n59906, n59907, n59908, n59909, n59910,
         n59911, n59912, n59913, n59914, n59915, n59916, n59917, n59918,
         n59919, n59920, n59921, n59922, n59923, n59924, n59925, n59926,
         n59927, n59928, n59929, n59930, n59931, n59932, n59933, n59934,
         n59935, n59936, n59937, n59938, n59939, n59940, n59941, n59942,
         n59943, n59944, n59945, n59946, n59947, n59948, n59949, n59950,
         n59951, n59952, n59953, n59954, n59955, n59956, n59957, n59958,
         n59959, n59960, n59961, n59962, n59963, n59964, n59965, n59966,
         n59967, n59968, n59969, n59970, n59971, n59972, n59973, n59974,
         n59975, n59976, n59977, n59978, n59979, n59980, n59981, n59982,
         n59983, n59984, n59985, n59986, n59987, n59988, n59989, n59990,
         n59991, n59992, n59993, n59994, n59995, n59996, n59997, n59998,
         n59999, n60000, n60001, n60002, n60003, n60004, n60005, n60006,
         n60007, n60008, n60009, n60010, n60011, n60012, n60013, n60014,
         n60015, n60016, n60017, n60018, n60019, n60020, n60021, n60022,
         n60023, n60024, n60025, n60026, n60027, n60028, n60029, n60030,
         n60031, n60032, n60033, n60034, n60035, n60036, n60037, n60038,
         n60039, n60040, n60041, n60042, n60043, n60044, n60045, n60046,
         n60047, n60048, n60049, n60050, n60051, n60052, n60053, n60054,
         n60055, n60056, n60057, n60058, n60059, n60060, n60061, n60062,
         n60063, n60064, n60065, n60066, n60067, n60068, n60069, n60070,
         n60071, n60072, n60073, n60074, n60075, n60076, n60077, n60078,
         n60079, n60080, n60081, n60082, n60083, n60084, n60085, n60086,
         n60087, n60088, n60089, n60090, n60091, n60092, n60093, n60094,
         n60095, n60096, n60097, n60098, n60099, n60100, n60101, n60102,
         n60103, n60104, n60105, n60106, n60107, n60108, n60109, n60110,
         n60111, n60112, n60113, n60114, n60115, n60116, n60117, n60118,
         n60119, n60120, n60121, n60122, n60123, n60124, n60125, n60126,
         n60127, n60128, n60129, n60130, n60131, n60132, n60133, n60134,
         n60135, n60136, n60137, n60138, n60139, n60140, n60141, n60142,
         n60143, n60144, n60145, n60146, n60147, n60148, n60149, n60150,
         n60151, n60152, n60153, n60154, n60155, n60156, n60157, n60158,
         n60159, n60160, n60161, n60162, n60163, n60164, n60165, n60166,
         n60167, n60168, n60169, n60170, n60171, n60172, n60173, n60174,
         n60175, n60176, n60177, n60178, n60179, n60180, n60181, n60182,
         n60183, n60184, n60185, n60186, n60187, n60188, n60189, n60190,
         n60191, n60192, n60193, n60194, n60195, n60196, n60197, n60198,
         n60199, n60200, n60201, n60202, n60203, n60204, n60205, n60206,
         n60207, n60208, n60209, n60210, n60211, n60212, n60213, n60214,
         n60215, n60216, n60217, n60218, n60219, n60220, n60221, n60222,
         n60223, n60224, n60225, n60226, n60227, n60228, n60229, n60230,
         n60231, n60232, n60233, n60234, n60235, n60236, n60237, n60238,
         n60239, n60240, n60241, n60242, n60243, n60244, n60245, n60246,
         n60247, n60248, n60249, n60250, n60251, n60252, n60253, n60254,
         n60255, n60256, n60257, n60258, n60259, n60260, n60261, n60262,
         n60263, n60264, n60265, n60266, n60267, n60268, n60269, n60270,
         n60271, n60272, n60273, n60274, n60275, n60276, n60277, n60278,
         n60279, n60280, n60281, n60282, n60283, n60284, n60285, n60286,
         n60287, n60288, n60289, n60290, n60291, n60292, n60293, n60294,
         n60295, n60296, n60297, n60298, n60299, n60300, n60301, n60302,
         n60303, n60304, n60305, n60306, n60307, n60308, n60309, n60310,
         n60311, n60312, n60313, n60314, n60315, n60316, n60317, n60318,
         n60319, n60320, n60321, n60322, n60323, n60324, n60325, n60326,
         n60327, n60328, n60329, n60330, n60331, n60332, n60333, n60334,
         n60335, n60336, n60337, n60338, n60339, n60340, n60341, n60342,
         n60343, n60344, n60345, n60346, n60347, n60348, n60349, n60350,
         n60351, n60352, n60353, n60354, n60355, n60356, n60357, n60358,
         n60359, n60360, n60361, n60362, n60363, n60364, n60365, n60366,
         n60367, n60368, n60369, n60370, n60371, n60372, n60373, n60374,
         n60375, n60376, n60377, n60378, n60379, n60380, n60381, n60382,
         n60383, n60384, n60385, n60386, n60387, n60388, n60389, n60390,
         n60391, n60392, n60393, n60394, n60395, n60396, n60397, n60398,
         n60399, n60400, n60401, n60402, n60403, n60404, n60405, n60406,
         n60407, n60408, n60409, n60410, n60411, n60412, n60413, n60414,
         n60415, n60416, n60417, n60418, n60419, n60420, n60421, n60422,
         n60423, n60424, n60425, n60426, n60427, n60428, n60429, n60430,
         n60431, n60432, n60433, n60434, n60435, n60436, n60437, n60438,
         n60439, n60440, n60441, n60442, n60443, n60444, n60445, n60446,
         n60447, n60448, n60449, n60450, n60451, n60452, n60453, n60454,
         n60455, n60456, n60457, n60458, n60459, n60460, n60461, n60462,
         n60463, n60464, n60465, n60466, n60467, n60468, n60469, n60470,
         n60471, n60472, n60473, n60474, n60475, n60476, n60477, n60478,
         n60479, n60480, n60481, n60482, n60483, n60484, n60485, n60486,
         n60487, n60488, n60489, n60490, n60491, n60492, n60493, n60494,
         n60495, n60496, n60497, n60498, n60499, n60500, n60501, n60502,
         n60503, n60504, n60505, n60506, n60507, n60508, n60509, n60510,
         n60511, n60512, n60513, n60514, n60515, n60516, n60517, n60518,
         n60519, n60520, n60521, n60522, n60523, n60524, n60525, n60526,
         n60527, n60528, n60529, n60530, n60531, n60532, n60533, n60534,
         n60535, n60536, n60537, n60538, n60539, n60540, n60541, n60542,
         n60543, n60544, n60545, n60546, n60547, n60548, n60549, n60550,
         n60551, n60552, n60553, n60554, n60555, n60556, n60557, n60558,
         n60559, n60560, n60561, n60562, n60563, n60564, n60565, n60566,
         n60567, n60568, n60569, n60570, n60571, n60572, n60573, n60574,
         n60575, n60576, n60577, n60578, n60579, n60580, n60581, n60582,
         n60583, n60584, n60585, n60586, n60587, n60588, n60589, n60590,
         n60591, n60592, n60593, n60594, n60595, n60596, n60597, n60598,
         n60599, n60600, n60601, n60602, n60603, n60604, n60605, n60606,
         n60607, n60608, n60609, n60610, n60611, n60612, n60613, n60614,
         n60615, n60616, n60617, n60618, n60619, n60620, n60621, n60622,
         n60623, n60624, n60625, n60626, n60627, n60628, n60629, n60630,
         n60631, n60632, n60633, n60634, n60635, n60636, n60637, n60638,
         n60639, n60640, n60641, n60642, n60643, n60644, n60645, n60646,
         n60647, n60648, n60649, n60650, n60651, n60652, n60653, n60654,
         n60655, n60656, n60657, n60658, n60659, n60660, n60661, n60662,
         n60663, n60664, n60665, n60666, n60667, n60668, n60669, n60670,
         n60671, n60672, n60673, n60674, n60675, n60676, n60677, n60678,
         n60679, n60680, n60681, n60682, n60683, n60684, n60685, n60686,
         n60687, n60688, n60689, n60690, n60691, n60692, n60693, n60694,
         n60695, n60696, n60697, n60698, n60699, n60700, n60701, n60702,
         n60703, n60704, n60705, n60706, n60707, n60708, n60709, n60710,
         n60711, n60712, n60713, n60714, n60715, n60716, n60717, n60718,
         n60719, n60720, n60721, n60722, n60723, n60724, n60725, n60726,
         n60727, n60728, n60729, n60730, n60731, n60732, n60733, n60734,
         n60735, n60736, n60737, n60738, n60739, n60740, n60741, n60742,
         n60743, n60744, n60745, n60746, n60747, n60748, n60749, n60750,
         n60751, n60752, n60753, n60754, n60755, n60756, n60757, n60758,
         n60759, n60760, n60761, n60762, n60763, n60764, n60765, n60766,
         n60767, n60768, n60769, n60770, n60771, n60772, n60773, n60774,
         n60775, n60776, n60777, n60778, n60779, n60780, n60781, n60782,
         n60783, n60784, n60785, n60786, n60787, n60788, n60789, n60790,
         n60791, n60792, n60793, n60794, n60795, n60796, n60797, n60798,
         n60799, n60800, n60801, n60802, n60803, n60804, n60805, n60806,
         n60807, n60808, n60809, n60810, n60811, n60812, n60813, n60814,
         n60815, n60816, n60817, n60818, n60819, n60820, n60821, n60822,
         n60823, n60824, n60825, n60826, n60827, n60828, n60829, n60830,
         n60831, n60832, n60833, n60834, n60835, n60836, n60837, n60838,
         n60839, n60840, n60841, n60842, n60843, n60844, n60845, n60846,
         n60847, n60848, n60849, n60850, n60851, n60852, n60853, n60854,
         n60855, n60856, n60857, n60858, n60859, n60860, n60861, n60862,
         n60863, n60864, n60865, n60866, n60867, n60868, n60869, n60870,
         n60871, n60872, n60873, n60874, n60875, n60876, n60877, n60878,
         n60879, n60880, n60881, n60882, n60883, n60884, n60885, n60886,
         n60887, n60888, n60889, n60890, n60891, n60892, n60893, n60894,
         n60895, n60896, n60897, n60898, n60899, n60900, n60901, n60902,
         n60903, n60904, n60905, n60906, n60907, n60908, n60909, n60910,
         n60911, n60912, n60913, n60914, n60915, n60916, n60917, n60918,
         n60919, n60920, n60921, n60922, n60923, n60924, n60925, n60926,
         n60927, n60928, n60929, n60930, n60931, n60932, n60933, n60934,
         n60935, n60936, n60937, n60938, n60939, n60940, n60941, n60942,
         n60943, n60944, n60945, n60946, n60947, n60948, n60949, n60950,
         n60951, n60952, n60953, n60954, n60955, n60956, n60957, n60958,
         n60959, n60960, n60961, n60962, n60963, n60964, n60965, n60966,
         n60967, n60968, n60969, n60970, n60971, n60972, n60973, n60974,
         n60975, n60976, n60977, n60978, n60979, n60980, n60981, n60982,
         n60983, n60984, n60985, n60986, n60987, n60988, n60989, n60990,
         n60991, n60992, n60993, n60994, n60995, n60996, n60997, n60998,
         n60999, n61000, n61001, n61002, n61003, n61004, n61005, n61006,
         n61007, n61008, n61009, n61010, n61011, n61012, n61013, n61014,
         n61015, n61016, n61017, n61018, n61019, n61020, n61021, n61022,
         n61023, n61024, n61025, n61026, n61027, n61028, n61029, n61030,
         n61031, n61032, n61033, n61034, n61035, n61036, n61037, n61038,
         n61039, n61040, n61041, n61042, n61043, n61044, n61045, n61046,
         n61047, n61048, n61049, n61050, n61051, n61052, n61053, n61054,
         n61055, n61056, n61057, n61058, n61059, n61060, n61061, n61062,
         n61063, n61064, n61065, n61066, n61067, n61068, n61069, n61070,
         n61071, n61072, n61073, n61074, n61075, n61076, n61077, n61078,
         n61079, n61080, n61081, n61082, n61083, n61084, n61085, n61086,
         n61087, n61088, n61089, n61090, n61091, n61092, n61093, n61094,
         n61095, n61096, n61097, n61098, n61099, n61100, n61101, n61102,
         n61103, n61104, n61105, n61106, n61107, n61108, n61109, n61110,
         n61111, n61112, n61113, n61114, n61115, n61116, n61117, n61118,
         n61119, n61120, n61121, n61122, n61123, n61124, n61125, n61126,
         n61127, n61128, n61129, n61130, n61131, n61132, n61133, n61134,
         n61135, n61136, n61137, n61138, n61139, n61140, n61141, n61142,
         n61143, n61144, n61145, n61146, n61147, n61148, n61149, n61150,
         n61151, n61152, n61153, n61154, n61155, n61156, n61157, n61158,
         n61159, n61160, n61161, n61162, n61163, n61164, n61165, n61166,
         n61167, n61168, n61169, n61170, n61171, n61172, n61173, n61174,
         n61175, n61176, n61177, n61178, n61179, n61180, n61181, n61182,
         n61183, n61184, n61185, n61186, n61187, n61188, n61189, n61190,
         n61191, n61192, n61193, n61194, n61195, n61196, n61197, n61198,
         n61199, n61200, n61201, n61202, n61203, n61204, n61205, n61206,
         n61207, n61208, n61209, n61210, n61211, n61212, n61213, n61214,
         n61215, n61216, n61217, n61218, n61219, n61220, n61221, n61222,
         n61223, n61224, n61225, n61226, n61227, n61228, n61229, n61230,
         n61231, n61232, n61233, n61234, n61235, n61236, n61237, n61238,
         n61239, n61240, n61241, n61242, n61243, n61244, n61245, n61246,
         n61247, n61248, n61249, n61250, n61251, n61252, n61253, n61254,
         n61255, n61256, n61257, n61258, n61259, n61260, n61261, n61262,
         n61263, n61264, n61265, n61266, n61267, n61268, n61269, n61270,
         n61271, n61272, n61273, n61274, n61275, n61276, n61277, n61278,
         n61279, n61280, n61281, n61282, n61283, n61284, n61285, n61286,
         n61287, n61288, n61289, n61290, n61291, n61292, n61293, n61294,
         n61295, n61296, n61297, n61298, n61299, n61300, n61301, n61302,
         n61303, n61304, n61305, n61306, n61307, n61308, n61309, n61310,
         n61311, n61312, n61313, n61314, n61315, n61316, n61317, n61318,
         n61319, n61320, n61321, n61322, n61323, n61324, n61325, n61326,
         n61327, n61328, n61329, n61330, n61331, n61332, n61333, n61334,
         n61335, n61336, n61337, n61338, n61339, n61340, n61341, n61342,
         n61343, n61344, n61345, n61346, n61347, n61348, n61349, n61350,
         n61351, n61352, n61353, n61354, n61355, n61356, n61357, n61358,
         n61359, n61360, n61361, n61362, n61363, n61364, n61365, n61366,
         n61367, n61368, n61369, n61370, n61371, n61372, n61373, n61374,
         n61375, n61376, n61377, n61378, n61379, n61380, n61381, n61382,
         n61383, n61384, n61385, n61386, n61387, n61388, n61389, n61390,
         n61391, n61392, n61393, n61394, n61395, n61396, n61397, n61398,
         n61399, n61400, n61401, n61402, n61403, n61404, n61405, n61406,
         n61407, n61408, n61409, n61410, n61411, n61412, n61413, n61414,
         n61415, n61416, n61417, n61418, n61419, n61420, n61421, n61422,
         n61423, n61424, n61425, n61426, n61427, n61428, n61429, n61430,
         n61431, n61432, n61433, n61434, n61435, n61436, n61437, n61438,
         n61439, n61440, n61441, n61442, n61443, n61444, n61445, n61446,
         n61447, n61448, n61449, n61450, n61451, n61452, n61453, n61454,
         n61455, n61456, n61457, n61458, n61459, n61460, n61461, n61462,
         n61463, n61464, n61465, n61466, n61467, n61468, n61469, n61470,
         n61471, n61472, n61473, n61474, n61475, n61476, n61477, n61478,
         n61479, n61480, n61481, n61482, n61483, n61484, n61485, n61486,
         n61487, n61488, n61489, n61490, n61491, n61492, n61493, n61494,
         n61495, n61496, n61497, n61498, n61499, n61500, n61501, n61502,
         n61503, n61504, n61505, n61506, n61507, n61508, n61509, n61510,
         n61511, n61512, n61513, n61514, n61515, n61516, n61517, n61518,
         n61519, n61520, n61521, n61522, n61523, n61524, n61525, n61526,
         n61527, n61528, n61529, n61530, n61531, n61532, n61533, n61534,
         n61535, n61536, n61537, n61538, n61539, n61540, n61541, n61542,
         n61543, n61544, n61545, n61546, n61547, n61548, n61549, n61550,
         n61551, n61552, n61553, n61554, n61555, n61556, n61557, n61558,
         n61559, n61560, n61561, n61562, n61563, n61564, n61565, n61566,
         n61567, n61568, n61569, n61570, n61571, n61572, n61573, n61574,
         n61575, n61576, n61577, n61578, n61579, n61580, n61581, n61582,
         n61583, n61584, n61585, n61586, n61587, n61588, n61589, n61590,
         n61591, n61592, n61593, n61594, n61595, n61596, n61597, n61598,
         n61599, n61600, n61601, n61602, n61603, n61604, n61605, n61606,
         n61607, n61608, n61609, n61610, n61611, n61612, n61613, n61614,
         n61615, n61616, n61617, n61618, n61619, n61620, n61621, n61622,
         n61623, n61624, n61625, n61626, n61627, n61628, n61629, n61630,
         n61631, n61632, n61633, n61634, n61635, n61636, n61637, n61638,
         n61639, n61640, n61641, n61642, n61643, n61644, n61645, n61646,
         n61647, n61648, n61649, n61650, n61651, n61652, n61653, n61654,
         n61655, n61656, n61657, n61658, n61659, n61660, n61661, n61662,
         n61663, n61664, n61665, n61666, n61667, n61668, n61669, n61670,
         n61671, n61672, n61673, n61674, n61675, n61676, n61677, n61678,
         n61679, n61680, n61681, n61682, n61683, n61684, n61685, n61686,
         n61687, n61688, n61689, n61690, n61691, n61692, n61693, n61694,
         n61695, n61696, n61697, n61698, n61699, n61700, n61701, n61702,
         n61703, n61704, n61705, n61706, n61707, n61708, n61709, n61710,
         n61711, n61712, n61713, n61714, n61715, n61716, n61717, n61718,
         n61719, n61720, n61721, n61722, n61723, n61724, n61725, n61726,
         n61727, n61728, n61729, n61730, n61731, n61732, n61733, n61734,
         n61735, n61736, n61737, n61738, n61739, n61740, n61741, n61742,
         n61743, n61744, n61745, n61746, n61747, n61748, n61749, n61750,
         n61751, n61752, n61753, n61754, n61755, n61756, n61757, n61758,
         n61759, n61760, n61761, n61762, n61763, n61764, n61765, n61766,
         n61767, n61768, n61769, n61770, n61771, n61772, n61773, n61774,
         n61775, n61776, n61777, n61778, n61779, n61780, n61781, n61782,
         n61783, n61784, n61785, n61786, n61787, n61788, n61789, n61790,
         n61791, n61792, n61793, n61794, n61795, n61796, n61797, n61798,
         n61799, n61800, n61801, n61802, n61803, n61804, n61805, n61806,
         n61807, n61808, n61809, n61810, n61811, n61812, n61813, n61814,
         n61815, n61816, n61817, n61818, n61819, n61820, n61821, n61822,
         n61823, n61824, n61825, n61826, n61827, n61828, n61829, n61830,
         n61831, n61832, n61833, n61834, n61835, n61836, n61837, n61838,
         n61839, n61840, n61841, n61842, n61843, n61844, n61845, n61846,
         n61847, n61848, n61849, n61850, n61851, n61852, n61853, n61854,
         n61855, n61856, n61857, n61858, n61859, n61860, n61861, n61862,
         n61863, n61864, n61865, n61866, n61867, n61868, n61869, n61870,
         n61871, n61872, n61873, n61874, n61875, n61876, n61877, n61878,
         n61879, n61880, n61881, n61882, n61883, n61884, n61885, n61886,
         n61887, n61888, n61889, n61890, n61891, n61892, n61893, n61894,
         n61895, n61896, n61897, n61898, n61899, n61900, n61901, n61902,
         n61903, n61904, n61905, n61906, n61907, n61908, n61909, n61910,
         n61911, n61912, n61913, n61914, n61915, n61916, n61917, n61918,
         n61919, n61920, n61921, n61922, n61923, n61924, n61925, n61926,
         n61927, n61928, n61929, n61930, n61931, n61932, n61933, n61934,
         n61935, n61936, n61937, n61938, n61939, n61940, n61941, n61942,
         n61943, n61944, n61945, n61946, n61947, n61948, n61949, n61950,
         n61951, n61952, n61953, n61954, n61955, n61956, n61957, n61958,
         n61959, n61960, n61961, n61962, n61963, n61964, n61965, n61966,
         n61967, n61968, n61969, n61970, n61971, n61972, n61973, n61974,
         n61975, n61976, n61977, n61978, n61979, n61980, n61981, n61982,
         n61983, n61984, n61985, n61986, n61987, n61988, n61989, n61990,
         n61991, n61992, n61993, n61994, n61995, n61996, n61997, n61998,
         n61999, n62000, n62001, n62002, n62003, n62004, n62005, n62006,
         n62007, n62008, n62009, n62010, n62011, n62012, n62013, n62014,
         n62015, n62016, n62017, n62018, n62019, n62020, n62021, n62022,
         n62023, n62024, n62025, n62026, n62027, n62028, n62029, n62030,
         n62031, n62032, n62033, n62034, n62035, n62036, n62037, n62038,
         n62039, n62040, n62041, n62042, n62043, n62044, n62045, n62046,
         n62047, n62048, n62049, n62050, n62051, n62052, n62053, n62054,
         n62055, n62056, n62057, n62058, n62059, n62060, n62061, n62062,
         n62063, n62064, n62065, n62066, n62067, n62068, n62069, n62070,
         n62071, n62072, n62073, n62074, n62075, n62076, n62077, n62078,
         n62079, n62080, n62081, n62082, n62083, n62084, n62085, n62086,
         n62087, n62088, n62089, n62090, n62091, n62092, n62093, n62094,
         n62095, n62096, n62097, n62098, n62099, n62100, n62101, n62102,
         n62103, n62104, n62105, n62106, n62107, n62108, n62109, n62110,
         n62111, n62112, n62113, n62114, n62115, n62116, n62117, n62118,
         n62119, n62120, n62121, n62122, n62123, n62124, n62125, n62126,
         n62127, n62128, n62129, n62130, n62131, n62132, n62133, n62134,
         n62135, n62136, n62137, n62138, n62139, n62140, n62141, n62142,
         n62143, n62144, n62145, n62146, n62147, n62148, n62149, n62150,
         n62151, n62152, n62153, n62154, n62155, n62156, n62157, n62158,
         n62159, n62160, n62161, n62162, n62163, n62164, n62165, n62166,
         n62167, n62168, n62169, n62170, n62171, n62172, n62173, n62174,
         n62175, n62176, n62177, n62178, n62179, n62180, n62181, n62182,
         n62183, n62184, n62185, n62186, n62187, n62188, n62189, n62190,
         n62191, n62192, n62193, n62194, n62195, n62196, n62197, n62198,
         n62199, n62200, n62201, n62202, n62203, n62204, n62205, n62206,
         n62207, n62208, n62209, n62210, n62211, n62212, n62213, n62214,
         n62215, n62216, n62217, n62218, n62219, n62220, n62221, n62222,
         n62223, n62224, n62225, n62226, n62227, n62228, n62229, n62230,
         n62231, n62232, n62233, n62234, n62235, n62236, n62237, n62238,
         n62239, n62240, n62241, n62242, n62243, n62244, n62245, n62246,
         n62247, n62248, n62249, n62250, n62251, n62252, n62253, n62254,
         n62255, n62256, n62257, n62258, n62259, n62260, n62261, n62262,
         n62263, n62264, n62265, n62266, n62267, n62268, n62269, n62270,
         n62271, n62272, n62273, n62274, n62275, n62276, n62277, n62278,
         n62279, n62280, n62281, n62282, n62283, n62284, n62285, n62286,
         n62287, n62288, n62289, n62290, n62291, n62292, n62293, n62294,
         n62295, n62296, n62297, n62298, n62299, n62300, n62301, n62302,
         n62303, n62304, n62305, n62306, n62307, n62308, n62309, n62310,
         n62311, n62312, n62313, n62314, n62315, n62316, n62317, n62318,
         n62319, n62320, n62321, n62322, n62323, n62324, n62325, n62326,
         n62327, n62328, n62329, n62330, n62331, n62332, n62333, n62334,
         n62335, n62336, n62337, n62338, n62339, n62340, n62341, n62342,
         n62343, n62344, n62345, n62346, n62347, n62348, n62349, n62350,
         n62351, n62352, n62353, n62354, n62355, n62356, n62357, n62358,
         n62359, n62360, n62361, n62362, n62363, n62364, n62365, n62366,
         n62367, n62368, n62369, n62370, n62371, n62372, n62373, n62374,
         n62375, n62376, n62377, n62378, n62379, n62380, n62381, n62382,
         n62383, n62384, n62385, n62386, n62387, n62388, n62389, n62390,
         n62391, n62392, n62393, n62394, n62395, n62396, n62397, n62398,
         n62399, n62400, n62401, n62402, n62403, n62404, n62405, n62406,
         n62407, n62408, n62409, n62410, n62411, n62412, n62413, n62414,
         n62415, n62416, n62417, n62418, n62419, n62420, n62421, n62422,
         n62423, n62424, n62425, n62426, n62427, n62428, n62429, n62430,
         n62431, n62432, n62433, n62434, n62435, n62436, n62437, n62438,
         n62439, n62440, n62441, n62442, n62443, n62444, n62445, n62446,
         n62447, n62448, n62449, n62450, n62451, n62452, n62453, n62454,
         n62455, n62456, n62457, n62458, n62459, n62460, n62461, n62462,
         n62463, n62464, n62465, n62466, n62467, n62468, n62469, n62470,
         n62471, n62472, n62473, n62474, n62475, n62476, n62477, n62478,
         n62479, n62480, n62481, n62482, n62483, n62484, n62485, n62486,
         n62487, n62488, n62489, n62490, n62491, n62492, n62493, n62494,
         n62495, n62496, n62497, n62498, n62499, n62500, n62501, n62502,
         n62503, n62504, n62505, n62506, n62507, n62508, n62509, n62510,
         n62511, n62512, n62513, n62514, n62515, n62516, n62517, n62518,
         n62519, n62520, n62521, n62522, n62523, n62524, n62525, n62526,
         n62527, n62528, n62529, n62530, n62531, n62532, n62533, n62534,
         n62535, n62536, n62537, n62538, n62539, n62540, n62541, n62542,
         n62543, n62544, n62545, n62546, n62547, n62548, n62549, n62550,
         n62551, n62552, n62553, n62554, n62555, n62556, n62557, n62558,
         n62559, n62560, n62561, n62562, n62563, n62564, n62565, n62566,
         n62567, n62568, n62569, n62570, n62571, n62572, n62573, n62574,
         n62575, n62576, n62577, n62578, n62579, n62580, n62581, n62582,
         n62583, n62584, n62585, n62586, n62587, n62588, n62589, n62590,
         n62591, n62592, n62593, n62594, n62595, n62596, n62597, n62598,
         n62599, n62600, n62601, n62602, n62603, n62604, n62605, n62606,
         n62607, n62608, n62609, n62610, n62611, n62612, n62613, n62614,
         n62615, n62616, n62617, n62618, n62619, n62620, n62621, n62622,
         n62623, n62624, n62625, n62626, n62627, n62628, n62629, n62630,
         n62631, n62632, n62633, n62634, n62635, n62636, n62637, n62638,
         n62639, n62640, n62641, n62642, n62643, n62644, n62645, n62646,
         n62647, n62648, n62649, n62650, n62651, n62652, n62653, n62654,
         n62655, n62656, n62657, n62658, n62659, n62660, n62661, n62662,
         n62663, n62664, n62665, n62666, n62667, n62668, n62669, n62670,
         n62671, n62672, n62673, n62674, n62675, n62676, n62677, n62678,
         n62679, n62680, n62681, n62682, n62683, n62684, n62685, n62686,
         n62687, n62688, n62689, n62690, n62691, n62692, n62693, n62694,
         n62695, n62696, n62697, n62698, n62699, n62700, n62701, n62702,
         n62703, n62704, n62705, n62706, n62707, n62708, n62709, n62710,
         n62711, n62712, n62713, n62714, n62715, n62716, n62717, n62718,
         n62719, n62720, n62721, n62722, n62723, n62724, n62725, n62726,
         n62727, n62728, n62729, n62730, n62731, n62732, n62733, n62734,
         n62735, n62736, n62737, n62738, n62739, n62740, n62741, n62742,
         n62743, n62744, n62745, n62746, n62747, n62748, n62749, n62750,
         n62751, n62752, n62753, n62754, n62755, n62756, n62757, n62758,
         n62759, n62760, n62761, n62762, n62763, n62764, n62765, n62766,
         n62767, n62768, n62769, n62770, n62771, n62772, n62773, n62774,
         n62775, n62776, n62777, n62778, n62779, n62780, n62781, n62782,
         n62783, n62784, n62785, n62786, n62787, n62788, n62789, n62790,
         n62791, n62792, n62793, n62794, n62795, n62796, n62797, n62798,
         n62799, n62800, n62801, n62802, n62803, n62804, n62805, n62806,
         n62807, n62808, n62809, n62810, n62811, n62812, n62813, n62814,
         n62815, n62816, n62817, n62818, n62819, n62820, n62821, n62822,
         n62823, n62824, n62825, n62826, n62827, n62828, n62829, n62830,
         n62831, n62832, n62833, n62834, n62835, n62836, n62837, n62838,
         n62839, n62840, n62841, n62842, n62843, n62844, n62845, n62846,
         n62847, n62848, n62849, n62850, n62851, n62852, n62853, n62854,
         n62855, n62856, n62857, n62858, n62859, n62860, n62861, n62862,
         n62863, n62864, n62865, n62866, n62867, n62868, n62869, n62870,
         n62871, n62872, n62873, n62874, n62875, n62876, n62877, n62878,
         n62879, n62880, n62881, n62882, n62883, n62884, n62885, n62886,
         n62887, n62888, n62889, n62890, n62891, n62892, n62893, n62894,
         n62895, n62896, n62897, n62898, n62899, n62900, n62901, n62902,
         n62903, n62904, n62905, n62906, n62907, n62908, n62909, n62910,
         n62911, n62912, n62913, n62914, n62915, n62916, n62917, n62918,
         n62919, n62920, n62921, n62922, n62923, n62924, n62925, n62926,
         n62927, n62928, n62929, n62930, n62931, n62932, n62933, n62934,
         n62935, n62936, n62937, n62938, n62939, n62940, n62941, n62942,
         n62943, n62944, n62945, n62946, n62947, n62948, n62949, n62950,
         n62951, n62952, n62953, n62954, n62955, n62956, n62957, n62958,
         n62959, n62960, n62961, n62962, n62963, n62964, n62965, n62966,
         n62967, n62968, n62969, n62970, n62971, n62972, n62973, n62974,
         n62975, n62976, n62977, n62978, n62979, n62980, n62981, n62982,
         n62983, n62984, n62985, n62986, n62987, n62988, n62989, n62990,
         n62991, n62992, n62993, n62994, n62995, n62996, n62997, n62998,
         n62999, n63000, n63001, n63002, n63003, n63004, n63005, n63006,
         n63007, n63008, n63009, n63010, n63011, n63012, n63013, n63014,
         n63015, n63016, n63017, n63018, n63019, n63020, n63021, n63022,
         n63023, n63024, n63025, n63026, n63027, n63028, n63029, n63030,
         n63031, n63032, n63033, n63034, n63035, n63036, n63037, n63038,
         n63039, n63040, n63041, n63042, n63043, n63044, n63045, n63046,
         n63047, n63048, n63049, n63050, n63051, n63052, n63053, n63054,
         n63055, n63056, n63057, n63058, n63059, n63060, n63061, n63062,
         n63063, n63064, n63065, n63066, n63067, n63068, n63069, n63070,
         n63071, n63072, n63073, n63074, n63075, n63076, n63077, n63078,
         n63079, n63080, n63081, n63082, n63083, n63084, n63085, n63086,
         n63087, n63088, n63089, n63090, n63091, n63092, n63093, n63094,
         n63095, n63096, n63097, n63098, n63099, n63100, n63101, n63102,
         n63103, n63104, n63105, n63106, n63107, n63108, n63109, n63110,
         n63111, n63112, n63113, n63114, n63115, n63116, n63117, n63118,
         n63119, n63120, n63121, n63122, n63123, n63124, n63125, n63126,
         n63127, n63128, n63129, n63130, n63131, n63132, n63133, n63134,
         n63135, n63136, n63137, n63138, n63139, n63140, n63141, n63142,
         n63143, n63144, n63145, n63146, n63147, n63148, n63149, n63150,
         n63151, n63152, n63153, n63154, n63155, n63156, n63157, n63158,
         n63159, n63160, n63161, n63162, n63163, n63164, n63165, n63166,
         n63167, n63168, n63169, n63170, n63171, n63172, n63173, n63174,
         n63175, n63176, n63177, n63178, n63179, n63180, n63181, n63182,
         n63183, n63184, n63185, n63186, n63187, n63188, n63189, n63190,
         n63191, n63192, n63193, n63194, n63195, n63196, n63197, n63198,
         n63199, n63200, n63201, n63202, n63203, n63204, n63205, n63206,
         n63207, n63208, n63209, n63210, n63211, n63212, n63213, n63214,
         n63215, n63216, n63217, n63218, n63219, n63220, n63221, n63222,
         n63223, n63224, n63225, n63226, n63227, n63228, n63229, n63230,
         n63231, n63232, n63233, n63234, n63235, n63236, n63237, n63238,
         n63239, n63240, n63241, n63242, n63243, n63244, n63245, n63246,
         n63247, n63248, n63249, n63250, n63251, n63252, n63253, n63254,
         n63255, n63256, n63257, n63258, n63259, n63260, n63261, n63262,
         n63263, n63264, n63265, n63266, n63267, n63268, n63269, n63270,
         n63271, n63272, n63273, n63274, n63275, n63276, n63277, n63278,
         n63279, n63280, n63281, n63282, n63283, n63284, n63285, n63286,
         n63287, n63288, n63289, n63290, n63291, n63292, n63293, n63294,
         n63295, n63296, n63297, n63298, n63299, n63300, n63301, n63302,
         n63303, n63304, n63305, n63306, n63307, n63308, n63309, n63310,
         n63311, n63312, n63313, n63314, n63315, n63316, n63317, n63318,
         n63319, n63320, n63321, n63322, n63323, n63324, n63325, n63326,
         n63327, n63328, n63329, n63330, n63331, n63332, n63333, n63334,
         n63335, n63336, n63337, n63338, n63339, n63340, n63341, n63342,
         n63343, n63344, n63345, n63346, n63347, n63348, n63349, n63350,
         n63351, n63352, n63353, n63354, n63355, n63356, n63357, n63358,
         n63359, n63360, n63361, n63362, n63363, n63364, n63365, n63366,
         n63367, n63368, n63369, n63370, n63371, n63372, n63373, n63374,
         n63375, n63376, n63377, n63378, n63379, n63380, n63381, n63382,
         n63383, n63384, n63385, n63386, n63387, n63388, n63389, n63390,
         n63391, n63392, n63393, n63394, n63395, n63396, n63397, n63398,
         n63399, n63400, n63401, n63402, n63403, n63404, n63405, n63406,
         n63407, n63408, n63409, n63410, n63411, n63412, n63413, n63414,
         n63415, n63416, n63417, n63418, n63419, n63420, n63421, n63422,
         n63423, n63424, n63425, n63426, n63427, n63428, n63429, n63430,
         n63431, n63432, n63433, n63434, n63435, n63436, n63437, n63438,
         n63439, n63440, n63441, n63442, n63443, n63444, n63445, n63446,
         n63447, n63448, n63449, n63450, n63451, n63452, n63453, n63454,
         n63455, n63456, n63457, n63458, n63459, n63460, n63461, n63462,
         n63463, n63464, n63465, n63466, n63467, n63468, n63469, n63470,
         n63471, n63472, n63473, n63474, n63475, n63476, n63477, n63478,
         n63479, n63480, n63481, n63482, n63483, n63484, n63485, n63486,
         n63487, n63488, n63489, n63490, n63491, n63492, n63493, n63494,
         n63495, n63496, n63497, n63498, n63499, n63500, n63501, n63502,
         n63503, n63504, n63505, n63506, n63507, n63508, n63509, n63510,
         n63511, n63512, n63513, n63514, n63515, n63516, n63517, n63518,
         n63519, n63520, n63521, n63522, n63523, n63524, n63525, n63526,
         n63527, n63528, n63529, n63530, n63531, n63532, n63533, n63534,
         n63535, n63536, n63537, n63538, n63539, n63540, n63541, n63542,
         n63543, n63544, n63545, n63546, n63547, n63548, n63549, n63550,
         n63551, n63552, n63553, n63554, n63555, n63556, n63557, n63558,
         n63559, n63560, n63561, n63562, n63563, n63564, n63565, n63566,
         n63567, n63568, n63569, n63570, n63571, n63572, n63573, n63574,
         n63575, n63576, n63577, n63578, n63579, n63580, n63581, n63582,
         n63583, n63584, n63585, n63586, n63587, n63588, n63589, n63590,
         n63591, n63592, n63593, n63594, n63595, n63596, n63597, n63598,
         n63599, n63600, n63601, n63602, n63603, n63604, n63605, n63606,
         n63607, n63608, n63609, n63610, n63611, n63612, n63613, n63614,
         n63615, n63616, n63617, n63618, n63619, n63620, n63621, n63622,
         n63623, n63624, n63625, n63626, n63627, n63628, n63629, n63630,
         n63631, n63632, n63633, n63634, n63635, n63636, n63637, n63638,
         n63639, n63640, n63641, n63642, n63643, n63644, n63645, n63646,
         n63647, n63648, n63649, n63650, n63651, n63652, n63653, n63654,
         n63655, n63656, n63657, n63658, n63659, n63660, n63661, n63662,
         n63663, n63664, n63665, n63666, n63667, n63668, n63669, n63670,
         n63671, n63672, n63673, n63674, n63675, n63676, n63677, n63678,
         n63679, n63680, n63681, n63682, n63683, n63684, n63685, n63686,
         n63687, n63688, n63689, n63690, n63691, n63692, n63693, n63694,
         n63695, n63696, n63697, n63698, n63699, n63700, n63701, n63702,
         n63703, n63704, n63705, n63706, n63707, n63708, n63709, n63710,
         n63711, n63712, n63713, n63714, n63715, n63716, n63717, n63718,
         n63719, n63720, n63721, n63722, n63723, n63724, n63725, n63726,
         n63727, n63728, n63729, n63730, n63731, n63732, n63733, n63734,
         n63735, n63736, n63737, n63738, n63739, n63740, n63741, n63742,
         n63743, n63744, n63745, n63746, n63747, n63748, n63749, n63750,
         n63751, n63752, n63753, n63754, n63755, n63756, n63757, n63758,
         n63759, n63760, n63761, n63762, n63763, n63764, n63765, n63766,
         n63767, n63768, n63769, n63770, n63771, n63772, n63773, n63774,
         n63775, n63776, n63777, n63778, n63779, n63780, n63781, n63782,
         n63783, n63784, n63785, n63786, n63787, n63788, n63789, n63790,
         n63791, n63792, n63793, n63794, n63795, n63796, n63797, n63798,
         n63799, n63800, n63801, n63802, n63803, n63804, n63805, n63806,
         n63807, n63808, n63809, n63810, n63811, n63812, n63813, n63814,
         n63815, n63816, n63817, n63818, n63819, n63820, n63821, n63822,
         n63823, n63824, n63825, n63826, n63827, n63828, n63829, n63830,
         n63831, n63832, n63833, n63834, n63835, n63836, n63837, n63838,
         n63839, n63840, n63841, n63842, n63843, n63844, n63845, n63846,
         n63847, n63848, n63849, n63850, n63851, n63852, n63853, n63854,
         n63855, n63856, n63857, n63858, n63859, n63860, n63861, n63862,
         n63863, n63864, n63865, n63866, n63867, n63868, n63869, n63870,
         n63871, n63872, n63873, n63874, n63875, n63876, n63877, n63878,
         n63879, n63880, n63881, n63882, n63883, n63884, n63885, n63886,
         n63887, n63888, n63889, n63890, n63891, n63892, n63893, n63894,
         n63895, n63896, n63897, n63898, n63899, n63900, n63901, n63902,
         n63903, n63904, n63905, n63906, n63907, n63908, n63909, n63910,
         n63911, n63912, n63913, n63914, n63915, n63916, n63917, n63918,
         n63919, n63920, n63921, n63922, n63923, n63924, n63925, n63926,
         n63927, n63928, n63929, n63930, n63931, n63932, n63933, n63934,
         n63935, n63936, n63937, n63938, n63939, n63940, n63941, n63942,
         n63943, n63944, n63945, n63946, n63947, n63948, n63949, n63950,
         n63951, n63952, n63953, n63954, n63955, n63956, n63957, n63958,
         n63959, n63960, n63961, n63962, n63963, n63964, n63965, n63966,
         n63967, n63968, n63969, n63970, n63971, n63972, n63973, n63974,
         n63975, n63976, n63977, n63978, n63979, n63980, n63981, n63982,
         n63983, n63984, n63985, n63986, n63987, n63988, n63989, n63990,
         n63991, n63992, n63993, n63994, n63995, n63996, n63997, n63998,
         n63999, n64000, n64001, n64002, n64003, n64004, n64005, n64006,
         n64007, n64008, n64009, n64010, n64011, n64012, n64013, n64014,
         n64015, n64016, n64017, n64018, n64019, n64020, n64021, n64022,
         n64023, n64024, n64025, n64026, n64027, n64028, n64029, n64030,
         n64031, n64032, n64033, n64034, n64035, n64036, n64037, n64038,
         n64039, n64040, n64041, n64042, n64043, n64044, n64045, n64046,
         n64047, n64048, n64049, n64050, n64051, n64052, n64053, n64054,
         n64055, n64056, n64057, n64058, n64059, n64060, n64061, n64062,
         n64063, n64064, n64065, n64066, n64067, n64068, n64069, n64070,
         n64071, n64072, n64073, n64074, n64075, n64076, n64077, n64078,
         n64079, n64080, n64081, n64082, n64083, n64084, n64085, n64086,
         n64087, n64088, n64089, n64090, n64091, n64092, n64093, n64094,
         n64095, n64096, n64097, n64098, n64099, n64100, n64101, n64102,
         n64103, n64104, n64105, n64106, n64107, n64108, n64109, n64110,
         n64111, n64112, n64113, n64114, n64115, n64116, n64117, n64118,
         n64119, n64120, n64121, n64122, n64123, n64124, n64125, n64126,
         n64127, n64128, n64129, n64130, n64131, n64132, n64133, n64134,
         n64135, n64136, n64137, n64138, n64139, n64140, n64141, n64142,
         n64143, n64144, n64145, n64146, n64147, n64148, n64149, n64150,
         n64151, n64152, n64153, n64154, n64155, n64156, n64157, n64158,
         n64159, n64160, n64161, n64162, n64163, n64164, n64165, n64166,
         n64167, n64168, n64169, n64170, n64171, n64172, n64173, n64174,
         n64175, n64176, n64177, n64178, n64179, n64180, n64181, n64182,
         n64183, n64184, n64185, n64186, n64187, n64188, n64189, n64190,
         n64191, n64192, n64193, n64194, n64195, n64196, n64197, n64198,
         n64199, n64200, n64201, n64202, n64203, n64204, n64205, n64206,
         n64207, n64208, n64209, n64210, n64211, n64212, n64213, n64214,
         n64215, n64216, n64217, n64218, n64219, n64220, n64221, n64222,
         n64223, n64224, n64225, n64226, n64227, n64228, n64229, n64230,
         n64231, n64232, n64233, n64234, n64235, n64236, n64237, n64238,
         n64239, n64240, n64241, n64242, n64243, n64244, n64245, n64246,
         n64247, n64248, n64249, n64250, n64251, n64252, n64253, n64254,
         n64255, n64256, n64257, n64258, n64259, n64260, n64261, n64262,
         n64263, n64264, n64265, n64266, n64267, n64268, n64269, n64270,
         n64271, n64272, n64273, n64274, n64275, n64276, n64277, n64278,
         n64279, n64280, n64281, n64282, n64283, n64284, n64285, n64286,
         n64287, n64288, n64289, n64290, n64291, n64292, n64293, n64294,
         n64295, n64296, n64297, n64298, n64299, n64300, n64301, n64302,
         n64303, n64304, n64305, n64306, n64307, n64308, n64309, n64310,
         n64311, n64312, n64313, n64314, n64315, n64316, n64317, n64318,
         n64319, n64320, n64321, n64322, n64323, n64324, n64325, n64326,
         n64327, n64328, n64329, n64330, n64331, n64332, n64333, n64334,
         n64335, n64336, n64337, n64338, n64339, n64340, n64341, n64342,
         n64343, n64344, n64345, n64346, n64347, n64348, n64349, n64350,
         n64351, n64352, n64353, n64354, n64355, n64356, n64357, n64358,
         n64359, n64360, n64361, n64362, n64363, n64364, n64365, n64366,
         n64367, n64368, n64369, n64370, n64371, n64372, n64373, n64374,
         n64375, n64376, n64377, n64378, n64379, n64380, n64381, n64382,
         n64383, n64384, n64385, n64386, n64387, n64388, n64389, n64390,
         n64391, n64392, n64393, n64394, n64395, n64396, n64397, n64398,
         n64399, n64400, n64401, n64402, n64403, n64404, n64405, n64406,
         n64407, n64408, n64409, n64410, n64411, n64412, n64413, n64414,
         n64415, n64416, n64417, n64418, n64419, n64420, n64421, n64422,
         n64423, n64424, n64425, n64426, n64427, n64428, n64429, n64430,
         n64431, n64432, n64433, n64434, n64435, n64436, n64437, n64438,
         n64439, n64440, n64441, n64442, n64443, n64444, n64445, n64446,
         n64447, n64448, n64449, n64450, n64451, n64452, n64453, n64454,
         n64455, n64456, n64457, n64458, n64459, n64460, n64461, n64462,
         n64463, n64464, n64465, n64466, n64467, n64468, n64469, n64470,
         n64471, n64472, n64473, n64474, n64475, n64476, n64477, n64478,
         n64479, n64480, n64481, n64482, n64483, n64484, n64485, n64486,
         n64487, n64488, n64489, n64490, n64491, n64492, n64493, n64494,
         n64495, n64496, n64497, n64498, n64499, n64500, n64501, n64502,
         n64503, n64504, n64505, n64506, n64507, n64508, n64509, n64510,
         n64511, n64512, n64513, n64514, n64515, n64516, n64517, n64518,
         n64519, n64520, n64521, n64522, n64523, n64524, n64525, n64526,
         n64527, n64528, n64529, n64530, n64531, n64532, n64533, n64534,
         n64535, n64536, n64537, n64538, n64539, n64540, n64541, n64542,
         n64543, n64544, n64545, n64546, n64547, n64548, n64549, n64550,
         n64551, n64552, n64553, n64554, n64555, n64556, n64557, n64558,
         n64559, n64560, n64561, n64562, n64563, n64564, n64565, n64566,
         n64567, n64568, n64569, n64570, n64571, n64572, n64573, n64574,
         n64575, n64576, n64577, n64578, n64579, n64580, n64581, n64582,
         n64583, n64584, n64585, n64586, n64587, n64588, n64589, n64590,
         n64591, n64592, n64593, n64594, n64595, n64596, n64597, n64598,
         n64599, n64600, n64601, n64602, n64603, n64604, n64605, n64606,
         n64607, n64608, n64609, n64610, n64611, n64612, n64613, n64614,
         n64615, n64616, n64617, n64618, n64619, n64620, n64621, n64622,
         n64623, n64624, n64625, n64626, n64627, n64628, n64629, n64630,
         n64631, n64632, n64633, n64634, n64635, n64636, n64637, n64638,
         n64639, n64640, n64641, n64642, n64643, n64644, n64645, n64646,
         n64647, n64648, n64649, n64650, n64651, n64652, n64653, n64654,
         n64655, n64656, n64657, n64658, n64659, n64660, n64661, n64662,
         n64663, n64664, n64665, n64666, n64667, n64668, n64669, n64670,
         n64671, n64672, n64673, n64674, n64675, n64676, n64677, n64678,
         n64679, n64680, n64681, n64682, n64683, n64684, n64685, n64686,
         n64687, n64688, n64689, n64690, n64691, n64692, n64693, n64694,
         n64695, n64696, n64697, n64698, n64699, n64700, n64701, n64702,
         n64703, n64704, n64705, n64706, n64707, n64708, n64709, n64710,
         n64711, n64712, n64713, n64714, n64715, n64716, n64717, n64718,
         n64719, n64720, n64721, n64722, n64723, n64724, n64725, n64726,
         n64727, n64728, n64729, n64730, n64731, n64732, n64733, n64734,
         n64735, n64736, n64737, n64738, n64739, n64740, n64741, n64742,
         n64743, n64744, n64745, n64746, n64747, n64748, n64749, n64750,
         n64751, n64752, n64753, n64754, n64755, n64756, n64757, n64758,
         n64759, n64760, n64761, n64762, n64763, n64764, n64765, n64766,
         n64767, n64768, n64769, n64770, n64771, n64772, n64773, n64774,
         n64775, n64776, n64777, n64778, n64779, n64780, n64781, n64782,
         n64783, n64784, n64785, n64786, n64787, n64788, n64789, n64790,
         n64791, n64792, n64793, n64794, n64795, n64796, n64797, n64798,
         n64799, n64800, n64801, n64802, n64803, n64804, n64805, n64806,
         n64807, n64808, n64809, n64810, n64811, n64812, n64813, n64814,
         n64815, n64816, n64817, n64818, n64819, n64820, n64821, n64822,
         n64823, n64824, n64825, n64826, n64827, n64828, n64829, n64830,
         n64831, n64832, n64833, n64834, n64835, n64836, n64837, n64838,
         n64839, n64840, n64841, n64842, n64843, n64844, n64845, n64846,
         n64847, n64848, n64849, n64850, n64851, n64852, n64853, n64854,
         n64855, n64856, n64857, n64858, n64859, n64860, n64861, n64862,
         n64863, n64864, n64865, n64866, n64867, n64868, n64869, n64870,
         n64871, n64872, n64873, n64874, n64875, n64876, n64877, n64878,
         n64879, n64880, n64881, n64882, n64883, n64884, n64885, n64886,
         n64887, n64888, n64889, n64890, n64891, n64892, n64893, n64894,
         n64895, n64896, n64897, n64898, n64899, n64900, n64901, n64902,
         n64903, n64904, n64905, n64906, n64907, n64908, n64909, n64910,
         n64911, n64912, n64913, n64914, n64915, n64916, n64917, n64918,
         n64919, n64920, n64921, n64922, n64923, n64924, n64925, n64926,
         n64927, n64928, n64929, n64930, n64931, n64932, n64933, n64934,
         n64935, n64936, n64937, n64938, n64939, n64940, n64941, n64942,
         n64943, n64944, n64945, n64946, n64947, n64948, n64949, n64950,
         n64951, n64952, n64953, n64954, n64955, n64956, n64957, n64958,
         n64959, n64960, n64961, n64962, n64963, n64964, n64965, n64966,
         n64967, n64968, n64969, n64970, n64971, n64972, n64973, n64974,
         n64975, n64976, n64977, n64978, n64979, n64980, n64981, n64982,
         n64983, n64984, n64985, n64986, n64987, n64988, n64989, n64990,
         n64991, n64992, n64993, n64994, n64995, n64996, n64997, n64998,
         n64999, n65000, n65001, n65002, n65003, n65004, n65005, n65006,
         n65007, n65008, n65009, n65010, n65011, n65012, n65013, n65014,
         n65015, n65016, n65017, n65018, n65019, n65020, n65021, n65022,
         n65023, n65024, n65025, n65026, n65027, n65028, n65029, n65030,
         n65031, n65032, n65033, n65034, n65035, n65036, n65037, n65038,
         n65039, n65040, n65041, n65042, n65043, n65044, n65045, n65046,
         n65047, n65048, n65049, n65050, n65051, n65052, n65053, n65054,
         n65055, n65056, n65057, n65058, n65059, n65060, n65061, n65062,
         n65063, n65064, n65065, n65066, n65067, n65068, n65069, n65070,
         n65071, n65072, n65073, n65074, n65075, n65076, n65077, n65078,
         n65079, n65080, n65081, n65082, n65083, n65084, n65085, n65086,
         n65087, n65088, n65089, n65090, n65091, n65092, n65093, n65094,
         n65095, n65096, n65097, n65098, n65099, n65100, n65101, n65102,
         n65103, n65104, n65105, n65106, n65107, n65108, n65109, n65110,
         n65111, n65112, n65113, n65114, n65115, n65116, n65117, n65118,
         n65119, n65120, n65121, n65122, n65123, n65124, n65125, n65126,
         n65127, n65128, n65129, n65130, n65131, n65132, n65133, n65134,
         n65135, n65136, n65137, n65138, n65139, n65140, n65141, n65142,
         n65143, n65144, n65145, n65146, n65147, n65148, n65149, n65150,
         n65151, n65152, n65153, n65154, n65155, n65156, n65157, n65158,
         n65159, n65160, n65161, n65162, n65163, n65164, n65165, n65166,
         n65167, n65168, n65169, n65170, n65171, n65172, n65173, n65174,
         n65175, n65176, n65177, n65178, n65179, n65180, n65181, n65182,
         n65183, n65184, n65185, n65186, n65187, n65188, n65189, n65190,
         n65191, n65192, n65193, n65194, n65195, n65196, n65197, n65198,
         n65199, n65200, n65201, n65202, n65203, n65204, n65205, n65206,
         n65207, n65208, n65209, n65210, n65211, n65212, n65213, n65214,
         n65215, n65216, n65217, n65218, n65219, n65220, n65221, n65222,
         n65223, n65224, n65225, n65226, n65227, n65228, n65229, n65230,
         n65231, n65232, n65233, n65234, n65235, n65236, n65237, n65238,
         n65239, n65240, n65241, n65242, n65243, n65244, n65245, n65246,
         n65247, n65248, n65249, n65250, n65251, n65252, n65253, n65254,
         n65255, n65256, n65257, n65258, n65259, n65260, n65261, n65262,
         n65263, n65264, n65265, n65266, n65267, n65268, n65269, n65270,
         n65271, n65272, n65273, n65274, n65275, n65276, n65277, n65278,
         n65279, n65280, n65281, n65282, n65283, n65284, n65285, n65286,
         n65287, n65288, n65289, n65290, n65291, n65292, n65293, n65294,
         n65295, n65296, n65297, n65298, n65299, n65300, n65301, n65302,
         n65303, n65304, n65305, n65306, n65307, n65308, n65309, n65310,
         n65311, n65312, n65313, n65314, n65315, n65316, n65317, n65318,
         n65319, n65320, n65321, n65322, n65323, n65324, n65325, n65326,
         n65327, n65328, n65329, n65330, n65331, n65332, n65333, n65334,
         n65335, n65336, n65337, n65338, n65339, n65340, n65341, n65342,
         n65343, n65344, n65345, n65346, n65347, n65348, n65349, n65350,
         n65351, n65352, n65353, n65354, n65355, n65356, n65357, n65358,
         n65359, n65360, n65361, n65362, n65363, n65364, n65365, n65366,
         n65367, n65368, n65369, n65370, n65371, n65372, n65373, n65374,
         n65375, n65376, n65377, n65378, n65379, n65380, n65381, n65382,
         n65383, n65384, n65385, n65386, n65387, n65388, n65389, n65390,
         n65391, n65392, n65393, n65394, n65395, n65396, n65397, n65398,
         n65399, n65400, n65401, n65402, n65403, n65404, n65405, n65406,
         n65407, n65408, n65409, n65410, n65411, n65412, n65413, n65414,
         n65415, n65416, n65417, n65418, n65419, n65420, n65421, n65422,
         n65423, n65424, n65425, n65426, n65427, n65428, n65429, n65430,
         n65431, n65432, n65433, n65434, n65435, n65436, n65437, n65438,
         n65439, n65440, n65441, n65442, n65443, n65444, n65445, n65446,
         n65447, n65448, n65449, n65450, n65451, n65452, n65453, n65454,
         n65455, n65456, n65457, n65458, n65459, n65460, n65461, n65462,
         n65463, n65464, n65465, n65466, n65467, n65468, n65469, n65470,
         n65471, n65472, n65473, n65474, n65475, n65476, n65477, n65478,
         n65479, n65480, n65481, n65482, n65483, n65484, n65485, n65486,
         n65487, n65488, n65489, n65490, n65491, n65492, n65493, n65494,
         n65495, n65496, n65497, n65498, n65499, n65500, n65501, n65502,
         n65503, n65504, n65505, n65506, n65507, n65508, n65509, n65510,
         n65511, n65512, n65513, n65514, n65515, n65516, n65517, n65518,
         n65519, n65520, n65521, n65522, n65523, n65524, n65525, n65526,
         n65527, n65528, n65529, n65530, n65531, n65532, n65533, n65534,
         n65535, n65536, n65537, n65538, n65539, n65540, n65541, n65542,
         n65543, n65544, n65545, n65546, n65547, n65548, n65549, n65550,
         n65551, n65552, n65553, n65554, n65555, n65556, n65557, n65558,
         n65559, n65560, n65561, n65562, n65563, n65564, n65565, n65566,
         n65567, n65568, n65569, n65570, n65571, n65572, n65573, n65574,
         n65575, n65576, n65577, n65578, n65579, n65580, n65581, n65582,
         n65583, n65584, n65585, n65586, n65587, n65588, n65589, n65590,
         n65591, n65592, n65593, n65594, n65595, n65596, n65597, n65598,
         n65599, n65600, n65601, n65602, n65603, n65604, n65605, n65606,
         n65607, n65608, n65609, n65610, n65611, n65612, n65613, n65614,
         n65615, n65616, n65617, n65618, n65619, n65620, n65621, n65622,
         n65623, n65624, n65625, n65626, n65627, n65628, n65629, n65630,
         n65631, n65632, n65633, n65634, n65635, n65636, n65637, n65638,
         n65639, n65640, n65641, n65642, n65643, n65644, n65645, n65646,
         n65647, n65648, n65649, n65650, n65651, n65652, n65653, n65654,
         n65655, n65656, n65657, n65658, n65659, n65660, n65661, n65662,
         n65663, n65664, n65665, n65666, n65667, n65668, n65669, n65670,
         n65671, n65672, n65673, n65674, n65675, n65676, n65677, n65678,
         n65679, n65680, n65681, n65682, n65683, n65684, n65685, n65686,
         n65687, n65688, n65689, n65690, n65691, n65692, n65693, n65694,
         n65695, n65696, n65697, n65698, n65699, n65700, n65701, n65702,
         n65703, n65704, n65705, n65706, n65707, n65708, n65709, n65710,
         n65711, n65712, n65713, n65714, n65715, n65716, n65717, n65718,
         n65719, n65720, n65721, n65722, n65723, n65724, n65725, n65726,
         n65727, n65728, n65729, n65730, n65731, n65732, n65733, n65734,
         n65735, n65736, n65737, n65738, n65739, n65740, n65741, n65742,
         n65743, n65744, n65745, n65746, n65747, n65748, n65749, n65750,
         n65751, n65752, n65753, n65754, n65755, n65756, n65757, n65758,
         n65759, n65760, n65761, n65762, n65763, n65764, n65765, n65766,
         n65767, n65768, n65769, n65770, n65771, n65772, n65773, n65774,
         n65775, n65776, n65777, n65778, n65779, n65780, n65781, n65782,
         n65783, n65784, n65785, n65786, n65787, n65788, n65789, n65790,
         n65791, n65792, n65793, n65794, n65795, n65796, n65797, n65798,
         n65799, n65800, n65801, n65802, n65803, n65804, n65805, n65806,
         n65807, n65808, n65809, n65810, n65811, n65812, n65813, n65814,
         n65815, n65816, n65817, n65818, n65819, n65820, n65821, n65822,
         n65823, n65824, n65825, n65826, n65827, n65828, n65829, n65830,
         n65831, n65832, n65833, n65834, n65835, n65836, n65837, n65838,
         n65839, n65840, n65841, n65842, n65843, n65844, n65845, n65846,
         n65847, n65848, n65849, n65850, n65851, n65852, n65853, n65854,
         n65855, n65856, n65857, n65858, n65859, n65860, n65861, n65862,
         n65863, n65864, n65865, n65866, n65867, n65868, n65869, n65870,
         n65871, n65872, n65873, n65874, n65875, n65876, n65877, n65878,
         n65879, n65880, n65881, n65882, n65883, n65884, n65885, n65886,
         n65887, n65888, n65889, n65890, n65891, n65892, n65893, n65894,
         n65895, n65896, n65897, n65898, n65899, n65900, n65901, n65902,
         n65903, n65904, n65905, n65906, n65907, n65908, n65909, n65910,
         n65911, n65912, n65913, n65914, n65915, n65916, n65917, n65918,
         n65919, n65920, n65921, n65922, n65923, n65924, n65925, n65926,
         n65927, n65928, n65929, n65930, n65931, n65932, n65933, n65934,
         n65935, n65936, n65937, n65938, n65939, n65940, n65941, n65942,
         n65943, n65944, n65945, n65946, n65947, n65948, n65949, n65950,
         n65951, n65952, n65953, n65954, n65955, n65956, n65957, n65958,
         n65959, n65960, n65961, n65962, n65963, n65964, n65965, n65966,
         n65967, n65968, n65969, n65970, n65971, n65972, n65973, n65974,
         n65975, n65976, n65977, n65978, n65979, n65980, n65981, n65982,
         n65983, n65984, n65985, n65986, n65987, n65988, n65989, n65990,
         n65991, n65992, n65993, n65994, n65995, n65996, n65997, n65998,
         n65999, n66000, n66001, n66002, n66003, n66004, n66005, n66006,
         n66007, n66008, n66009, n66010, n66011, n66012, n66013, n66014,
         n66015, n66016, n66017, n66018, n66019, n66020, n66021, n66022,
         n66023, n66024, n66025, n66026, n66027, n66028, n66029, n66030,
         n66031, n66032, n66033, n66034, n66035, n66036, n66037, n66038,
         n66039, n66040, n66041, n66042, n66043, n66044, n66045, n66046,
         n66047, n66048, n66049, n66050, n66051, n66052, n66053, n66054,
         n66055, n66056, n66057, n66058, n66059, n66060, n66061, n66062,
         n66063, n66064, n66065, n66066, n66067, n66068, n66069, n66070,
         n66071, n66072, n66073, n66074, n66075, n66076, n66077, n66078,
         n66079, n66080, n66081, n66082, n66083, n66084, n66085, n66086,
         n66087, n66088, n66089, n66090, n66091, n66092, n66093, n66094,
         n66095, n66096, n66097, n66098, n66099, n66100, n66101, n66102,
         n66103, n66104, n66105, n66106, n66107, n66108, n66109, n66110,
         n66111, n66112, n66113, n66114, n66115, n66116, n66117, n66118,
         n66119, n66120, n66121, n66122, n66123, n66124, n66125, n66126,
         n66127, n66128, n66129, n66130, n66131, n66132, n66133, n66134,
         n66135, n66136, n66137, n66138, n66139, n66140, n66141, n66142,
         n66143, n66144, n66145, n66146, n66147, n66148, n66149, n66150,
         n66151, n66152, n66153, n66154, n66155, n66156, n66157, n66158,
         n66159, n66160, n66161, n66162, n66163, n66164, n66165, n66166,
         n66167, n66168, n66169, n66170, n66171, n66172, n66173, n66174,
         n66175, n66176, n66177, n66178, n66179, n66180, n66181, n66182,
         n66183, n66184, n66185, n66186, n66187, n66188, n66189, n66190,
         n66191, n66192, n66193, n66194, n66195, n66196, n66197, n66198,
         n66199, n66200, n66201, n66202, n66203, n66204, n66205, n66206,
         n66207, n66208, n66209, n66210, n66211, n66212, n66213, n66214,
         n66215, n66216, n66217, n66218, n66219, n66220, n66221, n66222,
         n66223, n66224, n66225, n66226, n66227, n66228, n66229, n66230,
         n66231, n66232, n66233, n66234, n66235, n66236, n66237, n66238,
         n66239, n66240, n66241, n66242, n66243, n66244, n66245, n66246,
         n66247, n66248, n66249, n66250, n66251, n66252, n66253, n66254,
         n66255, n66256, n66257, n66258, n66259, n66260, n66261, n66262,
         n66263, n66264, n66265, n66266, n66267, n66268, n66269, n66270,
         n66271, n66272, n66273, n66274, n66275, n66276, n66277, n66278,
         n66279, n66280, n66281, n66282, n66283, n66284, n66285, n66286,
         n66287, n66288, n66289, n66290, n66291, n66292, n66293, n66294,
         n66295, n66296, n66297, n66298, n66299, n66300, n66301, n66302,
         n66303, n66304, n66305, n66306, n66307, n66308, n66309, n66310,
         n66311, n66312, n66313, n66314, n66315, n66316, n66317, n66318,
         n66319, n66320, n66321, n66322, n66323, n66324, n66325, n66326,
         n66327, n66328, n66329, n66330, n66331, n66332, n66333, n66334,
         n66335, n66336, n66337, n66338, n66339, n66340, n66341, n66342,
         n66343, n66344, n66345, n66346, n66347, n66348, n66349, n66350,
         n66351, n66352, n66353, n66354, n66355, n66356, n66357, n66358,
         n66359, n66360, n66361, n66362, n66363, n66364, n66365, n66366,
         n66367, n66368, n66369, n66370, n66371, n66372, n66373, n66374,
         n66375, n66376, n66377, n66378, n66379, n66380, n66381, n66382,
         n66383, n66384, n66385, n66386, n66387, n66388, n66389, n66390,
         n66391, n66392, n66393, n66394, n66395, n66396, n66397, n66398,
         n66399, n66400, n66401, n66402, n66403, n66404, n66405, n66406,
         n66407, n66408, n66409, n66410, n66411, n66412, n66413, n66414,
         n66415, n66416, n66417, n66418, n66419, n66420, n66421, n66422,
         n66423, n66424, n66425, n66426, n66427, n66428, n66429, n66430,
         n66431, n66432, n66433, n66434, n66435, n66436, n66437, n66438,
         n66439, n66440, n66441, n66442, n66443, n66444, n66445, n66446,
         n66447, n66448, n66449, n66450, n66451, n66452, n66453, n66454,
         n66455, n66456, n66457, n66458, n66459, n66460, n66461, n66462,
         n66463, n66464, n66465, n66466, n66467, n66468, n66469, n66470,
         n66471, n66472, n66473, n66474, n66475, n66476, n66477, n66478,
         n66479, n66480, n66481, n66482, n66483, n66484, n66485, n66486,
         n66487, n66488, n66489, n66490, n66491, n66492, n66493, n66494,
         n66495, n66496, n66497, n66498, n66499, n66500, n66501, n66502,
         n66503, n66504, n66505, n66506, n66507, n66508, n66509, n66510,
         n66511, n66512, n66513, n66514, n66515, n66516, n66517, n66518,
         n66519, n66520, n66521, n66522, n66523, n66524, n66525, n66526,
         n66527, n66528, n66529, n66530, n66531, n66532, n66533, n66534,
         n66535, n66536, n66537, n66538, n66539, n66540, n66541, n66542,
         n66543, n66544, n66545, n66546, n66547, n66548, n66549, n66550,
         n66551, n66552, n66553, n66554, n66555, n66556, n66557, n66558,
         n66559, n66560, n66561, n66562, n66563, n66564, n66565, n66566,
         n66567, n66568, n66569, n66570, n66571, n66572, n66573, n66574,
         n66575, n66576, n66577, n66578, n66579, n66580, n66581, n66582,
         n66583, n66584, n66585, n66586, n66587, n66588, n66589, n66590,
         n66591, n66592, n66593, n66594, n66595, n66596, n66597, n66598,
         n66599, n66600, n66601, n66602, n66603, n66604, n66605, n66606,
         n66607, n66608, n66609, n66610, n66611, n66612, n66613, n66614,
         n66615, n66616, n66617, n66618, n66619, n66620, n66621, n66622,
         n66623, n66624, n66625, n66626, n66627, n66628, n66629, n66630,
         n66631, n66632, n66633, n66634, n66635, n66636, n66637, n66638,
         n66639, n66640, n66641, n66642, n66643, n66644, n66645, n66646,
         n66647, n66648, n66649, n66650, n66651, n66652, n66653, n66654,
         n66655, n66656, n66657, n66658, n66659, n66660, n66661, n66662,
         n66663, n66664, n66665, n66666, n66667, n66668, n66669, n66670,
         n66671, n66672, n66673, n66674, n66675, n66676, n66677, n66678,
         n66679, n66680, n66681, n66682, n66683, n66684, n66685, n66686,
         n66687, n66688, n66689, n66690, n66691, n66692, n66693, n66694,
         n66695, n66696, n66697, n66698, n66699, n66700, n66701, n66702,
         n66703, n66704, n66705, n66706, n66707, n66708, n66709, n66710,
         n66711, n66712, n66713, n66714, n66715, n66716, n66717, n66718,
         n66719, n66720, n66721, n66722, n66723, n66724, n66725, n66726,
         n66727, n66728, n66729, n66730, n66731, n66732, n66733, n66734,
         n66735, n66736, n66737, n66738, n66739, n66740, n66741, n66742,
         n66743, n66744, n66745, n66746, n66747, n66748, n66749, n66750,
         n66751, n66752, n66753, n66754, n66755, n66756, n66757, n66758,
         n66759, n66760, n66761, n66762, n66763, n66764, n66765, n66766,
         n66767, n66768, n66769, n66770, n66771, n66772, n66773, n66774,
         n66775, n66776, n66777, n66778, n66779, n66780, n66781, n66782,
         n66783, n66784, n66785, n66786, n66787, n66788, n66789, n66790,
         n66791, n66792, n66793, n66794, n66795, n66796, n66797, n66798,
         n66799, n66800, n66801, n66802, n66803, n66804, n66805, n66806,
         n66807, n66808, n66809, n66810, n66811, n66812, n66813, n66814,
         n66815, n66816, n66817, n66818, n66819, n66820, n66821, n66822,
         n66823, n66824, n66825, n66826, n66827, n66828, n66829, n66830,
         n66831, n66832, n66833, n66834, n66835, n66836, n66837, n66838,
         n66839, n66840, n66841, n66842, n66843, n66844, n66845, n66846,
         n66847, n66848, n66849, n66850, n66851, n66852, n66853, n66854,
         n66855, n66856, n66857, n66858, n66859, n66860, n66861, n66862,
         n66863, n66864, n66865, n66866, n66867, n66868, n66869, n66870,
         n66871, n66872, n66873, n66874, n66875, n66876, n66877, n66878,
         n66879, n66880, n66881, n66882, n66883, n66884, n66885, n66886,
         n66887, n66888, n66889, n66890, n66891, n66892, n66893, n66894,
         n66895, n66896, n66897, n66898, n66899, n66900, n66901, n66902,
         n66903, n66904, n66905, n66906, n66907, n66908, n66909, n66910,
         n66911, n66912, n66913, n66914, n66915, n66916, n66917, n66918,
         n66919, n66920, n66921, n66922, n66923, n66924, n66925, n66926,
         n66927, n66928, n66929, n66930, n66931, n66932, n66933, n66934,
         n66935, n66936, n66937, n66938, n66939, n66940, n66941, n66942,
         n66943, n66944, n66945, n66946, n66947, n66948, n66949, n66950,
         n66951, n66952, n66953, n66954, n66955, n66956, n66957, n66958,
         n66959, n66960, n66961, n66962, n66963, n66964, n66965, n66966,
         n66967, n66968, n66969, n66970, n66971, n66972, n66973, n66974,
         n66975, n66976, n66977, n66978, n66979, n66980, n66981, n66982,
         n66983, n66984, n66985, n66986, n66987, n66988, n66989, n66990,
         n66991, n66992, n66993, n66994, n66995, n66996, n66997, n66998,
         n66999, n67000, n67001, n67002, n67003, n67004, n67005, n67006,
         n67007, n67008, n67009, n67010, n67011, n67012, n67013, n67014,
         n67015, n67016, n67017, n67018, n67019, n67020, n67021, n67022,
         n67023, n67024, n67025, n67026, n67027, n67028, n67029, n67030,
         n67031, n67032, n67033, n67034, n67035, n67036, n67037, n67038,
         n67039, n67040, n67041, n67042, n67043, n67044, n67045, n67046,
         n67047, n67048, n67049, n67050, n67051, n67052, n67053, n67054,
         n67055, n67056, n67057, n67058, n67059, n67060, n67061, n67062,
         n67063, n67064, n67065, n67066, n67067, n67068, n67069, n67070,
         n67071, n67072, n67073, n67074, n67075, n67076, n67077, n67078,
         n67079, n67080, n67081, n67082, n67083, n67084, n67085, n67086,
         n67087, n67088, n67089, n67090, n67091, n67092, n67093, n67094,
         n67095, n67096, n67097, n67098, n67099, n67100, n67101, n67102,
         n67103, n67104, n67105, n67106, n67107, n67108, n67109, n67110,
         n67111, n67112, n67113, n67114, n67115, n67116, n67117, n67118,
         n67119, n67120, n67121, n67122, n67123, n67124, n67125, n67126,
         n67127, n67128, n67129, n67130, n67131, n67132, n67133, n67134,
         n67135, n67136, n67137, n67138, n67139, n67140, n67141, n67142,
         n67143, n67144, n67145, n67146, n67147, n67148, n67149, n67150,
         n67151, n67152, n67153, n67154, n67155, n67156, n67157, n67158,
         n67159, n67160, n67161, n67162, n67163, n67164, n67165, n67166,
         n67167, n67168, n67169, n67170, n67171, n67172, n67173, n67174,
         n67175, n67176, n67177, n67178, n67179, n67180, n67181, n67182,
         n67183, n67184, n67185, n67186, n67187, n67188, n67189, n67190,
         n67191, n67192, n67193, n67194, n67195, n67196, n67197, n67198,
         n67199, n67200, n67201, n67202, n67203, n67204, n67205, n67206,
         n67207, n67208, n67209, n67210, n67211, n67212, n67213, n67214,
         n67215, n67216, n67217, n67218, n67219, n67220, n67221, n67222,
         n67223, n67224, n67225, n67226, n67227, n67228, n67229, n67230,
         n67231, n67232, n67233, n67234, n67235, n67236, n67237, n67238,
         n67239, n67240, n67241, n67242, n67243, n67244, n67245, n67246,
         n67247, n67248, n67249, n67250, n67251, n67252, n67253, n67254,
         n67255, n67256, n67257, n67258, n67259, n67260, n67261, n67262,
         n67263, n67264, n67265, n67266, n67267, n67268, n67269, n67270,
         n67271, n67272, n67273, n67274, n67275, n67276, n67277, n67278,
         n67279, n67280, n67281, n67282, n67283, n67284, n67285, n67286,
         n67287, n67288, n67289, n67290, n67291, n67292, n67293, n67294,
         n67295, n67296, n67297, n67298, n67299, n67300, n67301, n67302,
         n67303, n67304, n67305, n67306, n67307, n67308, n67309, n67310,
         n67311, n67312, n67313, n67314, n67315, n67316, n67317, n67318,
         n67319, n67320, n67321, n67322, n67323, n67324, n67325, n67326,
         n67327, n67328, n67329, n67330, n67331, n67332, n67333, n67334,
         n67335, n67336, n67337, n67338, n67339, n67340, n67341, n67342,
         n67343, n67344, n67345, n67346, n67347, n67348, n67349, n67350,
         n67351, n67352, n67353, n67354, n67355, n67356, n67357, n67358,
         n67359, n67360, n67361, n67362, n67363, n67364, n67365, n67366,
         n67367, n67368, n67369, n67370, n67371, n67372, n67373, n67374,
         n67375, n67376, n67377, n67378, n67379, n67380, n67381, n67382,
         n67383, n67384, n67385, n67386, n67387, n67388, n67389, n67390,
         n67391, n67392, n67393, n67394, n67395, n67396, n67397, n67398,
         n67399, n67400, n67401, n67402, n67403, n67404, n67405, n67406,
         n67407, n67408, n67409, n67410, n67411, n67412, n67413, n67414,
         n67415, n67416, n67417, n67418, n67419, n67420, n67421, n67422,
         n67423, n67424, n67425, n67426, n67427, n67428, n67429, n67430,
         n67431, n67432, n67433, n67434, n67435, n67436, n67437, n67438,
         n67439, n67440, n67441, n67442, n67443, n67444, n67445, n67446,
         n67447, n67448, n67449, n67450, n67451, n67452, n67453, n67454,
         n67455, n67456, n67457, n67458, n67459, n67460, n67461, n67462,
         n67463, n67464, n67465, n67466, n67467, n67468, n67469, n67470,
         n67471, n67472, n67473, n67474, n67475, n67476, n67477, n67478,
         n67479, n67480, n67481, n67482, n67483, n67484, n67485, n67486,
         n67487, n67488, n67489, n67490, n67491, n67492, n67493, n67494,
         n67495, n67496, n67497, n67498, n67499, n67500, n67501, n67502,
         n67503, n67504, n67505, n67506, n67507, n67508, n67509, n67510,
         n67511, n67512, n67513, n67514, n67515, n67516, n67517, n67518,
         n67519, n67520, n67521, n67522, n67523, n67524, n67525, n67526,
         n67527, n67528, n67529, n67530, n67531, n67532, n67533, n67534,
         n67535, n67536, n67537, n67538, n67539, n67540, n67541, n67542,
         n67543, n67544, n67545, n67546, n67547, n67548, n67549, n67550,
         n67551, n67552, n67553, n67554, n67555, n67556, n67557, n67558,
         n67559, n67560, n67561, n67562, n67563, n67564, n67565, n67566,
         n67567, n67568, n67569, n67570, n67571, n67572, n67573, n67574,
         n67575, n67576, n67577, n67578, n67579, n67580, n67581, n67582,
         n67583, n67584, n67585, n67586, n67587, n67588, n67589, n67590,
         n67591, n67592, n67593, n67594, n67595, n67596, n67597, n67598,
         n67599, n67600, n67601, n67602, n67603, n67604, n67605, n67606,
         n67607, n67608, n67609, n67610, n67611, n67612, n67613, n67614,
         n67615, n67616, n67617, n67618, n67619, n67620, n67621, n67622,
         n67623, n67624, n67625, n67626, n67627, n67628, n67629, n67630,
         n67631, n67632, n67633, n67634, n67635, n67636, n67637, n67638,
         n67639, n67640, n67641, n67642, n67643, n67644, n67645, n67646,
         n67647, n67648, n67649, n67650, n67651, n67652, n67653, n67654,
         n67655, n67656, n67657, n67658, n67659, n67660, n67661, n67662,
         n67663, n67664, n67665, n67666, n67667, n67668, n67669, n67670,
         n67671, n67672, n67673, n67674, n67675, n67676, n67677, n67678,
         n67679, n67680, n67681, n67682, n67683, n67684, n67685, n67686,
         n67687, n67688, n67689, n67690, n67691, n67692, n67693, n67694,
         n67695, n67696, n67697, n67698, n67699, n67700, n67701, n67702,
         n67703, n67704, n67705, n67706, n67707, n67708, n67709, n67710,
         n67711, n67712, n67713, n67714, n67715, n67716, n67717, n67718,
         n67719, n67720, n67721, n67722, n67723, n67724, n67725, n67726,
         n67727, n67728, n67729, n67730, n67731, n67732, n67733, n67734,
         n67735, n67736, n67737, n67738, n67739, n67740, n67741, n67742,
         n67743, n67744, n67745, n67746, n67747, n67748, n67749, n67750,
         n67751, n67752, n67753, n67754, n67755, n67756, n67757, n67758,
         n67759, n67760, n67761, n67762, n67763, n67764, n67765, n67766,
         n67767, n67768, n67769, n67770, n67771, n67772, n67773, n67774,
         n67775, n67776, n67777, n67778, n67779, n67780, n67781, n67782,
         n67783, n67784, n67785, n67786, n67787, n67788, n67789, n67790,
         n67791, n67792, n67793, n67794, n67795, n67796, n67797, n67798,
         n67799, n67800, n67801, n67802, n67803, n67804, n67805, n67806,
         n67807, n67808, n67809, n67810, n67811, n67812, n67813, n67814,
         n67815, n67816, n67817, n67818, n67819, n67820, n67821, n67822,
         n67823, n67824, n67825, n67826, n67827, n67828, n67829, n67830,
         n67831, n67832, n67833, n67834, n67835, n67836, n67837, n67838,
         n67839, n67840, n67841, n67842, n67843, n67844, n67845, n67846,
         n67847, n67848, n67849, n67850, n67851, n67852, n67853, n67854,
         n67855, n67856, n67857, n67858, n67859, n67860, n67861, n67862,
         n67863, n67864, n67865, n67866, n67867, n67868, n67869, n67870,
         n67871, n67872, n67873, n67874, n67875, n67876, n67877, n67878,
         n67879, n67880, n67881, n67882, n67883, n67884, n67885, n67886,
         n67887, n67888, n67889, n67890, n67891, n67892, n67893, n67894,
         n67895, n67896, n67897, n67898, n67899, n67900, n67901, n67902,
         n67903, n67904, n67905, n67906, n67907, n67908, n67909, n67910,
         n67911, n67912, n67913, n67914, n67915, n67916, n67917, n67918,
         n67919, n67920, n67921, n67922, n67923, n67924, n67925, n67926,
         n67927, n67928, n67929, n67930, n67931, n67932, n67933, n67934,
         n67935, n67936, n67937, n67938, n67939, n67940, n67941, n67942,
         n67943, n67944, n67945, n67946, n67947, n67948, n67949, n67950,
         n67951, n67952, n67953, n67954, n67955, n67956, n67957, n67958,
         n67959, n67960, n67961, n67962, n67963, n67964, n67965, n67966,
         n67967, n67968, n67969, n67970, n67971, n67972, n67973, n67974,
         n67975, n67976, n67977, n67978, n67979, n67980, n67981, n67982,
         n67983, n67984, n67985, n67986, n67987, n67988, n67989, n67990,
         n67991, n67992, n67993, n67994, n67995, n67996, n67997, n67998,
         n67999, n68000, n68001, n68002, n68003, n68004, n68005, n68006,
         n68007, n68008, n68009, n68010, n68011, n68012, n68013, n68014,
         n68015, n68016, n68017, n68018, n68019, n68020, n68021, n68022,
         n68023, n68024, n68025, n68026, n68027, n68028, n68029, n68030,
         n68031, n68032, n68033, n68034, n68035, n68036, n68037, n68038,
         n68039, n68040, n68041, n68042, n68043, n68044, n68045, n68046,
         n68047, n68048, n68049, n68050, n68051, n68052, n68053, n68054,
         n68055, n68056, n68057, n68058, n68059, n68060, n68061, n68062,
         n68063, n68064, n68065, n68066, n68067, n68068, n68069, n68070,
         n68071, n68072, n68073, n68074, n68075, n68076, n68077, n68078,
         n68079, n68080, n68081, n68082, n68083, n68084, n68085, n68086,
         n68087, n68088, n68089, n68090, n68091, n68092, n68093, n68094,
         n68095, n68096, n68097, n68098, n68099, n68100, n68101, n68102,
         n68103, n68104, n68105, n68106, n68107, n68108, n68109, n68110,
         n68111, n68112, n68113, n68114, n68115, n68116, n68117, n68118,
         n68119, n68120, n68121, n68122, n68123, n68124, n68125, n68126,
         n68127, n68128, n68129, n68130, n68131, n68132, n68133, n68134,
         n68135, n68136, n68137, n68138, n68139, n68140, n68141, n68142,
         n68143, n68144, n68145, n68146, n68147, n68148, n68149, n68150,
         n68151, n68152, n68153, n68154, n68155, n68156, n68157, n68158,
         n68159, n68160, n68161, n68162, n68163, n68164, n68165, n68166,
         n68167, n68168, n68169, n68170, n68171, n68172, n68173, n68174,
         n68175, n68176, n68177, n68178, n68179, n68180, n68181, n68182,
         n68183, n68184, n68185, n68186, n68187, n68188, n68189, n68190,
         n68191, n68192, n68193, n68194, n68195, n68196, n68197, n68198,
         n68199, n68200, n68201, n68202, n68203, n68204, n68205, n68206,
         n68207, n68208, n68209, n68210, n68211, n68212, n68213, n68214,
         n68215, n68216, n68217, n68218, n68219, n68220, n68221, n68222,
         n68223, n68224, n68225, n68226, n68227, n68228, n68229, n68230,
         n68231, n68232, n68233, n68234, n68235, n68236, n68237, n68238,
         n68239, n68240, n68241, n68242, n68243, n68244, n68245, n68246,
         n68247, n68248, n68249, n68250, n68251, n68252, n68253, n68254,
         n68255, n68256, n68257, n68258, n68259, n68260, n68261, n68262,
         n68263, n68264, n68265, n68266, n68267, n68268, n68269, n68270,
         n68271, n68272, n68273, n68274, n68275, n68276, n68277, n68278,
         n68279, n68280, n68281, n68282, n68283, n68284, n68285, n68286,
         n68287, n68288, n68289, n68290, n68291, n68292, n68293, n68294,
         n68295, n68296, n68297, n68298, n68299, n68300, n68301, n68302,
         n68303, n68304, n68305, n68306, n68307, n68308, n68309, n68310,
         n68311, n68312, n68313, n68314, n68315, n68316, n68317, n68318,
         n68319, n68320, n68321, n68322, n68323, n68324, n68325, n68326,
         n68327, n68328, n68329, n68330, n68331, n68332, n68333, n68334,
         n68335, n68336, n68337, n68338, n68339, n68340, n68341, n68342,
         n68343, n68344, n68345, n68346, n68347, n68348, n68349, n68350,
         n68351, n68352, n68353, n68354, n68355, n68356, n68357, n68358,
         n68359, n68360, n68361, n68362, n68363, n68364, n68365, n68366,
         n68367, n68368, n68369, n68370, n68371, n68372, n68373, n68374,
         n68375, n68376, n68377, n68378, n68379, n68380, n68381, n68382,
         n68383, n68384, n68385, n68386, n68387, n68388, n68389, n68390,
         n68391, n68392, n68393, n68394, n68395, n68396, n68397, n68398,
         n68399, n68400, n68401, n68402, n68403, n68404, n68405, n68406,
         n68407, n68408, n68409, n68410, n68411, n68412, n68413, n68414,
         n68415, n68416, n68417, n68418, n68419, n68420, n68421, n68422,
         n68423, n68424, n68425, n68426, n68427, n68428, n68429, n68430,
         n68431, n68432, n68433, n68434, n68435, n68436, n68437, n68438,
         n68439, n68440, n68441, n68442, n68443, n68444, n68445, n68446,
         n68447, n68448, n68449, n68450, n68451, n68452, n68453, n68454,
         n68455, n68456, n68457, n68458, n68459, n68460, n68461, n68462,
         n68463, n68464, n68465, n68466, n68467, n68468, n68469, n68470,
         n68471, n68472, n68473, n68474, n68475, n68476, n68477, n68478,
         n68479, n68480, n68481, n68482, n68483, n68484, n68485, n68486,
         n68487, n68488, n68489, n68490, n68491, n68492, n68493, n68494,
         n68495, n68496, n68497, n68498, n68499, n68500, n68501, n68502,
         n68503, n68504, n68505, n68506, n68507, n68508, n68509, n68510,
         n68511, n68512, n68513, n68514, n68515, n68516, n68517, n68518,
         n68519, n68520, n68521, n68522, n68523, n68524, n68525, n68526,
         n68527, n68528, n68529, n68530, n68531, n68532, n68533, n68534,
         n68535, n68536, n68537, n68538, n68539, n68540, n68541, n68542,
         n68543, n68544, n68545, n68546, n68547, n68548, n68549, n68550,
         n68551, n68552, n68553, n68554, n68555, n68556, n68557, n68558,
         n68559, n68560, n68561, n68562, n68563, n68564, n68565, n68566,
         n68567, n68568, n68569, n68570, n68571, n68572, n68573, n68574,
         n68575, n68576, n68577, n68578, n68579, n68580, n68581, n68582,
         n68583, n68584, n68585, n68586, n68587, n68588, n68589, n68590,
         n68591, n68592, n68593, n68594, n68595, n68596, n68597, n68598,
         n68599, n68600, n68601, n68602, n68603, n68604, n68605, n68606,
         n68607, n68608, n68609, n68610, n68611, n68612, n68613, n68614,
         n68615, n68616, n68617, n68618, n68619, n68620, n68621, n68622,
         n68623, n68624, n68625, n68626, n68627, n68628, n68629, n68630,
         n68631, n68632, n68633, n68634, n68635, n68636, n68637, n68638,
         n68639, n68640, n68641, n68642, n68643, n68644, n68645, n68646,
         n68647, n68648, n68649, n68650, n68651, n68652, n68653, n68654,
         n68655, n68656, n68657, n68658, n68659, n68660, n68661, n68662,
         n68663, n68664, n68665, n68666, n68667, n68668, n68669, n68670,
         n68671, n68672, n68673, n68674, n68675, n68676, n68677, n68678,
         n68679, n68680, n68681, n68682, n68683, n68684, n68685, n68686,
         n68687, n68688, n68689, n68690, n68691, n68692, n68693, n68694,
         n68695, n68696, n68697, n68698, n68699, n68700, n68701, n68702,
         n68703, n68704, n68705, n68706, n68707, n68708, n68709, n68710,
         n68711, n68712, n68713, n68714, n68715, n68716, n68717, n68718,
         n68719, n68720, n68721, n68722, n68723, n68724, n68725, n68726,
         n68727, n68728, n68729, n68730, n68731, n68732, n68733, n68734,
         n68735, n68736, n68737, n68738, n68739, n68740, n68741, n68742,
         n68743, n68744, n68745, n68746, n68747, n68748, n68749, n68750,
         n68751, n68752, n68753, n68754, n68755, n68756, n68757, n68758,
         n68759, n68760, n68761, n68762, n68763, n68764, n68765, n68766,
         n68767, n68768, n68769, n68770, n68771, n68772, n68773, n68774,
         n68775, n68776, n68777, n68778, n68779, n68780, n68781, n68782,
         n68783, n68784, n68785, n68786, n68787, n68788, n68789, n68790,
         n68791, n68792, n68793, n68794, n68795, n68796, n68797, n68798,
         n68799, n68800, n68801, n68802, n68803, n68804, n68805, n68806,
         n68807, n68808, n68809, n68810, n68811, n68812, n68813, n68814,
         n68815, n68816, n68817, n68818, n68819, n68820, n68821, n68822,
         n68823, n68824, n68825, n68826, n68827, n68828, n68829, n68830,
         n68831, n68832, n68833, n68834, n68835, n68836, n68837, n68838,
         n68839, n68840, n68841, n68842, n68843, n68844, n68845, n68846,
         n68847, n68848, n68849, n68850, n68851, n68852, n68853, n68854,
         n68855, n68856, n68857, n68858, n68859, n68860, n68861, n68862,
         n68863, n68864, n68865, n68866, n68867, n68868, n68869, n68870,
         n68871, n68872, n68873, n68874, n68875, n68876, n68877, n68878,
         n68879, n68880, n68881, n68882, n68883, n68884, n68885, n68886,
         n68887, n68888, n68889, n68890, n68891, n68892, n68893, n68894,
         n68895, n68896, n68897, n68898, n68899, n68900, n68901, n68902,
         n68903, n68904, n68905, n68906, n68907, n68908, n68909, n68910,
         n68911, n68912, n68913, n68914, n68915, n68916, n68917, n68918,
         n68919, n68920, n68921, n68922, n68923, n68924, n68925, n68926,
         n68927, n68928, n68929, n68930, n68931, n68932, n68933, n68934,
         n68935, n68936, n68937, n68938, n68939, n68940, n68941, n68942,
         n68943, n68944, n68945, n68946, n68947, n68948, n68949, n68950,
         n68951, n68952, n68953, n68954, n68955, n68956, n68957, n68958,
         n68959, n68960, n68961, n68962, n68963, n68964, n68965, n68966,
         n68967, n68968, n68969, n68970, n68971, n68972, n68973, n68974,
         n68975, n68976, n68977, n68978, n68979, n68980, n68981, n68982,
         n68983, n68984, n68985, n68986, n68987, n68988, n68989, n68990,
         n68991, n68992, n68993, n68994, n68995, n68996, n68997, n68998,
         n68999, n69000, n69001, n69002, n69003, n69004, n69005, n69006,
         n69007, n69008, n69009, n69010, n69011, n69012, n69013, n69014,
         n69015, n69016, n69017, n69018, n69019, n69020, n69021, n69022,
         n69023, n69024, n69025, n69026, n69027, n69028, n69029, n69030,
         n69031, n69032, n69033, n69034, n69035, n69036, n69037, n69038,
         n69039, n69040, n69041, n69042, n69043, n69044, n69045, n69046,
         n69047, n69048, n69049, n69050, n69051, n69052, n69053, n69054,
         n69055, n69056, n69057, n69058, n69059, n69060, n69061, n69062,
         n69063, n69064, n69065, n69066, n69067, n69068, n69069, n69070,
         n69071, n69072, n69073, n69074, n69075, n69076, n69077, n69078,
         n69079, n69080, n69081, n69082, n69083, n69084, n69085, n69086,
         n69087, n69088, n69089, n69090, n69091, n69092, n69093, n69094,
         n69095, n69096, n69097, n69098, n69099, n69100, n69101, n69102,
         n69103, n69104, n69105, n69106, n69107, n69108, n69109, n69110,
         n69111, n69112, n69113, n69114, n69115, n69116, n69117, n69118,
         n69119, n69120, n69121, n69122, n69123, n69124, n69125, n69126,
         n69127, n69128, n69129, n69130, n69131, n69132, n69133, n69134,
         n69135, n69136, n69137, n69138, n69139, n69140, n69141, n69142,
         n69143, n69144, n69145, n69146, n69147, n69148, n69149, n69150,
         n69151, n69152, n69153, n69154, n69155, n69156, n69157, n69158,
         n69159, n69160, n69161, n69162, n69163, n69164, n69165, n69166,
         n69167, n69168, n69169, n69170, n69171, n69172, n69173, n69174,
         n69175, n69176, n69177, n69178, n69179, n69180, n69181, n69182,
         n69183, n69184, n69185, n69186, n69187, n69188, n69189, n69190,
         n69191, n69192, n69193, n69194, n69195, n69196, n69197, n69198,
         n69199, n69200, n69201, n69202, n69203, n69204, n69205, n69206,
         n69207, n69208, n69209, n69210, n69211, n69212, n69213, n69214,
         n69215, n69216, n69217, n69218, n69219, n69220, n69221, n69222,
         n69223, n69224, n69225, n69226, n69227, n69228, n69229, n69230,
         n69231, n69232, n69233, n69234, n69235, n69236, n69237, n69238,
         n69239, n69240, n69241, n69242, n69243, n69244, n69245, n69246,
         n69247, n69248, n69249, n69250, n69251, n69252, n69253, n69254,
         n69255, n69256, n69257, n69258, n69259, n69260, n69261, n69262,
         n69263, n69264, n69265, n69266, n69267, n69268, n69269, n69270,
         n69271, n69272, n69273, n69274, n69275, n69276, n69277, n69278,
         n69279, n69280, n69281, n69282, n69283, n69284, n69285, n69286,
         n69287, n69288, n69289, n69290, n69291, n69292, n69293, n69294,
         n69295, n69296, n69297, n69298, n69299, n69300, n69301, n69302,
         n69303, n69304, n69305, n69306, n69307, n69308, n69309, n69310,
         n69311, n69312, n69313, n69314, n69315, n69316, n69317, n69318,
         n69319, n69320, n69321, n69322, n69323, n69324, n69325, n69326,
         n69327, n69328, n69329, n69330, n69331, n69332, n69333, n69334,
         n69335, n69336, n69337, n69338, n69339, n69340, n69341, n69342,
         n69343, n69344, n69345, n69346, n69347, n69348, n69349, n69350,
         n69351, n69352, n69353, n69354, n69355, n69356, n69357, n69358,
         n69359, n69360, n69361, n69362, n69363, n69364, n69365, n69366,
         n69367, n69368, n69369, n69370, n69371, n69372, n69373, n69374,
         n69375, n69376, n69377, n69378, n69379, n69380, n69381, n69382,
         n69383, n69384, n69385, n69386, n69387, n69388, n69389, n69390,
         n69391, n69392, n69393, n69394, n69395, n69396, n69397, n69398,
         n69399, n69400, n69401, n69402, n69403, n69404, n69405, n69406,
         n69407, n69408, n69409, n69410, n69411, n69412, n69413, n69414,
         n69415, n69416, n69417, n69418, n69419, n69420, n69421, n69422,
         n69423, n69424, n69425, n69426, n69427, n69428, n69429, n69430,
         n69431, n69432, n69433, n69434, n69435, n69436, n69437, n69438,
         n69439, n69440, n69441, n69442, n69443, n69444, n69445, n69446,
         n69447, n69448, n69449, n69450, n69451, n69452, n69453, n69454,
         n69455, n69456, n69457, n69458, n69459, n69460, n69461, n69462,
         n69463, n69464, n69465, n69466, n69467, n69468, n69469, n69470,
         n69471, n69472, n69473, n69474, n69475, n69476, n69477, n69478,
         n69479, n69480, n69481, n69482, n69483, n69484, n69485, n69486,
         n69487, n69488, n69489, n69490, n69491, n69492, n69493, n69494,
         n69495, n69496, n69497, n69498, n69499, n69500, n69501, n69502,
         n69503, n69504, n69505, n69506, n69507, n69508, n69509, n69510,
         n69511, n69512, n69513, n69514, n69515, n69516, n69517, n69518,
         n69519, n69520, n69521, n69522, n69523, n69524, n69525, n69526,
         n69527, n69528, n69529, n69530, n69531, n69532, n69533, n69534,
         n69535, n69536, n69537, n69538, n69539, n69540, n69541, n69542,
         n69543, n69544, n69545, n69546, n69547, n69548, n69549, n69550,
         n69551, n69552, n69553, n69554, n69555, n69556, n69557, n69558,
         n69559, n69560, n69561, n69562, n69563, n69564, n69565, n69566,
         n69567, n69568, n69569, n69570, n69571, n69572, n69573, n69574,
         n69575, n69576, n69577, n69578, n69579, n69580, n69581, n69582,
         n69583, n69584, n69585, n69586, n69587, n69588, n69589, n69590,
         n69591, n69592, n69593, n69594, n69595, n69596, n69597, n69598,
         n69599, n69600, n69601, n69602, n69603, n69604, n69605, n69606,
         n69607, n69608, n69609, n69610, n69611, n69612, n69613, n69614,
         n69615, n69616, n69617, n69618, n69619, n69620, n69621, n69622,
         n69623, n69624, n69625, n69626, n69627, n69628, n69629, n69630,
         n69631, n69632, n69633, n69634, n69635, n69636, n69637, n69638,
         n69639, n69640, n69641, n69642, n69643, n69644, n69645, n69646,
         n69647, n69648, n69649, n69650, n69651, n69652, n69653, n69654,
         n69655, n69656, n69657, n69658, n69659, n69660, n69661, n69662,
         n69663, n69664, n69665, n69666, n69667, n69668, n69669, n69670,
         n69671, n69672, n69673, n69674, n69675, n69676, n69677, n69678,
         n69679, n69680, n69681, n69682, n69683, n69684, n69685, n69686,
         n69687, n69688, n69689, n69690, n69691, n69692, n69693, n69694,
         n69695, n69696, n69697, n69698, n69699, n69700, n69701, n69702,
         n69703, n69704, n69705, n69706, n69707, n69708, n69709, n69710,
         n69711, n69712, n69713, n69714, n69715, n69716, n69717, n69718,
         n69719, n69720, n69721, n69722, n69723, n69724, n69725, n69726,
         n69727, n69728, n69729, n69730, n69731, n69732, n69733, n69734,
         n69735, n69736, n69737, n69738, n69739, n69740, n69741, n69742,
         n69743, n69744, n69745, n69746, n69747, n69748, n69749, n69750,
         n69751, n69752, n69753, n69754, n69755, n69756, n69757, n69758,
         n69759, n69760, n69761, n69762, n69763, n69764, n69765, n69766,
         n69767, n69768, n69769, n69770, n69771, n69772, n69773, n69774,
         n69775, n69776, n69777, n69778, n69779, n69780, n69781, n69782,
         n69783, n69784, n69785, n69786, n69787, n69788, n69789, n69790,
         n69791, n69792, n69793, n69794, n69795, n69796, n69797, n69798,
         n69799, n69800, n69801, n69802, n69803, n69804, n69805, n69806,
         n69807, n69808, n69809, n69810, n69811, n69812, n69813, n69814,
         n69815, n69816, n69817, n69818, n69819, n69820, n69821, n69822,
         n69823, n69824, n69825, n69826, n69827, n69828, n69829, n69830,
         n69831, n69832, n69833, n69834, n69835, n69836, n69837, n69838,
         n69839, n69840, n69841, n69842, n69843, n69844, n69845, n69846,
         n69847, n69848, n69849, n69850, n69851, n69852, n69853, n69854,
         n69855, n69856, n69857, n69858, n69859, n69860, n69861, n69862,
         n69863, n69864, n69865, n69866, n69867, n69868, n69869, n69870,
         n69871, n69872, n69873, n69874, n69875, n69876, n69877, n69878,
         n69879, n69880, n69881, n69882, n69883, n69884, n69885, n69886,
         n69887, n69888, n69889, n69890, n69891, n69892, n69893, n69894,
         n69895, n69896, n69897, n69898, n69899, n69900, n69901, n69902,
         n69903, n69904, n69905, n69906, n69907, n69908, n69909, n69910,
         n69911, n69912, n69913, n69914, n69915, n69916, n69917, n69918,
         n69919, n69920, n69921, n69922, n69923, n69924, n69925, n69926,
         n69927, n69928, n69929, n69930, n69931, n69932, n69933, n69934,
         n69935, n69936, n69937, n69938, n69939, n69940, n69941, n69942,
         n69943, n69944, n69945, n69946, n69947, n69948, n69949, n69950,
         n69951, n69952, n69953, n69954, n69955, n69956, n69957, n69958,
         n69959, n69960, n69961, n69962, n69963, n69964, n69965, n69966,
         n69967, n69968, n69969, n69970, n69971, n69972, n69973, n69974,
         n69975, n69976, n69977, n69978, n69979, n69980, n69981, n69982,
         n69983, n69984, n69985, n69986, n69987, n69988, n69989, n69990,
         n69991, n69992, n69993, n69994, n69995, n69996, n69997, n69998,
         n69999, n70000, n70001, n70002, n70003, n70004, n70005, n70006,
         n70007, n70008, n70009, n70010, n70011, n70012, n70013, n70014,
         n70015, n70016, n70017, n70018, n70019, n70020, n70021, n70022,
         n70023, n70024, n70025, n70026, n70027, n70028, n70029, n70030,
         n70031, n70032, n70033, n70034, n70035, n70036, n70037, n70038,
         n70039, n70040, n70041, n70042, n70043, n70044, n70045, n70046,
         n70047, n70048, n70049, n70050, n70051, n70052, n70053, n70054,
         n70055, n70056, n70057, n70058, n70059, n70060, n70061, n70062,
         n70063, n70064, n70065, n70066, n70067, n70068, n70069, n70070,
         n70071, n70072, n70073, n70074, n70075, n70076, n70077, n70078,
         n70079, n70080, n70081, n70082, n70083, n70084, n70085, n70086,
         n70087, n70088, n70089, n70090, n70091, n70092, n70093, n70094,
         n70095, n70096, n70097, n70098, n70099, n70100, n70101, n70102,
         n70103, n70104, n70105, n70106, n70107, n70108, n70109, n70110,
         n70111, n70112, n70113, n70114, n70115, n70116, n70117, n70118,
         n70119, n70120, n70121, n70122, n70123, n70124, n70125, n70126,
         n70127, n70128, n70129, n70130, n70131, n70132, n70133, n70134,
         n70135, n70136, n70137, n70138, n70139, n70140, n70141, n70142,
         n70143, n70144, n70145, n70146, n70147, n70148, n70149, n70150,
         n70151, n70152, n70153, n70154, n70155, n70156, n70157, n70158,
         n70159, n70160, n70161, n70162, n70163, n70164, n70165, n70166,
         n70167, n70168, n70169, n70170, n70171, n70172, n70173, n70174,
         n70175, n70176, n70177, n70178, n70179, n70180, n70181, n70182,
         n70183, n70184, n70185, n70186, n70187, n70188, n70189, n70190,
         n70191, n70192, n70193, n70194, n70195, n70196, n70197, n70198,
         n70199, n70200, n70201, n70202, n70203, n70204, n70205, n70206,
         n70207, n70208, n70209, n70210, n70211, n70212, n70213, n70214,
         n70215, n70216, n70217, n70218, n70219, n70220, n70221, n70222,
         n70223, n70224, n70225, n70226, n70227, n70228, n70229, n70230,
         n70231, n70232, n70233, n70234, n70235, n70236, n70237, n70238,
         n70239, n70240, n70241, n70242, n70243, n70244, n70245, n70246,
         n70247, n70248, n70249, n70250, n70251, n70252, n70253, n70254,
         n70255, n70256, n70257, n70258, n70259, n70260, n70261, n70262,
         n70263, n70264, n70265, n70266, n70267, n70268, n70269, n70270,
         n70271, n70272, n70273, n70274, n70275, n70276, n70277, n70278,
         n70279, n70280, n70281, n70282, n70283, n70284, n70285, n70286,
         n70287, n70288, n70289, n70290, n70291, n70292, n70293, n70294,
         n70295, n70296, n70297, n70298, n70299, n70300, n70301, n70302,
         n70303, n70304, n70305, n70306, n70307, n70308, n70309, n70310,
         n70311, n70312, n70313, n70314, n70315, n70316, n70317, n70318,
         n70319, n70320, n70321, n70322, n70323, n70324, n70325, n70326,
         n70327, n70328, n70329, n70330, n70331, n70332, n70333, n70334,
         n70335, n70336, n70337, n70338, n70339, n70340, n70341, n70342,
         n70343, n70344, n70345, n70346, n70347, n70348, n70349, n70350,
         n70351, n70352, n70353, n70354, n70355, n70356, n70357, n70358,
         n70359, n70360, n70361, n70362, n70363, n70364, n70365, n70366,
         n70367, n70368, n70369, n70370, n70371, n70372, n70373, n70374,
         n70375, n70376, n70377, n70378, n70379, n70380, n70381, n70382,
         n70383, n70384, n70385, n70386, n70387, n70388, n70389, n70390,
         n70391, n70392, n70393, n70394, n70395, n70396, n70397, n70398,
         n70399, n70400, n70401, n70402, n70403, n70404, n70405, n70406,
         n70407, n70408, n70409, n70410, n70411, n70412, n70413, n70414,
         n70415, n70416, n70417, n70418, n70419, n70420, n70421, n70422,
         n70423, n70424, n70425, n70426, n70427, n70428, n70429, n70430,
         n70431, n70432, n70433, n70434, n70435, n70436, n70437, n70438,
         n70439, n70440, n70441, n70442, n70443, n70444, n70445, n70446,
         n70447, n70448, n70449, n70450, n70451, n70452, n70453, n70454,
         n70455, n70456, n70457, n70458, n70459, n70460, n70461, n70462,
         n70463, n70464, n70465, n70466, n70467, n70468, n70469, n70470,
         n70471, n70472, n70473, n70474, n70475, n70476, n70477, n70478,
         n70479, n70480, n70481, n70482, n70483, n70484, n70485, n70486,
         n70487, n70488, n70489, n70490, n70491, n70492, n70493, n70494,
         n70495, n70496, n70497, n70498, n70499, n70500, n70501, n70502,
         n70503, n70504, n70505, n70506, n70507, n70508, n70509, n70510,
         n70511, n70512, n70513, n70514, n70515, n70516, n70517, n70518,
         n70519, n70520, n70521, n70522, n70523, n70524, n70525, n70526,
         n70527, n70528, n70529, n70530, n70531, n70532, n70533, n70534,
         n70535, n70536, n70537, n70538, n70539, n70540, n70541, n70542,
         n70543, n70544, n70545, n70546, n70547, n70548, n70549, n70550,
         n70551, n70552, n70553, n70554, n70555, n70556, n70557, n70558,
         n70559, n70560, n70561, n70562, n70563, n70564, n70565, n70566,
         n70567, n70568, n70569, n70570, n70571, n70572, n70573, n70574,
         n70575, n70576, n70577, n70578, n70579, n70580, n70581, n70582,
         n70583, n70584, n70585, n70586, n70587, n70588, n70589, n70590,
         n70591, n70592, n70593, n70594, n70595, n70596, n70597, n70598,
         n70599, n70600, n70601, n70602, n70603, n70604, n70605, n70606,
         n70607, n70608, n70609, n70610, n70611, n70612, n70613, n70614,
         n70615, n70616, n70617, n70618, n70619, n70620, n70621, n70622,
         n70623, n70624, n70625, n70626, n70627, n70628, n70629, n70630,
         n70631, n70632, n70633, n70634, n70635, n70636, n70637, n70638,
         n70639, n70640, n70641, n70642, n70643, n70644, n70645, n70646,
         n70647, n70648, n70649, n70650, n70651, n70652, n70653, n70654,
         n70655, n70656, n70657, n70658, n70659, n70660, n70661, n70662,
         n70663, n70664, n70665, n70666, n70667, n70668, n70669, n70670,
         n70671, n70672, n70673, n70674, n70675, n70676, n70677, n70678,
         n70679, n70680, n70681, n70682, n70683, n70684, n70685, n70686,
         n70687, n70688, n70689, n70690, n70691, n70692, n70693, n70694,
         n70695, n70696, n70697, n70698, n70699, n70700, n70701, n70702,
         n70703, n70704, n70705, n70706, n70707, n70708, n70709, n70710,
         n70711, n70712, n70713, n70714, n70715, n70716, n70717, n70718,
         n70719, n70720, n70721, n70722, n70723, n70724, n70725, n70726,
         n70727, n70728, n70729, n70730, n70731, n70732, n70733, n70734,
         n70735, n70736, n70737, n70738, n70739, n70740, n70741, n70742,
         n70743, n70744, n70745, n70746, n70747, n70748, n70749, n70750,
         n70751, n70752, n70753, n70754, n70755, n70756, n70757, n70758,
         n70759, n70760, n70761, n70762, n70763, n70764, n70765, n70766,
         n70767, n70768, n70769, n70770, n70771, n70772, n70773, n70774,
         n70775, n70776, n70777, n70778, n70779, n70780, n70781, n70782,
         n70783, n70784, n70785, n70786, n70787, n70788, n70789, n70790,
         n70791, n70792, n70793, n70794, n70795, n70796, n70797, n70798,
         n70799, n70800, n70801, n70802, n70803, n70804, n70805, n70806,
         n70807, n70808, n70809, n70810, n70811, n70812, n70813, n70814,
         n70815, n70816, n70817, n70818, n70819, n70820, n70821, n70822,
         n70823, n70824, n70825, n70826, n70827, n70828, n70829, n70830,
         n70831, n70832, n70833, n70834, n70835, n70836, n70837, n70838,
         n70839, n70840, n70841, n70842, n70843, n70844, n70845, n70846,
         n70847, n70848, n70849, n70850, n70851, n70852, n70853, n70854,
         n70855, n70856, n70857, n70858, n70859, n70860, n70861, n70862,
         n70863, n70864, n70865, n70866, n70867, n70868, n70869, n70870,
         n70871, n70872, n70873, n70874, n70875, n70876, n70877, n70878,
         n70879, n70880, n70881, n70882, n70883, n70884, n70885, n70886,
         n70887, n70888, n70889, n70890, n70891, n70892, n70893, n70894,
         n70895, n70896, n70897, n70898, n70899, n70900, n70901, n70902,
         n70903, n70904, n70905, n70906, n70907, n70908, n70909, n70910,
         n70911, n70912, n70913, n70914, n70915, n70916, n70917, n70918,
         n70919, n70920, n70921, n70922, n70923, n70924, n70925, n70926,
         n70927, n70928, n70929, n70930, n70931, n70932, n70933, n70934,
         n70935, n70936, n70937, n70938, n70939, n70940, n70941, n70942,
         n70943, n70944, n70945, n70946, n70947, n70948, n70949, n70950,
         n70951, n70952, n70953, n70954, n70955, n70956, n70957, n70958,
         n70959, n70960, n70961, n70962, n70963, n70964, n70965, n70966,
         n70967, n70968, n70969, n70970, n70971, n70972, n70973, n70974,
         n70975, n70976, n70977, n70978, n70979, n70980, n70981, n70982,
         n70983, n70984, n70985, n70986, n70987, n70988, n70989, n70990,
         n70991, n70992, n70993, n70994, n70995, n70996, n70997, n70998,
         n70999, n71000, n71001, n71002, n71003, n71004, n71005, n71006,
         n71007, n71008, n71009, n71010, n71011, n71012, n71013, n71014,
         n71015, n71016, n71017, n71018, n71019, n71020, n71021, n71022,
         n71023, n71024, n71025, n71026, n71027, n71028, n71029, n71030,
         n71031, n71032, n71033, n71034, n71035, n71036, n71037, n71038,
         n71039, n71040, n71041, n71042, n71043, n71044, n71045, n71046,
         n71047, n71048, n71049, n71050, n71051, n71052, n71053, n71054,
         n71055, n71056, n71057, n71058, n71059, n71060, n71061, n71062,
         n71063, n71064, n71065, n71066, n71067, n71068, n71069, n71070,
         n71071, n71072, n71073, n71074, n71075, n71076, n71077, n71078,
         n71079, n71080, n71081, n71082, n71083, n71084, n71085, n71086,
         n71087, n71088, n71089, n71090, n71091, n71092, n71093, n71094,
         n71095, n71096, n71097, n71098, n71099, n71100, n71101, n71102,
         n71103, n71104, n71105, n71106, n71107, n71108, n71109, n71110,
         n71111, n71112, n71113, n71114, n71115, n71116, n71117, n71118,
         n71119, n71120, n71121, n71122, n71123, n71124, n71125, n71126,
         n71127, n71128, n71129, n71130, n71131, n71132, n71133, n71134,
         n71135, n71136, n71137, n71138, n71139, n71140, n71141, n71142,
         n71143, n71144, n71145, n71146, n71147, n71148, n71149, n71150,
         n71151, n71152, n71153, n71154, n71155, n71156, n71157, n71158,
         n71159, n71160, n71161, n71162, n71163, n71164, n71165, n71166,
         n71167, n71168, n71169, n71170, n71171, n71172, n71173, n71174,
         n71175, n71176, n71177, n71178, n71179, n71180, n71181, n71182,
         n71183, n71184, n71185, n71186, n71187, n71188, n71189, n71190,
         n71191, n71192, n71193, n71194, n71195, n71196, n71197, n71198,
         n71199, n71200, n71201, n71202, n71203, n71204, n71205, n71206,
         n71207, n71208, n71209, n71210, n71211, n71212, n71213, n71214,
         n71215, n71216, n71217, n71218, n71219, n71220, n71221, n71222,
         n71223, n71224, n71225, n71226, n71227, n71228, n71229, n71230,
         n71231, n71232, n71233, n71234, n71235, n71236, n71237, n71238,
         n71239, n71240, n71241, n71242, n71243, n71244, n71245, n71246,
         n71247, n71248, n71249, n71250, n71251, n71252, n71253, n71254,
         n71255, n71256, n71257, n71258, n71259, n71260, n71261, n71262,
         n71263, n71264, n71265, n71266, n71267, n71268, n71269, n71270,
         n71271, n71272, n71273, n71274, n71275, n71276, n71277, n71278,
         n71279, n71280, n71281, n71282, n71283, n71284, n71285, n71286,
         n71287, n71288, n71289, n71290, n71291, n71292, n71293, n71294,
         n71295, n71296, n71297, n71298, n71299, n71300, n71301, n71302,
         n71303, n71304, n71305, n71306, n71307, n71308, n71309, n71310,
         n71311, n71312, n71313, n71314, n71315, n71316, n71317, n71318,
         n71319, n71320, n71321, n71322, n71323, n71324, n71325, n71326,
         n71327, n71328, n71329, n71330, n71331, n71332, n71333, n71334,
         n71335, n71336, n71337, n71338, n71339, n71340, n71341, n71342,
         n71343, n71344, n71345, n71346, n71347, n71348, n71349, n71350,
         n71351, n71352, n71353, n71354, n71355, n71356, n71357, n71358,
         n71359, n71360, n71361, n71362, n71363, n71364, n71365, n71366,
         n71367, n71368, n71369, n71370, n71371, n71372, n71373, n71374,
         n71375, n71376, n71377, n71378, n71379, n71380, n71381, n71382,
         n71383, n71384, n71385, n71386, n71387, n71388, n71389, n71390,
         n71391, n71392, n71393, n71394, n71395, n71396, n71397, n71398,
         n71399, n71400, n71401, n71402, n71403, n71404, n71405, n71406,
         n71407, n71408, n71409, n71410, n71411, n71412, n71413, n71414,
         n71415, n71416, n71417, n71418, n71419, n71420, n71421, n71422,
         n71423, n71424, n71425, n71426, n71427, n71428, n71429, n71430,
         n71431, n71432, n71433, n71434, n71435, n71436, n71437, n71438,
         n71439, n71440, n71441, n71442, n71443, n71444, n71445, n71446,
         n71447, n71448, n71449, n71450, n71451, n71452, n71453, n71454,
         n71455, n71456, n71457, n71458, n71459, n71460, n71461, n71462,
         n71463, n71464, n71465, n71466, n71467, n71468, n71469, n71470,
         n71471, n71472, n71473, n71474, n71475, n71476, n71477, n71478,
         n71479, n71480, n71481, n71482, n71483, n71484, n71485, n71486,
         n71487, n71488, n71489, n71490, n71491, n71492, n71493, n71494,
         n71495, n71496, n71497, n71498, n71499, n71500, n71501, n71502,
         n71503, n71504, n71505, n71506, n71507, n71508, n71509, n71510,
         n71511, n71512, n71513, n71514, n71515, n71516, n71517, n71518,
         n71519, n71520, n71521, n71522, n71523, n71524, n71525, n71526,
         n71527, n71528, n71529, n71530, n71531, n71532, n71533, n71534,
         n71535, n71536, n71537, n71538, n71539, n71540, n71541, n71542,
         n71543, n71544, n71545, n71546, n71547, n71548, n71549, n71550,
         n71551, n71552, n71553, n71554, n71555, n71556, n71557, n71558,
         n71559, n71560, n71561, n71562, n71563, n71564, n71565, n71566,
         n71567, n71568, n71569, n71570, n71571, n71572, n71573, n71574,
         n71575, n71576, n71577, n71578, n71579, n71580, n71581, n71582,
         n71583, n71584, n71585, n71586, n71587, n71588, n71589, n71590,
         n71591, n71592, n71593, n71594, n71595, n71596, n71597, n71598,
         n71599, n71600, n71601, n71602, n71603, n71604, n71605, n71606,
         n71607, n71608, n71609, n71610, n71611, n71612, n71613, n71614,
         n71615, n71616, n71617, n71618, n71619, n71620, n71621, n71622,
         n71623, n71624, n71625, n71626, n71627, n71628, n71629, n71630,
         n71631, n71632, n71633, n71634, n71635, n71636, n71637, n71638,
         n71639, n71640, n71641, n71642, n71643, n71644, n71645, n71646,
         n71647, n71648, n71649, n71650, n71651, n71652, n71653, n71654,
         n71655, n71656, n71657, n71658, n71659, n71660, n71661, n71662,
         n71663, n71664, n71665, n71666, n71667, n71668, n71669, n71670,
         n71671, n71672, n71673, n71674, n71675, n71676, n71677, n71678,
         n71679, n71680, n71681, n71682, n71683, n71684, n71685, n71686,
         n71687, n71688, n71689, n71690, n71691, n71692, n71693, n71694,
         n71695, n71696, n71697, n71698, n71699, n71700, n71701, n71702,
         n71703, n71704, n71705, n71706, n71707, n71708, n71709, n71710,
         n71711, n71712, n71713, n71714, n71715, n71716, n71717, n71718,
         n71719, n71720, n71721, n71722, n71723, n71724, n71725, n71726,
         n71727, n71728, n71729, n71730, n71731, n71732, n71733, n71734,
         n71735, n71736, n71737, n71738, n71739, n71740, n71741, n71742,
         n71743, n71744, n71745, n71746, n71747, n71748, n71749, n71750,
         n71751, n71752, n71753, n71754, n71755, n71756, n71757, n71758,
         n71759, n71760, n71761, n71762, n71763, n71764, n71765, n71766,
         n71767, n71768, n71769, n71770, n71771, n71772, n71773, n71774,
         n71775, n71776, n71777, n71778, n71779, n71780, n71781, n71782,
         n71783, n71784, n71785, n71786, n71787, n71788, n71789, n71790,
         n71791, n71792, n71793, n71794, n71795, n71796, n71797, n71798,
         n71799, n71800, n71801, n71802, n71803, n71804, n71805, n71806,
         n71807, n71808, n71809, n71810, n71811, n71812, n71813, n71814,
         n71815, n71816, n71817, n71818, n71819, n71820, n71821, n71822,
         n71823, n71824, n71825, n71826, n71827, n71828, n71829, n71830,
         n71831, n71832, n71833, n71834, n71835, n71836, n71837, n71838,
         n71839, n71840, n71841, n71842, n71843, n71844, n71845, n71846,
         n71847, n71848, n71849, n71850, n71851, n71852, n71853, n71854,
         n71855, n71856, n71857, n71858, n71859, n71860, n71861, n71862,
         n71863, n71864, n71865, n71866, n71867, n71868, n71869, n71870,
         n71871, n71872, n71873, n71874, n71875, n71876, n71877, n71878,
         n71879, n71880, n71881, n71882, n71883, n71884, n71885, n71886,
         n71887, n71888, n71889, n71890, n71891, n71892, n71893, n71894,
         n71895, n71896, n71897, n71898, n71899, n71900, n71901, n71902,
         n71903, n71904, n71905, n71906, n71907, n71908, n71909, n71910,
         n71911, n71912, n71913, n71914, n71915, n71916, n71917, n71918,
         n71919, n71920, n71921, n71922, n71923, n71924, n71925, n71926,
         n71927, n71928, n71929, n71930, n71931, n71932, n71933, n71934,
         n71935, n71936, n71937, n71938, n71939, n71940, n71941, n71942,
         n71943, n71944, n71945, n71946, n71947, n71948, n71949, n71950,
         n71951, n71952, n71953, n71954, n71955, n71956, n71957, n71958,
         n71959, n71960, n71961, n71962, n71963, n71964, n71965, n71966,
         n71967, n71968, n71969, n71970, n71971, n71972, n71973, n71974,
         n71975, n71976, n71977, n71978, n71979, n71980, n71981, n71982,
         n71983, n71984, n71985, n71986, n71987, n71988, n71989, n71990,
         n71991, n71992, n71993, n71994, n71995, n71996, n71997, n71998,
         n71999, n72000, n72001, n72002, n72003, n72004, n72005, n72006,
         n72007, n72008, n72009, n72010, n72011, n72012, n72013, n72014,
         n72015, n72016, n72017, n72018, n72019, n72020, n72021, n72022,
         n72023, n72024, n72025, n72026, n72027, n72028, n72029, n72030,
         n72031, n72032, n72033, n72034, n72035, n72036, n72037, n72038,
         n72039, n72040, n72041, n72042, n72043, n72044, n72045, n72046,
         n72047, n72048, n72049, n72050, n72051, n72052, n72053, n72054,
         n72055, n72056, n72057, n72058, n72059, n72060, n72061, n72062,
         n72063, n72064, n72065, n72066, n72067, n72068, n72069, n72070,
         n72071, n72072, n72073, n72074, n72075, n72076, n72077, n72078,
         n72079, n72080, n72081, n72082, n72083, n72084, n72085, n72086,
         n72087, n72088, n72089, n72090, n72091, n72092, n72093, n72094,
         n72095, n72096, n72097, n72098, n72099, n72100, n72101, n72102,
         n72103, n72104, n72105, n72106, n72107, n72108, n72109, n72110,
         n72111, n72112, n72113, n72114, n72115, n72116, n72117, n72118,
         n72119, n72120, n72121, n72122, n72123, n72124, n72125, n72126,
         n72127, n72128, n72129, n72130, n72131, n72132, n72133, n72134,
         n72135, n72136, n72137, n72138, n72139, n72140, n72141, n72142,
         n72143, n72144, n72145, n72146, n72147, n72148, n72149, n72150,
         n72151, n72152, n72153, n72154, n72155, n72156, n72157, n72158,
         n72159, n72160, n72161, n72162, n72163, n72164, n72165, n72166,
         n72167, n72168, n72169, n72170, n72171, n72172, n72173, n72174,
         n72175, n72176, n72177, n72178, n72179, n72180, n72181, n72182,
         n72183, n72184, n72185, n72186, n72187, n72188, n72189, n72190,
         n72191, n72192, n72193, n72194, n72195, n72196, n72197, n72198,
         n72199, n72200, n72201, n72202, n72203, n72204, n72205, n72206,
         n72207, n72208, n72209, n72210, n72211, n72212, n72213, n72214,
         n72215, n72216, n72217, n72218, n72219, n72220, n72221, n72222,
         n72223, n72224, n72225, n72226, n72227, n72228, n72229, n72230,
         n72231, n72232, n72233, n72234, n72235, n72236, n72237, n72238,
         n72239, n72240, n72241, n72242, n72243, n72244, n72245, n72246,
         n72247, n72248, n72249, n72250, n72251, n72252, n72253, n72254,
         n72255, n72256, n72257, n72258, n72259, n72260, n72261, n72262,
         n72263, n72264, n72265, n72266, n72267, n72268, n72269, n72270,
         n72271, n72272, n72273, n72274, n72275, n72276, n72277, n72278,
         n72279, n72280, n72281, n72282, n72283, n72284, n72285, n72286,
         n72287, n72288, n72289, n72290, n72291, n72292, n72293, n72294,
         n72295, n72296, n72297, n72298, n72299, n72300, n72301, n72302,
         n72303, n72304, n72305, n72306, n72307, n72308, n72309, n72310,
         n72311, n72312, n72313, n72314, n72315, n72316, n72317, n72318,
         n72319, n72320, n72321, n72322, n72323, n72324, n72325, n72326,
         n72327, n72328, n72329, n72330, n72331, n72332, n72333, n72334,
         n72335, n72336, n72337, n72338, n72339, n72340, n72341, n72342,
         n72343, n72344, n72345, n72346, n72347, n72348, n72349, n72350,
         n72351, n72352, n72353, n72354, n72355, n72356, n72357, n72358,
         n72359, n72360, n72361, n72362, n72363, n72364, n72365, n72366,
         n72367, n72368, n72369, n72370, n72371, n72372, n72373, n72374,
         n72375, n72376, n72377, n72378, n72379, n72380, n72381, n72382,
         n72383, n72384, n72385, n72386, n72387, n72388, n72389, n72390,
         n72391, n72392, n72393, n72394, n72395, n72396, n72397, n72398,
         n72399, n72400, n72401, n72402, n72403, n72404, n72405, n72406,
         n72407, n72408, n72409, n72410, n72411, n72412, n72413, n72414,
         n72415, n72416, n72417, n72418, n72419, n72420, n72421, n72422,
         n72423, n72424, n72425, n72426, n72427, n72428, n72429, n72430,
         n72431, n72432, n72433, n72434, n72435, n72436, n72437, n72438,
         n72439, n72440, n72441, n72442, n72443, n72444, n72445, n72446,
         n72447, n72448, n72449, n72450, n72451, n72452, n72453, n72454,
         n72455, n72456, n72457, n72458, n72459, n72460, n72461, n72462,
         n72463, n72464, n72465, n72466, n72467, n72468, n72469, n72470,
         n72471, n72472, n72473, n72474, n72475, n72476, n72477, n72478,
         n72479, n72480, n72481, n72482, n72483, n72484, n72485, n72486,
         n72487, n72488, n72489, n72490, n72491, n72492, n72493, n72494,
         n72495, n72496, n72497, n72498, n72499, n72500, n72501, n72502,
         n72503, n72504, n72505, n72506, n72507, n72508, n72509, n72510,
         n72511, n72512, n72513, n72514, n72515, n72516, n72517, n72518,
         n72519, n72520, n72521, n72522, n72523, n72524, n72525, n72526,
         n72527, n72528, n72529, n72530, n72531, n72532, n72533, n72534,
         n72535, n72536, n72537, n72538, n72539, n72540, n72541, n72542,
         n72543, n72544, n72545, n72546, n72547, n72548, n72549, n72550,
         n72551, n72552, n72553, n72554, n72555, n72556, n72557, n72558,
         n72559, n72560, n72561, n72562, n72563, n72564, n72565, n72566,
         n72567, n72568, n72569, n72570, n72571, n72572, n72573, n72574,
         n72575, n72576, n72577, n72578, n72579, n72580, n72581, n72582,
         n72583, n72584, n72585, n72586, n72587, n72588, n72589, n72590,
         n72591, n72592, n72593, n72594, n72595, n72596, n72597, n72598,
         n72599, n72600, n72601, n72602, n72603, n72604, n72605, n72606,
         n72607, n72608, n72609, n72610, n72611, n72612, n72613, n72614,
         n72615, n72616, n72617, n72618, n72619, n72620, n72621, n72622,
         n72623, n72624, n72625, n72626, n72627, n72628, n72629, n72630,
         n72631, n72632, n72633, n72634, n72635, n72636, n72637, n72638,
         n72639, n72640, n72641, n72642, n72643, n72644, n72645, n72646,
         n72647, n72648, n72649, n72650, n72651, n72652, n72653, n72654,
         n72655, n72656, n72657, n72658, n72659, n72660, n72661, n72662,
         n72663, n72664, n72665, n72666, n72667, n72668, n72669, n72670,
         n72671, n72672, n72673, n72674, n72675, n72676, n72677, n72678,
         n72679, n72680, n72681, n72682, n72683, n72684, n72685, n72686,
         n72687, n72688, n72689, n72690, n72691, n72692, n72693, n72694,
         n72695, n72696, n72697, n72698, n72699, n72700, n72701, n72702,
         n72703, n72704, n72705, n72706, n72707, n72708, n72709, n72710,
         n72711, n72712, n72713, n72714, n72715, n72716, n72717, n72718,
         n72719, n72720, n72721, n72722, n72723, n72724, n72725, n72726,
         n72727, n72728, n72729, n72730, n72731, n72732, n72733, n72734,
         n72735, n72736, n72737, n72738, n72739, n72740, n72741, n72742,
         n72743, n72744, n72745, n72746, n72747, n72748, n72749, n72750,
         n72751, n72752, n72753, n72754, n72755, n72756, n72757, n72758,
         n72759, n72760, n72761, n72762, n72763, n72764, n72765, n72766,
         n72767, n72768, n72769, n72770, n72771, n72772, n72773, n72774,
         n72775, n72776, n72777, n72778, n72779, n72780, n72781, n72782,
         n72783, n72784, n72785, n72786, n72787, n72788, n72789, n72790,
         n72791, n72792, n72793, n72794, n72795, n72796, n72797, n72798,
         n72799, n72800, n72801, n72802, n72803, n72804, n72805, n72806,
         n72807, n72808, n72809, n72810, n72811, n72812, n72813, n72814,
         n72815, n72816, n72817, n72818, n72819, n72820, n72821, n72822,
         n72823, n72824, n72825, n72826, n72827, n72828, n72829, n72830,
         n72831, n72832, n72833, n72834, n72835, n72836, n72837, n72838,
         n72839, n72840, n72841, n72842, n72843, n72844, n72845, n72846,
         n72847, n72848, n72849, n72850, n72851, n72852, n72853, n72854,
         n72855, n72856, n72857, n72858, n72859, n72860, n72861, n72862,
         n72863, n72864, n72865, n72866, n72867, n72868, n72869, n72870,
         n72871, n72872, n72873, n72874, n72875, n72876, n72877, n72878,
         n72879, n72880, n72881, n72882, n72883, n72884, n72885, n72886,
         n72887, n72888, n72889, n72890, n72891, n72892, n72893, n72894,
         n72895, n72896, n72897, n72898, n72899, n72900, n72901, n72902,
         n72903, n72904, n72905, n72906, n72907, n72908, n72909, n72910,
         n72911, n72912, n72913, n72914, n72915, n72916, n72917, n72918,
         n72919, n72920, n72921, n72922, n72923, n72924, n72925, n72926,
         n72927, n72928, n72929, n72930, n72931, n72932, n72933, n72934,
         n72935, n72936, n72937, n72938, n72939, n72940, n72941, n72942,
         n72943, n72944, n72945, n72946, n72947, n72948, n72949, n72950,
         n72951, n72952, n72953, n72954, n72955, n72956, n72957, n72958,
         n72959, n72960, n72961, n72962, n72963, n72964, n72965, n72966,
         n72967, n72968, n72969, n72970, n72971, n72972, n72973, n72974,
         n72975, n72976, n72977, n72978, n72979, n72980, n72981, n72982,
         n72983, n72984, n72985, n72986, n72987, n72988, n72989, n72990,
         n72991, n72992, n72993, n72994, n72995, n72996, n72997, n72998,
         n72999, n73000, n73001, n73002, n73003, n73004, n73005, n73006,
         n73007, n73008, n73009, n73010, n73011, n73012, n73013, n73014,
         n73015, n73016, n73017, n73018, n73019, n73020, n73021, n73022,
         n73023, n73024, n73025, n73026, n73027, n73028, n73029, n73030,
         n73031, n73032, n73033, n73034, n73035, n73036, n73037, n73038,
         n73039, n73040, n73041, n73042, n73043, n73044, n73045, n73046,
         n73047, n73048, n73049, n73050, n73051, n73052, n73053, n73054,
         n73055, n73056, n73057, n73058, n73059, n73060, n73061, n73062,
         n73063, n73064, n73065, n73066, n73067, n73068, n73069, n73070,
         n73071, n73072, n73073, n73074, n73075, n73076, n73077, n73078,
         n73079, n73080, n73081, n73082, n73083, n73084, n73085, n73086,
         n73087, n73088, n73089, n73090, n73091, n73092, n73093, n73094,
         n73095, n73096, n73097, n73098, n73099, n73100, n73101, n73102,
         n73103, n73104, n73105, n73106, n73107, n73108, n73109, n73110,
         n73111, n73112, n73113, n73114, n73115, n73116, n73117, n73118,
         n73119, n73120, n73121, n73122, n73123, n73124, n73125, n73126,
         n73127, n73128, n73129, n73130, n73131, n73132, n73133, n73134,
         n73135, n73136, n73137, n73138, n73139, n73140, n73141, n73142,
         n73143, n73144, n73145, n73146, n73147, n73148, n73149, n73150,
         n73151, n73152, n73153, n73154, n73155, n73156, n73157, n73158,
         n73159, n73160, n73161, n73162, n73163, n73164, n73165, n73166,
         n73167, n73168, n73169, n73170, n73171, n73172, n73173, n73174,
         n73175, n73176, n73177, n73178, n73179, n73180, n73181, n73182,
         n73183, n73184, n73185, n73186, n73187, n73188, n73189, n73190,
         n73191, n73192, n73193, n73194, n73195, n73196, n73197, n73198,
         n73199, n73200, n73201, n73202, n73203, n73204, n73205, n73206,
         n73207, n73208, n73209, n73210, n73211, n73212, n73213, n73214,
         n73215, n73216, n73217, n73218, n73219, n73220, n73221, n73222,
         n73223, n73224, n73225, n73226, n73227, n73228, n73229, n73230,
         n73231, n73232, n73233, n73234, n73235, n73236, n73237, n73238,
         n73239, n73240, n73241, n73242, n73243, n73244, n73245, n73246,
         n73247, n73248, n73249, n73250, n73251, n73252, n73253, n73254,
         n73255, n73256, n73257, n73258, n73259, n73260, n73261, n73262,
         n73263, n73264, n73265, n73266, n73267, n73268, n73269, n73270,
         n73271, n73272, n73273, n73274, n73275, n73276, n73277, n73278,
         n73279, n73280, n73281, n73282, n73283, n73284, n73285, n73286,
         n73287, n73288, n73289, n73290, n73291, n73292, n73293, n73294,
         n73295, n73296, n73297, n73298, n73299, n73300, n73301, n73302,
         n73303, n73304, n73305, n73306, n73307, n73308, n73309, n73310,
         n73311, n73312, n73313, n73314, n73315, n73316, n73317, n73318,
         n73319, n73320, n73321, n73322, n73323, n73324, n73325, n73326,
         n73327, n73328, n73329, n73330, n73331, n73332, n73333, n73334,
         n73335, n73336, n73337, n73338, n73339, n73340, n73341, n73342,
         n73343, n73344, n73345, n73346, n73347, n73348, n73349, n73350,
         n73351, n73352, n73353, n73354, n73355, n73356, n73357, n73358,
         n73359, n73360, n73361, n73362, n73363, n73364, n73365, n73366,
         n73367, n73368, n73369, n73370, n73371, n73372, n73373, n73374,
         n73375, n73376, n73377, n73378, n73379, n73380, n73381, n73382,
         n73383, n73384, n73385, n73386, n73387, n73388, n73389, n73390,
         n73391, n73392, n73393, n73394, n73395, n73396, n73397, n73398,
         n73399, n73400, n73401, n73402, n73403, n73404, n73405, n73406,
         n73407, n73408, n73409, n73410, n73411, n73412, n73413, n73414,
         n73415, n73416, n73417, n73418, n73419, n73420, n73421, n73422,
         n73423, n73424, n73425, n73426, n73427, n73428, n73429, n73430,
         n73431, n73432, n73433, n73434, n73435, n73436, n73437, n73438,
         n73439, n73440, n73441, n73442, n73443, n73444, n73445, n73446,
         n73447, n73448, n73449, n73450, n73451, n73452, n73453, n73454,
         n73455, n73456, n73457, n73458, n73459, n73460, n73461, n73462,
         n73463, n73464, n73465, n73466, n73467, n73468, n73469, n73470,
         n73471, n73472, n73473, n73474, n73475, n73476, n73477, n73478,
         n73479, n73480, n73481, n73482, n73483, n73484, n73485, n73486,
         n73487, n73488, n73489, n73490, n73491, n73492, n73493, n73494,
         n73495, n73496, n73497, n73498, n73499, n73500, n73501, n73502,
         n73503, n73504, n73505, n73506, n73507, n73508, n73509, n73510,
         n73511, n73512, n73513, n73514, n73515, n73516, n73517, n73518,
         n73519, n73520, n73521, n73522, n73523, n73524, n73525, n73526,
         n73527, n73528, n73529, n73530, n73531, n73532, n73533, n73534,
         n73535, n73536, n73537, n73538, n73539, n73540, n73541, n73542,
         n73543, n73544, n73545, n73546, n73547, n73548, n73549, n73550,
         n73551, n73552, n73553, n73554, n73555, n73556, n73557, n73558,
         n73559, n73560, n73561, n73562, n73563, n73564, n73565, n73566,
         n73567, n73568, n73569, n73570, n73571, n73572, n73573, n73574,
         n73575, n73576, n73577, n73578, n73579, n73580, n73581, n73582,
         n73583, n73584, n73585, n73586, n73587, n73588, n73589, n73590,
         n73591, n73592, n73593, n73594, n73595, n73596, n73597, n73598,
         n73599, n73600, n73601, n73602, n73603, n73604, n73605, n73606,
         n73607, n73608, n73609, n73610, n73611, n73612, n73613, n73614,
         n73615, n73616, n73617, n73618, n73619, n73620, n73621, n73622,
         n73623, n73624, n73625, n73626, n73627, n73628, n73629, n73630,
         n73631, n73632, n73633, n73634, n73635, n73636, n73637, n73638,
         n73639, n73640, n73641, n73642, n73643, n73644, n73645, n73646,
         n73647, n73648, n73649, n73650, n73651, n73652, n73653, n73654,
         n73655, n73656, n73657, n73658, n73659, n73660, n73661, n73662,
         n73663, n73664, n73665, n73666, n73667, n73668, n73669, n73670,
         n73671, n73672, n73673, n73674, n73675, n73676, n73677, n73678,
         n73679, n73680, n73681, n73682, n73683, n73684, n73685, n73686,
         n73687, n73688, n73689, n73690, n73691, n73692, n73693, n73694,
         n73695, n73696, n73697, n73698, n73699, n73700, n73701, n73702,
         n73703, n73704, n73705, n73706, n73707, n73708, n73709, n73710,
         n73711, n73712, n73713, n73714, n73715, n73716, n73717, n73718,
         n73719, n73720, n73721, n73722, n73723, n73724, n73725, n73726,
         n73727, n73728, n73729, n73730, n73731, n73732, n73733, n73734,
         n73735, n73736, n73737, n73738, n73739, n73740, n73741, n73742,
         n73743, n73744, n73745, n73746, n73747, n73748, n73749, n73750,
         n73751, n73752, n73753, n73754, n73755, n73756, n73757, n73758,
         n73759, n73760, n73761, n73762, n73763, n73764, n73765, n73766,
         n73767, n73768, n73769, n73770, n73771, n73772, n73773, n73774,
         n73775, n73776, n73777, n73778, n73779, n73780, n73781, n73782,
         n73783, n73784, n73785, n73786, n73787, n73788, n73789, n73790,
         n73791, n73792, n73793, n73794, n73795, n73796, n73797, n73798,
         n73799, n73800, n73801, n73802, n73803, n73804, n73805, n73806,
         n73807, n73808, n73809, n73810, n73811, n73812, n73813, n73814,
         n73815, n73816, n73817, n73818, n73819, n73820, n73821, n73822,
         n73823, n73824, n73825, n73826, n73827, n73828, n73829, n73830,
         n73831, n73832, n73833, n73834, n73835, n73836, n73837, n73838,
         n73839, n73840, n73841, n73842, n73843, n73844, n73845, n73846,
         n73847, n73848, n73849, n73850, n73851, n73852, n73853, n73854,
         n73855, n73856, n73857, n73858, n73859, n73860, n73861, n73862,
         n73863, n73864, n73865, n73866, n73867, n73868, n73869, n73870,
         n73871, n73872, n73873, n73874, n73875, n73876, n73877, n73878,
         n73879, n73880, n73881, n73882, n73883, n73884, n73885, n73886,
         n73887, n73888, n73889, n73890, n73891, n73892, n73893, n73894,
         n73895, n73896, n73897, n73898, n73899, n73900, n73901, n73902,
         n73903, n73904, n73905, n73906, n73907, n73908, n73909, n73910,
         n73911, n73912, n73913, n73914, n73915, n73916, n73917, n73918,
         n73919, n73920, n73921, n73922, n73923, n73924, n73925, n73926,
         n73927, n73928, n73929, n73930, n73931, n73932, n73933, n73934,
         n73935, n73936, n73937, n73938, n73939, n73940, n73941, n73942,
         n73943, n73944, n73945, n73946, n73947, n73948, n73949, n73950,
         n73951, n73952, n73953, n73954, n73955, n73956, n73957, n73958,
         n73959, n73960, n73961, n73962, n73963, n73964, n73965, n73966,
         n73967, n73968, n73969, n73970, n73971, n73972, n73973, n73974,
         n73975, n73976, n73977, n73978, n73979, n73980, n73981, n73982,
         n73983, n73984, n73985, n73986, n73987, n73988, n73989, n73990,
         n73991, n73992, n73993, n73994, n73995, n73996, n73997, n73998,
         n73999, n74000, n74001, n74002, n74003, n74004, n74005, n74006,
         n74007, n74008, n74009, n74010, n74011, n74012, n74013, n74014,
         n74015, n74016, n74017, n74018, n74019, n74020, n74021, n74022,
         n74023, n74024, n74025, n74026, n74027, n74028, n74029, n74030,
         n74031, n74032, n74033, n74034, n74035, n74036, n74037, n74038,
         n74039, n74040, n74041, n74042, n74043, n74044, n74045, n74046,
         n74047, n74048, n74049, n74050, n74051, n74052, n74053, n74054,
         n74055, n74056, n74057, n74058, n74059, n74060, n74061, n74062,
         n74063, n74064, n74065, n74066, n74067, n74068, n74069, n74070,
         n74071, n74072, n74073, n74074, n74075, n74076, n74077, n74078,
         n74079, n74080, n74081, n74082, n74083, n74084, n74085, n74086,
         n74087, n74088, n74089, n74090, n74091, n74092, n74093, n74094,
         n74095, n74096, n74097, n74098, n74099, n74100, n74101, n74102,
         n74103, n74104, n74105, n74106, n74107, n74108, n74109, n74110,
         n74111, n74112, n74113, n74114, n74115, n74116, n74117, n74118,
         n74119, n74120, n74121, n74122, n74123, n74124, n74125, n74126,
         n74127, n74128, n74129, n74130, n74131, n74132, n74133, n74134,
         n74135, n74136, n74137, n74138, n74139, n74140, n74141, n74142,
         n74143, n74144, n74145, n74146, n74147, n74148, n74149, n74150,
         n74151, n74152, n74153, n74154, n74155, n74156, n74157, n74158,
         n74159, n74160, n74161, n74162, n74163, n74164, n74165, n74166,
         n74167, n74168, n74169, n74170, n74171, n74172, n74173, n74174,
         n74175, n74176, n74177, n74178, n74179, n74180, n74181, n74182,
         n74183, n74184, n74185, n74186, n74187, n74188, n74189, n74190,
         n74191, n74192, n74193, n74194, n74195, n74196, n74197, n74198,
         n74199, n74200, n74201, n74202, n74203, n74204, n74205, n74206,
         n74207, n74208, n74209, n74210, n74211, n74212, n74213, n74214,
         n74215, n74216, n74217, n74218, n74219, n74220, n74221, n74222,
         n74223, n74224, n74225, n74226, n74227, n74228, n74229, n74230,
         n74231, n74232, n74233, n74234, n74235, n74236, n74237, n74238,
         n74239, n74240, n74241, n74242, n74243, n74244, n74245, n74246,
         n74247, n74248, n74249, n74250, n74251, n74252, n74253, n74254,
         n74255, n74256, n74257, n74258, n74259, n74260, n74261, n74262,
         n74263, n74264, n74265, n74266, n74267, n74268, n74269, n74270,
         n74271, n74272, n74273, n74274, n74275, n74276, n74277, n74278,
         n74279, n74280, n74281, n74282, n74283, n74284, n74285, n74286,
         n74287, n74288, n74289, n74290, n74291, n74292, n74293, n74294,
         n74295, n74296, n74297, n74298, n74299, n74300, n74301, n74302,
         n74303, n74304, n74305, n74306, n74307, n74308, n74309, n74310,
         n74311, n74312, n74313, n74314, n74315, n74316, n74317, n74318,
         n74319, n74320, n74321, n74322, n74323, n74324, n74325, n74326,
         n74327, n74328, n74329, n74330, n74331, n74332, n74333, n74334,
         n74335, n74336, n74337, n74338, n74339, n74340, n74341, n74342,
         n74343, n74344, n74345, n74346, n74347, n74348, n74349, n74350,
         n74351, n74352, n74353, n74354, n74355, n74356, n74357, n74358,
         n74359, n74360, n74361, n74362, n74363, n74364, n74365, n74366,
         n74367, n74368, n74369, n74370, n74371, n74372, n74373, n74374,
         n74375, n74376, n74377, n74378, n74379, n74380, n74381, n74382,
         n74383, n74384, n74385, n74386, n74387, n74388, n74389, n74390,
         n74391, n74392, n74393, n74394, n74395, n74396, n74397, n74398,
         n74399, n74400, n74401, n74402, n74403, n74404, n74405, n74406,
         n74407, n74408, n74409, n74410, n74411, n74412, n74413, n74414,
         n74415, n74416, n74417, n74418, n74419, n74420, n74421, n74422,
         n74423, n74424, n74425, n74426, n74427, n74428, n74429, n74430,
         n74431, n74432, n74433, n74434, n74435, n74436, n74437, n74438,
         n74439, n74440, n74441, n74442, n74443, n74444, n74445, n74446,
         n74447, n74448, n74449, n74450, n74451, n74452, n74453, n74454,
         n74455, n74456, n74457, n74458, n74459, n74460, n74461, n74462,
         n74463, n74464, n74465, n74466, n74467, n74468, n74469, n74470,
         n74471, n74472, n74473, n74474, n74475, n74476, n74477, n74478,
         n74479, n74480, n74481, n74482, n74483, n74484, n74485, n74486,
         n74487, n74488, n74489, n74490, n74491, n74492, n74493, n74494,
         n74495, n74496, n74497, n74498, n74499, n74500, n74501, n74502,
         n74503, n74504, n74505, n74506, n74507, n74508, n74509, n74510,
         n74511, n74512, n74513, n74514, n74515, n74516, n74517, n74518,
         n74519, n74520, n74521, n74522, n74523, n74524, n74525, n74526,
         n74527, n74528, n74529, n74530, n74531, n74532, n74533, n74534,
         n74535, n74536, n74537, n74538, n74539, n74540, n74541, n74542,
         n74543, n74544, n74545, n74546, n74547, n74548, n74549, n74550,
         n74551, n74552, n74553, n74554, n74555, n74556, n74557, n74558,
         n74559, n74560, n74561, n74562, n74563, n74564, n74565, n74566,
         n74567, n74568, n74569, n74570, n74571, n74572, n74573, n74574,
         n74575, n74576, n74577, n74578, n74579, n74580, n74581, n74582,
         n74583, n74584, n74585, n74586, n74587, n74588, n74589, n74590,
         n74591, n74592, n74593, n74594, n74595, n74596, n74597, n74598,
         n74599, n74600, n74601, n74602, n74603, n74604, n74605, n74606,
         n74607, n74608, n74609, n74610, n74611, n74612, n74613, n74614,
         n74615, n74616, n74617, n74618, n74619, n74620, n74621, n74622,
         n74623, n74624, n74625, n74626, n74627, n74628, n74629, n74630,
         n74631, n74632, n74633, n74634, n74635, n74636, n74637, n74638,
         n74639, n74640, n74641, n74642, n74643, n74644, n74645, n74646,
         n74647, n74648, n74649, n74650, n74651, n74652, n74653, n74654,
         n74655, n74656, n74657, n74658, n74659, n74660, n74661, n74662,
         n74663, n74664, n74665, n74666, n74667, n74668, n74669, n74670,
         n74671, n74672, n74673, n74674, n74675, n74676, n74677, n74678,
         n74679, n74680, n74681, n74682, n74683, n74684, n74685, n74686,
         n74687, n74688, n74689, n74690, n74691, n74692, n74693, n74694,
         n74695, n74696, n74697, n74698, n74699, n74700, n74701, n74702,
         n74703, n74704, n74705, n74706, n74707, n74708, n74709, n74710,
         n74711, n74712, n74713, n74714, n74715, n74716, n74717, n74718,
         n74719, n74720, n74721, n74722, n74723, n74724, n74725, n74726,
         n74727, n74728, n74729, n74730, n74731, n74732, n74733, n74734,
         n74735, n74736, n74737, n74738, n74739, n74740, n74741, n74742,
         n74743, n74744, n74745, n74746, n74747, n74748, n74749, n74750,
         n74751, n74752, n74753, n74754, n74755, n74756, n74757, n74758,
         n74759, n74760, n74761, n74762, n74763, n74764, n74765, n74766,
         n74767, n74768, n74769, n74770, n74771, n74772, n74773, n74774,
         n74775, n74776, n74777, n74778, n74779, n74780, n74781, n74782,
         n74783, n74784, n74785, n74786, n74787, n74788, n74789, n74790,
         n74791, n74792, n74793, n74794, n74795, n74796, n74797, n74798,
         n74799, n74800, n74801, n74802, n74803, n74804, n74805, n74806,
         n74807, n74808, n74809, n74810, n74811, n74812, n74813, n74814,
         n74815, n74816, n74817, n74818, n74819, n74820, n74821, n74822,
         n74823, n74824, n74825, n74826, n74827, n74828, n74829, n74830,
         n74831, n74832, n74833, n74834, n74835, n74836, n74837, n74838,
         n74839, n74840, n74841, n74842, n74843, n74844, n74845, n74846,
         n74847, n74848, n74849, n74850, n74851, n74852, n74853, n74854,
         n74855, n74856, n74857, n74858, n74859, n74860, n74861, n74862,
         n74863, n74864, n74865, n74866, n74867, n74868, n74869, n74870,
         n74871, n74872, n74873, n74874, n74875, n74876, n74877, n74878,
         n74879, n74880, n74881, n74882, n74883, n74884, n74885, n74886,
         n74887, n74888, n74889, n74890, n74891, n74892, n74893, n74894,
         n74895, n74896, n74897, n74898, n74899, n74900, n74901, n74902,
         n74903, n74904, n74905, n74906, n74907, n74908, n74909, n74910,
         n74911, n74912, n74913, n74914, n74915, n74916, n74917, n74918,
         n74919, n74920, n74921, n74922, n74923, n74924, n74925, n74926,
         n74927, n74928, n74929, n74930, n74931, n74932, n74933, n74934,
         n74935, n74936, n74937, n74938, n74939, n74940, n74941, n74942,
         n74943, n74944, n74945, n74946, n74947, n74948, n74949, n74950,
         n74951, n74952, n74953, n74954, n74955, n74956, n74957, n74958,
         n74959, n74960, n74961, n74962, n74963, n74964, n74965, n74966,
         n74967, n74968, n74969, n74970, n74971, n74972, n74973, n74974,
         n74975, n74976, n74977, n74978, n74979, n74980, n74981, n74982,
         n74983, n74984, n74985, n74986, n74987, n74988, n74989, n74990,
         n74991, n74992, n74993, n74994, n74995, n74996, n74997, n74998,
         n74999, n75000, n75001, n75002, n75003, n75004, n75005, n75006,
         n75007, n75008, n75009, n75010, n75011, n75012, n75013, n75014,
         n75015, n75016, n75017, n75018, n75019, n75020, n75021, n75022,
         n75023, n75024, n75025, n75026, n75027, n75028, n75029, n75030,
         n75031, n75032, n75033, n75034, n75035, n75036, n75037, n75038,
         n75039, n75040, n75041, n75042, n75043, n75044, n75045, n75046,
         n75047, n75048, n75049, n75050, n75051, n75052, n75053, n75054,
         n75055, n75056, n75057, n75058, n75059, n75060, n75061, n75062,
         n75063, n75064, n75065, n75066, n75067, n75068, n75069, n75070,
         n75071, n75072, n75073, n75074, n75075, n75076, n75077, n75078,
         n75079, n75080, n75081, n75082, n75083, n75084, n75085, n75086,
         n75087, n75088, n75089, n75090, n75091, n75092, n75093, n75094,
         n75095, n75096, n75097, n75098, n75099, n75100, n75101, n75102,
         n75103, n75104, n75105, n75106, n75107, n75108, n75109, n75110,
         n75111, n75112, n75113, n75114, n75115, n75116, n75117, n75118,
         n75119, n75120, n75121, n75122, n75123, n75124, n75125, n75126,
         n75127, n75128, n75129, n75130, n75131, n75132, n75133, n75134,
         n75135, n75136, n75137, n75138, n75139, n75140, n75141, n75142,
         n75143, n75144, n75145, n75146, n75147, n75148, n75149, n75150,
         n75151, n75152, n75153, n75154, n75155, n75156, n75157, n75158,
         n75159, n75160, n75161, n75162, n75163, n75164, n75165, n75166,
         n75167, n75168, n75169, n75170, n75171, n75172, n75173, n75174,
         n75175, n75176, n75177, n75178, n75179, n75180, n75181, n75182,
         n75183, n75184, n75185, n75186, n75187, n75188, n75189, n75190,
         n75191, n75192, n75193, n75194, n75195, n75196, n75197, n75198,
         n75199, n75200, n75201, n75202, n75203, n75204, n75205, n75206,
         n75207, n75208, n75209, n75210, n75211, n75212, n75213, n75214,
         n75215, n75216, n75217, n75218, n75219, n75220, n75221, n75222,
         n75223, n75224, n75225, n75226, n75227, n75228, n75229, n75230,
         n75231, n75232, n75233, n75234, n75235, n75236, n75237, n75238,
         n75239, n75240, n75241, n75242, n75243, n75244, n75245, n75246,
         n75247, n75248, n75249, n75250, n75251, n75252, n75253, n75254,
         n75255, n75256, n75257, n75258, n75259, n75260, n75261, n75262,
         n75263, n75264, n75265, n75266, n75267, n75268, n75269, n75270,
         n75271, n75272, n75273, n75274, n75275, n75276, n75277, n75278,
         n75279, n75280, n75281, n75282, n75283, n75284, n75285, n75286,
         n75287, n75288, n75289, n75290, n75291, n75292, n75293, n75294,
         n75295, n75296, n75297, n75298, n75299, n75300, n75301, n75302,
         n75303, n75304, n75305, n75306, n75307, n75308, n75309, n75310,
         n75311, n75312, n75313, n75314, n75315, n75316, n75317, n75318,
         n75319, n75320, n75321, n75322, n75323, n75324, n75325, n75326,
         n75327, n75328, n75329, n75330, n75331, n75332, n75333, n75334,
         n75335, n75336, n75337, n75338, n75339, n75340, n75341, n75342,
         n75343, n75344, n75345, n75346, n75347, n75348, n75349, n75350,
         n75351, n75352, n75353, n75354, n75355, n75356, n75357, n75358,
         n75359, n75360, n75361, n75362, n75363, n75364, n75365, n75366,
         n75367, n75368, n75369, n75370, n75371, n75372, n75373, n75374,
         n75375, n75376, n75377, n75378, n75379, n75380, n75381, n75382,
         n75383, n75384, n75385, n75386, n75387, n75388, n75389, n75390,
         n75391, n75392, n75393, n75394, n75395, n75396, n75397, n75398,
         n75399, n75400, n75401, n75402, n75403, n75404, n75405, n75406,
         n75407, n75408, n75409, n75410, n75411, n75412, n75413, n75414,
         n75415, n75416, n75417, n75418, n75419, n75420, n75421, n75422,
         n75423, n75424, n75425, n75426, n75427, n75428, n75429, n75430,
         n75431, n75432, n75433, n75434, n75435, n75436, n75437, n75438,
         n75439, n75440, n75441, n75442, n75443, n75444, n75445, n75446,
         n75447, n75448, n75449, n75450, n75451, n75452, n75453, n75454,
         n75455, n75456, n75457, n75458, n75459, n75460, n75461, n75462,
         n75463, n75464, n75465, n75466, n75467, n75468, n75469, n75470,
         n75471, n75472, n75473, n75474, n75475, n75476, n75477, n75478,
         n75479, n75480, n75481, n75482, n75483, n75484, n75485, n75486,
         n75487, n75488, n75489, n75490, n75491, n75492, n75493, n75494,
         n75495, n75496, n75497, n75498, n75499, n75500, n75501, n75502,
         n75503, n75504, n75505, n75506, n75507, n75508, n75509, n75510,
         n75511, n75512, n75513, n75514, n75515, n75516, n75517, n75518,
         n75519, n75520, n75521, n75522, n75523, n75524, n75525, n75526,
         n75527, n75528, n75529, n75530, n75531, n75532, n75533, n75534,
         n75535, n75536, n75537, n75538, n75539, n75540, n75541, n75542,
         n75543, n75544, n75545, n75546, n75547, n75548, n75549, n75550,
         n75551, n75552, n75553, n75554, n75555, n75556, n75557, n75558,
         n75559, n75560, n75561, n75562, n75563, n75564, n75565, n75566,
         n75567, n75568, n75569, n75570, n75571, n75572, n75573, n75574,
         n75575, n75576, n75577, n75578, n75579, n75580, n75581, n75582,
         n75583, n75584, n75585, n75586, n75587, n75588, n75589, n75590,
         n75591, n75592, n75593, n75594, n75595, n75596, n75597, n75598,
         n75599, n75600, n75601, n75602, n75603, n75604, n75605, n75606,
         n75607, n75608, n75609, n75610, n75611, n75612, n75613, n75614,
         n75615, n75616, n75617, n75618, n75619, n75620, n75621, n75622,
         n75623, n75624, n75625, n75626, n75627, n75628, n75629, n75630,
         n75631, n75632, n75633, n75634, n75635, n75636, n75637, n75638,
         n75639, n75640, n75641, n75642, n75643, n75644, n75645, n75646,
         n75647, n75648, n75649, n75650, n75651, n75652, n75653, n75654,
         n75655, n75656, n75657, n75658, n75659, n75660, n75661, n75662,
         n75663, n75664, n75665, n75666, n75667, n75668, n75669, n75670,
         n75671, n75672, n75673, n75674, n75675, n75676, n75677, n75678,
         n75679, n75680, n75681, n75682, n75683, n75684, n75685, n75686,
         n75687, n75688, n75689, n75690, n75691, n75692, n75693, n75694,
         n75695, n75696, n75697, n75698, n75699, n75700, n75701, n75702,
         n75703, n75704, n75705, n75706, n75707, n75708, n75709, n75710,
         n75711, n75712, n75713, n75714, n75715, n75716, n75717, n75718,
         n75719, n75720, n75721, n75722, n75723, n75724, n75725, n75726,
         n75727, n75728, n75729, n75730, n75731, n75732, n75733, n75734,
         n75735, n75736, n75737, n75738, n75739, n75740, n75741, n75742,
         n75743, n75744, n75745, n75746, n75747, n75748, n75749, n75750,
         n75751, n75752, n75753, n75754, n75755, n75756, n75757, n75758,
         n75759, n75760, n75761, n75762, n75763, n75764, n75765, n75766,
         n75767, n75768, n75769, n75770, n75771, n75772, n75773, n75774,
         n75775, n75776, n75777, n75778, n75779, n75780, n75781, n75782,
         n75783, n75784, n75785, n75786, n75787, n75788, n75789, n75790,
         n75791, n75792, n75793, n75794, n75795, n75796, n75797, n75798,
         n75799, n75800, n75801, n75802, n75803, n75804, n75805, n75806,
         n75807, n75808, n75809, n75810, n75811, n75812, n75813, n75814,
         n75815, n75816, n75817, n75818, n75819, n75820, n75821, n75822,
         n75823, n75824, n75825, n75826, n75827, n75828, n75829, n75830,
         n75831, n75832, n75833, n75834, n75835, n75836, n75837, n75838,
         n75839, n75840, n75841, n75842, n75843, n75844, n75845, n75846,
         n75847, n75848, n75849, n75850, n75851, n75852, n75853, n75854,
         n75855, n75856, n75857, n75858, n75859, n75860, n75861, n75862,
         n75863, n75864, n75865, n75866, n75867, n75868, n75869, n75870,
         n75871, n75872, n75873, n75874, n75875, n75876, n75877, n75878,
         n75879, n75880, n75881, n75882, n75883, n75884, n75885, n75886,
         n75887, n75888, n75889, n75890, n75891, n75892, n75893, n75894,
         n75895, n75896, n75897, n75898, n75899, n75900, n75901, n75902,
         n75903, n75904, n75905, n75906, n75907, n75908, n75909, n75910,
         n75911, n75912, n75913, n75914, n75915, n75916, n75917, n75918,
         n75919, n75920, n75921, n75922, n75923, n75924, n75925, n75926,
         n75927, n75928, n75929, n75930, n75931, n75932, n75933, n75934,
         n75935, n75936, n75937, n75938, n75939, n75940, n75941, n75942,
         n75943, n75944, n75945, n75946, n75947, n75948, n75949, n75950,
         n75951, n75952, n75953, n75954, n75955, n75956, n75957, n75958,
         n75959, n75960, n75961, n75962, n75963, n75964, n75965, n75966,
         n75967, n75968, n75969, n75970, n75971, n75972, n75973, n75974,
         n75975, n75976, n75977, n75978, n75979, n75980, n75981, n75982,
         n75983, n75984, n75985, n75986, n75987, n75988, n75989, n75990,
         n75991, n75992, n75993, n75994, n75995, n75996, n75997, n75998,
         n75999, n76000, n76001, n76002, n76003, n76004, n76005, n76006,
         n76007, n76008, n76009, n76010, n76011, n76012, n76013, n76014,
         n76015, n76016, n76017, n76018, n76019, n76020, n76021, n76022,
         n76023, n76024, n76025, n76026, n76027, n76028, n76029, n76030,
         n76031, n76032, n76033, n76034, n76035, n76036, n76037, n76038,
         n76039, n76040, n76041, n76042, n76043, n76044, n76045, n76046,
         n76047, n76048, n76049, n76050, n76051, n76052, n76053, n76054,
         n76055, n76056, n76057, n76058, n76059, n76060, n76061, n76062,
         n76063, n76064, n76065, n76066, n76067, n76068, n76069, n76070,
         n76071, n76072, n76073, n76074, n76075, n76076, n76077, n76078,
         n76079, n76080, n76081, n76082, n76083, n76084, n76085, n76086,
         n76087, n76088, n76089, n76090, n76091, n76092, n76093, n76094,
         n76095, n76096, n76097, n76098, n76099, n76100, n76101, n76102,
         n76103, n76104, n76105, n76106, n76107, n76108, n76109, n76110,
         n76111, n76112, n76113, n76114, n76115, n76116, n76117, n76118,
         n76119, n76120, n76121, n76122, n76123, n76124, n76125, n76126,
         n76127, n76128, n76129, n76130, n76131, n76132, n76133, n76134,
         n76135, n76136, n76137, n76138, n76139, n76140, n76141, n76142,
         n76143, n76144, n76145, n76146, n76147, n76148, n76149, n76150,
         n76151, n76152, n76153, n76154, n76155, n76156, n76157, n76158,
         n76159, n76160, n76161, n76162, n76163, n76164, n76165, n76166,
         n76167, n76168, n76169, n76170, n76171, n76172, n76173, n76174,
         n76175, n76176, n76177, n76178, n76179, n76180, n76181, n76182,
         n76183, n76184, n76185, n76186, n76187, n76188, n76189, n76190,
         n76191, n76192, n76193, n76194, n76195, n76196, n76197, n76198,
         n76199, n76200, n76201, n76202, n76203, n76204, n76205, n76206,
         n76207, n76208, n76209, n76210, n76211, n76212, n76213, n76214,
         n76215, n76216, n76217, n76218, n76219, n76220, n76221, n76222,
         n76223, n76224, n76225, n76226, n76227, n76228, n76229, n76230,
         n76231, n76232, n76233, n76234, n76235, n76236, n76237, n76238,
         n76239, n76240, n76241, n76242, n76243, n76244, n76245, n76246,
         n76247, n76248, n76249, n76250, n76251, n76252, n76253, n76254,
         n76255, n76256, n76257, n76258, n76259, n76260, n76261, n76262,
         n76263, n76264, n76265, n76266, n76267, n76268, n76269, n76270,
         n76271, n76272, n76273, n76274, n76275, n76276, n76277, n76278,
         n76279, n76280, n76281, n76282, n76283, n76284, n76285, n76286,
         n76287, n76288, n76289, n76290, n76291, n76292, n76293, n76294,
         n76295, n76296, n76297, n76298, n76299, n76300, n76301, n76302,
         n76303, n76304, n76305, n76306, n76307, n76308, n76309, n76310,
         n76311, n76312, n76313, n76314, n76315, n76316, n76317, n76318,
         n76319, n76320, n76321, n76322, n76323, n76324, n76325, n76326,
         n76327, n76328, n76329, n76330, n76331, n76332, n76333, n76334,
         n76335, n76336, n76337, n76338, n76339, n76340, n76341, n76342,
         n76343, n76344, n76345, n76346, n76347, n76348, n76349, n76350,
         n76351, n76352, n76353, n76354, n76355, n76356, n76357, n76358,
         n76359, n76360, n76361, n76362, n76363, n76364, n76365, n76366,
         n76367, n76368, n76369, n76370, n76371, n76372, n76373, n76374,
         n76375, n76376, n76377, n76378, n76379, n76380, n76381, n76382,
         n76383, n76384, n76385, n76386, n76387, n76388, n76389, n76390,
         n76391, n76392, n76393, n76394, n76395, n76396, n76397, n76398,
         n76399, n76400, n76401, n76402, n76403, n76404, n76405, n76406,
         n76407, n76408, n76409, n76410, n76411, n76412, n76413, n76414,
         n76415, n76416, n76417, n76418, n76419, n76420, n76421, n76422,
         n76423, n76424, n76425, n76426, n76427, n76428, n76429, n76430,
         n76431, n76432, n76433, n76434, n76435, n76436, n76437, n76438,
         n76439, n76440, n76441, n76442, n76443, n76444, n76445, n76446,
         n76447, n76448, n76449, n76450, n76451, n76452, n76453, n76454,
         n76455, n76456, n76457, n76458, n76459, n76460, n76461, n76462,
         n76463, n76464, n76465, n76466, n76467, n76468, n76469, n76470,
         n76471, n76472, n76473, n76474, n76475, n76476, n76477, n76478,
         n76479, n76480, n76481, n76482, n76483, n76484, n76485, n76486,
         n76487, n76488, n76489, n76490, n76491, n76492, n76493, n76494,
         n76495, n76496, n76497, n76498, n76499, n76500, n76501, n76502,
         n76503, n76504, n76505, n76506, n76507, n76508, n76509, n76510,
         n76511, n76512, n76513, n76514, n76515, n76516, n76517, n76518,
         n76519, n76520, n76521, n76522, n76523, n76524, n76525, n76526,
         n76527, n76528, n76529, n76530, n76531, n76532, n76533, n76534,
         n76535, n76536, n76537, n76538, n76539, n76540, n76541, n76542,
         n76543, n76544, n76545, n76546, n76547, n76548, n76549, n76550,
         n76551, n76552, n76553, n76554, n76555, n76556, n76557, n76558,
         n76559, n76560, n76561, n76562, n76563, n76564, n76565, n76566,
         n76567, n76568, n76569, n76570, n76571, n76572, n76573, n76574,
         n76575, n76576, n76577, n76578, n76579, n76580, n76581, n76582,
         n76583, n76584, n76585, n76586, n76587, n76588, n76589, n76590,
         n76591, n76592, n76593, n76594, n76595, n76596, n76597, n76598,
         n76599, n76600, n76601, n76602, n76603, n76604, n76605, n76606,
         n76607, n76608, n76609, n76610, n76611, n76612, n76613, n76614,
         n76615, n76616, n76617, n76618, n76619, n76620, n76621, n76622,
         n76623, n76624, n76625, n76626, n76627, n76628, n76629, n76630,
         n76631, n76632, n76633, n76634, n76635, n76636, n76637, n76638,
         n76639, n76640, n76641, n76642, n76643, n76644, n76645, n76646,
         n76647, n76648, n76649, n76650, n76651, n76652, n76653, n76654,
         n76655, n76656, n76657, n76658, n76659, n76660, n76661, n76662,
         n76663, n76664, n76665, n76666, n76667, n76668, n76669, n76670,
         n76671, n76672, n76673, n76674, n76675, n76676, n76677, n76678,
         n76679, n76680, n76681, n76682, n76683, n76684, n76685, n76686,
         n76687, n76688, n76689, n76690, n76691, n76692, n76693, n76694,
         n76695, n76696, n76697, n76698, n76699, n76700, n76701, n76702,
         n76703, n76704, n76705, n76706, n76707, n76708, n76709, n76710,
         n76711, n76712, n76713, n76714, n76715, n76716, n76717, n76718,
         n76719, n76720, n76721, n76722, n76723, n76724, n76725, n76726,
         n76727, n76728, n76729, n76730, n76731, n76732, n76733, n76734,
         n76735, n76736, n76737, n76738, n76739, n76740, n76741, n76742,
         n76743, n76744, n76745, n76746, n76747, n76748, n76749, n76750,
         n76751, n76752, n76753, n76754, n76755, n76756, n76757, n76758,
         n76759, n76760, n76761, n76762, n76763, n76764, n76765, n76766,
         n76767, n76768, n76769, n76770, n76771, n76772, n76773, n76774,
         n76775, n76776, n76777, n76778, n76779, n76780, n76781, n76782,
         n76783, n76784, n76785, n76786, n76787, n76788, n76789, n76790,
         n76791, n76792, n76793, n76794, n76795, n76796, n76797, n76798,
         n76799, n76800, n76801, n76802, n76803, n76804, n76805, n76806,
         n76807, n76808, n76809, n76810, n76811, n76812, n76813, n76814,
         n76815, n76816, n76817, n76818, n76819, n76820, n76821, n76822,
         n76823, n76824, n76825, n76826, n76827, n76828, n76829, n76830,
         n76831, n76832, n76833, n76834, n76835, n76836, n76837, n76838,
         n76839, n76840, n76841, n76842, n76843, n76844, n76845, n76846,
         n76847, n76848, n76849, n76850, n76851, n76852, n76853, n76854,
         n76855, n76856, n76857, n76858, n76859, n76860, n76861, n76862,
         n76863, n76864, n76865, n76866, n76867, n76868, n76869, n76870,
         n76871, n76872, n76873, n76874, n76875, n76876, n76877, n76878,
         n76879, n76880, n76881, n76882, n76883, n76884, n76885, n76886,
         n76887, n76888, n76889, n76890, n76891, n76892, n76893, n76894,
         n76895, n76896, n76897, n76898, n76899, n76900, n76901, n76902,
         n76903, n76904, n76905, n76906, n76907, n76908, n76909, n76910,
         n76911, n76912, n76913, n76914, n76915, n76916, n76917, n76918,
         n76919, n76920, n76921, n76922, n76923, n76924, n76925, n76926,
         n76927, n76928, n76929, n76930, n76931, n76932, n76933, n76934,
         n76935, n76936, n76937, n76938, n76939, n76940, n76941, n76942,
         n76943, n76944, n76945, n76946, n76947, n76948, n76949, n76950,
         n76951, n76952, n76953, n76954, n76955, n76956, n76957, n76958,
         n76959, n76960, n76961, n76962, n76963, n76964, n76965, n76966,
         n76967, n76968, n76969, n76970, n76971, n76972, n76973, n76974,
         n76975, n76976, n76977, n76978, n76979, n76980, n76981, n76982,
         n76983, n76984, n76985, n76986, n76987, n76988, n76989, n76990,
         n76991, n76992, n76993, n76994, n76995, n76996, n76997, n76998,
         n76999, n77000, n77001, n77002, n77003, n77004, n77005, n77006,
         n77007, n77008, n77009, n77010, n77011, n77012, n77013, n77014,
         n77015, n77016, n77017, n77018, n77019, n77020, n77021, n77022,
         n77023, n77024, n77025, n77026, n77027, n77028, n77029, n77030,
         n77031, n77032, n77033, n77034, n77035, n77036, n77037, n77038,
         n77039, n77040, n77041, n77042, n77043, n77044, n77045, n77046,
         n77047, n77048, n77049, n77050, n77051, n77052, n77053, n77054,
         n77055, n77056, n77057, n77058, n77059, n77060, n77061, n77062,
         n77063, n77064, n77065, n77066, n77067, n77068, n77069, n77070,
         n77071, n77072, n77073, n77074, n77075, n77076, n77077, n77078,
         n77079, n77080, n77081, n77082, n77083, n77084, n77085, n77086,
         n77087, n77088, n77089, n77090, n77091, n77092, n77093, n77094,
         n77095, n77096, n77097, n77098, n77099, n77100, n77101, n77102,
         n77103, n77104, n77105, n77106, n77107, n77108, n77109, n77110,
         n77111, n77112, n77113, n77114, n77115, n77116, n77117, n77118,
         n77119, n77120, n77121, n77122, n77123, n77124, n77125, n77126,
         n77127, n77128, n77129, n77130, n77131, n77132, n77133, n77134,
         n77135, n77136, n77137, n77138, n77139, n77140, n77141, n77142,
         n77143, n77144, n77145, n77146, n77147, n77148, n77149, n77150,
         n77151, n77152, n77153, n77154, n77155, n77156, n77157, n77158,
         n77159, n77160, n77161, n77162, n77163, n77164, n77165, n77166,
         n77167, n77168, n77169, n77170, n77171, n77172, n77173, n77174,
         n77175, n77176, n77177, n77178, n77179, n77180, n77181, n77182,
         n77183, n77184, n77185, n77186, n77187, n77188, n77189, n77190,
         n77191, n77192, n77193, n77194, n77195, n77196, n77197, n77198,
         n77199, n77200, n77201, n77202, n77203, n77204, n77205, n77206,
         n77207, n77208, n77209, n77210, n77211, n77212, n77213, n77214,
         n77215, n77216, n77217, n77218, n77219, n77220, n77221, n77222,
         n77223, n77224, n77225, n77226, n77227, n77228, n77229, n77230,
         n77231, n77232, n77233, n77234, n77235, n77236, n77237, n77238,
         n77239, n77240, n77241, n77242, n77243, n77244, n77245, n77246,
         n77247, n77248, n77249, n77250, n77251, n77252, n77253, n77254,
         n77255, n77256, n77257, n77258, n77259, n77260, n77261, n77262,
         n77263, n77264, n77265, n77266, n77267, n77268, n77269, n77270,
         n77271, n77272, n77273, n77274, n77275, n77276, n77277, n77278,
         n77279, n77280, n77281, n77282, n77283, n77284, n77285, n77286,
         n77287, n77288, n77289, n77290, n77291, n77292, n77293, n77294,
         n77295, n77296, n77297, n77298, n77299, n77300, n77301, n77302,
         n77303, n77304, n77305, n77306, n77307, n77308, n77309, n77310,
         n77311, n77312, n77313, n77314, n77315, n77316, n77317, n77318,
         n77319, n77320, n77321, n77322, n77323, n77324, n77325, n77326,
         n77327, n77328, n77329, n77330, n77331, n77332, n77333, n77334,
         n77335, n77336, n77337, n77338, n77339, n77340, n77341, n77342,
         n77343, n77344, n77345, n77346, n77347, n77348, n77349, n77350,
         n77351, n77352, n77353, n77354, n77355, n77356, n77357, n77358,
         n77359, n77360, n77361, n77362, n77363, n77364, n77365, n77366,
         n77367, n77368, n77369, n77370, n77371, n77372, n77373, n77374,
         n77375, n77376, n77377, n77378, n77379, n77380, n77381, n77382,
         n77383, n77384, n77385, n77386, n77387, n77388, n77389, n77390,
         n77391, n77392, n77393, n77394, n77395, n77396, n77397, n77398,
         n77399, n77400, n77401, n77402, n77403, n77404, n77405, n77406,
         n77407, n77408, n77409, n77410, n77411, n77412, n77413, n77414,
         n77415, n77416, n77417, n77418, n77419, n77420, n77421, n77422,
         n77423, n77424, n77425, n77426, n77427, n77428, n77429, n77430,
         n77431, n77432, n77433, n77434, n77435, n77436, n77437, n77438,
         n77439, n77440, n77441, n77442, n77443, n77444, n77445, n77446,
         n77447, n77448, n77449, n77450, n77451, n77452, n77453, n77454,
         n77455, n77456, n77457, n77458, n77459, n77460, n77461, n77462,
         n77463, n77464, n77465, n77466, n77467, n77468, n77469, n77470,
         n77471, n77472, n77473, n77474, n77475, n77476, n77477, n77478,
         n77479, n77480, n77481, n77482, n77483, n77484, n77485, n77486,
         n77487, n77488, n77489, n77490, n77491, n77492, n77493, n77494,
         n77495, n77496, n77497, n77498, n77499, n77500, n77501, n77502,
         n77503, n77504, n77505, n77506, n77507, n77508, n77509, n77510,
         n77511, n77512, n77513, n77514, n77515, n77516, n77517, n77518,
         n77519, n77520, n77521, n77522, n77523, n77524, n77525, n77526,
         n77527, n77528, n77529, n77530, n77531, n77532, n77533, n77534,
         n77535, n77536, n77537, n77538, n77539, n77540, n77541, n77542,
         n77543, n77544, n77545, n77546, n77547, n77548, n77549, n77550,
         n77551, n77552, n77553, n77554, n77555, n77556, n77557, n77558,
         n77559, n77560, n77561, n77562, n77563, n77564, n77565, n77566,
         n77567, n77568, n77569, n77570, n77571, n77572, n77573, n77574,
         n77575, n77576, n77577, n77578, n77579, n77581, n77582, n77583,
         n77584, n77585, n77586, n77587, n77588, n77589, n77590, n77591,
         n77592, n77593, n77594, n77595, n77596, n77597, n77598, n77599,
         n77600, n77601, n77602, n77603, n77604, n77605, n77606, n77607,
         n77608, n77609, n77610, n77611, n77612, n77613, n77614, n77615,
         n77616, n77617, n77618, n77619, n77620, n77621, n77622, n77623,
         n77624, n77625, n77626, n77627, n77628, n77629, n77630, n77631,
         n77632, n77633, n77634, n77635, n77636, n77637, n77638, n77639,
         n77640, n77641, n77642, n77643, n77644, n77645, n77646, n77647,
         n77648, n77649, n77650, n77651, n77652, n77653, n77654, n77655,
         n77656, n77657, n77658, n77659, n77660, n77661, n77662, n77663,
         n77664, n77665, n77666, n77667, n77668, n77669, n77670, n77671,
         n77672, n77673, n77674, n77675, n77676, n77677, n77678, n77679,
         n77680, n77681, n77682, n77683, n77684, n77685, n77686, n77687,
         n77688, n77689, n77690, n77691, n77692, n77693, n77694, n77695,
         n77696, n77697, n77698, n77699, n77700, n77701, n77702, n77703,
         n77704, n77705, n77706, n77707, n77708, n77709, n77710, n77711,
         n77712, n77713, n77714, n77715, n77716, n77717, n77718, n77719,
         n77720, n77721, n77722, n77723, n77724, n77725, n77726, n77727,
         n77728, n77729, n77730, n77731, n77732, n77733, n77734, n77735,
         n77736, n77737, n77738, n77739, n77740, n77741, n77742, n77743,
         n77744, n77745, n77746, n77747, n77748, n77749, n77750, n77751,
         n77752, n77753, n77754, n77755, n77756, n77757, n77758, n77759,
         n77760, n77761, n77762, n77763, n77764, n77765, n77766, n77767,
         n77768, n77769, n77770, n77771, n77772, n77773, n77774, n77775,
         n77776, n77777, n77778, n77779, n77780, n77781, n77782, n77783,
         n77784, n77785, n77786, n77787, n77788, n77789, n77790, n77791,
         n77792, n77793, n77794, n77795, n77796, n77797, n77798, n77799,
         n77800, n77801, n77802, n77803, n77804, n77805, n77806, n77807,
         n77808, n77809, n77810, n77811, n77812, n77813, n77814, n77815,
         n77816, n77817, n77818, n77819, n77820, n77821, n77822, n77823,
         n77824, n77825, n77826, n77827, n77828, n77829, n77830, n77831,
         n77832, n77833, n77834, n77835, n77836, n77837, n77838, n77839,
         n77840, n77841, n77842, n77843, n77844, n77845, n77846, n77847,
         n77848, n77849, n77850, n77851, n77852, n77853, n77854, n77855,
         n77856, n77857, n77858, n77859, n77860, n77861, n77862, n77863,
         n77864, n77865, n77866, n77867, n77868, n77869, n77870, n77871,
         n77872, n77873, n77874, n77875, n77876, n77877, n77878, n77879,
         n77880, n77881, n77882, n77883, n77884, n77885, n77886, n77887,
         n77888, n77889, n77890, n77891, n77892, n77893, n77894, n77895,
         n77896, n77897, n77898, n77899, n77900, n77901, n77902, n77903,
         n77904, n77905, n77906, n77907, n77908, n77909, n77910, n77911,
         n77912, n77913, n77914, n77915, n77916, n77917, n77918, n77919,
         n77920, n77921, n77922, n77923, n77924, n77925, n77926, n77927,
         n77928, n77929, n77930, n77931, n77932, n77933, n77934, n77935,
         n77936, n77937, n77938, n77939, n77940, n77941, n77942, n77943,
         n77944, n77945, n77946, n77947, n77948, n77949, n77950, n77951,
         n77952, n77953, n77954, n77955, n77956, n77957, n77958, n77959,
         n77960, n77961, n77962, n77963, n77964, n77965, n77966, n77967,
         n77968, n77969, n77970, n77971, n77972, n77973, n77974, n77975,
         n77976, n77977, n77978, n77979, n77980, n77981, n77982, n77983,
         n77984, n77985, n77986, n77987, n77988, n77989, n77990, n77991,
         n77992, n77993, n77994, n77995, n77996, n77997, n77998, n77999,
         n78000, n78001, n78002, n78003, n78004, n78005, n78006, n78007,
         n78008, n78009, n78010, n78011, n78012, n78013, n78014, n78015,
         n78016, n78017, n78018, n78019, n78020, n78021, n78022, n78023,
         n78024, n78025, n78026, n78027, n78028, n78029, n78030, n78031,
         n78032, n78033, n78034, n78035, n78036, n78037, n78038, n78039,
         n78040, n78041, n78042, n78043, n78044, n78045, n78046, n78047,
         n78048, n78049, n78050, n78051, n78052, n78053, n78054, n78055,
         n78056, n78057, n78058, n78059, n78060, n78061, n78062, n78063,
         n78064, n78065, n78066, n78067, n78068, n78069, n78070, n78071,
         n78072, n78073, n78074, n78075, n78076, n78077, n78078, n78079,
         n78080, n78081, n78082, n78083, n78084, n78085, n78086, n78087,
         n78088, n78089, n78090, n78091, n78092, n78093, n78094, n78095,
         n78096, n78097, n78098, n78099, n78100, n78101, n78102, n78103,
         n78104, n78105, n78106, n78107, n78108, n78109, n78110, n78111,
         n78112, n78113, n78114, n78115, n78116, n78117, n78118, n78119,
         n78120, n78121, n78122, n78123, n78124, n78125, n78126, n78127,
         n78128, n78129, n78130, n78131, n78132, n78133, n78134, n78135,
         n78136, n78137, n78138, n78139, n78140, n78141, n78142, n78143,
         n78144, n78145, n78146, n78147, n78148, n78149, n78150, n78151,
         n78152, n78153, n78154, n78155, n78156, n78157, n78158, n78159,
         n78160, n78161, n78162, n78163, n78164, n78165, n78166, n78167,
         n78168, n78169, n78170, n78171, n78172, n78173, n78174, n78175,
         n78176, n78177, n78181, n78182, n78183, n78184, n78185, n78187,
         n78188, n78189, n78190, n78191, n78192, n78193, n78194, n78195,
         n78196, n78197, n78198, n78199, n78200, n78201, n78202, n78203,
         n78204, n78205, n78206, n78207, n78208, n78209, n78210, n78211,
         n78212, n78213, n78214, n78215, n78216, n78217, n78218, n78219,
         n78220, n78221, n78222, n78223, n78224, n78225, n78226, n78227,
         n78228, n78229, n78230, n78231, n78232, n78233, n78234, n78235,
         n78236, n78237, n78238, n78239, n78240, n78241, n78242, n78243,
         n78244, n78245, n78246, n78247, n78248, n78249, n78250, n78251,
         n78252, n78253, n78254, n78255, n78256, n78257, n78258, n78259,
         n78260, n78261, n78262, n78263, n78264, n78265, n78326, n78327,
         n78328, n78329, n78330, n78331, n78332, n78333, n78334, n78335,
         n78336, n78337, n78338, n78339, n78340, n78341, n78342, n78343,
         n78344, n78345, n78346, n78347, n78348, n78349, n78350, n78351,
         n78352, n78353, n78354, n78355, n78356, n78357, n78358, n78359,
         n78360, n78361, n78362, n78363, n78364, n78365, n78366, n78367,
         n78368, n78369, n78370, n78371, n78372, n78373, n78374, n78375,
         n78376, n78377, n78378, n78379, n78380, n78381, n78382, n78383,
         n78384, n78385, n78386, n78387, n78388, n78389, n78390, n78391,
         n78392, n78393, n78394, n78395, n78396, n78397, n78398, n78399,
         n78400, n78401, n78402, n78403, n78404, n78405, n78406, n78407,
         n78408, n78409, n78410, n78411, n78412, n78413, n78414, n78415,
         n78416, n78417, n78418, n78419, n78420, n78421, n78422, n78423,
         n78424, n78425, n78426, n78427, n78428, n78429, n78430, n78431,
         n78432, n78433, n78434, n78435, n78436, n78437, n78438, n78439,
         n78440, n78441, n78442, n78443, n78444, n78445, n78446, n78447,
         n78448, n78449, n78450;
  wire   [31:2] icbiu_adr_ic_word;
  wire   [31:2] sbbiu_adr_sb;
  wire   [31:13] icqmem_adr_qmem;
  wire   [28:16] ex_insn;
  wire   [28:16] wb_insn;
  wire   [19:0] or1200_ic_top_tag;
  wire   [31:0] or1200_ic_top_from_icram;
  wire   [11:4] or1200_ic_top_ictag_addr;
  wire   [13:1] or1200_cpu_to_sr;
  wire   [15:0] or1200_cpu_esr;
  wire   [31:17] or1200_cpu_spr_dat_ppc;
  wire   [31:1] or1200_cpu_spr_dat_rf;
  wire   [31:0] or1200_cpu_rf_datab;
  wire   [4:0] or1200_cpu_rf_addrb;
  wire   [3:0] or1200_dc_top_dcram_we;
  wire   [31:0] or1200_dc_top_to_dcram;
  wire   [11:4] or1200_dc_top_dctag_addr;
  wire   [7:2] or1200_cpu_or1200_genpc_pcreg_default;
  wire   [28:16] or1200_cpu_or1200_if_insn_saved;
  wire   [6:0] or1200_cpu_or1200_fpu_fpu_conv_shr;
  wire   [31:0] or1200_cpu_or1200_fpu_result_arith;
  wire   [31:0] or1200_cpu_or1200_fpu_result_conv;
  wire   [30:24] or1200_cpu_or1200_fpu_fpu_arith_s_output_o;
  wire   [31:0] or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output;
  wire   [26:0] or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr;
  wire   [26:0] or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt;
  wire   [23:0] or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor;
  wire   [49:42] or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd;
  wire   [9:0] or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp;
  wire   [31:0] or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output;
  wire   [47:0] or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48;
  wire   [22:0] or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24;
  wire   [9:0] or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10;
  wire   [31:0] or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o;
  wire   [26:1] or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o;
  wire   [7:0] or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o;
  wire   [26:0] or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o;
  wire   [26:0] or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o;
  wire   [47:0] or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f;
  wire   [7:0] or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r;
  wire   [2:0] or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1;
  wire   [1:0] or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3;
  wire   [1:0] or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1;
  wire   [7:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o;
  wire   [4:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1;
  wire   [7:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1;
  wire   [7:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in;
  wire   [7:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in;
  wire   [9:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o;
  wire   [26:1] or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd;
  wire   [22:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2;
  wire   [8:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1;
  wire   [9:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i;
  wire   [31:0] or1200_cpu_or1200_rf_rf_dataw;
  wire   [4:0] or1200_cpu_or1200_rf_rf_addrw;
  wire   [4:0] or1200_cpu_or1200_rf_rf_addra;
  wire   [63:0] or1200_cpu_or1200_mult_mac_mul_prod;
  wire   [2:1] or1200_cpu_or1200_except_delayed_tee;
  wire   [2:1] or1200_cpu_or1200_except_delayed_iee;
  wire   [23:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i;
  wire   [23:0] or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i;

  OR2x2_ASAP7_75t_SL or1200_dc_top_C234 ( .A(or1200_dc_top_dcfsm_tag_we), .B(
        n78176), .Y(or1200_dc_top_dctag_we) );
  OR2x2_ASAP7_75t_SL or1200_dc_top_C238 ( .A(n78176), .B(dc_en), .Y(
        or1200_dc_top_dctag_en) );
  OR2x2_ASAP7_75t_SL or1200_ic_top_C174 ( .A(or1200_ic_top_icram_we_3_), .B(
        n78175), .Y(or1200_ic_top_ictag_we) );
  OR2x2_ASAP7_75t_SL or1200_ic_top_C178 ( .A(n78175), .B(ic_en), .Y(
        or1200_ic_top_ictag_en) );
  INVx1_ASAP7_75t_SL or1200_ic_top_I_1 ( .A(n78175), .Y(or1200_ic_top_ictag_v)
         );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dbg_ack_reg ( .D(n78439), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(or1200_du_dbg_ack) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dbg_ack_o_reg ( .D(n4183), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(dbg_ack_o) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_bit_eph_select_reg ( 
        .D(n53192), .CLK(clk_i), .RESET(rst_i), .SET(n53192), .QN(n3351) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_reg_4_ ( 
        .D(n27979), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_reg_5_ ( 
        .D(n27978), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_reg_6_ ( 
        .D(n27977), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_reg_7_ ( 
        .D(n12855), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_1_ ( 
        .D(n3341), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_2_ ( 
        .D(n3340), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_1_ ( 
        .D(n3339), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_2_ ( 
        .D(n3338), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_0_), .CLK(
        clk_i), .QN(n3337) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_1_ ( 
        .D(n12864), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_2_ ( 
        .D(n12827), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_3_ ( 
        .D(n21879), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_4_ ( 
        .D(n12863), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_5_ ( 
        .D(n12861), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_6_), .CLK(
        clk_i), .QN(n3331) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_7_ ( 
        .D(n53191), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_8_ ( 
        .D(n53190), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_9_ ( 
        .D(n53189), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_10_ ( 
        .D(n51955), .CLK(clk_i), .QN(n3327) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_11_ ( 
        .D(n78213), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_12_ ( 
        .D(n78214), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_13_ ( 
        .D(n78215), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_14_ ( 
        .D(n78216), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_15_ ( 
        .D(n78212), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_16_ ( 
        .D(n51956), .CLK(clk_i), .QN(n3321) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_17_ ( 
        .D(n78211), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_18_ ( 
        .D(n78210), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_19_ ( 
        .D(n78220), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_20_ ( 
        .D(n78221), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_21_ ( 
        .D(n78219), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_22_ ( 
        .D(n78222), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_23_ ( 
        .D(n78217), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_24_ ( 
        .D(n51957), .CLK(clk_i), .QN(n3313) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_25_ ( 
        .D(n78218), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_26_ ( 
        .D(n53176), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_fract_o_reg_27_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_27_), .CLK(
        clk_i), .QN(n3310) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_27_ ( 
        .D(n5349), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_27_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_26_ ( 
        .D(n3308), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_26_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_25_ ( 
        .D(n3307), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_25_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_24_ ( 
        .D(n3306), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_24_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_23_ ( 
        .D(n3305), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_23_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_22_ ( 
        .D(n3304), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_22_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_21_ ( 
        .D(n3303), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_21_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_20_ ( 
        .D(n3302), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_20_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_19_ ( 
        .D(n3301), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_19_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_18_ ( 
        .D(n3300), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_18_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_17_ ( 
        .D(n3299), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_17_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_16_ ( 
        .D(n3298), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_16_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_15_ ( 
        .D(n3297), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_15_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_14_ ( 
        .D(n3296), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_14_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_13_ ( 
        .D(n3295), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_13_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_12_ ( 
        .D(n3294), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_12_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_11_ ( 
        .D(n3293), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_11_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_10_ ( 
        .D(n3292), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_10_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_9_ ( 
        .D(n3291), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_9_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_8_ ( 
        .D(n3290), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_8_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_7_ ( 
        .D(n3289), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_7_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_6_ ( 
        .D(n3288), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_6_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_5_ ( 
        .D(n3287), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_5_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_4_ ( 
        .D(n3286), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_4_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_3_ ( 
        .D(n3285), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_3_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_2_ ( 
        .D(n3284), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_2_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_1_ ( 
        .D(n3283), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_1_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_reg_0_ ( 
        .D(n3282), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_0_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1_reg_0_ ( 
        .D(n3281), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1_reg_1_ ( 
        .D(n3280), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1_reg_2_ ( 
        .D(n3279), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1_reg_3_ ( 
        .D(n3278), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1_reg_4_ ( 
        .D(n3277), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1_reg_5_ ( 
        .D(n3276), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1_reg_6_ ( 
        .D(n3275), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1_reg_7_ ( 
        .D(n3274), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_0_ ( 
        .D(n12876), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_1_ ( 
        .D(n12875), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_2_ ( 
        .D(n3271), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_3_ ( 
        .D(n12873), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_4_ ( 
        .D(n12871), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_5_ ( 
        .D(n52545), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_6_ ( 
        .D(n52546), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_7_ ( 
        .D(n3266), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_8_ ( 
        .D(n3265), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_exp_10_o_reg_9_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_s_exp_10_o_9_), 
        .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_0_ ( 
        .D(n12874), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_1_ ( 
        .D(n3262), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_2_ ( 
        .D(n27047), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_3_ ( 
        .D(n3260), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_4_ ( 
        .D(n3259), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_5_ ( 
        .D(n3258), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_6_ ( 
        .D(n3257), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_7_ ( 
        .D(n3256), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_8_ ( 
        .D(n51958), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o_reg_9_ ( 
        .D(n3254), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in_reg_0_ ( 
        .D(n52547), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in_reg_1_ ( 
        .D(n78376), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in_reg_2_ ( 
        .D(n78379), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in_reg_3_ ( 
        .D(n78370), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in_reg_4_ ( 
        .D(n78381), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in_reg_5_ ( 
        .D(n78361), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in_reg_6_ ( 
        .D(n78363), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in_reg_7_ ( 
        .D(n78383), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in_reg_0_ ( 
        .D(n52549), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in_reg_1_ ( 
        .D(n78375), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in_reg_2_ ( 
        .D(n78378), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in_reg_3_ ( 
        .D(n78371), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in_reg_4_ ( 
        .D(n78380), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in_reg_6_ ( 
        .D(n78362), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in_reg_7_ ( 
        .D(n78382), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_0_ ( 
        .D(n27037), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_1_ ( 
        .D(n27038), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_2_ ( 
        .D(n27039), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_3_ ( 
        .D(n27040), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_4_ ( 
        .D(n27041), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_5_ ( 
        .D(n27042), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_6_ ( 
        .D(n27043), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_7_ ( 
        .D(n27044), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_8_ ( 
        .D(n27045), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_exp_10_o_reg_9_ ( 
        .D(n27046), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[0]), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[1]), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[2]), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[3]), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[4]), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[5]), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[6]), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_7_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[7]), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_8_ ( 
        .D(n3217), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_9_ ( 
        .D(n3216), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_10_ ( 
        .D(n3215), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_11_ ( 
        .D(n3214), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_12_ ( 
        .D(n3213), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_13_ ( 
        .D(n3212), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_14_ ( 
        .D(n3211), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_15_ ( 
        .D(n3210), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_16_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[16]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_17_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[17]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[18]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_19_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[19]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_20_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[20]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_21_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[21]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[22]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_reg_23_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[23]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_26_ ( 
        .D(n17036), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_26_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_27_ ( 
        .D(n17034), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_27_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_28_ ( 
        .D(n17035), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_28_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_29_ ( 
        .D(n17033), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_29_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_30_ ( 
        .D(n17032), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_30_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_31_ ( 
        .D(n17031), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_31_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_32_ ( 
        .D(n17027), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_32_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_33_ ( 
        .D(n17028), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_33_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_34_ ( 
        .D(n52521), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_34_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_35_ ( 
        .D(n52522), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_35_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_36_ ( 
        .D(n52518), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_36_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_37_ ( 
        .D(n52524), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_37_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_38_ ( 
        .D(n52520), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_38_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_39_ ( 
        .D(n52523), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_39_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_40_ ( 
        .D(n52517), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_40_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_41_ ( 
        .D(n52519), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_41_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_42_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[42]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_42_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_43_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[43]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_43_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_44_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[44]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_44_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_45_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[45]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_45_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_46_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[46]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_46_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_47_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[47]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_47_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_48_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[48]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_48_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_reg_49_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[49]), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_49_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_N586), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_1_ ( 
        .D(n3176), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_2_ ( 
        .D(n51978), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_3_ ( 
        .D(n3174), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_4_ ( 
        .D(n51979), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_5_ ( 
        .D(n51980), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_6_ ( 
        .D(n51981), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_7_ ( 
        .D(n12856), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_reg_8_ ( 
        .D(n53175), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_reg_1_ ( 
        .D(n3167), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_reg_5_ ( 
        .D(n3163), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_0_ ( 
        .D(n3162), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_1_ ( 
        .D(n3161), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_2_ ( 
        .D(n3160), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_3_ ( 
        .D(n3159), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_4_ ( 
        .D(n3158), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_5_ ( 
        .D(n3157), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_6_ ( 
        .D(n3156), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_7_ ( 
        .D(n3155), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1_reg_8_ ( 
        .D(n3154), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_0_ ( 
        .D(n27066), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_1_ ( 
        .D(n27067), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_2_ ( 
        .D(n27068), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_3_ ( 
        .D(n27069), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_4_ ( 
        .D(n27070), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_5_ ( 
        .D(n27071), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_6_ ( 
        .D(n27072), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_7_ ( 
        .D(n27073), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_8_ ( 
        .D(n27074), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i_reg_9_ ( 
        .D(n27075), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_expa_ff_reg ( 
        .D(n3143), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_expa_ff) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_reg ( 
        .D(n4743), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_qnan_d) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_ine_reg ( .D(
        n3142), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_ine_conv) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_8_ ( .D(n9485), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3141) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_freeze_flushpipe_r_reg ( .D(
        n9468), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3426) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_11_ ( 
        .D(n9698), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3138) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_load_reg ( .D(n9474), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3136) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_31_ ( .D(n9423), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3134) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_sel_imm_reg ( .D(n9195), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3132) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_31_ ( 
        .D(n9676), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3130) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_31_ ( .D(
        n78327), .CLK(clk_i), .QN(n3128) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_7_ ( 
        .D(n9632), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3127) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_7_ ( .D(
        n59581), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_7_ ( 
        .D(n78340), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_10_ ( 
        .D(n3124), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[10]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_9_ ( .D(
        or1200_cpu_to_sr[9]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n3123) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_0_ ( .D(
        or1200_immu_top_N3), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n3121) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_21_ ( .D(n9584), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3117) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_11_ ( 
        .D(n9628), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3115) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_11_ ( .D(
        n59580), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_11_ ( 
        .D(n78346), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_14_ ( 
        .D(n3112), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[14]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_cache_dirty_needs_writeback_reg ( 
        .D(n9391), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3111) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_cnt_reg_3_ ( .D(n9384), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3109) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_cnt_reg_2_ ( .D(n9378), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3107) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_load_reg ( .D(n9344), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3105) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_fsm_state_cur_reg_0_ ( .D(n78265), 
        .CLK(clk_i), .RESET(n53192), .SET(dwb_rst_i), .QN(n3103) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_stb_o_reg ( .D(dwb_biu_N36), .CLK(clk_i), .RESET(n53192), .SET(dwb_rst_i), .QN(n3100) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_ack_cnt_reg ( .D(n52473), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n3376) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_biu_ack_cnt_reg ( .D(n52472), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n3097) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_err_cnt_reg ( .D(n9388), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n3095) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_biu_err_cnt_reg ( .D(n9387), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n3375) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_state_reg_1_ ( .D(
        n9383), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3092) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_state_reg_2_ ( .D(
        n9390), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3090) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_hitmiss_eval_reg ( .D(
        n9382), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3088) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_state_reg_0_ ( .D(
        n9381), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3086) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_did_early_load_ack_reg ( 
        .D(n9389), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3084) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_cache_inhibit_reg ( 
        .D(n9347), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3082) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_lsu_except_align_reg ( .D(n9458), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3080) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_31_ ( .D(n9677), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3078) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_lsu_ex_lsu_op_reg_3_ ( .D(n9459), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3076) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_store_reg ( .D(n52470), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3074) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_0_ ( .D(n3072), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3071) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_7_ ( .D(n3069), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3068) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_lsu_dcpu_adr_r_reg_0_ ( .D(n3066), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3419) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_2_ ( 
        .D(n3064), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3063) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_3_ ( 
        .D(n3061), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3060) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_4_ ( 
        .D(n3058), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3057) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_5_ ( 
        .D(n3055), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3054) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_6_ ( 
        .D(n3052), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3051) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_7_ ( 
        .D(n3049), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3048) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_8_ ( 
        .D(n3046), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3045) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_9_ ( 
        .D(n3043), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3042) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_10_ ( 
        .D(n3040), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3039) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_11_ ( 
        .D(n3037), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3036) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_12_ ( 
        .D(n3034), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3033) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_13_ ( 
        .D(n3031), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3030) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_14_ ( 
        .D(n3028), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3027) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_15_ ( 
        .D(n3025), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3024) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_16_ ( 
        .D(n3022), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3021) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_17_ ( 
        .D(n3019), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3018) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_18_ ( 
        .D(n3016), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3015) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_19_ ( 
        .D(n3013), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3012) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_20_ ( 
        .D(n3010), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3009) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_21_ ( 
        .D(n3007), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3006) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_22_ ( 
        .D(n3004), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3003) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_23_ ( 
        .D(n3001), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3000) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_24_ ( 
        .D(n2998), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2997) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_25_ ( 
        .D(n2995), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2994) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_26_ ( 
        .D(n2992), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2991) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_27_ ( 
        .D(n2989), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2988) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_28_ ( 
        .D(n2986), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2985) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_29_ ( 
        .D(n2983), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2982) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_30_ ( 
        .D(n2980), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2979) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_addrtarget_reg_31_ ( 
        .D(n2977), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2976) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_30_ ( .D(n9424), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2974) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_branch_op_reg_1_ ( .D(
        n9456), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2972) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_op_reg_1_ ( .D(
        n9606), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2970) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_0_ ( .D(n2967), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(supv) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dmr1_reg_23_ ( .D(n9326), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n2966) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_23_ ( .D(n2964), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2963) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_10_ ( .D(
        or1200_cpu_to_sr[10]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n2961) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_31_ ( .D(n2959), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2958) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_31_ ( 
        .D(n9673), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2956) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_31_ ( 
        .D(n59579), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_31_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2_reg ( 
        .D(n78435), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_sign_i_reg ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n254), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_output_o_31_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_31_ ( 
        .D(n27324), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[31]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_22_ ( 
        .D(n2953), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_22_ ( 
        .D(n2952), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N105), .CLK(clk_i), .QN(n2951) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_22_ ( .D(
        n2950), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[22]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_22_ ( 
        .D(n9617), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2949) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_22_ ( .D(
        n59578), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_22_ ( 
        .D(n78364), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_25_ ( 
        .D(n2946), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_31_ ( 
        .D(n2945), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[31]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_31_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N114), .CLK(clk_i), .QN(n2944) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_21_ ( .D(
        n51976), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[21]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_21_ ( .D(n2942), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2941) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_21_ ( 
        .D(n9649), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2939) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_21_ ( 
        .D(n59577), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_21_ ( 
        .D(n78367), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_24_ ( 
        .D(n2936), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_infa_f_r_reg ( 
        .D(n2935), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_infa_f_r) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_inf_reg ( 
        .D(n4747), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_inf_d) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_opa_nan_reg ( 
        .D(n2934), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_nan) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_0_ ( 
        .D(n52486), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_1_ ( 
        .D(n52499), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_2_ ( 
        .D(n52498), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_3_ ( 
        .D(n78190), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_4_ ( 
        .D(n52492), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_5_ ( 
        .D(n52493), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_6_ ( 
        .D(n52489), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_7_ ( 
        .D(n52494), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_8_ ( 
        .D(n78189), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_9_ ( 
        .D(n52505), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_10_ ( 
        .D(n52496), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_11_ ( 
        .D(n52506), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_12_ ( 
        .D(n52507), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_13_ ( 
        .D(n52508), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_14_ ( 
        .D(n52490), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_15_ ( 
        .D(n52503), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_16_ ( 
        .D(n52502), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_17_ ( 
        .D(n52501), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_18_ ( 
        .D(n52500), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_19_ ( 
        .D(n52491), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_20_ ( 
        .D(n52509), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_21_ ( 
        .D(n52497), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_22_ ( 
        .D(n52504), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_24_ ( 
        .D(n78199), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_25_ ( 
        .D(n78200), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_26_ ( 
        .D(n78197), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_27_ ( 
        .D(n78201), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[27]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_28_ ( 
        .D(n78202), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[28]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_29_ ( 
        .D(n78246), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[29]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_30_ ( 
        .D(n78203), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[30]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_30_ ( 
        .D(n9640), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2902) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_30_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_30_), .CLK(clk_i), 
        .QN(n2900) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_ine_o_reg ( 
        .D(n2899), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_ine_o) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_0_ ( 
        .D(n2898), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_1_ ( 
        .D(n2897), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_2_ ( 
        .D(n2896), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_3_ ( 
        .D(n2895), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_4_ ( 
        .D(n2894), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_5_ ( 
        .D(n2893), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_6_ ( 
        .D(n2892), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_7_ ( 
        .D(n2891), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_8_ ( 
        .D(n2890), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_9_ ( 
        .D(n2889), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_10_ ( 
        .D(n2888), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_11_ ( 
        .D(n2887), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_12_ ( 
        .D(n2886), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_13_ ( 
        .D(n2885), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_14_ ( 
        .D(n2884), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_15_ ( 
        .D(n2883), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_16_ ( 
        .D(n2882), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_17_ ( 
        .D(n2881), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_18_ ( 
        .D(n2880), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_19_ ( 
        .D(n2879), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_20_ ( 
        .D(n2878), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_21_ ( 
        .D(n2877), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_23_ ( 
        .D(n2876), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_24_ ( 
        .D(n2875), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_25_ ( 
        .D(n2874), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_26_ ( 
        .D(n2873), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_27_ ( 
        .D(n2872), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[27]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_28_ ( 
        .D(n2871), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[28]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_29_ ( 
        .D(n2870), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[29]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_29_ ( 
        .D(n2869), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[29]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_29_ ( .D(
        n78209), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[29]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_29_ ( 
        .D(n9641), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2867) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_29_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_), .CLK(clk_i), 
        .QN(n2865) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_28_ ( 
        .D(n2864), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[28]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_28_ ( .D(
        n78196), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[28]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_28_ ( 
        .D(n9642), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2862) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_28_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_), .CLK(clk_i), 
        .QN(n2860) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_27_ ( 
        .D(n2859), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[27]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_27_ ( 
        .D(n2858), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[27]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_27_ ( .D(
        n78195), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[27]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_27_ ( 
        .D(n9643), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2856) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_27_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_), .CLK(clk_i), 
        .QN(n2854) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_15_ ( 
        .D(n5544), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_15_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N98), .CLK(clk_i), .QN(n2853) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_15_ ( .D(
        n2852), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[15]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_15_ ( .D(n77129), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2850) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_15_ ( 
        .D(n9655), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2848) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_15_ ( 
        .D(n59572), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_15_ ( 
        .D(n78353), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_18_ ( 
        .D(n2845), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[18]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_lsu_dcpu_adr_r_reg_1_ ( .D(n2844), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2843) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_7_ ( 
        .D(n9663), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2841) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_7_ ( 
        .D(n59571), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_10_ ( 
        .D(n2838), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[10]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_12_ ( .D(or1200_du_N107), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n2837) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_12_ ( 
        .D(n9658), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2835) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_12_ ( 
        .D(n78351), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_15_ ( 
        .D(n2832), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[15]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_3_ ( .D(
        or1200_cpu_to_sr[3]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n3418) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_8_ ( 
        .D(n9662), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2830) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_8_ ( 
        .D(n78343), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_11_ ( 
        .D(n2827), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[11]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_comp_op_reg_0_ ( .D(n9580), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2826) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_21_ ( .D(n9212), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2824) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_21_ ( .D(n2822), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2821) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_31_ ( .D(n9202), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2819) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_31_ ( .D(n2817), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2816) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_28_ ( .D(n51945), .CLK(clk_i), .RESET(rst_i), .SET(n53192), .QN(n2814) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_28_ ( .D(n2811), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(ex_insn[28]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_28_ ( .D(n2808), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(wb_insn[28]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rfwb_op_reg_1_ ( .D(n9465), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2807) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_2_ ( .D(n2805), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2804) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_2_ ( 
        .D(n9668), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2802) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_2_ ( 
        .D(n78433), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_5_ ( 
        .D(n2799), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[5]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_7_ ( .D(n9334), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n2798) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_11_ ( .D(n9330), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n2796) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_4_ ( .D(n76992), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n2794) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_4_ ( .D(n2792), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2791) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_4_ ( 
        .D(n9635), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2789) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_4_ ( .D(
        n59567), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_4_ ( 
        .D(n78334), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_7_ ( 
        .D(n2786), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[7]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_4_ ( .D(n9337), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n2785) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_4_ ( .D(
        or1200_cpu_to_sr[4]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n2783) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_hitmiss_eval_reg ( .D(
        n9471), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2781) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_state_reg_1_ ( .D(
        n77355), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2779) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_state_reg_0_ ( .D(
        n9477), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2777) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_biu_stb_reg_reg ( .D(iwb_biu_N62), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n2775) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_stb_o_reg ( .D(iwb_biu_N36), .CLK(clk_i), .RESET(n53192), .SET(iwb_rst_i), .QN(n2773) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_fsm_state_cur_reg_0_ ( .D(n78181), 
        .CLK(clk_i), .RESET(n53192), .SET(iwb_rst_i), .QN(n3374) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_11_ ( .D(n2770), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n2769) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_cyc_o_reg ( .D(n78181), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n2767) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_err_cnt_reg ( .D(n9481), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n2765) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_biu_err_cnt_reg ( .D(n9480), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n2763) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_ack_cnt_reg ( .D(n9482), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n2761) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_biu_ack_cnt_reg ( .D(n9479), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n2759) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_saved_reg ( .D(n9455), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n2757) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_err_saved_reg_2_ ( .D(n9392), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2755) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_0_ ( .D(n9454), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2753) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_1_ ( .D(n9453), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2751) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_2_ ( .D(n9452), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2749) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_3_ ( .D(n9451), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2747) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_4_ ( .D(n9450), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2745) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_5_ ( .D(n9449), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2743) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_6_ ( .D(n9448), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2741) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_7_ ( .D(n9447), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2739) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_8_ ( .D(n9446), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2737) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_9_ ( .D(n9445), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2735) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_10_ ( .D(n9444), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2733) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_11_ ( .D(n9443), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2731) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_12_ ( .D(n9442), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2729) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_13_ ( .D(n9441), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2727) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_14_ ( .D(n9440), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2725) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_15_ ( .D(n9439), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2723) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_17_ ( .D(n9437), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2721) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_18_ ( .D(n9436), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2719) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_19_ ( .D(n9435), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2717) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_20_ ( .D(n9434), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2715) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_21_ ( .D(n9433), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2713) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_23_ ( .D(n9431), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2711) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_24_ ( .D(n9430), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2709) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_25_ ( .D(n9429), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2707) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_27_ ( .D(n9427), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2705) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_29_ ( .D(n9425), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2703) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_16_ ( .D(n2700), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_if_insn_saved[16]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_22_ ( .D(n2698), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_if_insn_saved[22]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_26_ ( .D(n2696), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_if_insn_saved[26]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_insn_saved_reg_28_ ( .D(n2694), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_if_insn_saved[28]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_branch_op_reg_2_ ( .D(
        n9675), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2693) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_op_reg_2_ ( .D(
        n9674), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2691) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_7_ ( .D(
        or1200_cpu_to_sr[7]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n2687) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_20_ ( .D(n9585), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2685) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_20_ ( .D(n9213), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2683) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_20_ ( .D(n2681), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2680) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_19_ ( .D(n9586), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2678) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_19_ ( .D(n9214), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2676) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_19_ ( .D(n2674), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2673) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_18_ ( .D(n9587), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2671) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_18_ ( .D(n9215), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2669) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_18_ ( .D(n2667), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2666) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_17_ ( .D(n9588), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2664) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_17_ ( .D(n9216), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2662) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_17_ ( .D(n2660), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2659) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_16_ ( .D(n9589), 
        .CLK(clk_i), .RESET(rst_i), .SET(n53192), .QN(n2657) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_16_ ( .D(n2654), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(ex_insn[16]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_16_ ( .D(n2651), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(wb_insn[16]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_15_ ( .D(n9590), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3392) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_15_ ( .D(n9218), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2649) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_15_ ( .D(n2647), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2646) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_14_ ( .D(n9591), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2644) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_14_ ( .D(n9219), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2642) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_14_ ( .D(n2640), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2639) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_13_ ( .D(n9592), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2637) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_13_ ( .D(n9220), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2635) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_13_ ( .D(n2633), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2632) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_12_ ( .D(n9593), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2630) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_12_ ( .D(n9221), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2628) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_12_ ( .D(n2626), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2625) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_11_ ( .D(n9594), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2623) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_11_ ( .D(n9222), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2621) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_11_ ( .D(n2619), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2618) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_30_ ( .D(n9571), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2616) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_30_ ( .D(n9203), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2614) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_30_ ( .D(n2612), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2611) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_26_ ( .D(n9575), 
        .CLK(clk_i), .RESET(rst_i), .SET(n53192), .QN(n2609) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_lsu_ex_lsu_op_reg_0_ ( .D(n60727), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2607) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_26_ ( .D(n2604), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(ex_insn[26]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_26_ ( .D(n2601), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(wb_insn[26]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_branch_op_reg_0_ ( .D(
        n9457), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2600) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_branch_op_reg_0_ ( .D(
        n9607), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2598) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_27_ ( .D(n9574), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2596) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_27_ ( .D(n9206), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2594) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_27_ ( .D(n2592), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2591) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_29_ ( .D(n9572), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2589) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_macrc_op_reg ( .D(n9196), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2587) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_spr_read_reg ( .D(n9608), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2585) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_freeze_multicycle_cnt_reg_0_ ( 
        .D(n9495), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2583) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rfwb_op_reg_3_ ( .D(n9463), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2581) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_valid_re_reg ( .D(
        n9565), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2579) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_valid_re_r_reg ( .D(n2579), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_op_valid_re_r) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_spr_write_reg ( .D(n9494), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2577) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rf_addrw_reg_0_ ( .D(n9201), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2575) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_rfaddrw_reg_0_ ( .D(
        n2573), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2572) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_lsu_ex_lsu_op_reg_2_ ( .D(n9460), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3423) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_lsu_ex_lsu_op_reg_1_ ( .D(n9461), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2569) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rfwb_op_reg_2_ ( .D(n9464), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2567) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_22_ ( .D(n2565), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2564) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_1_ ( .D(n2562), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2561) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_30_ ( .D(n2559), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2558) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_29_ ( .D(n2556), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2555) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_28_ ( .D(n75887), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2552) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_27_ ( .D(n2550), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2549) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op_reg_4_ ( .D(n9235), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2547) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_11_ ( .D(n2545), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2544) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_29_ ( .D(n9204), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2542) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_29_ ( .D(n2540), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2539) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dbg_is_o_reg_1_ ( .D(n52471), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2536) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_0_ ( .D(n9605), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3390) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_0_ ( .D(n2533), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2532) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1_reg_0_ ( 
        .D(n78438), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_reg_0_ ( 
        .D(n27420), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_reg_0_ ( 
        .D(n27421), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_sign_o_reg ( 
        .D(n2527), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_sign_o) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_mac_op_reg_0_ ( .D(n9568), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2526) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_0_ ( .D(n9233), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2524) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_0_ ( .D(n2522), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2521) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op_reg_0_ ( .D(n9239), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2519) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_1_ ( .D(n9604), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2517) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_1_ ( .D(n2515), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2514) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1_reg_1_ ( 
        .D(n78437), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_reg_1_ ( 
        .D(n78251), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_reg_1_ ( 
        .D(n78250), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_1_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op_reg_1_ ( .D(n9238), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2508) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_1_ ( .D(n9232), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2506) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_1_ ( .D(n2504), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2503) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_mac_op_reg_1_ ( .D(n9567), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2501) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_2_ ( .D(n9603), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2499) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_2_ ( .D(n2497), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2496) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_r_reg_2_ ( .D(n2493), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_op_r_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1_reg_2_ ( 
        .D(n78436), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_reg_2_ ( 
        .D(n27433), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_2_), .CLK(clk_i), 
        .QN(n2491) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_31_ ( 
        .D(n2490), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[31]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_24_ ( 
        .D(n2489), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_25_ ( 
        .D(n2488), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_29_ ( 
        .D(n2487), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[29]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_32_ ( 
        .D(n52485), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[32]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_38_ ( 
        .D(n2485), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[38]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_44_ ( 
        .D(n2484), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[44]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_45_ ( 
        .D(n2483), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[45]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_46_ ( 
        .D(n2482), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[46]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_47_ ( 
        .D(n2481), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[47]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_2_ ( 
        .D(n2480), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_7_ ( 
        .D(n2479), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_8_ ( 
        .D(n2478), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_12_ ( 
        .D(n2477), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_15_ ( 
        .D(n2476), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r_reg_7_ ( 
        .D(n2474), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_mac_op_reg_2_ ( .D(n9566), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2473) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op_reg_2_ ( .D(n2470), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(or1200_cpu_alu_op_2_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_2_ ( .D(n9231), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2469) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_2_ ( .D(n2467), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2466) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_3_ ( .D(n9602), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2464) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_3_ ( .D(n2462), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2461) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_r_reg_3_ ( .D(n2458), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_op_r_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_start_i_reg ( .D(
        n2457), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_start_i) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_state_reg ( 
        .D(n9559), .CLK(clk_i), .QN(n2455) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_reg_0_ ( 
        .D(n2454), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_reg_2_ ( 
        .D(n2453), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_reg_4_ ( 
        .D(n2452), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_reg_1_ ( 
        .D(n9562), .CLK(clk_i), .QN(n2451) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_0_ ( 
        .D(n2449), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[0]), .CLK(clk_i), 
        .QN(n2448) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_2_ ( 
        .D(n2447), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_2_ ( 
        .D(n27447), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_8_ ( 
        .D(n2445), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_8_ ( 
        .D(n27448), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_10_ ( 
        .D(n2443), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_10_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[10]), .CLK(clk_i), 
        .QN(n2442) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_18_ ( 
        .D(n2441), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[18]), .CLK(clk_i), 
        .QN(n2440) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_26_ ( 
        .D(n2439), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shl1_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_v_shl_0_), .CLK(
        clk_i), .QN(n2437) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_0_ ( 
        .D(n2436), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_1_ ( 
        .D(n2435), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_1_ ( 
        .D(n78229), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_1_ ( 
        .D(n2433), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_2_ ( 
        .D(n2432), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_9_ ( 
        .D(n2431), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_9_ ( 
        .D(n78233), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_9_ ( 
        .D(n2429), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_6_ ( 
        .D(n2428), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_6_ ( 
        .D(n5507), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_6_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N89), .CLK(clk_i), .QN(n2427) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_6_ ( .D(
        n51959), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_10_ ( 
        .D(n2425), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_7_ ( 
        .D(n2424), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_7_ ( 
        .D(n5506), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_7_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N90), .CLK(clk_i), .QN(n2423) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_7_ ( .D(
        n2422), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_17_ ( 
        .D(n2421), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_17_ ( 
        .D(n78237), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_18_ ( 
        .D(n2419), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_15_ ( 
        .D(n2418), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_25_ ( 
        .D(n2417), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_25_ ( 
        .D(n27456), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_26_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_N139), .CLK(clk_i), .QN(DP_OP_742J1_130_9702_n59) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_3_ ( 
        .D(n2414), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_3_ ( 
        .D(n78230), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_3_ ( 
        .D(n2412), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_0_ ( 
        .D(n2411), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_0_ ( 
        .D(n5550), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_0_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N83), .CLK(clk_i), .QN(n2410) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_0_ ( .D(
        n2409), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_11_ ( 
        .D(n2408), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_11_ ( 
        .D(n78234), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_11_ ( 
        .D(n2406), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_8_ ( 
        .D(n2405), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_8_ ( 
        .D(n5505), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_8_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N91), .CLK(clk_i), .QN(n2404) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_8_ ( .D(
        n51975), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_19_ ( 
        .D(n2402), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_19_ ( 
        .D(n78238), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_19_ ( 
        .D(n2400), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_16_ ( 
        .D(n2399), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_4_ ( 
        .D(n2398), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[4]), .CLK(clk_i), 
        .QN(n2397) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_4_ ( 
        .D(n2396), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_1_ ( 
        .D(n2395), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_1_ ( 
        .D(n5539), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_1_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N84), .CLK(clk_i), .QN(n2394) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_1_ ( .D(
        n51974), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_12_ ( 
        .D(n2392), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_12_ ( 
        .D(n78235), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_12_ ( 
        .D(n2390), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_9_ ( 
        .D(n2389), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_9_ ( 
        .D(n5503), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_9_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N92), .CLK(clk_i), .QN(n2388) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_9_ ( .D(
        n51973), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_20_ ( 
        .D(n2386), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_20_ ( 
        .D(n2384), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_17_ ( 
        .D(n2383), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_5_ ( 
        .D(n2382), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_5_ ( 
        .D(n27472), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_5_ ( 
        .D(n2380), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_2_ ( 
        .D(n2379), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_2_ ( 
        .D(n5513), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_2_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N85), .CLK(clk_i), .QN(n2378) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_2_ ( .D(
        n2377), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_21_ ( 
        .D(n2376), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_21_ ( 
        .D(n2374), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_18_ ( 
        .D(n2373), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_13_ ( 
        .D(n2372), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_13_ ( 
        .D(n2370), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_10_ ( 
        .D(n2369), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_10_ ( 
        .D(n5549), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_10_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N93), .CLK(clk_i), .QN(n2368) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_10_ ( .D(
        n51972), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_7_ ( 
        .D(n2366), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_7_ ( 
        .D(n78232), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_8_ ( 
        .D(n2364), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_5_ ( 
        .D(n2363), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_5_ ( 
        .D(n5508), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_5_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N88), .CLK(clk_i), .QN(n2362) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_5_ ( .D(
        n51971), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_23_ ( 
        .D(n2360), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_23_ ( 
        .D(n78241), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_15_ ( 
        .D(n2358), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_15_ ( 
        .D(n78236), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_6_ ( 
        .D(n2356), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_6_ ( 
        .D(n78231), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_6_ ( 
        .D(n2354), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_3_ ( 
        .D(n2353), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_3_ ( 
        .D(n5510), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_3_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N86), .CLK(clk_i), .QN(n2352) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_3_ ( .D(
        n51970), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_7_ ( 
        .D(n2350), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_4_ ( 
        .D(n2349), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_4_ ( 
        .D(n5509), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_4_ ( .D(
        or1200_cpu_or1200_fpu_fpu_arith_N87), .CLK(clk_i), .QN(n2348) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_4_ ( .D(
        n51960), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_14_ ( 
        .D(n2346), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_14_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[14]), .CLK(clk_i), 
        .QN(n2345) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_14_ ( 
        .D(n2344), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_11_ ( 
        .D(n2343), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_11_ ( 
        .D(n5548), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_11_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N94), .CLK(clk_i), .QN(n2342) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_11_ ( .D(
        n51969), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_15_ ( 
        .D(n2340), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_12_ ( 
        .D(n2339), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_12_ ( 
        .D(n5547), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_12_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N95), .CLK(clk_i), .QN(n2338) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_12_ ( .D(
        n51968), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_22_ ( 
        .D(n2336), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[22]), .CLK(clk_i), 
        .QN(n2335) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_22_ ( 
        .D(n2334), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_19_ ( 
        .D(n2333), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_23_ ( 
        .D(n2332), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_20_ ( 
        .D(n2331), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_16_ ( 
        .D(n2330), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_16_ ( 
        .D(n27495), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_16_ ( 
        .D(n2328), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_13_ ( 
        .D(n2327), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_13_ ( 
        .D(n5546), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_13_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N96), .CLK(clk_i), .QN(n2326) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_13_ ( .D(
        n51967), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_17_ ( 
        .D(n2324), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_14_ ( 
        .D(n2323), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_14_ ( 
        .D(n5545), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_14_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N97), .CLK(clk_i), .QN(n2322) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_14_ ( .D(
        n51966), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_qutnt_o_reg_24_ ( 
        .D(n2320), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_24_ ( 
        .D(n78242), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_24_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_24_ ( 
        .D(n2318), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_24_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2_reg_21_ ( 
        .D(n2317), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_reg_25_ ( 
        .D(n2316), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_25_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_1_ ( 
        .D(n2313), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_2_ ( 
        .D(n2311), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_3_ ( 
        .D(n2309), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_4_ ( 
        .D(n2307), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_5_ ( 
        .D(n2305), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_6_ ( 
        .D(n2303), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_7_ ( 
        .D(n2301), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_8_ ( 
        .D(n2299), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_9_ ( 
        .D(n2297), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_10_ ( 
        .D(n2295), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_11_ ( 
        .D(n2293), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_12_ ( 
        .D(n2291), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_13_ ( 
        .D(n2289), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_14_ ( 
        .D(n2287), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_15_ ( 
        .D(n2285), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_16_ ( 
        .D(n2283), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_17_ ( 
        .D(n2281), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_18_ ( 
        .D(n2279), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_19_ ( 
        .D(n2277), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_20_ ( 
        .D(n2275), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_21_ ( 
        .D(n2273), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_22_ ( 
        .D(n2271), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_23_ ( 
        .D(n2269), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_24_ ( 
        .D(n2267), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_25_ ( 
        .D(n2265), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd_reg_26_ ( 
        .D(n2263), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_26_ ( 
        .D(n2262), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_26_ ( 
        .D(n27499), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_26_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_25_ ( 
        .D(n2260), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_25_ ( 
        .D(n27500), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_25_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_24_ ( 
        .D(n2258), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_24_ ( 
        .D(n27501), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_24_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_23_ ( 
        .D(n70499), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_23_ ( 
        .D(n27502), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_22_ ( 
        .D(n2254), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_22_ ( 
        .D(n27503), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_21_ ( 
        .D(n70523), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_21_ ( 
        .D(n27504), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_20_ ( 
        .D(n2250), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_20_ ( 
        .D(n27505), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_19_ ( 
        .D(n2248), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_19_ ( 
        .D(n27506), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_18_ ( 
        .D(n2246), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_18_ ( 
        .D(n27507), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_17_ ( 
        .D(n2244), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_17_ ( 
        .D(n27508), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_16_ ( 
        .D(n2242), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_16_ ( 
        .D(n27509), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_15_ ( 
        .D(n2240), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_15_ ( 
        .D(n27510), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_14_ ( 
        .D(n2238), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_14_ ( 
        .D(n27511), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_13_ ( 
        .D(n2236), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_13_ ( 
        .D(n27512), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_12_ ( 
        .D(n2234), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_12_ ( 
        .D(n27513), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_11_ ( 
        .D(n2232), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_11_ ( 
        .D(n27514), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_10_ ( 
        .D(n2230), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_10_ ( 
        .D(n27515), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_9_ ( 
        .D(n2228), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_9_ ( 
        .D(n27516), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_8_ ( 
        .D(n2226), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_8_ ( 
        .D(n27517), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_7_ ( 
        .D(n70514), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_7_ ( 
        .D(n27518), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_6_ ( 
        .D(n70512), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_6_ ( 
        .D(n27519), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_5_ ( 
        .D(n2220), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_5_ ( 
        .D(n27520), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_4_ ( 
        .D(n2218), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_4_ ( 
        .D(n27521), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_3_ ( 
        .D(n2216), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_3_ ( 
        .D(n27522), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_2_ ( 
        .D(n70507), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_2_ ( 
        .D(n27523), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_1_ ( 
        .D(n70505), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_1_ ( 
        .D(n27524), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_rmndr_o_reg_0_ ( 
        .D(n2210), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_reg_0_ ( 
        .D(n27525), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_state_reg ( .D(n2208), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_state) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_count_reg_5_ ( .D(
        n2207), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_count_5_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_count_reg_0_ ( .D(
        n2206), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_count_0_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_count_reg_1_ ( .D(
        n2205), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_count_1_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_count_reg_2_ ( .D(
        n2204), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_count_2_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_count_reg_3_ ( .D(
        n2203), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_count_3_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_count_reg_4_ ( .D(
        n2202), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_count_4_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_ready_o_reg ( .D(n2201), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_done) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_14_ ( .D(n2200), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2199) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_12_ ( .D(n2197), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2196) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_8_ ( .D(n2194), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2193) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rfwb_op_reg_0_ ( .D(n9466), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2191) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_valid_reg ( .D(
        n2189), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2188) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op_reg_3_ ( .D(n9236), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2186) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_3_ ( .D(n9230), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2184) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_3_ ( .D(n2182), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2181) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_conv_shr_reg_0_ ( .D(n2179), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_conv_shr[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_conv_shr_reg_1_ ( .D(n27531), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_conv_shr[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_conv_shr_reg_2_ ( .D(n27532), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_conv_shr[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_conv_shr_reg_3_ ( .D(n27533), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_conv_shr[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_conv_shr_reg_4_ ( .D(n27534), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_conv_shr[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_conv_shr_reg_5_ ( .D(n27535), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_conv_shr[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_conv_shr_reg_6_ ( .D(n27536), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_conv_shr[6]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_4_ ( .D(n9601), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2172) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_4_ ( .D(n2170), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2169) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_r_reg_4_ ( .D(n2166), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_op_r_4_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_4_ ( .D(n9229), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2165) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_4_ ( .D(n2163), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2162) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_5_ ( .D(n9600), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2160) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_5_ ( .D(n2158), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2157) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_r_reg_5_ ( .D(n2154), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_op_r_5_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_5_ ( .D(n9228), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2153) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_5_ ( .D(n2151), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2150) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_6_ ( .D(n9599), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2148) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_6_ ( .D(n2146), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2145) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_r_reg_6_ ( .D(n2142), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_op_r_6_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op2_reg_0_ ( .D(n9243), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2141) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_6_ ( .D(n9227), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2139) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_6_ ( .D(n2137), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2136) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_7_ ( .D(n9598), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2134) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_7_ ( .D(n2132), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2131) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op2_reg_1_ ( .D(n9242), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2129) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_7_ ( .D(n9226), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2127) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_7_ ( .D(n2125), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2124) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_8_ ( .D(n9597), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2122) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_8_ ( .D(n2120), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2119) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op2_reg_2_ ( .D(n9241), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2117) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_8_ ( .D(n9225), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2115) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_8_ ( .D(n2113), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2112) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_9_ ( .D(n9596), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2110) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_9_ ( .D(n2108), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2107) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_alu_op2_reg_3_ ( .D(n9240), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2105) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_9_ ( .D(n9224), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2103) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_9_ ( .D(n2101), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2100) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_10_ ( .D(n9595), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2098) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_10_ ( .D(n2096), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2095) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_10_ ( .D(n9223), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2093) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_10_ ( .D(n2091), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2090) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_22_ ( .D(n2087), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(id_insn_22_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_comp_op_reg_1_ ( .D(n9579), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2086) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_22_ ( .D(n2083), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(ex_insn[22]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_22_ ( .D(n2080), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(wb_insn[22]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rf_addrw_reg_1_ ( .D(n9200), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2079) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_rfaddrw_reg_1_ ( .D(
        n2077), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2076) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_12_ ( .D(n2074), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2073) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_23_ ( .D(n9582), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2071) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_comp_op_reg_2_ ( .D(n9578), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2069) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_23_ ( .D(n9210), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2067) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_23_ ( .D(n2065), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2064) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rf_addrw_reg_2_ ( .D(n9199), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2062) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_rfaddrw_reg_2_ ( .D(
        n2060), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2059) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_13_ ( .D(n2057), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2056) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_24_ ( .D(n9581), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2054) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_comp_op_reg_3_ ( .D(n9577), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2052) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_24_ ( .D(n9209), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2050) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_24_ ( .D(n2048), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2047) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rf_addrw_reg_3_ ( .D(n9198), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2045) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_rfaddrw_reg_3_ ( .D(
        n2043), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2042) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_14_ ( .D(n2040), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2039) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_id_insn_reg_25_ ( .D(n9576), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2037) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_sig_trap_reg ( .D(n9570), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2035) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_sig_syscall_reg ( .D(n9569), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2033) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_insn_reg_25_ ( .D(n9208), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2031) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_insn_reg_25_ ( .D(n2029), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2028) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_rf_addrw_reg_4_ ( .D(n9197), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2026) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_wb_rfaddrw_reg_4_ ( .D(
        n2024), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2023) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_0_ ( 
        .D(n9670), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2021) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_0_ ( 
        .D(n2018), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_3_ ( 
        .D(n2017), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[3]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_1_ ( 
        .D(n9669), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2016) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_1_ ( 
        .D(n2013), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_4_ ( 
        .D(n2012), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[4]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_23_ ( 
        .D(n9647), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2011) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_23_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .CLK(clk_i), 
        .QN(n2009) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_40_ ( 
        .D(n2008), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r_reg_0_ ( 
        .D(n2007), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_22_ ( 
        .D(n9648), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2006) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_22_ ( 
        .D(n59561), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_r_a_reg ( 
        .D(n78365), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_r_a) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_39_ ( 
        .D(n2003), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[39]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_25_ ( 
        .D(n2002), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[25]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_14_ ( 
        .D(n9656), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n2001) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_14_ ( 
        .D(n78432), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_14_ ( 
        .D(n1998), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_31_ ( 
        .D(n1997), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[31]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_17_ ( 
        .D(n1996), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[17]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_4_ ( 
        .D(n9666), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1995) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_4_ ( 
        .D(n59559), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_4_ ( 
        .D(n78335), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_4_ ( 
        .D(n1992), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_7_ ( 
        .D(n1990), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[7]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_1_ ( 
        .D(n9638), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1989) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_1_ ( .D(
        n59442), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_1_ ( 
        .D(n78330), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_4_ ( 
        .D(n1986), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[4]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_1_ ( .D(or1200_du_N96), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1985) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_1_ ( .D(n9340), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1983) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_3_ ( 
        .D(n9636), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1981) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_3_ ( .D(
        n59558), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_3_ ( 
        .D(n78332), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_6_ ( 
        .D(n1979), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[6]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_3_ ( .D(n9338), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1978) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_3_ ( .D(or1200_du_N98), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1976) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_3_ ( .D(n1974), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1973) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_3_ ( 
        .D(n9667), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1971) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_3_ ( 
        .D(n59557), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_3_ ( 
        .D(n78333), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_3_ ( 
        .D(n1969), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_6_ ( 
        .D(n1968), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[6]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_6_ ( 
        .D(n9633), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1967) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_6_ ( .D(
        n59556), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_6_ ( 
        .D(n78338), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_9_ ( 
        .D(n1964), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[9]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_6_ ( .D(n18256), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1963) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_6_ ( .D(n9335), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1961) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_6_ ( .D(n1959), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1958) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_6_ ( 
        .D(n9664), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1956) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_6_ ( 
        .D(n78339), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_6_ ( 
        .D(n1953), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_9_ ( 
        .D(n1952), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[9]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_6_ ( .D(
        or1200_cpu_to_sr[6]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1951) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_8_ ( 
        .D(n9631), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1949) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_8_ ( .D(
        n59554), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_8_ ( 
        .D(n78342), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_11_ ( 
        .D(n1946), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[11]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_8_ ( .D(n9333), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1945) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_8_ ( .D(
        or1200_cpu_to_sr[8]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1943) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_12_ ( 
        .D(n9627), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1941) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_12_ ( .D(
        n59553), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_12_ ( 
        .D(n78350), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_15_ ( 
        .D(n1939), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[15]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_12_ ( .D(n9329), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1938) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_12_ ( .D(
        or1200_cpu_to_sr[12]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1936) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_14_ ( 
        .D(n9625), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1934) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_14_ ( 
        .D(n78427), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_17_ ( 
        .D(n1931), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[17]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_bit_eph_reg ( .D(
        n9467), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n3417) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_15_ ( 
        .D(n9624), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1929) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_15_ ( .D(
        n59551), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_15_ ( 
        .D(n78426), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_18_ ( 
        .D(n1926), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[18]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_15_ ( .D(n1925), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1924) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_31_ ( .D(n1922), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1921) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_29_ ( .D(n1919), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1918) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_27_ ( .D(n1916), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1915) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_25_ ( .D(n1913), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1912) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_23_ ( .D(n1910), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1909) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_21_ ( .D(n1907), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1906) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_19_ ( .D(n1904), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1903) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_17_ ( .D(n1901), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1900) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_16_ ( .D(n1898), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1897) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_18_ ( .D(n1895), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1894) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_20_ ( .D(n1892), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1891) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_22_ ( .D(n1889), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1888) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_24_ ( .D(n1886), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1885) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_26_ ( .D(n1883), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1882) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_28_ ( .D(n1880), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1879) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_ex_simm_reg_30_ ( .D(n1877), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1876) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_30_ ( 
        .D(n9609), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1874) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_30_ ( 
        .D(n78383), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_30_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_29_ ( 
        .D(n9610), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1871) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_29_ ( 
        .D(n78363), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_29_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_28_ ( 
        .D(n9611), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1868) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_28_ ( 
        .D(n78361), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_28_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_27_ ( 
        .D(n9612), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1865) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_27_ ( 
        .D(n78381), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_27_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_23_ ( 
        .D(n9616), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1862) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_23_ ( 
        .D(n78372), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o_reg_0_ ( 
        .D(n1859), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_exp_o_reg_0_ ( 
        .D(n27627), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_21_ ( 
        .D(n9618), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1857) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_21_ ( .D(
        n59546), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_21_ ( 
        .D(n78366), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_24_ ( 
        .D(n1854), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[24]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_last_eval_miss_reg ( 
        .D(n9164), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1853) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_cnt_reg_3_ ( .D(n9476), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1851) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_cnt_reg_2_ ( .D(n9475), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1849) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_5_ ( .D(n18405), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1847) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_5_ ( .D(n61667), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1844) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_5_ ( 
        .D(n9665), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1842) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_5_ ( 
        .D(n59545), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_5_ ( 
        .D(n78337), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_5_ ( 
        .D(n1839), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_22_ ( 
        .D(n1838), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_8_ ( 
        .D(n1837), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[8]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_5_ ( 
        .D(n9634), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1836) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_5_ ( .D(
        n59544), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_5_ ( 
        .D(n78336), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_8_ ( 
        .D(n1833), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[8]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_5_ ( .D(n9336), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1832) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_5_ ( .D(
        or1200_cpu_to_sr[5]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1830) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_7_ ( .D(n58417), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1828) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_8_ ( .D(or1200_du_N103), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1826) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_9_ ( .D(or1200_du_N104), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1824) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_9_ ( .D(n1822), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1821) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_9_ ( 
        .D(n9630), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1819) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_9_ ( .D(
        n59543), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_9_ ( 
        .D(n78344), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_12_ ( 
        .D(n1816), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[12]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_9_ ( .D(n9332), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1815) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_9_ ( 
        .D(n9661), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1813) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_9_ ( 
        .D(n59542), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_9_ ( 
        .D(n78345), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_9_ ( 
        .D(n1810), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_26_ ( 
        .D(n1809), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_12_ ( 
        .D(n1808), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[12]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_10_ ( .D(or1200_du_N105), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1807) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_10_ ( .D(n1805), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1804) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_10_ ( 
        .D(n9629), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1802) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_10_ ( 
        .D(n78348), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_13_ ( 
        .D(n1799), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[13]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_10_ ( .D(n9331), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1798) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_10_ ( 
        .D(n9660), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1796) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_10_ ( 
        .D(n59541), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_10_ ( 
        .D(n78349), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_10_ ( 
        .D(n1793), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_27_ ( 
        .D(n1792), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[27]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_13_ ( 
        .D(n1791), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[13]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_11_ ( .D(or1200_du_N106), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1790) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_11_ ( .D(n1788), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1787) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_11_ ( 
        .D(n9659), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1785) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_11_ ( 
        .D(n59540), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_11_ ( 
        .D(n78347), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_11_ ( 
        .D(n1782), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_14_ ( 
        .D(n1780), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[14]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_13_ ( .D(or1200_du_N108), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1779) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_13_ ( .D(n1777), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1776) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_13_ ( 
        .D(n9626), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1774) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_13_ ( .D(
        n59539), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_13_ ( 
        .D(n78428), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_16_ ( 
        .D(n1771), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[16]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_13_ ( .D(n9328), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1770) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_13_ ( .D(
        or1200_cpu_to_sr[13]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1768) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_13_ ( 
        .D(n9657), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1766) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_13_ ( 
        .D(n59538), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_13_ ( 
        .D(n78352), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_13_ ( 
        .D(n1764), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_16_ ( 
        .D(n1762), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[16]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_2_ ( 
        .D(n9637), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1761) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_2_ ( .D(
        n59708), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_2_ ( 
        .D(n78331), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_5_ ( 
        .D(n1758), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[5]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_2_ ( .D(or1200_du_N97), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1757) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_2_ ( .D(n9339), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1755) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_ctrl_except_illegal_reg ( .D(
        n51982), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1753) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_sel_o_reg_0_ ( .D(n1749), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(dwb_sel_o[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_sel_o_reg_1_ ( .D(n1746), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(dwb_sel_o[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_sel_o_reg_2_ ( .D(n1743), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(dwb_sel_o[2]) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_sel_o_reg_3_ ( .D(n1740), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(dwb_sel_o[3]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_2_ ( .D(
        or1200_cpu_to_sr[2]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1739) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_1_ ( .D(
        or1200_cpu_to_sr[1]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1737) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_1_ ( .D(n9492), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1735) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1_reg_0_ ( 
        .D(n1735), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_reg_0_ ( 
        .D(n78248), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3_reg_0_ ( 
        .D(n78247), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_2_ ( .D(n9493), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1733) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1_reg_1_ ( 
        .D(n1733), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_reg_1_ ( 
        .D(n78249), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3_reg_1_ ( 
        .D(n78326), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_sign_reg ( .D(
        n1729), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_intfloat_conv_sign)
         );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_lsu_dcpu_adr_r_reg_2_ ( .D(n1728), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1727) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_0_ ( 
        .D(n9639), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1725) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_0_ ( 
        .D(n78329), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_3_ ( 
        .D(n1722), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[3]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_drr_reg_0_ ( .D(or1200_du_N95), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1721) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dsr_reg_0_ ( .D(n9341), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1719) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_0_ ( .D(n9491), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1717) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_0_ ( .D(n1715), .CLK(clk_i), 
        .QN(dbg_dat_o[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_1_ ( .D(n1714), .CLK(clk_i), 
        .QN(dbg_dat_o[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_2_ ( .D(n1713), .CLK(clk_i), 
        .QN(dbg_dat_o[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_3_ ( .D(n1712), .CLK(clk_i), 
        .QN(dbg_dat_o[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_4_ ( .D(n1711), .CLK(clk_i), 
        .QN(dbg_dat_o[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_5_ ( .D(n1710), .CLK(clk_i), 
        .QN(dbg_dat_o[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_6_ ( .D(n1709), .CLK(clk_i), 
        .QN(dbg_dat_o[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_8_ ( .D(n1708), .CLK(clk_i), 
        .QN(dbg_dat_o[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_9_ ( .D(n1707), .CLK(clk_i), 
        .QN(dbg_dat_o[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_10_ ( .D(n1706), .CLK(clk_i), 
        .QN(dbg_dat_o[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_12_ ( .D(n1705), .CLK(clk_i), 
        .QN(dbg_dat_o[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_13_ ( .D(n1704), .CLK(clk_i), 
        .QN(dbg_dat_o[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_14_ ( .D(n1703), .CLK(clk_i), 
        .QN(dbg_dat_o[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_15_ ( .D(n1702), .CLK(clk_i), 
        .QN(dbg_dat_o[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_21_ ( .D(n1701), .CLK(clk_i), 
        .QN(dbg_dat_o[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_27_ ( .D(n1700), .CLK(clk_i), 
        .QN(dbg_dat_o[27]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_28_ ( .D(n1699), .CLK(clk_i), 
        .QN(dbg_dat_o[28]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_29_ ( .D(n52475), .CLK(clk_i), 
        .QN(dbg_dat_o[29]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_30_ ( .D(n1697), .CLK(clk_i), 
        .QN(dbg_dat_o[30]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_31_ ( .D(n1696), .CLK(clk_i), 
        .QN(dbg_dat_o[31]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_16_ ( 
        .D(n5543), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_16_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N99), .CLK(clk_i), .QN(n1695) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_16_ ( .D(
        n51965), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[16]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_16_ ( .D(n1693), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1692) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_16_ ( 
        .D(n9623), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1690) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_16_ ( .D(
        n57312), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_16_ ( 
        .D(n78425), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_19_ ( 
        .D(n1687), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[19]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_16_ ( .D(n78187), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1686) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_16_ ( .D(n1684), .CLK(clk_i), 
        .QN(dbg_dat_o[16]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_16_ ( 
        .D(n9654), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1683) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_16_ ( 
        .D(n59486), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_16_ ( 
        .D(n78431), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_16_ ( 
        .D(n1680), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_33_ ( 
        .D(n1679), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[33]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_19_ ( 
        .D(n1678), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_17_ ( 
        .D(n5542), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_17_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N100), .CLK(clk_i), .QN(n1677) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_17_ ( .D(
        n51964), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[17]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_17_ ( .D(n75375), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1674) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_17_ ( 
        .D(n9622), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1672) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_17_ ( 
        .D(n78424), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_20_ ( 
        .D(n1669), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_17_ ( .D(n1668), .CLK(clk_i), 
        .QN(dbg_dat_o[17]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_17_ ( 
        .D(n9653), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1667) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_17_ ( 
        .D(n59535), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_17_ ( 
        .D(n1664), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_34_ ( 
        .D(n1663), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[34]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_20_ ( 
        .D(n1662), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_18_ ( 
        .D(n5541), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N101), .CLK(clk_i), .QN(n1661) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_18_ ( .D(
        n51963), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[18]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_18_ ( .D(n1659), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1658) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_18_ ( 
        .D(n9621), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1656) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_18_ ( .D(
        n59534), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_18_ ( 
        .D(n78354), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_21_ ( 
        .D(n1653), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_18_ ( .D(n1652), .CLK(clk_i), 
        .QN(dbg_dat_o[18]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_18_ ( 
        .D(n9652), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1651) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_18_ ( 
        .D(n59533), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_18_ ( 
        .D(n78355), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_18_ ( 
        .D(n1648), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_35_ ( 
        .D(n1647), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[35]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_21_ ( 
        .D(n1646), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_19_ ( 
        .D(n5540), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_19_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N102), .CLK(clk_i), .QN(n1645) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_19_ ( .D(
        n51962), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[19]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_19_ ( .D(n1643), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1642) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_19_ ( 
        .D(n9620), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1640) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_19_ ( .D(
        n59532), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_19_ ( 
        .D(n78356), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_22_ ( 
        .D(n1638), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_19_ ( .D(n1637), .CLK(clk_i), 
        .QN(dbg_dat_o[19]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_19_ ( 
        .D(n9651), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1636) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_19_ ( 
        .D(n59531), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_19_ ( 
        .D(n78357), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_36_ ( 
        .D(n1633), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[36]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_22_ ( 
        .D(n1632), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_20_ ( 
        .D(n5538), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_20_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N103), .CLK(clk_i), .QN(n1631) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_20_ ( .D(
        n51961), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[20]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_20_ ( .D(n1629), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1628) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_20_ ( 
        .D(n9619), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1626) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_20_ ( .D(
        n1626), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_20_ ( 
        .D(n78368), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_23_ ( 
        .D(n1623), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_20_ ( .D(n1622), .CLK(clk_i), 
        .QN(dbg_dat_o[20]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_20_ ( 
        .D(n9650), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1621) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_20_ ( 
        .D(n57377), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_20_ ( 
        .D(n78369), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_20_ ( 
        .D(n1618), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_37_ ( 
        .D(n1617), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[37]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_23_ ( 
        .D(n1616), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_21_ ( 
        .D(n5537), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_21_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_N104), .CLK(clk_i), .QN(n1615) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_23_ ( 
        .D(n1614), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_23_ ( 
        .D(n1613), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_output1_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_24_ ( 
        .D(n1612), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_24_ ( 
        .D(n1611), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_24_ ( .D(
        n78194), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[24]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_24_ ( .D(n1609), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1608) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_24_ ( 
        .D(n9615), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1606) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_24_ ( 
        .D(n78376), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_24_) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_24_ ( .D(n1603), .CLK(clk_i), 
        .QN(dbg_dat_o[24]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_24_ ( 
        .D(n9646), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1602) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_24_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_), .CLK(clk_i), 
        .QN(n1600) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_div_zero_o_reg ( .D(
        n1597), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_dbz) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o_reg_1_ ( 
        .D(n78374), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_exp_o_reg_1_ ( 
        .D(n27713), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_25_ ( 
        .D(n1594), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_25_ ( 
        .D(n1593), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_25_ ( .D(
        n78193), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[25]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_25_ ( .D(n1591), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1590) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_25_ ( 
        .D(n9614), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1588) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_25_ ( 
        .D(n78379), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_25_) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_25_ ( .D(n52474), .CLK(clk_i), 
        .QN(dbg_dat_o[25]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_25_ ( 
        .D(n9645), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1584) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_25_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_), .CLK(clk_i), 
        .QN(n1582) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r_reg_2_ ( 
        .D(n1580), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o_reg_2_ ( 
        .D(n78377), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_exp_o_reg_2_ ( 
        .D(n27721), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_26_ ( 
        .D(n1577), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_26_ ( 
        .D(n1576), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_26_ ( .D(
        n78192), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[26]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_wbmux_muxreg_reg_26_ ( .D(n1574), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1573) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_b_reg_26_ ( 
        .D(n9613), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1571) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_reg_26_ ( 
        .D(n78370), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_26_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_26_ ( 
        .D(n1568), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_26_ ( .D(n1567), .CLK(clk_i), 
        .QN(dbg_dat_o[26]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_operandmuxes_operand_a_reg_26_ ( 
        .D(n9644), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1566) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_26_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_), .CLK(clk_i), 
        .QN(n1564) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_ine_o_reg ( 
        .D(n1562), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_ine) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_ine_o_reg ( .D(n1561), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_ine_o) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_ine_o_reg ( .D(n27728), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_ine) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o_reg_3_ ( 
        .D(n1558), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_exp_o_reg_3_ ( 
        .D(n27729), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o_reg_4_ ( 
        .D(n78358), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_exp_o_reg_4_ ( 
        .D(n27731), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_28_ ( 
        .D(n1553), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[28]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_29_ ( 
        .D(n1552), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[29]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_output_o_reg_30_ ( 
        .D(n1551), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[30]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o_reg_5_ ( 
        .D(n78359), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_exp_o_reg_5_ ( 
        .D(n27733), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fractb_28_o_reg_0_ ( 
        .D(n1547), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_0_ ( 
        .D(n1546), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_fracta_28_o_reg_26_ ( 
        .D(n1543), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o_reg_6_ ( 
        .D(n78223), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_exp_o_reg_6_ ( 
        .D(n27735), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_30_ ( 
        .D(n1540), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[30]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_output1_reg_30_ ( 
        .D(n1539), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[30]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_30_ ( .D(
        n78191), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[30]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_qnan_o_reg ( .D(n1537), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_qnan) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_6_ ( .D(n9487), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1536) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_overflow_o_reg ( .D(
        n1534), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_overflow) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_3_ ( .D(n9490), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1533) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_underflow_o_reg ( .D(
        n1531), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_underflow) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o_reg_7_ ( 
        .D(n78224), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_exp_o_reg_7_ ( 
        .D(n27738), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_a_is_qnan_reg ( .D(n1523), .CLK(
        clk_i), .QN(or1200_cpu_or1200_fpu_a_is_qnan) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_output_o_reg_22_ ( 
        .D(n1522), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_snan_r_a_reg ( 
        .D(n1521), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_snan_r_a) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_snan_reg ( 
        .D(n27100), .CLK(clk_i), .QN(n1520) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_4_ ( .D(n9489), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1519) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_zero_reg ( .D(
        n1517), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_zero_conv) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_snan_reg ( .D(
        n1516), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_snan_conv) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_a_is_zero_reg ( .D(n53614), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_a_is_zero) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_a_is_snan_reg ( .D(n1514), .CLK(
        clk_i), .QN(or1200_cpu_or1200_fpu_a_is_snan) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_a_is_inf_reg ( .D(n58420), .CLK(
        clk_i), .QN(or1200_cpu_or1200_fpu_a_is_inf) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_b_is_inf_reg ( .D(n1512), .CLK(
        clk_i), .QN(or1200_cpu_or1200_fpu_b_is_inf) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_23_ ( .D(
        n1511), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[23]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dmr1_reg_22_ ( .D(n9327), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1510) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_du_dbg_bp_r_reg ( .D(or1200_du_N76), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1508) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_b_is_snan_reg ( .D(n1506), .CLK(
        clk_i), .QN(or1200_cpu_or1200_fpu_b_is_snan) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_22_ ( .D(n1505), .CLK(clk_i), 
        .QN(dbg_dat_o[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_b_is_qnan_reg ( .D(n1504), .CLK(
        clk_i), .QN(or1200_cpu_or1200_fpu_b_is_qnan) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_b_is_zero_reg ( .D(n78170), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_b_is_zero) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_zero_o_reg ( .D(n1502), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_zero) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_output_o_reg_31_ ( .D(
        n1501), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_arith[31]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_snan_o_reg ( .D(n74772), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_snan) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_5_ ( .D(n9488), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1499) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_inf_o_reg ( .D(n1497), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_inf) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_10_ ( .D(n52469), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1496) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_freeze_waiting_on_reg_0_ ( .D(
        n9671), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1494) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_freeze_waiting_on_reg_1_ ( .D(
        n9672), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1492) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_a_b_sign_xor_reg ( .D(n78182), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_a_b_sign_xor) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_9_ ( .D(n9484), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1489) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_23_ ( .D(n1487), .CLK(clk_i), 
        .QN(dbg_dat_o[23]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_0_ ( .D(n9307), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1486) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_1_ ( .D(n9306), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1484) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_2_ ( .D(n9305), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1482) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_3_ ( .D(n9304), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1480) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_4_ ( .D(n9303), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1478) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_5_ ( .D(n9302), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1476) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_6_ ( .D(n9301), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1474) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_7_ ( .D(n9300), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1472) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_8_ ( .D(n9299), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1470) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_9_ ( .D(n9298), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1468) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_10_ ( .D(n9297), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1466) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_11_ ( .D(n9296), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1464) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_12_ ( .D(n9295), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1462) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_13_ ( .D(n9294), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1460) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_14_ ( .D(n9293), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1458) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_15_ ( .D(n9292), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1456) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_16_ ( .D(n9291), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1454) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_17_ ( .D(n9290), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1452) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_18_ ( .D(n9289), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1450) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_19_ ( .D(n9288), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1448) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_20_ ( .D(n9287), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1446) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_21_ ( .D(n9286), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1444) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_22_ ( .D(n9285), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1442) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_23_ ( .D(n9284), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1440) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_24_ ( .D(n9283), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1438) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_25_ ( .D(n9282), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1436) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_26_ ( .D(n9281), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1434) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_27_ ( .D(n9280), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1432) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_29_ ( .D(n9279), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1430) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_30_ ( .D(n9278), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1428) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_31_ ( .D(n9277), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1426) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_0_ ( .D(or1200_pic_N47), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1424) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_1_ ( .D(or1200_pic_N48), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1422) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_2_ ( .D(n9325), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1420) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_2_ ( .D(or1200_pic_N49), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1418) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_3_ ( .D(n9324), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1416) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_3_ ( .D(or1200_pic_N50), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1414) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_4_ ( .D(n9323), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1412) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_4_ ( .D(or1200_pic_N51), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1410) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_5_ ( .D(n9322), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1408) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_5_ ( .D(or1200_pic_N52), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1406) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_6_ ( .D(n9321), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1404) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_6_ ( .D(or1200_pic_N53), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1402) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_7_ ( .D(n9320), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1400) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_7_ ( .D(or1200_pic_N54), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1398) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_8_ ( .D(n9319), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1396) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_8_ ( .D(or1200_pic_N55), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1394) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_9_ ( .D(n9318), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1392) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_9_ ( .D(or1200_pic_N56), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1390) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_10_ ( .D(n9317), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1388) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_10_ ( .D(or1200_pic_N57), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1386) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_11_ ( .D(n9316), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1384) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_12_ ( .D(n9315), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1382) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_12_ ( .D(or1200_pic_N59), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1380) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_13_ ( .D(n9314), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1378) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_13_ ( .D(or1200_pic_N60), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1376) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_14_ ( .D(n9313), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1374) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_14_ ( .D(or1200_pic_N61), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1372) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_15_ ( .D(n9312), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1370) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_15_ ( .D(or1200_pic_N62), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1368) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_16_ ( .D(n9311), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1366) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_16_ ( .D(or1200_pic_N63), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1364) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_17_ ( .D(n9310), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1362) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_17_ ( .D(or1200_pic_N64), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1360) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_18_ ( .D(n9309), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1358) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_18_ ( .D(or1200_pic_N65), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1356) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picmr_reg_19_ ( .D(n1353), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(or1200_pic_picmr_19_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_19_ ( .D(or1200_pic_N66), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1352) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_we_o_reg ( .D(n1350), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1349) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_biu_stb_reg_reg ( .D(dwb_biu_N62), .CLK(
        clk_i), .RESET(n53192), .SET(rst_i), .QN(n1347) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_2_ ( .D(
        n9346), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1345) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_3_ ( .D(
        n9345), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1343) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_cyc_o_reg ( .D(n78265), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1341) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_2_ ( .D(n9343), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1339) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_3_ ( .D(n9342), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1337) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_4_ ( .D(
        n9348), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1335) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_4_ ( .D(n1333), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1332) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_5_ ( .D(
        n9355), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1330) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_5_ ( .D(n1328), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1327) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_6_ ( .D(
        n9354), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1325) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_6_ ( .D(n1323), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1322) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_7_ ( .D(
        n9353), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1320) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_7_ ( .D(n1318), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1317) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_8_ ( .D(
        n9352), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1315) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_8_ ( .D(n1313), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1312) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_9_ ( .D(
        n9351), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1310) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_9_ ( .D(n1308), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1307) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_10_ ( .D(
        n9350), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1305) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_10_ ( .D(n1303), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1302) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_11_ ( .D(
        n9349), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1300) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_11_ ( .D(n1298), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1297) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_0_ ( .D(
        n9377), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1295) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_0_ ( .D(n1293), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1292) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_1_ ( .D(
        n9376), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1290) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_1_ ( .D(n1288), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1287) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_12_ ( .D(
        n9375), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1285) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_12_ ( .D(n58610), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1282) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_13_ ( .D(
        n9374), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1280) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_13_ ( .D(n1278), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1277) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_14_ ( .D(
        n9373), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1275) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_14_ ( .D(n58602), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1272) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_15_ ( .D(
        n9372), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1270) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_15_ ( .D(n58594), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1267) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_16_ ( .D(
        n9371), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1265) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_16_ ( .D(n1263), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1262) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_17_ ( .D(
        n9370), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1260) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_17_ ( .D(n58596), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1257) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_18_ ( .D(
        n9369), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1255) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_18_ ( .D(n1253), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1252) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_19_ ( .D(
        n9368), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1250) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_19_ ( .D(n58590), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1247) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_20_ ( .D(
        n9367), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1245) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_20_ ( .D(n58586), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1242) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_21_ ( .D(
        n9366), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1240) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_21_ ( .D(n1238), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1237) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_22_ ( .D(
        n9365), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1235) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_22_ ( .D(n58605), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1232) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_23_ ( .D(
        n9364), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1230) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_23_ ( .D(n58603), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1227) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_24_ ( .D(
        n9363), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1225) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_24_ ( .D(n1223), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1222) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_25_ ( .D(
        n9362), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1220) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_25_ ( .D(n58593), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1217) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_26_ ( .D(
        n9361), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1215) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_26_ ( .D(n58580), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1212) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_27_ ( .D(
        n9360), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1210) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_27_ ( .D(n58584), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1207) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_28_ ( .D(
        n9359), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1205) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_28_ ( .D(n58581), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1202) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_29_ ( .D(
        n9358), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1200) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_29_ ( .D(n58585), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1197) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_30_ ( .D(
        n9357), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1195) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_30_ ( .D(n1193), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1192) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_addr_r_reg_31_ ( .D(
        n9356), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1190) );
  ASYNC_DFFHx1_ASAP7_75t_SL dwb_biu_wb_adr_o_reg_31_ ( .D(n1188), .CLK(clk_i), 
        .RESET(n53192), .SET(dwb_rst_i), .QN(n1187) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_dc_top_or1200_dc_fsm_cache_miss_reg ( .D(
        n9380), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1185) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_11_ ( .D(n9264), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1183) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttmr_reg_28_ ( .D(n9244), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1181) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_0_ ( .D(n9275), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1179) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_1_ ( .D(n9274), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1177) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_2_ ( .D(n9273), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1175) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_3_ ( .D(n9272), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1173) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_4_ ( .D(n9271), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1171) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_5_ ( .D(n9270), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1169) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_6_ ( .D(n9269), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1167) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_7_ ( .D(n9268), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1165) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_8_ ( .D(n9267), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1163) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_9_ ( .D(n9266), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1161) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_10_ ( .D(n9265), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1159) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_12_ ( .D(n9263), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1157) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_13_ ( .D(n9262), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1155) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_14_ ( .D(n9261), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1153) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_15_ ( .D(n9260), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1151) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_16_ ( .D(n9259), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1149) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_17_ ( .D(n9258), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1147) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_18_ ( .D(n9257), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1145) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_19_ ( .D(n9256), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1143) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_20_ ( .D(n9255), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1141) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_21_ ( .D(n9254), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1139) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_22_ ( .D(n9253), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1137) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_23_ ( .D(n9252), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1135) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_24_ ( .D(n9251), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1133) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_25_ ( .D(n9250), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1131) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_26_ ( .D(n9249), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1129) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_27_ ( .D(n9276), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1127) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_28_ ( .D(n9248), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1125) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_29_ ( .D(n9247), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1123) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_30_ ( .D(n9246), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1121) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_tt_ttcr_reg_31_ ( .D(n9245), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(n1119) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_sprs_sr_reg_reg_11_ ( .D(
        or1200_cpu_to_sr[11]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1117) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_pic_picsr_reg_11_ ( .D(or1200_pic_N58), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1115) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_11_ ( .D(n1113), .CLK(clk_i), 
        .QN(dbg_dat_o[11]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_11_ ( .D(n9706), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1112) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_11_ ( .D(
        or1200_immu_top_N14), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1110) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_11_ ( .D(n9413), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1108) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_11_ ( 
        .D(n9185), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1106) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_10_ ( 
        .D(n9699), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1104) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_10_ ( .D(n1102), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1101) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_10_ ( .D(
        or1200_immu_top_N13), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1099) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_10_ ( .D(n9414), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1097) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_10_ ( 
        .D(n9186), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1095) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_9_ ( 
        .D(n9700), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1093) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_9_ ( .D(n1091), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1090) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_9_ ( .D(
        or1200_immu_top_N12), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1088) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_9_ ( .D(n9415), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1086) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_9_ ( .D(
        n9187), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1084) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_8_ ( 
        .D(n9701), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1082) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_8_ ( .D(n1080), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1079) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_8_ ( .D(n1076), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_immu_top_icpu_adr_default_8_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_8_ ( .D(n9416), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1075) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_8_ ( .D(
        n9188), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1073) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_7_ ( 
        .D(n9702), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1071) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_7_ ( .D(n1069), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1068) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_7_ ( .D(
        or1200_immu_top_N10), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1066) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_7_ ( .D(n9417), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1064) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_7_ ( .D(
        n1061), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_genpc_pcreg_default[7]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_6_ ( 
        .D(n9703), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1060) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_6_ ( .D(n1058), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1057) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_6_ ( .D(
        or1200_immu_top_N9), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1055) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_6_ ( .D(n9418), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1053) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_6_ ( .D(
        n1050), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_genpc_pcreg_default[6]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_5_ ( 
        .D(n9704), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1049) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_5_ ( .D(n1047), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1046) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_5_ ( .D(
        or1200_immu_top_N8), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1044) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_5_ ( .D(n9419), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1042) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_5_ ( .D(
        n1039), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_genpc_pcreg_default[5]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_4_ ( 
        .D(n9705), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1038) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_4_ ( .D(n1036), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1035) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_4_ ( .D(
        or1200_immu_top_N7), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1033) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_4_ ( .D(n9420), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1031) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_4_ ( .D(
        n1028), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_genpc_pcreg_default[4]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_31_ ( .D(
        or1200_immu_top_N34), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1027) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_31_ ( 
        .D(n9678), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1025) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_31_ ( .D(n1023), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1022) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_31_ ( .D(n9393), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1020) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_30_ ( .D(
        or1200_immu_top_N33), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n1018) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_30_ ( 
        .D(n9679), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1016) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_30_ ( .D(n1014), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1013) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_30_ ( .D(n9394), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1011) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_29_ ( .D(
        n51954), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1009) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_29_ ( 
        .D(n9680), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1007) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_29_ ( .D(n58562), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n1004) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_29_ ( .D(n9395), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1002) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_28_ ( .D(
        n51953), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n1000) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_28_ ( 
        .D(n9681), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n998) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_28_ ( .D(n58564), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n995) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_28_ ( .D(n9396), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n993) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_27_ ( .D(
        or1200_immu_top_N30), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n991) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_27_ ( 
        .D(n9682), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n989) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_27_ ( .D(n58563), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n986) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_27_ ( .D(n9397), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n984) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_26_ ( .D(
        or1200_immu_top_N29), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n982) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_26_ ( 
        .D(n9683), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n980) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_26_ ( .D(n978), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n977) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_26_ ( .D(n9398), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n975) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_25_ ( .D(
        n51952), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n973) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_25_ ( 
        .D(n9684), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n971) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_25_ ( .D(n58561), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n968) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_25_ ( .D(n9399), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n966) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_24_ ( .D(
        or1200_immu_top_N27), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n964) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_24_ ( 
        .D(n9685), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n962) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_24_ ( .D(n960), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n959) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_24_ ( .D(n9400), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n957) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_23_ ( .D(
        or1200_immu_top_N26), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n955) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_23_ ( 
        .D(n9686), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n953) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_23_ ( .D(n951), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n950) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_23_ ( .D(n9401), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n948) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_22_ ( .D(
        or1200_immu_top_N25), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n946) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_22_ ( 
        .D(n9687), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n944) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_22_ ( .D(n942), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n941) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_22_ ( .D(n9402), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n939) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_21_ ( .D(
        or1200_immu_top_N24), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n937) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_21_ ( 
        .D(n9688), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n935) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_21_ ( .D(n933), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n932) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_21_ ( .D(n9403), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n930) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_20_ ( .D(
        n51951), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n928) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_20_ ( 
        .D(n9689), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n926) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_20_ ( .D(n924), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n923) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_20_ ( .D(n9404), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n921) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_19_ ( .D(
        n51950), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n919) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_19_ ( 
        .D(n9690), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n917) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_19_ ( .D(n915), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n914) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_19_ ( .D(n9405), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n912) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_18_ ( .D(
        or1200_immu_top_N21), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n910) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_18_ ( 
        .D(n9691), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n908) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_18_ ( .D(n906), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n905) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_18_ ( .D(n9406), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n903) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_17_ ( .D(
        or1200_immu_top_N20), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n901) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_17_ ( 
        .D(n9692), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n899) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_17_ ( .D(n897), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n896) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_17_ ( .D(n9407), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n894) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_16_ ( .D(
        n51949), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n892) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_16_ ( 
        .D(n9693), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n890) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_16_ ( .D(n888), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n887) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_16_ ( .D(n9408), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n885) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_15_ ( .D(
        n51948), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n883) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_15_ ( 
        .D(n9694), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n881) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_15_ ( .D(n879), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n878) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_15_ ( .D(n9409), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n876) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_14_ ( .D(
        n51947), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n874) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_14_ ( 
        .D(n9695), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n872) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_14_ ( .D(n870), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n869) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_14_ ( .D(n9410), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n867) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_13_ ( .D(
        n51946), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n865) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_13_ ( 
        .D(n9696), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n863) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_13_ ( .D(n861), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n860) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_13_ ( .D(n9411), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n858) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_12_ ( .D(
        or1200_immu_top_N15), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n856) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_12_ ( .D(n9412), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n854) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_12_ ( 
        .D(n9697), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n852) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_12_ ( .D(n850), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n849) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_12_ ( 
        .D(n9184), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n847) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_3_ ( .D(
        or1200_immu_top_N6), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n845) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_3_ ( .D(n9421), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n843) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_3_ ( .D(
        n840), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_genpc_pcreg_default[3]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_adr_default_reg_2_ ( .D(
        or1200_immu_top_N5), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n839) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_if_addr_saved_reg_2_ ( .D(n9422), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n837) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_2_ ( 
        .D(n9473), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n835) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_2_ ( .D(n9469), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n833) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_ic_top_or1200_ic_fsm_saved_addr_r_reg_3_ ( 
        .D(n9472), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n831) );
  ASYNC_DFFHx1_ASAP7_75t_SL iwb_biu_wb_adr_o_reg_3_ ( .D(n77806), .CLK(clk_i), 
        .RESET(n53192), .SET(iwb_rst_i), .QN(n829) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_2_ ( .D(
        n826), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_genpc_pcreg_default[2]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_13_ ( 
        .D(n9183), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n823) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_14_ ( .D(
        icqmem_adr_qmem[14]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n821) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_14_ ( 
        .D(n9182), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n819) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_15_ ( .D(
        icqmem_adr_qmem[15]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n817) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_15_ ( 
        .D(n9181), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n815) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_16_ ( .D(
        icqmem_adr_qmem[16]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n813) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_16_ ( 
        .D(n9180), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n811) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_17_ ( .D(
        icqmem_adr_qmem[17]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n809) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_17_ ( 
        .D(n9179), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n807) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_18_ ( .D(
        icqmem_adr_qmem[18]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n805) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_18_ ( 
        .D(n9178), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n803) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_19_ ( .D(
        icqmem_adr_qmem[19]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n801) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_19_ ( 
        .D(n9177), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n799) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_20_ ( .D(
        icqmem_adr_qmem[20]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n797) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_20_ ( 
        .D(n9176), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n795) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_21_ ( 
        .D(n9175), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n791) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_22_ ( .D(
        icqmem_adr_qmem[22]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n789) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_22_ ( 
        .D(n9174), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n787) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_23_ ( .D(
        icqmem_adr_qmem[23]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n785) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_23_ ( 
        .D(n9173), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n783) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_24_ ( .D(
        icqmem_adr_qmem[24]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n781) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_24_ ( 
        .D(n9172), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n779) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_25_ ( .D(
        icqmem_adr_qmem[25]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n777) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_25_ ( 
        .D(n9171), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n775) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_26_ ( .D(
        icqmem_adr_qmem[26]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n773) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_26_ ( 
        .D(n9170), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n771) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_27_ ( 
        .D(n9169), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n767) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_28_ ( .D(
        icqmem_adr_qmem[28]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n765) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_28_ ( 
        .D(n9168), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n763) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_29_ ( 
        .D(n9167), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n759) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_30_ ( .D(
        icqmem_adr_qmem[30]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n757) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_30_ ( 
        .D(n9166), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n755) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_immu_top_icpu_vpn_r_reg_31_ ( .D(
        icqmem_adr_qmem[31]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n753) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_genpc_pcreg_default_reg_31_ ( 
        .D(n9165), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n751) );
  DFFHQNx1_ASAP7_75t_SL or1200_du_dbg_dat_o_reg_7_ ( .D(n749), .CLK(clk_i), 
        .QN(dbg_dat_o[7]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpcsr_r_reg_7_ ( .D(n9486), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(n748) );
  INVx1_ASAP7_75t_SL U150 ( .A(n3418), .Y(dc_en) );
  A2O1A1Ixp33_ASAP7_75t_SL U464 ( .A1(n57189), .A2(n53628), .B(n4134), .C(n235), .Y(icbiu_adr_ic_word[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1102 ( .A1(n3918), .A2(n3917), .B(n53192), .C(
        n53628), .Y(sbbiu_adr_sb[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1109 ( .A1(n3916), .A2(n3915), .B(n53192), .C(
        n53628), .Y(sbbiu_adr_sb[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1116 ( .A1(n3914), .A2(n3913), .B(n53192), .C(
        n53628), .Y(sbbiu_adr_sb[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1123 ( .A1(n3912), .A2(n3911), .B(n53192), .C(
        n53628), .Y(sbbiu_adr_sb[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1130 ( .A1(n3910), .A2(n3909), .B(n53192), .C(
        n53628), .Y(sbbiu_adr_sb[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1137 ( .A1(n3908), .A2(n3907), .B(n53192), .C(
        n53628), .Y(sbbiu_adr_sb[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1144 ( .A1(n3923), .A2(n3922), .B(n53192), .C(
        n53628), .Y(sbbiu_adr_sb[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1151 ( .A1(n3921), .A2(n3920), .B(n53192), .C(
        n53628), .Y(sbbiu_adr_sb[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1166 ( .A1(n4317), .A2(n4318), .B(n1285), .C(n527), 
        .Y(sbbiu_adr_sb[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1172 ( .A1(n4317), .A2(n4318), .B(n1280), .C(n529), 
        .Y(sbbiu_adr_sb[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1178 ( .A1(n4317), .A2(n4318), .B(n1275), .C(n531), 
        .Y(sbbiu_adr_sb[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1184 ( .A1(n4317), .A2(n4318), .B(n1270), .C(n533), 
        .Y(sbbiu_adr_sb[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1190 ( .A1(n4317), .A2(n4318), .B(n1265), .C(n535), 
        .Y(sbbiu_adr_sb[16]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1196 ( .A1(n4317), .A2(n4318), .B(n1260), .C(n537), 
        .Y(sbbiu_adr_sb[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1202 ( .A1(n4317), .A2(n4318), .B(n1255), .C(n539), 
        .Y(sbbiu_adr_sb[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1208 ( .A1(n4317), .A2(n4318), .B(n1250), .C(n541), 
        .Y(sbbiu_adr_sb[19]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1214 ( .A1(n4317), .A2(n4318), .B(n1245), .C(n543), 
        .Y(sbbiu_adr_sb[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1220 ( .A1(n4317), .A2(n4318), .B(n1240), .C(n545), 
        .Y(sbbiu_adr_sb[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1226 ( .A1(n4317), .A2(n4318), .B(n1235), .C(n547), 
        .Y(sbbiu_adr_sb[22]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1232 ( .A1(n4317), .A2(n4318), .B(n1230), .C(n549), 
        .Y(sbbiu_adr_sb[23]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1238 ( .A1(n4317), .A2(n4318), .B(n1225), .C(n551), 
        .Y(sbbiu_adr_sb[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1244 ( .A1(n4317), .A2(n4318), .B(n1220), .C(n553), 
        .Y(sbbiu_adr_sb[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1250 ( .A1(n4317), .A2(n4318), .B(n1215), .C(n555), 
        .Y(sbbiu_adr_sb[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1256 ( .A1(n4317), .A2(n4318), .B(n1210), .C(n557), 
        .Y(sbbiu_adr_sb[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1262 ( .A1(n4317), .A2(n4318), .B(n1205), .C(n559), 
        .Y(sbbiu_adr_sb[28]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1268 ( .A1(n4317), .A2(n4318), .B(n1200), .C(n561), 
        .Y(sbbiu_adr_sb[29]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1274 ( .A1(n4317), .A2(n4318), .B(n1195), .C(n563), 
        .Y(sbbiu_adr_sb[30]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1280 ( .A1(n4317), .A2(n4318), .B(n1190), .C(n565), 
        .Y(sbbiu_adr_sb[31]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1295 ( .A1(n57189), .A2(n53628), .B(n4135), .C(
        n572), .Y(icbiu_adr_ic_word[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1309 ( .A1(n57189), .A2(n53628), .B(n4136), .C(
        n579), .Y(icbiu_adr_ic_word[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1329 ( .A1(n57189), .A2(n53628), .B(n78056), .C(
        n589), .Y(icbiu_adr_ic_word[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1343 ( .A1(n57189), .A2(n53628), .B(n4138), .C(
        n596), .Y(icbiu_adr_ic_word[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1357 ( .A1(n57189), .A2(n53628), .B(n4089), .C(
        n603), .Y(icbiu_adr_ic_word[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1371 ( .A1(n57189), .A2(n53628), .B(n4090), .C(
        n610), .Y(icbiu_adr_ic_word[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1385 ( .A1(n57189), .A2(n53628), .B(n4091), .C(
        n617), .Y(icbiu_adr_ic_word[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1407 ( .A1(n4095), .A2(n78183), .B(n57189), .C(
        n626), .Y(icbiu_adr_ic_word[31]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1422 ( .A1(n4097), .A2(n78185), .B(n57189), .C(
        n631), .Y(icbiu_adr_ic_word[30]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1438 ( .A1(n78208), .A2(n4099), .B(n57189), .C(
        n636), .Y(icbiu_adr_ic_word[29]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1453 ( .A1(n4101), .A2(n78262), .B(n57189), .C(
        n643), .Y(icbiu_adr_ic_word[28]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1468 ( .A1(n4103), .A2(n78204), .B(n57189), .C(
        n648), .Y(icbiu_adr_ic_word[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1483 ( .A1(n4106), .A2(n78207), .B(n57189), .C(
        n653), .Y(icbiu_adr_ic_word[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1498 ( .A1(n4108), .A2(n78206), .B(n57189), .C(
        n658), .Y(icbiu_adr_ic_word[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1513 ( .A1(n4110), .A2(n78205), .B(n57189), .C(
        n663), .Y(icbiu_adr_ic_word[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1528 ( .A1(n4112), .A2(n78263), .B(n57189), .C(
        n668), .Y(icbiu_adr_ic_word[23]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1543 ( .A1(n4114), .A2(n78252), .B(n57189), .C(
        n673), .Y(icbiu_adr_ic_word[22]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1558 ( .A1(n4116), .A2(n78259), .B(n57189), .C(
        n678), .Y(icbiu_adr_ic_word[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1573 ( .A1(n4118), .A2(n78258), .B(n57189), .C(
        n683), .Y(icbiu_adr_ic_word[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1588 ( .A1(n4120), .A2(n78188), .B(n57189), .C(
        n688), .Y(icbiu_adr_ic_word[19]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1603 ( .A1(n4122), .A2(n78257), .B(n57189), .C(
        n693), .Y(icbiu_adr_ic_word[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1618 ( .A1(n4124), .A2(n78256), .B(n57189), .C(
        n698), .Y(icbiu_adr_ic_word[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1633 ( .A1(n4126), .A2(n78255), .B(n57189), .C(
        n703), .Y(icbiu_adr_ic_word[16]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1648 ( .A1(n4128), .A2(n78254), .B(n57189), .C(
        n708), .Y(icbiu_adr_ic_word[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1663 ( .A1(n4130), .A2(n78261), .B(n57189), .C(
        n713), .Y(icbiu_adr_ic_word[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1678 ( .A1(n4132), .A2(n78264), .B(n57189), .C(
        n720), .Y(icbiu_adr_ic_word[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U1692 ( .A1(n57189), .A2(n53628), .B(n4133), .C(
        n727), .Y(icbiu_adr_ic_word[12]) );
  NAND3xp33_ASAP7_75t_SL U8647 ( .A(n7636), .B(n7637), .C(n7635), .Y(
        or1200_cpu_rf_addrb[0]) );
  NAND3xp33_ASAP7_75t_SL U8651 ( .A(n7631), .B(n7632), .C(n7630), .Y(
        or1200_cpu_rf_addrb[1]) );
  NAND3xp33_ASAP7_75t_SL U8655 ( .A(n7626), .B(n7627), .C(n7625), .Y(
        or1200_cpu_rf_addrb[2]) );
  NAND3xp33_ASAP7_75t_SL U8659 ( .A(n7621), .B(n7622), .C(n7620), .Y(
        or1200_cpu_rf_addrb[3]) );
  NAND3xp33_ASAP7_75t_SL U8663 ( .A(n7616), .B(n7617), .C(n7615), .Y(
        or1200_cpu_rf_addrb[4]) );
  OAI21xp33_ASAP7_75t_SL U8699 ( .A1(n4092), .A2(n57189), .B(n7192), .Y(
        icbiu_adr_ic_word[3]) );
  NAND2xp33_ASAP7_75t_SL U9405 ( .A(n4304), .B(n4305), .Y(
        or1200_dc_top_to_dcram[0]) );
  NAND2xp33_ASAP7_75t_SL U9408 ( .A(n4273), .B(n4274), .Y(
        or1200_dc_top_to_dcram[1]) );
  NAND2xp33_ASAP7_75t_SL U9411 ( .A(n4244), .B(n4245), .Y(
        or1200_dc_top_to_dcram[2]) );
  NAND2xp33_ASAP7_75t_SL U9414 ( .A(n4238), .B(n4239), .Y(
        or1200_dc_top_to_dcram[3]) );
  NAND2xp33_ASAP7_75t_SL U9417 ( .A(n4236), .B(n4237), .Y(
        or1200_dc_top_to_dcram[4]) );
  NAND2xp33_ASAP7_75t_SL U9420 ( .A(n4234), .B(n4235), .Y(
        or1200_dc_top_to_dcram[5]) );
  NAND2xp33_ASAP7_75t_SL U9423 ( .A(n4232), .B(n4233), .Y(
        or1200_dc_top_to_dcram[6]) );
  NAND2xp33_ASAP7_75t_SL U9426 ( .A(n4230), .B(n4231), .Y(
        or1200_dc_top_to_dcram[7]) );
  OAI21xp33_ASAP7_75t_SL U9435 ( .A1(n59696), .A2(n4302), .B(n4303), .Y(
        or1200_dc_top_to_dcram[10]) );
  OAI21xp33_ASAP7_75t_SL U9475 ( .A1(n59696), .A2(n4265), .B(n4266), .Y(
        or1200_dc_top_to_dcram[22]) );
  OAI21xp33_ASAP7_75t_SL U9482 ( .A1(n59696), .A2(n4256), .B(n4257), .Y(
        or1200_dc_top_to_dcram[24]) );
  OAI21xp33_ASAP7_75t_SL U9488 ( .A1(n59696), .A2(n4254), .B(n4255), .Y(
        or1200_dc_top_to_dcram[25]) );
  OAI21xp33_ASAP7_75t_SL U9494 ( .A1(n59696), .A2(n4252), .B(n4253), .Y(
        or1200_dc_top_to_dcram[26]) );
  OAI21xp33_ASAP7_75t_SL U9500 ( .A1(n59696), .A2(n4250), .B(n4251), .Y(
        or1200_dc_top_to_dcram[27]) );
  OAI21xp33_ASAP7_75t_SL U9506 ( .A1(n59696), .A2(n4248), .B(n4249), .Y(
        or1200_dc_top_to_dcram[28]) );
  OAI21xp33_ASAP7_75t_SL U9512 ( .A1(n59696), .A2(n4246), .B(n4247), .Y(
        or1200_dc_top_to_dcram[29]) );
  OAI21xp33_ASAP7_75t_SL U9518 ( .A1(n59696), .A2(n4242), .B(n4243), .Y(
        or1200_dc_top_to_dcram[30]) );
  OAI21xp33_ASAP7_75t_SL U9525 ( .A1(n59696), .A2(n4240), .B(n4241), .Y(
        or1200_dc_top_to_dcram[31]) );
  OAI21xp33_ASAP7_75t_SL U9536 ( .A1(n78174), .A2(n3906), .B(n4320), .Y(
        or1200_dc_top_dcram_we[0]) );
  OAI21xp33_ASAP7_75t_SL U9540 ( .A1(n78174), .A2(n3905), .B(n4320), .Y(
        or1200_dc_top_dcram_we[1]) );
  OAI21xp33_ASAP7_75t_SL U9547 ( .A1(n78174), .A2(n3904), .B(n4320), .Y(
        or1200_dc_top_dcram_we[2]) );
  OAI21xp33_ASAP7_75t_SL U9550 ( .A1(n78174), .A2(n3903), .B(n4320), .Y(
        or1200_dc_top_dcram_we[3]) );
  NOR2xp33_ASAP7_75t_SL U9971 ( .A(n78176), .B(n4306), .Y(
        or1200_dc_top_dctag_v) );
  A2O1A1Ixp33_ASAP7_75t_SL U10143 ( .A1(n4049), .A2(n4050), .B(n4139), .C(
        n4140), .Y(or1200_ic_top_ictag_addr[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10144 ( .A1(n4053), .A2(n4054), .B(n4139), .C(
        n4141), .Y(or1200_ic_top_ictag_addr[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10145 ( .A1(n4057), .A2(n4058), .B(n4139), .C(
        n4142), .Y(or1200_ic_top_ictag_addr[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10146 ( .A1(n4061), .A2(n4062), .B(n4139), .C(
        n4143), .Y(or1200_ic_top_ictag_addr[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10147 ( .A1(n4066), .A2(n4067), .B(n4139), .C(
        n4144), .Y(or1200_ic_top_ictag_addr[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10148 ( .A1(n4070), .A2(n4071), .B(n4139), .C(
        n4145), .Y(or1200_ic_top_ictag_addr[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10149 ( .A1(n4041), .A2(n4042), .B(n4139), .C(
        n4146), .Y(or1200_ic_top_ictag_addr[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10150 ( .A1(n4045), .A2(n4046), .B(n4139), .C(
        n4147), .Y(or1200_ic_top_ictag_addr[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10159 ( .A1(n4224), .A2(n4225), .B(n59696), .C(
        n4226), .Y(or1200_dc_top_to_dcram[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10160 ( .A1(n4227), .A2(n4228), .B(n59696), .C(
        n4229), .Y(or1200_dc_top_to_dcram[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10161 ( .A1(n4262), .A2(n4263), .B(n59696), .C(
        n4264), .Y(or1200_dc_top_to_dcram[23]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10162 ( .A1(n4267), .A2(n4268), .B(n59696), .C(
        n4269), .Y(or1200_dc_top_to_dcram[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10163 ( .A1(n4270), .A2(n4271), .B(n59696), .C(
        n4272), .Y(or1200_dc_top_to_dcram[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10164 ( .A1(n4275), .A2(n4276), .B(n59696), .C(
        n4277), .Y(or1200_dc_top_to_dcram[19]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10165 ( .A1(n4278), .A2(n4279), .B(n59696), .C(
        n4280), .Y(or1200_dc_top_to_dcram[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10166 ( .A1(n4281), .A2(n4282), .B(n59696), .C(
        n4283), .Y(or1200_dc_top_to_dcram[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10167 ( .A1(n4284), .A2(n4285), .B(n59696), .C(
        n4286), .Y(or1200_dc_top_to_dcram[16]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10168 ( .A1(n4287), .A2(n4288), .B(n59696), .C(
        n4289), .Y(or1200_dc_top_to_dcram[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10169 ( .A1(n4290), .A2(n4291), .B(n59696), .C(
        n4292), .Y(or1200_dc_top_to_dcram[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10170 ( .A1(n4293), .A2(n4294), .B(n59696), .C(
        n4295), .Y(or1200_dc_top_to_dcram[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10171 ( .A1(n4296), .A2(n4297), .B(n59696), .C(
        n4298), .Y(or1200_dc_top_to_dcram[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10172 ( .A1(n4299), .A2(n4300), .B(n59696), .C(
        n4301), .Y(or1200_dc_top_to_dcram[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10173 ( .A1(n3907), .A2(n3908), .B(n78176), .C(
        n4309), .Y(or1200_dc_top_dctag_addr[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10174 ( .A1(n3909), .A2(n3910), .B(n78176), .C(
        n4310), .Y(or1200_dc_top_dctag_addr[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10175 ( .A1(n3911), .A2(n3912), .B(n78176), .C(
        n4311), .Y(or1200_dc_top_dctag_addr[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10176 ( .A1(n3913), .A2(n3914), .B(n78176), .C(
        n4312), .Y(or1200_dc_top_dctag_addr[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10177 ( .A1(n3915), .A2(n3916), .B(n78176), .C(
        n4313), .Y(or1200_dc_top_dctag_addr[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10178 ( .A1(n3917), .A2(n3918), .B(n78176), .C(
        n4314), .Y(or1200_dc_top_dctag_addr[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10179 ( .A1(n3920), .A2(n3921), .B(n78176), .C(
        n4315), .Y(or1200_dc_top_dctag_addr[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL U10180 ( .A1(n3922), .A2(n3923), .B(n78176), .C(
        n4316), .Y(or1200_dc_top_dctag_addr[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U195 ( .A1(
        or1200_cpu_or1200_rf_n145), .A2(or1200_cpu_or1200_rf_n144), .B(n53192), 
        .C(or1200_cpu_or1200_rf_n142), .Y(or1200_cpu_or1200_rf_rf_addra[0]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U194 ( .A1(
        or1200_cpu_or1200_rf_n141), .A2(or1200_cpu_or1200_rf_n140), .B(n53192), 
        .C(or1200_cpu_or1200_rf_n139), .Y(or1200_cpu_or1200_rf_rf_addra[1]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U193 ( .A1(
        or1200_cpu_or1200_rf_n138), .A2(or1200_cpu_or1200_rf_n137), .B(n53192), 
        .C(or1200_cpu_or1200_rf_n136), .Y(or1200_cpu_or1200_rf_rf_addra[2]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U192 ( .A1(
        or1200_cpu_or1200_rf_n135), .A2(or1200_cpu_or1200_rf_n134), .B(n53192), 
        .C(or1200_cpu_or1200_rf_n133), .Y(or1200_cpu_or1200_rf_rf_addra[3]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U191 ( .A1(
        or1200_cpu_or1200_rf_n132), .A2(or1200_cpu_or1200_rf_n131), .B(n53192), 
        .C(or1200_cpu_or1200_rf_n130), .Y(or1200_cpu_or1200_rf_rf_addra[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U189 ( .A1(
        or1200_cpu_or1200_rf_n129), .A2(or1200_cpu_or1200_rf_n128), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_addrw[0]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U188 ( .A1(
        or1200_cpu_or1200_rf_n125), .A2(or1200_cpu_or1200_rf_n124), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_addrw[1]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U187 ( .A1(
        or1200_cpu_or1200_rf_n123), .A2(or1200_cpu_or1200_rf_n122), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_addrw[2]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U186 ( .A1(
        or1200_cpu_or1200_rf_n121), .A2(or1200_cpu_or1200_rf_n120), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_addrw[3]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U185 ( .A1(
        or1200_cpu_or1200_rf_n119), .A2(or1200_cpu_or1200_rf_n118), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_addrw[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U182 ( .A1(
        or1200_cpu_or1200_rf_n117), .A2(or1200_cpu_or1200_rf_n116), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[0]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U181 ( .A1(
        or1200_cpu_or1200_rf_n113), .A2(or1200_cpu_or1200_rf_n112), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[1]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U180 ( .A1(
        or1200_cpu_or1200_rf_n111), .A2(or1200_cpu_or1200_rf_n110), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[2]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U179 ( .A1(
        or1200_cpu_or1200_rf_n109), .A2(or1200_cpu_or1200_rf_n108), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[3]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U178 ( .A1(
        or1200_cpu_or1200_rf_n107), .A2(or1200_cpu_or1200_rf_n106), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[4]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U177 ( .A1(
        or1200_cpu_or1200_rf_n105), .A2(or1200_cpu_or1200_rf_n104), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[5]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U176 ( .A1(
        or1200_cpu_or1200_rf_n103), .A2(or1200_cpu_or1200_rf_n102), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U175 ( .A1(
        or1200_cpu_or1200_rf_n101), .A2(or1200_cpu_or1200_rf_n100), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U174 ( .A1(
        or1200_cpu_or1200_rf_n99), .A2(or1200_cpu_or1200_rf_n98), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U173 ( .A1(
        or1200_cpu_or1200_rf_n97), .A2(or1200_cpu_or1200_rf_n96), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U172 ( .A1(
        or1200_cpu_or1200_rf_n95), .A2(or1200_cpu_or1200_rf_n94), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[10]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U171 ( .A1(
        or1200_cpu_or1200_rf_n93), .A2(or1200_cpu_or1200_rf_n92), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U170 ( .A1(
        or1200_cpu_or1200_rf_n91), .A2(or1200_cpu_or1200_rf_n90), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U169 ( .A1(
        or1200_cpu_or1200_rf_n89), .A2(or1200_cpu_or1200_rf_n88), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U168 ( .A1(
        or1200_cpu_or1200_rf_n87), .A2(or1200_cpu_or1200_rf_n86), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U167 ( .A1(
        or1200_cpu_or1200_rf_n85), .A2(or1200_cpu_or1200_rf_n84), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U166 ( .A1(
        or1200_cpu_or1200_rf_n83), .A2(or1200_cpu_or1200_rf_n82), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[16]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U165 ( .A1(
        or1200_cpu_or1200_rf_n81), .A2(or1200_cpu_or1200_rf_n80), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U164 ( .A1(
        or1200_cpu_or1200_rf_n79), .A2(or1200_cpu_or1200_rf_n78), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U163 ( .A1(
        or1200_cpu_or1200_rf_n77), .A2(or1200_cpu_or1200_rf_n76), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[19]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U162 ( .A1(
        or1200_cpu_or1200_rf_n75), .A2(or1200_cpu_or1200_rf_n74), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U161 ( .A1(
        or1200_cpu_or1200_rf_n73), .A2(or1200_cpu_or1200_rf_n72), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U160 ( .A1(
        or1200_cpu_or1200_rf_n71), .A2(or1200_cpu_or1200_rf_n70), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[22]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U159 ( .A1(
        or1200_cpu_or1200_rf_n69), .A2(or1200_cpu_or1200_rf_n68), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[23]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U158 ( .A1(
        or1200_cpu_or1200_rf_n67), .A2(or1200_cpu_or1200_rf_n66), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[24]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U157 ( .A1(
        or1200_cpu_or1200_rf_n65), .A2(or1200_cpu_or1200_rf_n64), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[25]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U156 ( .A1(
        or1200_cpu_or1200_rf_n63), .A2(or1200_cpu_or1200_rf_n62), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[26]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U155 ( .A1(
        or1200_cpu_or1200_rf_n61), .A2(or1200_cpu_or1200_rf_n60), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[27]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U154 ( .A1(
        or1200_cpu_or1200_rf_n59), .A2(or1200_cpu_or1200_rf_n58), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[28]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U153 ( .A1(
        or1200_cpu_or1200_rf_n57), .A2(or1200_cpu_or1200_rf_n56), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[29]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U152 ( .A1(
        or1200_cpu_or1200_rf_n55), .A2(or1200_cpu_or1200_rf_n54), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[30]) );
  A2O1A1Ixp33_ASAP7_75t_SL or1200_cpu_or1200_rf_U151 ( .A1(
        or1200_cpu_or1200_rf_n53), .A2(or1200_cpu_or1200_rf_n52), .B(n53192), 
        .C(n53628), .Y(or1200_cpu_or1200_rf_rf_dataw[31]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_rf_addra_last_reg_0_ ( .D(
        or1200_cpu_or1200_rf_n11), .CLK(clk_i), .QN(
        or1200_cpu_or1200_rf_addra_last_0_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_rf_rf_we_allow_reg ( .D(
        or1200_cpu_or1200_rf_n12), .CLK(clk_i), .RESET(n53192), .SET(rst_i), 
        .QN(or1200_cpu_or1200_rf_rf_we_allow) );
  AND2x2_ASAP7_75t_SL or1200_cpu_or1200_rf_C150 ( .A(or1200_cpu_or1200_rf_N31), 
        .B(or1200_cpu_or1200_rf_rf_we_allow), .Y(or1200_cpu_or1200_rf_rf_we)
         );
  OR2x2_ASAP7_75t_SL or1200_cpu_or1200_rf_C158 ( .A(or1200_cpu_or1200_rf_N36), 
        .B(n78177), .Y(or1200_cpu_or1200_rf_rf_ena) );
  tpram or1200_cpu_or1200_rf_rf_a ( .clock(clk_i), .rst(rst_i), .ce_a(
        or1200_cpu_or1200_rf_rf_ena), .addr_a(or1200_cpu_or1200_rf_rf_addra), 
        .do_a({or1200_cpu_spr_dat_rf, or1200_cpu_rf_dataa_0_}), .ce_b(
        or1200_cpu_or1200_rf_rf_enb), .addr_b(or1200_cpu_rf_addrb), .do_b(
        or1200_cpu_rf_datab), .ce_w(or1200_cpu_or1200_rf_rf_we), .we_w(
        or1200_cpu_or1200_rf_rf_we), .addr_w(or1200_cpu_or1200_rf_rf_addrw), 
        .di_w(or1200_cpu_or1200_rf_rf_dataw) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_63_ ( 
        .D(n78169), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n192) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_62_ ( 
        .D(n78172), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n190) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_61_ ( 
        .D(n78168), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n188) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_60_ ( 
        .D(n51985), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n186) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_59_ ( 
        .D(n51986), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n184) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_58_ ( 
        .D(n51987), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n182) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_57_ ( 
        .D(n51988), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n180) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_53_ ( 
        .D(n51999), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n172) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_52_ ( 
        .D(n52000), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n170) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_51_ ( 
        .D(n52008), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n168) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_50_ ( 
        .D(n52003), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n166) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_49_ ( 
        .D(n78171), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n164) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_48_ ( 
        .D(n52006), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n162) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_47_ ( 
        .D(n52011), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n160) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_46_ ( 
        .D(n52012), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n158) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_45_ ( 
        .D(n52004), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n156) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_43_ ( 
        .D(n52009), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n152) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_42_ ( 
        .D(n51998), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n150) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_41_ ( 
        .D(n51997), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n148) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_40_ ( 
        .D(n51990), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n146) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_39_ ( 
        .D(n51993), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n144) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_38_ ( 
        .D(n51996), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n142) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_37_ ( 
        .D(n51994), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n140) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_36_ ( 
        .D(n51995), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n138) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_35_ ( 
        .D(n51991), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n136) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_34_ ( 
        .D(n51992), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n134) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_33_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N34), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n132) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_32_ ( 
        .D(n52013), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n130) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_31_ ( 
        .D(n52014), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n128) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_30_ ( 
        .D(n52061), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n126) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_29_ ( 
        .D(n52060), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n124) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_28_ ( 
        .D(n52059), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n122) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_27_ ( 
        .D(n52058), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n120) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_26_ ( 
        .D(n52057), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n118) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_25_ ( 
        .D(n52056), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n116) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_24_ ( 
        .D(n52055), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n114) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_23_ ( 
        .D(n52053), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n112) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_22_ ( 
        .D(n52054), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n110) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_21_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N22), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n108) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_20_ ( 
        .D(n52052), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n106) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_19_ ( 
        .D(n52051), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n104) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_18_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N19), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n102) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_17_ ( 
        .D(n52050), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n100) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_16_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N17), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n98) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_15_ ( 
        .D(n52049), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n96) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_14_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N15), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n94) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_13_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N14), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n92) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_12_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N13), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n90) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_11_ ( 
        .D(n52048), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n88) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_10_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N11), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n86) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_9_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N10), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n84) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_8_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N9), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n82) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_7_ ( 
        .D(n63349), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n80) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_6_ ( 
        .D(n63295), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n78) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_5_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N6), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n76) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_4_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N5), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n74) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_3_ ( 
        .D(n58577), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n72) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_2_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N3), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n70) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_1_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_mult_x_1_n211), 
        .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n68) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_0_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N1), .CLK(clk_i), 
        .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n66) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_63_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n192), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[63]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_62_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n190), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[62]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_61_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n188), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[61]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_60_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n186), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[60]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_59_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n184), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[59]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_58_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n182), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[58]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_57_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n180), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[57]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_56_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n178), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[56]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_55_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n176), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[55]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_54_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n174), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[54]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_53_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n172), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[53]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_52_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n170), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[52]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_51_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n168), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[51]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_50_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n166), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[50]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_49_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n164), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[49]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_48_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n162), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[48]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_47_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n160), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[47]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_46_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n158), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[46]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_45_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n156), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[45]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_44_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n154), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[44]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_43_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n152), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[43]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_42_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n150), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[42]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_41_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n148), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[41]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_40_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n146), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[40]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_39_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n144), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[39]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_38_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n142), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[38]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_37_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n140), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[37]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_36_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n138), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[36]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_35_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n136), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[35]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_34_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n134), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[34]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_33_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n132), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[33]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_32_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n130), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[32]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_31_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n128), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[31]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_30_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n126), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[30]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_29_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n124), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[29]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_28_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n122), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[28]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_27_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n120), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[27]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_26_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n118), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[26]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_25_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n116), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[25]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_24_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n114), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[24]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_23_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n112), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[23]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_22_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n110), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[22]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_21_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n108), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[21]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_20_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n106), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[20]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_19_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n104), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[19]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_18_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n102), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[18]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_17_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n100), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[17]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_16_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n98), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[16]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_15_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n96), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[15]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_14_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n94), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[14]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_13_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n92), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[13]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_12_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n90), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[12]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_11_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n88), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[11]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_10_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n86), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[10]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_9_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n84), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[9]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_8_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n82), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[8]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_7_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n80), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[7]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_6_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n78), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[6]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_5_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n76), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[5]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_4_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n74), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[4]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_3_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n72), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[3]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_2_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n70), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[2]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_1_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n68), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p1_reg_0_ ( 
        .D(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n66), .CLK(clk_i), 
        .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_mult_mac_mul_prod[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_63_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1496), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n2) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_62_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1497), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n4) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_61_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1498), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n6) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_60_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1499), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n8) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_59_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1500), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n10) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_58_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1501), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n12) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_57_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1502), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n14) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_56_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1503), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n16) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_55_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1504), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n18) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_54_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1505), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n20) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_53_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1506), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n22) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_52_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1507), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n24) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_51_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1508), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n26) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_50_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1509), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n28) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_49_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1510), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n30) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_48_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1511), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n32) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_47_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1512), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n34) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_46_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1513), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n36) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_45_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1514), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n38) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_44_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1515), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n40) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_43_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1516), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n42) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_42_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1517), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n44) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_41_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1518), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n46) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_40_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1519), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n48) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_39_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1520), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n50) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_38_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1521), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n52) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_37_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1522), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n54) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_36_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1523), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n56) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_35_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1524), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n58) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_34_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1525), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n60) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_33_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1526), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n62) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_32_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1528), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n64) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_31_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1529), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n66) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_30_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1530), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n68) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_29_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1531), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n70) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_28_ ( 
        .D(n14253), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n72) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_27_ ( 
        .D(n14494), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n74) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_26_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1534), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n76) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_25_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1535), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n78) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_24_ ( 
        .D(n12980), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n80) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_23_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1537), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n82) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_22_ ( 
        .D(n12981), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n84) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_21_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1539), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n86) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_20_ ( 
        .D(n12986), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n88) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_19_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1541), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n90) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_18_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1542), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n92) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_17_ ( 
        .D(n14251), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n94) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_16_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1544), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n96) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_15_ ( 
        .D(n12970), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n98) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_14_ ( 
        .D(n14249), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n100) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_13_ ( 
        .D(n52047), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_n102) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_12_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1548), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n104) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_11_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1549), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n106) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_10_ ( 
        .D(or1200_cpu_or1200_mult_mac_n1550), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n108) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_9_ ( .D(
        or1200_cpu_or1200_mult_mac_n1551), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n110) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_8_ ( .D(
        or1200_cpu_or1200_mult_mac_n1552), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n112) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_7_ ( .D(
        or1200_cpu_or1200_mult_mac_n1553), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n114) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_6_ ( .D(
        or1200_cpu_or1200_mult_mac_n1554), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n116) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_5_ ( .D(
        or1200_cpu_or1200_mult_mac_n1555), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n118) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_4_ ( .D(
        or1200_cpu_or1200_mult_mac_n1556), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n120) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_3_ ( .D(
        or1200_cpu_or1200_mult_mac_n1557), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n122) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_2_ ( .D(
        or1200_cpu_or1200_mult_mac_n1558), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n124) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_1_ ( .D(
        or1200_cpu_or1200_mult_mac_n1559), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n126) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_quot_r_reg_0_ ( .D(
        or1200_cpu_or1200_mult_mac_n1527), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n128) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_cntr_reg_0_ ( .D(
        or1200_cpu_or1200_mult_mac_n1106), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_div_cntr_0_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_cntr_reg_1_ ( .D(
        or1200_cpu_or1200_mult_mac_n1105), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_div_cntr_1_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_cntr_reg_2_ ( .D(
        or1200_cpu_or1200_mult_mac_n1104), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_div_cntr_2_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_cntr_reg_3_ ( .D(
        or1200_cpu_or1200_mult_mac_n1103), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_div_cntr_3_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_cntr_reg_4_ ( .D(
        or1200_cpu_or1200_mult_mac_n1107), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_div_cntr_4_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_cntr_reg_5_ ( .D(
        or1200_cpu_or1200_mult_mac_n1560), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n135) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_div_free_reg ( .D(
        or1200_cpu_or1200_mult_mac_n136), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_div_free) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_stall_r_reg ( .D(
        or1200_cpu_or1200_mult_mac_N503), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n139) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_0_ ( .D(
        or1200_cpu_or1200_mult_mac_n1625), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n141) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_1_ ( .D(
        or1200_cpu_or1200_mult_mac_n1592), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n143) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_2_ ( .D(
        or1200_cpu_or1200_mult_mac_n1591), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n145) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_3_ ( .D(
        or1200_cpu_or1200_mult_mac_n1590), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n147) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_4_ ( .D(
        or1200_cpu_or1200_mult_mac_n1589), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n149) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_5_ ( .D(
        or1200_cpu_or1200_mult_mac_n1588), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n151) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_6_ ( .D(
        or1200_cpu_or1200_mult_mac_n1587), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n153) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_7_ ( .D(
        or1200_cpu_or1200_mult_mac_n1586), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n155) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_8_ ( .D(
        or1200_cpu_or1200_mult_mac_n1585), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n157) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_9_ ( .D(
        or1200_cpu_or1200_mult_mac_n1584), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n159) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_10_ ( .D(
        or1200_cpu_or1200_mult_mac_n1583), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n161) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_11_ ( .D(
        or1200_cpu_or1200_mult_mac_n1582), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n163) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_12_ ( .D(
        or1200_cpu_or1200_mult_mac_n1581), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n165) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_13_ ( .D(
        or1200_cpu_or1200_mult_mac_n1580), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n167) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_14_ ( .D(
        or1200_cpu_or1200_mult_mac_n1579), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n169) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_15_ ( .D(
        or1200_cpu_or1200_mult_mac_n1578), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n171) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_16_ ( .D(
        or1200_cpu_or1200_mult_mac_n1577), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n173) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_17_ ( .D(
        or1200_cpu_or1200_mult_mac_n1576), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n175) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_18_ ( .D(
        or1200_cpu_or1200_mult_mac_n1575), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n177) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_19_ ( .D(
        or1200_cpu_or1200_mult_mac_n1574), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n179) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_20_ ( .D(
        or1200_cpu_or1200_mult_mac_n1573), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n181) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_21_ ( .D(
        or1200_cpu_or1200_mult_mac_n1572), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n183) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_22_ ( .D(
        or1200_cpu_or1200_mult_mac_n1571), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n185) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_23_ ( .D(
        or1200_cpu_or1200_mult_mac_n1570), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n187) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_24_ ( .D(
        or1200_cpu_or1200_mult_mac_n1569), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n189) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_25_ ( .D(
        or1200_cpu_or1200_mult_mac_n1568), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n191) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_26_ ( .D(
        or1200_cpu_or1200_mult_mac_n1567), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n193) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_27_ ( .D(
        or1200_cpu_or1200_mult_mac_n1566), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n195) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_28_ ( .D(
        or1200_cpu_or1200_mult_mac_n1565), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n197) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_29_ ( .D(
        or1200_cpu_or1200_mult_mac_n1564), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n199) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_30_ ( .D(
        or1200_cpu_or1200_mult_mac_n1563), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n201) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_31_ ( .D(
        or1200_cpu_or1200_mult_mac_n1562), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n203) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_32_ ( .D(
        or1200_cpu_or1200_mult_mac_n1624), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n205) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_33_ ( .D(
        or1200_cpu_or1200_mult_mac_n1623), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n207) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_34_ ( .D(
        or1200_cpu_or1200_mult_mac_n1622), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n209) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_35_ ( .D(
        or1200_cpu_or1200_mult_mac_n1621), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n211) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_36_ ( .D(
        or1200_cpu_or1200_mult_mac_n1620), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n213) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_37_ ( .D(
        or1200_cpu_or1200_mult_mac_n1619), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n215) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_38_ ( .D(
        or1200_cpu_or1200_mult_mac_n1618), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n217) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_39_ ( .D(
        or1200_cpu_or1200_mult_mac_n1617), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n219) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_40_ ( .D(
        or1200_cpu_or1200_mult_mac_n1616), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n221) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_41_ ( .D(
        or1200_cpu_or1200_mult_mac_n1615), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n223) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_42_ ( .D(
        or1200_cpu_or1200_mult_mac_n1614), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n225) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_43_ ( .D(
        or1200_cpu_or1200_mult_mac_n1613), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n227) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_44_ ( .D(
        or1200_cpu_or1200_mult_mac_n1612), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n229) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_45_ ( .D(
        or1200_cpu_or1200_mult_mac_n1611), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n231) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_46_ ( .D(
        or1200_cpu_or1200_mult_mac_n1610), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n233) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_47_ ( .D(
        or1200_cpu_or1200_mult_mac_n1609), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n235) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_48_ ( .D(
        or1200_cpu_or1200_mult_mac_n1608), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n237) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_49_ ( .D(
        or1200_cpu_or1200_mult_mac_n1607), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n239) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_50_ ( .D(
        or1200_cpu_or1200_mult_mac_n1606), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n241) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_51_ ( .D(
        or1200_cpu_or1200_mult_mac_n1605), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n243) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_52_ ( .D(
        or1200_cpu_or1200_mult_mac_n1604), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n245) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_53_ ( .D(
        or1200_cpu_or1200_mult_mac_n1603), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n247) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_54_ ( .D(
        or1200_cpu_or1200_mult_mac_n1602), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n249) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_55_ ( .D(
        or1200_cpu_or1200_mult_mac_n1601), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n251) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_56_ ( .D(
        or1200_cpu_or1200_mult_mac_n1600), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n253) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_57_ ( .D(
        or1200_cpu_or1200_mult_mac_n1599), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n255) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_58_ ( .D(
        or1200_cpu_or1200_mult_mac_n1598), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n257) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_59_ ( .D(
        or1200_cpu_or1200_mult_mac_n1597), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n259) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_60_ ( .D(
        or1200_cpu_or1200_mult_mac_n1596), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n261) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_61_ ( .D(
        or1200_cpu_or1200_mult_mac_n1595), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n263) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_62_ ( .D(
        or1200_cpu_or1200_mult_mac_n1594), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n265) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_r_reg_63_ ( .D(
        or1200_cpu_or1200_mult_mac_n1593), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n267) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r3_reg_0_ ( .D(
        or1200_cpu_or1200_mult_mac_mac_op_r2_0_), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n269) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r3_reg_1_ ( .D(
        or1200_cpu_or1200_mult_mac_mac_op_r2_1_), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n271) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r3_reg_2_ ( .D(
        or1200_cpu_or1200_mult_mac_mac_op_r2_2_), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n273) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r2_reg_0_ ( .D(
        or1200_cpu_or1200_mult_mac_n278), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_mac_op_r2_0_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r2_reg_1_ ( .D(
        or1200_cpu_or1200_mult_mac_n280), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_mac_op_r2_1_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r2_reg_2_ ( .D(
        or1200_cpu_or1200_mult_mac_n282), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_mac_op_r2_2_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r1_reg_0_ ( .D(
        or1200_cpu_or1200_mult_mac_N292), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n278) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r1_reg_1_ ( .D(
        or1200_cpu_or1200_mult_mac_N293), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n280) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mac_op_r1_reg_2_ ( .D(
        or1200_cpu_or1200_mult_mac_N294), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_mult_mac_n282) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_stall_count_reg_1_ ( 
        .D(or1200_cpu_or1200_mult_mac_n285), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_mult_mac_mul_stall_count_1_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_stall_count_reg_0_ ( 
        .D(or1200_cpu_or1200_mult_mac_N290), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n285) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_0_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[0]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n287) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_1_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[1]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n289) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_2_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[2]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n291) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_3_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[3]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n293) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_4_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[4]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n295) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_5_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[5]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n297) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_6_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[6]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n299) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_7_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[7]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n301) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_8_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[8]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n303) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_9_ ( .D(
        or1200_cpu_or1200_mult_mac_mul_prod[9]), .CLK(clk_i), .RESET(n53192), 
        .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n305) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_10_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[10]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n307) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_11_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[11]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n309) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_12_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[12]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n311) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_13_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[13]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n313) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_14_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[14]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n315) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_15_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[15]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n317) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_16_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[16]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n319) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_17_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[17]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n321) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_18_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[18]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n323) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_19_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[19]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n325) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_20_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[20]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n327) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_21_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[21]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n329) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_22_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[22]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n331) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_23_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[23]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n333) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_24_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[24]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n335) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_25_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[25]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n337) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_26_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[26]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n339) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_27_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[27]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n341) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_28_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[28]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n343) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_29_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[29]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n345) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_30_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[30]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n347) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_31_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[31]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n349) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_32_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[32]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n351) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_33_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[33]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n353) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_34_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[34]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n355) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_35_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[35]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n357) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_36_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[36]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n359) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_37_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[37]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n361) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_38_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[38]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n363) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_39_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[39]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n365) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_40_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[40]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n367) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_41_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[41]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n369) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_42_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[42]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n371) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_43_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[43]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n373) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_44_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[44]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n375) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_45_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[45]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n377) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_46_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[46]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n379) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_47_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[47]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n381) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_48_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[48]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n383) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_49_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[49]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n385) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_50_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[50]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n387) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_51_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[51]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n389) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_52_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[52]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n391) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_53_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[53]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n393) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_54_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[54]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n395) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_55_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[55]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n397) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_56_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[56]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n399) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_57_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[57]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n401) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_58_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[58]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n403) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_59_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[59]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n405) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_60_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[60]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n407) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_61_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[61]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n409) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_62_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[62]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n411) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_mul_prod_r_reg_63_ ( 
        .D(or1200_cpu_or1200_mult_mac_mul_prod[63]), .CLK(clk_i), .RESET(
        n53192), .SET(rst_i), .QN(or1200_cpu_or1200_mult_mac_n413) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_ex_freeze_r_reg ( .D(
        n57073), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_ex_freeze_r) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_14_ ( 
        .D(n59560), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_14_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_0_ ( 
        .D(n59565), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_30_ ( 
        .D(n59576), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_30_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_2_ ( 
        .D(n59568), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_6_ ( 
        .D(n59555), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_24_ ( .D(
        n57068), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_28_ ( .D(
        n1868), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_23_ ( .D(
        n59547), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_29_ ( .D(
        n59549), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_29_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_27_ ( .D(
        n59548), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_27_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r_reg_1_ ( 
        .D(n1598), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SRAM or1200_immu_top_icpu_vpn_r_reg_27_ ( .D(
        icqmem_adr_qmem[27]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n769) );
  ASYNC_DFFHx1_ASAP7_75t_SRAM or1200_immu_top_icpu_vpn_r_reg_21_ ( .D(
        icqmem_adr_qmem[21]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n793) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_17_ ( .D(
        n59536), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_14_ ( .D(
        n59552), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[14]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_44_ ( 
        .D(n52005), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n154) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_1_ ( 
        .D(n59564), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_56_ ( 
        .D(n52010), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n178) );
  OAI31xp33_ASAP7_75t_SRAM U9857 ( .A1(n22057), .A2(n4152), .A3(n53192), .B(
        n3645), .Y(or1200_ic_top_icram_we_3_) );
  INVx1_ASAP7_75t_SL U3307 ( .A(n2783), .Y(ic_en) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_rf_spr_du_cs_reg ( .D(
        or1200_cpu_or1200_rf_n44), .CLK(clk_i), .QN(
        or1200_cpu_or1200_rf_spr_du_cs) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_12_ ( 
        .D(n59570), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_12_) );
  ASYNC_DFFHx1_ASAP7_75t_SRAM or1200_cpu_or1200_sprs_sr_reg_reg_15_ ( .D(n2688), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(or1200_cpu_sr_15_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r_reg_5_ ( 
        .D(n1550), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r_reg_4_ ( 
        .D(n1556), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]) );
  ASYNC_DFFHx1_ASAP7_75t_SRAM or1200_immu_top_icpu_vpn_r_reg_29_ ( .D(
        icqmem_adr_qmem[29]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n761) );
  TIELOx1_ASAP7_75t_SL U27514 ( .L(n78441) );
  spram or1200_ic_top_or1200_ic_tag_ic_tag0 ( .clock(clk_i), .ce(
        or1200_ic_top_ictag_en), .wren(or1200_ic_top_ictag_we), .address(
        or1200_ic_top_ictag_addr), .data({icbiu_adr_ic_word[31:12], 
        or1200_ic_top_ictag_v}), .q({or1200_ic_top_tag, or1200_ic_top_tag_v})
         );
  spram or1200_ic_top_or1200_ic_ram_ic_ram0 ( .clock(clk_i), .ce(ic_en), 
        .wren(or1200_ic_top_icram_we_3_), .address(icbiu_adr_ic_word[11:2]), 
        .data(iwb_dat_i), .q(or1200_ic_top_from_icram) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_extend_flush_reg ( .D(
        or1200_cpu_or1200_except_n1731), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n116) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_except_type_reg_1_ ( .D(
        or1200_cpu_or1200_except_n1733), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_except_type_1_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_except_type_reg_0_ ( .D(
        or1200_cpu_or1200_except_n1734), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n120) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dsx_reg ( .D(
        or1200_cpu_or1200_except_n1735), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n122) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_31_ ( .D(
        or1200_cpu_or1200_except_n1699), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n124) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_30_ ( .D(
        or1200_cpu_or1200_except_n1700), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n126) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_29_ ( .D(
        or1200_cpu_or1200_except_n1701), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n128) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_28_ ( .D(
        or1200_cpu_or1200_except_n1702), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n130) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_27_ ( .D(
        or1200_cpu_or1200_except_n1703), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n132) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_26_ ( .D(
        or1200_cpu_or1200_except_n1704), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n134) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_25_ ( .D(
        or1200_cpu_or1200_except_n1705), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n136) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_24_ ( .D(
        or1200_cpu_or1200_except_n1706), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n138) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_23_ ( .D(
        or1200_cpu_or1200_except_n1707), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n140) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_22_ ( .D(
        or1200_cpu_or1200_except_n1708), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n142) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_21_ ( .D(
        or1200_cpu_or1200_except_n1709), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n144) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_20_ ( .D(
        or1200_cpu_or1200_except_n1710), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n146) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_19_ ( .D(
        or1200_cpu_or1200_except_n1711), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n148) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_18_ ( .D(
        or1200_cpu_or1200_except_n1712), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n150) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_17_ ( .D(
        or1200_cpu_or1200_except_n1713), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n152) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_16_ ( .D(
        or1200_cpu_or1200_except_n1714), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n154) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_15_ ( .D(
        or1200_cpu_or1200_except_n1715), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n156) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_14_ ( .D(
        or1200_cpu_or1200_except_n1716), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n158) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_13_ ( .D(
        or1200_cpu_or1200_except_n1717), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n160) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_12_ ( .D(
        or1200_cpu_or1200_except_n1718), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n162) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_11_ ( .D(
        or1200_cpu_or1200_except_n1719), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n164) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_10_ ( .D(
        or1200_cpu_or1200_except_n1720), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n166) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_9_ ( .D(
        or1200_cpu_or1200_except_n1721), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n168) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_8_ ( .D(
        or1200_cpu_or1200_except_n1722), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n170) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_7_ ( .D(
        or1200_cpu_or1200_except_n1723), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n172) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_6_ ( .D(
        or1200_cpu_or1200_except_n1724), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n174) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_5_ ( .D(
        or1200_cpu_or1200_except_n1725), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n176) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_4_ ( .D(
        or1200_cpu_or1200_except_n1726), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n178) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_3_ ( .D(
        or1200_cpu_or1200_except_n1727), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n180) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_2_ ( .D(
        or1200_cpu_or1200_except_n1728), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n182) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_1_ ( .D(
        or1200_cpu_or1200_except_n1729), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n184) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_eear_reg_0_ ( .D(
        or1200_cpu_or1200_except_n1730), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n186) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_0_ ( .D(
        or1200_cpu_or1200_except_n1784), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n188) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_1_ ( .D(
        or1200_cpu_or1200_except_n1783), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_epcr_1_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_2_ ( .D(
        or1200_cpu_or1200_except_n1782), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n192) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_3_ ( .D(
        or1200_cpu_or1200_except_n1781), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n194) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_4_ ( .D(
        or1200_cpu_or1200_except_n1780), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n196) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_5_ ( .D(
        or1200_cpu_or1200_except_n1779), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n198) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_6_ ( .D(
        or1200_cpu_or1200_except_n1778), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n200) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_7_ ( .D(
        or1200_cpu_or1200_except_n1777), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n202) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_8_ ( .D(
        or1200_cpu_or1200_except_n1776), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n204) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_9_ ( .D(
        or1200_cpu_or1200_except_n1775), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n206) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_10_ ( .D(
        or1200_cpu_or1200_except_n1774), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n208) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_11_ ( .D(
        or1200_cpu_or1200_except_n1773), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n210) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_12_ ( .D(
        or1200_cpu_or1200_except_n1772), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n212) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_13_ ( .D(
        or1200_cpu_or1200_except_n1771), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n214) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_14_ ( .D(
        or1200_cpu_or1200_except_n1770), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n216) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_15_ ( .D(
        or1200_cpu_or1200_except_n1769), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n218) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_16_ ( .D(
        or1200_cpu_or1200_except_n1768), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n220) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_17_ ( .D(
        or1200_cpu_or1200_except_n1767), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n222) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_18_ ( .D(
        or1200_cpu_or1200_except_n1766), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n224) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_19_ ( .D(
        or1200_cpu_or1200_except_n1765), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n226) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_20_ ( .D(
        or1200_cpu_or1200_except_n1764), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n228) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_21_ ( .D(
        or1200_cpu_or1200_except_n1763), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n230) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_22_ ( .D(
        or1200_cpu_or1200_except_n1762), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n232) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_23_ ( .D(
        or1200_cpu_or1200_except_n1761), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n234) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_24_ ( .D(
        or1200_cpu_or1200_except_n1760), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n236) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_25_ ( .D(
        or1200_cpu_or1200_except_n1759), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n238) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_26_ ( .D(
        or1200_cpu_or1200_except_n1758), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n240) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_27_ ( .D(
        or1200_cpu_or1200_except_n1757), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n242) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_28_ ( .D(
        or1200_cpu_or1200_except_n1756), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n244) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_29_ ( .D(
        or1200_cpu_or1200_except_n1755), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n246) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_30_ ( .D(
        or1200_cpu_or1200_except_n1754), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n248) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_epcr_reg_31_ ( .D(
        or1200_cpu_or1200_except_n1753), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_epcr_31_) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_16_ ( .D(
        or1200_cpu_or1200_except_n1736), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n252) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_15_ ( .D(
        or1200_cpu_or1200_except_n253), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_esr[15]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_14_ ( .D(
        or1200_cpu_or1200_except_n1738), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n256) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_13_ ( .D(
        or1200_cpu_or1200_except_n1739), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n258) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_12_ ( .D(
        or1200_cpu_or1200_except_n1740), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n260) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_11_ ( .D(
        or1200_cpu_or1200_except_n1741), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n262) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_10_ ( .D(
        or1200_cpu_or1200_except_n1742), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n264) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_9_ ( .D(
        or1200_cpu_or1200_except_n1743), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n266) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_8_ ( .D(
        or1200_cpu_or1200_except_n1744), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n268) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_7_ ( .D(
        or1200_cpu_or1200_except_n1745), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n270) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_6_ ( .D(
        or1200_cpu_or1200_except_n1746), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n272) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_5_ ( .D(
        or1200_cpu_or1200_except_n1747), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n274) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_4_ ( .D(
        or1200_cpu_or1200_except_n1748), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n276) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_3_ ( .D(
        or1200_cpu_or1200_except_n1749), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n278) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_2_ ( .D(
        or1200_cpu_or1200_except_n1750), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n280) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_1_ ( .D(
        or1200_cpu_or1200_except_n1751), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n282) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_esr_reg_0_ ( .D(
        or1200_cpu_or1200_except_n283), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_esr[0]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_except_type_reg_3_ ( .D(
        or1200_cpu_or1200_except_n1787), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n286) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_state_reg_2_ ( .D(
        or1200_cpu_or1200_except_n1785), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n288) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_state_reg_1_ ( .D(
        or1200_cpu_or1200_except_n1786), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n290) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_except_type_reg_2_ ( .D(
        or1200_cpu_or1200_except_n1732), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n292) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_state_reg_0_ ( .D(
        or1200_cpu_or1200_except_n1788), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n294) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_2_ ( .D(
        or1200_cpu_or1200_except_n303), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n302) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_3_ ( .D(
        or1200_cpu_or1200_except_n306), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n305) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_4_ ( .D(
        or1200_cpu_or1200_except_n309), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n308) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_5_ ( .D(
        or1200_cpu_or1200_except_n312), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n311) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_6_ ( .D(
        or1200_cpu_or1200_except_n315), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n314) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_7_ ( .D(
        or1200_cpu_or1200_except_n318), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n317) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_8_ ( .D(
        or1200_cpu_or1200_except_n321), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n320) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_9_ ( .D(
        or1200_cpu_or1200_except_n324), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n323) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_10_ ( .D(
        or1200_cpu_or1200_except_n327), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n326) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_11_ ( .D(
        or1200_cpu_or1200_except_n330), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n329) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_12_ ( .D(
        or1200_cpu_or1200_except_n333), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n332) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_13_ ( .D(
        or1200_cpu_or1200_except_n336), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n335) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_14_ ( .D(
        or1200_cpu_or1200_except_n339), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n338) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_15_ ( .D(
        or1200_cpu_or1200_except_n342), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n341) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_16_ ( .D(
        or1200_cpu_or1200_except_n345), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n344) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_17_ ( .D(
        or1200_cpu_or1200_except_n348), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n347) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_18_ ( .D(
        or1200_cpu_or1200_except_n351), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n350) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_19_ ( .D(
        or1200_cpu_or1200_except_n354), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n353) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_20_ ( .D(
        or1200_cpu_or1200_except_n357), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n356) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_21_ ( .D(
        or1200_cpu_or1200_except_n360), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n359) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_22_ ( .D(
        or1200_cpu_or1200_except_n363), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n362) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_23_ ( .D(
        or1200_cpu_or1200_except_n366), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n365) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_24_ ( .D(
        or1200_cpu_or1200_except_n369), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n368) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_25_ ( .D(
        or1200_cpu_or1200_except_n372), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n371) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_26_ ( .D(
        or1200_cpu_or1200_except_n375), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n374) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_27_ ( .D(
        or1200_cpu_or1200_except_n378), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n377) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_28_ ( .D(
        or1200_cpu_or1200_except_n381), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n380) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_29_ ( .D(
        or1200_cpu_or1200_except_n384), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n383) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_30_ ( .D(
        or1200_cpu_or1200_except_n387), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n386) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dl_pc_reg_31_ ( .D(
        or1200_cpu_or1200_except_n390), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n389) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_2_ ( .D(
        or1200_cpu_or1200_except_n399), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n398) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_3_ ( .D(
        or1200_cpu_or1200_except_n402), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n401) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_4_ ( .D(
        or1200_cpu_or1200_except_n405), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n404) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_5_ ( .D(
        or1200_cpu_or1200_except_n408), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n407) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_6_ ( .D(
        or1200_cpu_or1200_except_n411), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n410) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_7_ ( .D(
        or1200_cpu_or1200_except_n414), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n413) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_8_ ( .D(
        or1200_cpu_or1200_except_n417), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n416) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_9_ ( .D(
        or1200_cpu_or1200_except_n420), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n419) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_10_ ( .D(
        or1200_cpu_or1200_except_n423), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n422) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_11_ ( .D(
        or1200_cpu_or1200_except_n426), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n425) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_12_ ( .D(
        or1200_cpu_or1200_except_n429), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n428) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_13_ ( .D(
        or1200_cpu_or1200_except_n432), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n431) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_14_ ( .D(
        or1200_cpu_or1200_except_n435), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n434) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_15_ ( .D(
        or1200_cpu_or1200_except_n438), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n437) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_16_ ( .D(
        or1200_cpu_or1200_except_n441), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n440) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_17_ ( .D(
        or1200_cpu_or1200_except_n444), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[17]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_18_ ( .D(
        or1200_cpu_or1200_except_n447), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n446) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_19_ ( .D(
        or1200_cpu_or1200_except_n450), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[19]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_20_ ( .D(
        or1200_cpu_or1200_except_n453), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[20]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_21_ ( .D(
        or1200_cpu_or1200_except_n456), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[21]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_22_ ( .D(
        or1200_cpu_or1200_except_n459), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[22]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_23_ ( .D(
        or1200_cpu_or1200_except_n462), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n461) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_24_ ( .D(
        or1200_cpu_or1200_except_n465), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[24]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_25_ ( .D(
        or1200_cpu_or1200_except_n468), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n467) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_26_ ( .D(
        or1200_cpu_or1200_except_n471), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[26]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_27_ ( .D(
        or1200_cpu_or1200_except_n474), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[27]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_28_ ( .D(
        or1200_cpu_or1200_except_n477), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n476) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_29_ ( .D(
        or1200_cpu_or1200_except_n480), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[29]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_30_ ( .D(
        or1200_cpu_or1200_except_n483), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n482) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_wb_pc_reg_31_ ( .D(
        or1200_cpu_or1200_except_n486), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_spr_dat_ppc[31]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_2_ ( .D(
        or1200_cpu_or1200_except_n1791), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n492) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_3_ ( .D(
        or1200_cpu_or1200_except_n1792), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n494) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_4_ ( .D(
        or1200_cpu_or1200_except_n1793), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n496) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_5_ ( .D(
        or1200_cpu_or1200_except_n1794), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n498) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_6_ ( .D(
        or1200_cpu_or1200_except_n1795), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n500) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_7_ ( .D(
        or1200_cpu_or1200_except_n1796), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n502) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_8_ ( .D(
        or1200_cpu_or1200_except_n1797), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n504) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_9_ ( .D(
        or1200_cpu_or1200_except_n1798), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n506) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_10_ ( .D(
        or1200_cpu_or1200_except_n1799), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n508) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_11_ ( .D(
        or1200_cpu_or1200_except_n1800), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n510) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_12_ ( .D(
        or1200_cpu_or1200_except_n1801), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n512) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_13_ ( .D(
        or1200_cpu_or1200_except_n1802), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n514) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_14_ ( .D(
        or1200_cpu_or1200_except_n1803), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n516) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_15_ ( .D(
        or1200_cpu_or1200_except_n1804), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n518) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_16_ ( .D(
        or1200_cpu_or1200_except_n1805), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n520) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_17_ ( .D(
        or1200_cpu_or1200_except_n1806), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n522) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_18_ ( .D(
        or1200_cpu_or1200_except_n1807), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n524) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_19_ ( .D(
        or1200_cpu_or1200_except_n1808), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n526) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_20_ ( .D(
        or1200_cpu_or1200_except_n1809), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n528) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_21_ ( .D(
        or1200_cpu_or1200_except_n1810), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n530) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_22_ ( .D(
        or1200_cpu_or1200_except_n1811), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n532) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_23_ ( .D(
        or1200_cpu_or1200_except_n1812), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n534) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_24_ ( .D(
        or1200_cpu_or1200_except_n1813), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n536) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_25_ ( .D(
        or1200_cpu_or1200_except_n1814), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n538) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_26_ ( .D(
        or1200_cpu_or1200_except_n1815), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n540) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_27_ ( .D(
        or1200_cpu_or1200_except_n1816), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n542) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_28_ ( .D(
        or1200_cpu_or1200_except_n1817), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n544) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_29_ ( .D(
        or1200_cpu_or1200_except_n1818), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n546) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_30_ ( .D(
        or1200_cpu_or1200_except_n1819), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n548) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_reg_31_ ( .D(
        or1200_cpu_or1200_except_n1820), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n550) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_trace_trap_reg ( .D(
        or1200_cpu_or1200_except_n553), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n552) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_pc_val_reg ( .D(
        or1200_cpu_or1200_except_n1821), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n555) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_exceptflags_reg_2_ ( 
        .D(or1200_cpu_or1200_except_n1824), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n561) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_delayed2_ex_dslot_reg ( 
        .D(or1200_cpu_or1200_except_n1825), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n563) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_delayed1_ex_dslot_reg ( 
        .D(or1200_cpu_or1200_except_n1826), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n565) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_dslot_reg ( .D(
        or1200_cpu_or1200_except_n1827), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n567) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_delayed_tee_reg_2_ ( .D(
        or1200_cpu_or1200_except_n1694), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_except_delayed_tee[2]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_delayed_tee_reg_1_ ( .D(
        n58626), .CLK(clk_i), .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_except_delayed_tee[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_delayed_tee_reg_0_ ( .D(
        n78260), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_except_n571) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_delayed_iee_reg_2_ ( .D(
        or1200_cpu_or1200_except_n1696), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_except_delayed_iee[2]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_delayed_iee_reg_1_ ( .D(
        or1200_cpu_or1200_except_n1697), .CLK(clk_i), .RESET(rst_i), .SET(
        n53192), .QN(or1200_cpu_or1200_except_delayed_iee[1]) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_delayed_iee_reg_0_ ( .D(
        n78253), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_except_n575) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_2_ ( .D(
        or1200_cpu_or1200_except_n584), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n583) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_3_ ( .D(
        or1200_cpu_or1200_except_n587), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n586) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_4_ ( .D(
        or1200_cpu_or1200_except_n590), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n589) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_5_ ( .D(
        or1200_cpu_or1200_except_n593), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n592) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_6_ ( .D(
        or1200_cpu_or1200_except_n596), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n595) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_7_ ( .D(
        or1200_cpu_or1200_except_n599), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n598) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_8_ ( .D(
        or1200_cpu_or1200_except_n602), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n601) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_9_ ( .D(
        or1200_cpu_or1200_except_n605), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n604) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_10_ ( .D(
        or1200_cpu_or1200_except_n608), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n607) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_11_ ( .D(
        or1200_cpu_or1200_except_n611), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n610) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_12_ ( .D(
        or1200_cpu_or1200_except_n614), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n613) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_13_ ( .D(
        or1200_cpu_or1200_except_n617), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n616) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_14_ ( .D(
        or1200_cpu_or1200_except_n620), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n619) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_15_ ( .D(
        or1200_cpu_or1200_except_n623), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n622) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_16_ ( .D(
        or1200_cpu_or1200_except_n626), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n625) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_17_ ( .D(
        or1200_cpu_or1200_except_n629), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n628) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_18_ ( .D(
        or1200_cpu_or1200_except_n632), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n631) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_19_ ( .D(
        or1200_cpu_or1200_except_n635), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n634) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_20_ ( .D(
        or1200_cpu_or1200_except_n638), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n637) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_21_ ( .D(
        or1200_cpu_or1200_except_n641), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n640) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_22_ ( .D(
        or1200_cpu_or1200_except_n644), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n643) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_23_ ( .D(
        or1200_cpu_or1200_except_n647), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n646) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_24_ ( .D(
        or1200_cpu_or1200_except_n650), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n649) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_25_ ( .D(
        or1200_cpu_or1200_except_n653), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n652) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_26_ ( .D(
        or1200_cpu_or1200_except_n656), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n655) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_27_ ( .D(
        or1200_cpu_or1200_except_n659), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n658) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_28_ ( .D(
        or1200_cpu_or1200_except_n662), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n661) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_29_ ( .D(
        or1200_cpu_or1200_except_n665), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n664) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_30_ ( .D(
        or1200_cpu_or1200_except_n668), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n667) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_reg_31_ ( .D(
        or1200_cpu_or1200_except_n671), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n670) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_exceptflags_reg_2_ ( 
        .D(or1200_cpu_or1200_except_n1830), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n677) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_id_pc_val_reg ( .D(
        or1200_cpu_or1200_except_n1831), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n679) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_sr_ted_prev_reg ( .D(
        or1200_cpu_or1200_except_n682), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n681) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dmr1_bt_prev_reg ( .D(
        or1200_cpu_or1200_except_n685), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n684) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dmr1_st_prev_reg ( .D(
        n76670), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_except_n687) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_dsr_te_prev_reg ( .D(
        or1200_cpu_or1200_except_n691), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(or1200_cpu_or1200_except_n690) );
  ASYNC_DFFHx1_ASAP7_75t_SL or1200_cpu_or1200_except_ex_freeze_prev_reg ( .D(
        n57073), .CLK(clk_i), .RESET(rst_i), .SET(n53192), .QN(
        or1200_cpu_or1200_except_ex_freeze_prev) );
  spram or1200_dc_top_or1200_dc_tag_dc_tag0 ( .clock(clk_i), .ce(
        or1200_dc_top_dctag_en), .wren(or1200_dc_top_dctag_we), .address(
        or1200_dc_top_dctag_addr), .data({sbbiu_adr_sb[31:12], 
        or1200_dc_top_dctag_v, n78441}), .q({or1200_dc_top_tag_19_, 
        or1200_dc_top_tag_18_, or1200_dc_top_tag_17_, or1200_dc_top_tag_16_, 
        or1200_dc_top_tag_15_, or1200_dc_top_tag_14_, or1200_dc_top_tag_13_, 
        or1200_dc_top_tag_12_, or1200_dc_top_tag_11_, or1200_dc_top_tag_10_, 
        or1200_dc_top_tag_9_, or1200_dc_top_tag_8_, or1200_dc_top_tag_7_, 
        or1200_dc_top_tag_6_, or1200_dc_top_tag_5_, or1200_dc_top_tag_4_, 
        or1200_dc_top_tag_3_, or1200_dc_top_tag_2_, or1200_dc_top_tag_1_, 
        or1200_dc_top_tag_0_, or1200_dc_top_tag_v, or1200_dc_top_dirty}) );
  spram or1200_dc_top_or1200_dc_ram_dc_ram3 ( .clock(clk_i), .ce(dc_en), 
        .wren(or1200_dc_top_dcram_we[3]), .address(sbbiu_adr_sb[11:2]), .data(
        or1200_dc_top_to_dcram[31:24]), .q({or1200_dc_top_from_dcram_31_, 
        or1200_dc_top_from_dcram_30_, or1200_dc_top_from_dcram_29_, 
        or1200_dc_top_from_dcram_28_, or1200_dc_top_from_dcram_27_, 
        or1200_dc_top_from_dcram_26_, or1200_dc_top_from_dcram_25_, 
        or1200_dc_top_from_dcram_24_}) );
  spram or1200_dc_top_or1200_dc_ram_dc_ram2 ( .clock(clk_i), .ce(dc_en), 
        .wren(or1200_dc_top_dcram_we[2]), .address(sbbiu_adr_sb[11:2]), .data(
        or1200_dc_top_to_dcram[23:16]), .q({or1200_dc_top_from_dcram_23_, 
        or1200_dc_top_from_dcram_22_, or1200_dc_top_from_dcram_21_, 
        or1200_dc_top_from_dcram_20_, or1200_dc_top_from_dcram_19_, 
        or1200_dc_top_from_dcram_18_, or1200_dc_top_from_dcram_17_, 
        or1200_dc_top_from_dcram_16_}) );
  spram or1200_dc_top_or1200_dc_ram_dc_ram1 ( .clock(clk_i), .ce(dc_en), 
        .wren(or1200_dc_top_dcram_we[1]), .address(sbbiu_adr_sb[11:2]), .data(
        or1200_dc_top_to_dcram[15:8]), .q({or1200_dc_top_from_dcram_15_, 
        or1200_dc_top_from_dcram_14_, or1200_dc_top_from_dcram_13_, 
        or1200_dc_top_from_dcram_12_, or1200_dc_top_from_dcram_11_, 
        or1200_dc_top_from_dcram_10_, or1200_dc_top_from_dcram_9_, 
        or1200_dc_top_from_dcram_8_}) );
  spram or1200_dc_top_or1200_dc_ram_dc_ram0 ( .clock(clk_i), .ce(dc_en), 
        .wren(or1200_dc_top_dcram_we[0]), .address(sbbiu_adr_sb[11:2]), .data(
        or1200_dc_top_to_dcram[7:0]), .q({or1200_dc_top_from_dcram_7_, 
        or1200_dc_top_from_dcram_6_, or1200_dc_top_from_dcram_5_, 
        or1200_dc_top_from_dcram_4_, or1200_dc_top_from_dcram_3_, 
        or1200_dc_top_from_dcram_2_, or1200_dc_top_from_dcram_1_, 
        or1200_dc_top_from_dcram_0_}) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_6_ ( 
        .D(n27033), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_6_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_reg_5_ ( 
        .D(n78361), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_5_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_reg_6_ ( 
        .D(n78363), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_6_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_reg_0_ ( 
        .D(n78372), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_0_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_0_ ( 
        .D(n78429), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_0_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_2_ ( 
        .D(n78433), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_2_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_6_ ( 
        .D(n78339), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_6_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_31_ ( 
        .D(n28158), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[31]) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_47_ ( 
        .D(n28207), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n120), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n1), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n2), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_0_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n3), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n4), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_1_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n5), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n6), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_2_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n7), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_3_ ( 
        .D(n74344), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n9), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n10), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_4_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n11), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_5_ ( 
        .D(n74357), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n13), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n14), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_6_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_7_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n15), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_7_ ( 
        .D(n74316), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_8_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n17), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_8_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n18), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_8_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_9_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n19), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_9_ ( 
        .D(n74327), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_10_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n21), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_10_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n22), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_10_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_11_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n23), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_11_ ( 
        .D(n74349), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_12_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n25), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_12_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n26), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_12_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_13_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n27), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_13_ ( 
        .D(n74393), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_14_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n29), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_14_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n30), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_14_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_15_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n31), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_15_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n32), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_15_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_16_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n33), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_16_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n34), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_16_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_17_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n35), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_17_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n36), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_17_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n37), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n38), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_18_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_19_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n39), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_19_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n40), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_19_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_20_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n41), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_20_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n42), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_20_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_21_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n43), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_21_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n44), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_21_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n45), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n46), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_22_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_23_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n47), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_23_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_30_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n48), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[30]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_29_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n49), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[29]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_28_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n50), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[28]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_27_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n51), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[27]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_26_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n52), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[26]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_25_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n53), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[25]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_24_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n54), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[24]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_output_o_reg_23_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n55), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_ine_o_reg ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n56), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_ine) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_reg_24_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n57), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n58), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n59), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n60), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n61), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n62), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n63), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n64), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_7_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n65), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_8_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n66), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_9_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n67), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_10_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n68), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_11_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n69), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_12_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n70), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_13_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n71), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_14_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n72), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_15_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n73), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_16_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n74), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_17_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n75), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n76), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_19_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n77), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_20_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n78), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_21_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n79), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n80), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_23_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n81), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_24_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n82), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_24_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_25_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n83), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_25_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_26_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n84), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_26_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_27_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n85), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_27_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_28_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n86), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_28_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_29_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n87), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_29_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_30_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n88), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_30_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_31_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n89), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_31_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_32_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n90), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_32_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_33_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n91), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_33_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_34_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n92), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_34_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_35_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n93), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_35_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_36_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n94), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_36_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_37_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n95), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_37_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_38_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n96), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_38_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_39_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n97), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_39_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_40_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n98), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_40_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_41_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n99), .CLK(clk_i), 
        .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_41_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_42_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n100), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_42_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_43_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n101), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_43_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_44_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n102), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_44_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_45_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n103), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_45_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_46_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_N2648), .CLK(
        clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_reg_47_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n105), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_47_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n106), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_reg_1_ ( 
        .D(n28105), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n108), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n109), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n110), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n111), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n112), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_reg_7_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n113), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n126), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n127), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n128), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n129), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n130), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_N2435), .CLK(
        clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n131) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n132), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n133), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n134), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n135), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n136), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n137), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_0_ ( 
        .D(n28198), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_1_ ( 
        .D(n28199), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_2_ ( 
        .D(n28200), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_4_ ( 
        .D(n28202), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_5_ ( 
        .D(n28203), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_6_ ( 
        .D(n28204), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_7_ ( 
        .D(n28161), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_8_ ( 
        .D(n28162), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_9_ ( 
        .D(n28163), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_10_ ( 
        .D(n28164), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_11_ ( 
        .D(n28165), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_13_ ( 
        .D(n28167), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_14_ ( 
        .D(n28168), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_15_ ( 
        .D(n28169), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_16_ ( 
        .D(n28170), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_17_ ( 
        .D(n28171), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_18_ ( 
        .D(n28172), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_20_ ( 
        .D(n28174), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_21_ ( 
        .D(n28175), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_22_ ( 
        .D(n28176), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_23_ ( 
        .D(n28177), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_24_ ( 
        .D(n28178), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_24_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_25_ ( 
        .D(n28179), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_25_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_27_ ( 
        .D(n28181), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_28_ ( 
        .D(n28182), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_29_ ( 
        .D(n28183), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_30_ ( 
        .D(n28184), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_31_ ( 
        .D(n28185), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_32_ ( 
        .D(n28186), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_32_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_33_ ( 
        .D(n28187), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_33_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_34_ ( 
        .D(n28188), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_35_ ( 
        .D(n28189), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_35_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_36_ ( 
        .D(n28190), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_36_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_37_ ( 
        .D(n28191), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_37_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_38_ ( 
        .D(n28208), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_40_ ( 
        .D(n28193), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_41_ ( 
        .D(n28194), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_42_ ( 
        .D(n28195), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_44_ ( 
        .D(n28196), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_46_ ( 
        .D(n28206), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_1_ ( 
        .D(n27028), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_2_ ( 
        .D(n27029), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_3_ ( 
        .D(n27030), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_4_ ( 
        .D(n27031), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_5_ ( 
        .D(n27032), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_7_ ( 
        .D(n27034), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_8_ ( 
        .D(n27035), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_9_ ( 
        .D(n27036), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_reg_1_ ( 
        .D(n78376), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_reg_2_ ( 
        .D(n78379), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_reg_3_ ( 
        .D(n78370), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_reg_4_ ( 
        .D(n78381), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_reg_7_ ( 
        .D(n78383), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_reg_0_ ( 
        .D(n78373), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_reg_1_ ( 
        .D(n78375), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_reg_2_ ( 
        .D(n78378), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_reg_3_ ( 
        .D(n78371), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_reg_4_ ( 
        .D(n78380), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_reg_5_ ( 
        .D(n78360), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_reg_6_ ( 
        .D(n78362), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_reg_7_ ( 
        .D(n78382), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_0_ ( 
        .D(n78329), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_1_ ( 
        .D(n78330), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_2_ ( 
        .D(n78331), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_3_ ( 
        .D(n78332), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_4_ ( 
        .D(n78334), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_5_ ( 
        .D(n78336), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_6_ ( 
        .D(n78338), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_7_ ( 
        .D(n78340), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_8_ ( 
        .D(n78342), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_9_ ( 
        .D(n78344), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_10_ ( 
        .D(n78348), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_11_ ( 
        .D(n78346), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_12_ ( 
        .D(n78350), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_13_ ( 
        .D(n78428), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_14_ ( 
        .D(n78427), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_15_ ( 
        .D(n78426), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_16_ ( 
        .D(n78425), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_17_ ( 
        .D(n78424), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_18_ ( 
        .D(n78354), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_19_ ( 
        .D(n78356), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_20_ ( 
        .D(n78368), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_21_ ( 
        .D(n78366), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_reg_22_ ( 
        .D(n78364), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_1_ ( 
        .D(n78434), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_3_ ( 
        .D(n78333), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_4_ ( 
        .D(n78335), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_5_ ( 
        .D(n78337), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_7_ ( 
        .D(n78341), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_8_ ( 
        .D(n78343), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_9_ ( 
        .D(n78345), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_10_ ( 
        .D(n78349), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_11_ ( 
        .D(n78347), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_12_ ( 
        .D(n78351), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_13_ ( 
        .D(n78352), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_14_ ( 
        .D(n78432), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_15_ ( 
        .D(n78353), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_16_ ( 
        .D(n78431), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_17_ ( 
        .D(n78430), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_18_ ( 
        .D(n78355), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_19_ ( 
        .D(n78357), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_20_ ( 
        .D(n78369), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_21_ ( 
        .D(n78367), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_reg_22_ ( 
        .D(n78365), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_sign_i_reg ( 
        .D(n28160), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_output_o_31_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_reg_0_ ( 
        .D(n78248), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_reg_1_ ( 
        .D(n78249), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_1_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_sign_o_reg ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n254), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_sign) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_7_ ( 
        .D(n78419), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[7]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_8_ ( 
        .D(n78418), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[8]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_9_ ( 
        .D(n78417), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[9]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_10_ ( 
        .D(n78416), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[10]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_11_ ( 
        .D(n78415), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[11]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_12_ ( 
        .D(n78414), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[12]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_13_ ( 
        .D(n78413), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[13]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_14_ ( 
        .D(n78412), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[14]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_15_ ( 
        .D(n78411), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[15]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_16_ ( 
        .D(n78410), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[16]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_17_ ( 
        .D(n78409), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[17]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_18_ ( 
        .D(n78408), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[18]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_19_ ( 
        .D(n78407), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[19]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_20_ ( 
        .D(n78406), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[20]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_21_ ( 
        .D(n78405), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[21]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_22_ ( 
        .D(n78404), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[22]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_23_ ( 
        .D(n78403), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[23]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_24_ ( 
        .D(n78402), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[24]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_25_ ( 
        .D(n78401), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[25]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_26_ ( 
        .D(n78400), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[26]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_27_ ( 
        .D(n78227), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[27]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_28_ ( 
        .D(n78399), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[28]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_29_ ( 
        .D(n78398), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[29]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_30_ ( 
        .D(n78397), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[30]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_31_ ( 
        .D(n78226), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[31]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_32_ ( 
        .D(n78396), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[32]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_33_ ( 
        .D(n78395), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[33]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_34_ ( 
        .D(n78225), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[34]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_35_ ( 
        .D(n78394), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[35]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_36_ ( 
        .D(n78393), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[36]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_37_ ( 
        .D(n78392), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[37]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_40_ ( 
        .D(n78390), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[40]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_41_ ( 
        .D(n78389), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[41]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_42_ ( 
        .D(n78388), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[42]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_44_ ( 
        .D(n78386), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[44]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_45_ ( 
        .D(n78385), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[45]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_0_ ( 
        .D(n78421), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[0]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_1_ ( 
        .D(n28210), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[1]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_2_ ( 
        .D(n78228), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[2]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_3_ ( 
        .D(n78423), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[3]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_4_ ( 
        .D(n28213), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[4]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_5_ ( 
        .D(n78422), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[5]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_6_ ( 
        .D(n78420), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[6]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_43_ ( 
        .D(n78387), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[43]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_46_ ( 
        .D(n78384), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[46]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_47_ ( 
        .D(n28256), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[47]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_38_ ( 
        .D(n78391), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[38]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n103), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n106), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n109), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n112), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n115), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n118), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n121), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_7_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n124), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_8_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n127), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_9_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n130), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_10_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n133), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_11_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n136), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_12_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n139), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_13_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n142), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_14_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n145), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_15_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n148), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_16_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n151), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_17_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n154), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n157), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_19_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n160), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_20_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n163), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_21_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n166), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n169), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_23_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n172), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_24_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n175), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_24_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_25_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n178), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_25_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_26_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n181), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_26_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_27_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n184), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_27_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_28_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n187), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_28_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_29_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n190), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_29_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_31_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n196), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_31_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_32_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n199), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_32_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_33_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n202), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_33_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_34_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n205), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_34_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_35_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n208), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_35_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_36_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n211), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_36_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_37_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n214), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_37_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_38_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n217), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_38_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_40_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n223), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_40_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_41_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n226), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_41_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_42_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n229), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_42_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_43_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n232), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_43_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_44_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n235), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_44_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_45_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n238), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_45_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_46_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n241), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_46_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_47_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n244), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_47_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n249), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_start_i_reg ( 
        .D(n78245), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_start_i) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_0_ ( 
        .D(n78329), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_1_ ( 
        .D(n78330), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_2_ ( 
        .D(n78331), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_3_ ( 
        .D(n78332), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_4_ ( 
        .D(n78334), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_5_ ( 
        .D(n78336), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_6_ ( 
        .D(n78338), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_7_ ( 
        .D(n78340), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_8_ ( 
        .D(n78342), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_9_ ( 
        .D(n78344), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_10_ ( 
        .D(n78348), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_11_ ( 
        .D(n78346), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_12_ ( 
        .D(n78350), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_13_ ( 
        .D(n78428), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_14_ ( 
        .D(n78427), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_15_ ( 
        .D(n78426), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_16_ ( 
        .D(n78425), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_17_ ( 
        .D(n78424), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_18_ ( 
        .D(n78354), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_19_ ( 
        .D(n78356), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_20_ ( 
        .D(n78368), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_21_ ( 
        .D(n78366), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_22_ ( 
        .D(n78364), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i_reg_23_ ( 
        .D(n78243), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_0_ ( 
        .D(n78429), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_1_ ( 
        .D(n78434), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_2_ ( 
        .D(n78433), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[2]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_3_ ( 
        .D(n78333), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[3]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_4_ ( 
        .D(n78335), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_5_ ( 
        .D(n78337), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_6_ ( 
        .D(n78339), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[6]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_7_ ( 
        .D(n78341), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[7]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_8_ ( 
        .D(n78343), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[8]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_9_ ( 
        .D(n78345), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[9]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_10_ ( 
        .D(n78349), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[10]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_11_ ( 
        .D(n78347), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[11]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_12_ ( 
        .D(n78351), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[12]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_13_ ( 
        .D(n78352), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[13]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_14_ ( 
        .D(n78432), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[14]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_15_ ( 
        .D(n78353), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[15]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_16_ ( 
        .D(n78431), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[16]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_17_ ( 
        .D(n78430), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[17]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_18_ ( 
        .D(n78355), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[18]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_19_ ( 
        .D(n78357), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[19]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_20_ ( 
        .D(n78369), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[20]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_21_ ( 
        .D(n78367), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_22_ ( 
        .D(n78365), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[22]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i_reg_23_ ( 
        .D(n78244), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[23]) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n1), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n2), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n3), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n4), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n5), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n6), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n7), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_reg_7_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n8), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n11), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n12), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n13), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n14), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n15), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_7_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n16), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_8_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n17), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_9_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n18), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_10_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n19), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_11_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n20), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_12_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n21), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_13_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n22), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_14_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n23), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_15_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n24), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_16_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n25), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_17_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n26), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n27), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_19_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n28), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_20_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n29), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_21_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n30), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n31), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n32), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n33), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n34), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n35), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n36), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n37), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_6_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n38), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_6_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_7_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n39), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_7_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_8_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n40), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_8_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_9_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n41), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_9_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_10_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n42), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_10_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_11_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n43), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_11_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_12_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n44), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_12_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_13_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n45), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_13_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_14_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n46), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_14_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_15_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n47), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_15_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_16_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n48), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_16_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_17_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n49), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_18_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n50), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_18_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_19_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n51), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_19_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_20_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n52), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_20_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_21_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n53), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_21_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_22_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n54), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_22_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_23_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n55), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_reg_24_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n56), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_24_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_in_00_reg ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n57), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_in_00) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n58), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_N398) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n59), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n60), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n61), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n62), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n63), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_5_) );
  OAI21xp33_ASAP7_75t_SL U8688 ( .A1(n4093), .A2(n57189), .B(n8750), .Y(
        icbiu_adr_ic_word[2]) );
  OAI21xp33_ASAP7_75t_SL U9557 ( .A1(n4317), .A2(n1345), .B(n6739), .Y(
        sbbiu_adr_sb[2]) );
  OAI21xp33_ASAP7_75t_SL U9560 ( .A1(n4317), .A2(n1343), .B(n6731), .Y(
        sbbiu_adr_sb[3]) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1_reg ( 
        .D(n78328), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_start_i_reg ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_s_start_i), .CLK(clk_i), .QN(n2456)
         );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_20_ ( 
        .D(n78239), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_21_ ( 
        .D(n78240), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_13_ ( 
        .D(n27477), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_19_ ( 
        .D(n1634), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n123), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n121), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n122), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n124), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_3_ ( 
        .D(n28201), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_12_ ( 
        .D(n28166), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_19_ ( 
        .D(n28173), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_26_ ( 
        .D(n28180), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_39_ ( 
        .D(n28192), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_43_ ( 
        .D(n28205), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_reg_45_ ( 
        .D(n28197), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n250), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1_reg_3_ ( 
        .D(n1525), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shr1_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_N190), .CLK(
        clk_i), .QN(n3309) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1_reg_0_ ( 
        .D(n1528), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[0]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1_reg_1_ ( 
        .D(n1527), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[1]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1_reg_4_ ( 
        .D(n1524), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n119), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_reg_3_ ( 
        .D(n27980), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_r_reg_0_ ( .D(n2529), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_op_r_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_reg_4_ ( 
        .D(n3164), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_op_r_reg_1_ ( .D(n2511), 
        .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_op_r_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n116), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_reg_0_ ( 
        .D(n3168), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n117), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in_reg_5_ ( 
        .D(n78360), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_reg_0_ ( 
        .D(n52526), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_28_ ( 
        .D(n52484), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n114), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n115), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_reg_1_ ( 
        .D(n27982), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_30_ ( 
        .D(n1763), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_17_ ( 
        .D(n78430), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_17_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_43_ ( 
        .D(n1560), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_42_ ( 
        .D(n1581), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_41_ ( 
        .D(n1599), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_reg_0_ ( 
        .D(n27027), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_0_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_24_ ( 
        .D(n59530), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_28_ ( 
        .D(n59574), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_26_ ( 
        .D(n59528), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_29_ ( 
        .D(n59575), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_27_ ( 
        .D(n59573), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_23_ ( 
        .D(n1563), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r_reg_6_ ( 
        .D(n2475), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[6]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_23_ ( 
        .D(n59563), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f_reg_21_ ( 
        .D(n1991), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r_reg_3_ ( 
        .D(n1559), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[3]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_8_ ( 
        .D(n59569), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_8_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_30_ ( 
        .D(n59550), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_30_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_26_ ( 
        .D(n1571), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_0_ ( .D(
        n59710), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[0]) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_reg_25_ ( 
        .D(n59529), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_7_ ( 
        .D(n78341), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_7_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_10_ ( 
        .D(n57500), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[10]) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_reg_5_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n125), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_1_ ( 
        .D(n78434), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_1_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_reg_0_ ( 
        .D(n78429), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_0_) );
  ASYNC_DFFHx1_ASAP7_75t_SRAM or1200_cpu_or1200_if_if_bypass_reg_reg ( .D(
        or1200_cpu_or1200_if_if_bypass), .CLK(clk_i), .RESET(n53192), .SET(
        rst_i), .QN(n3119) );
  DFFHQNx3_ASAP7_75t_SL or1200_cpu_or1200_rf_addra_last_reg_2_ ( .D(
        or1200_cpu_or1200_rf_n9), .CLK(clk_i), .QN(
        or1200_cpu_or1200_rf_addra_last_2_) );
  DFFHQNx3_ASAP7_75t_SL or1200_cpu_or1200_rf_addra_last_reg_4_ ( .D(
        or1200_cpu_or1200_rf_n7), .CLK(clk_i), .QN(
        or1200_cpu_or1200_rf_addra_last_4_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n251), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_) );
  DFFHQNx3_ASAP7_75t_SL or1200_cpu_or1200_rf_addra_last_reg_1_ ( .D(
        or1200_cpu_or1200_rf_n10), .CLK(clk_i), .QN(
        or1200_cpu_or1200_rf_addra_last_1_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_reg_2_ ( 
        .D(n27981), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_reg_3_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n252), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_3_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_0_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n9), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_0_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_reg_1_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n10), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_1_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_reg_3_ ( 
        .D(n9560), .CLK(clk_i), .QN(n2450) );
  ASYNC_DFFHx1_ASAP7_75t_SRAM or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_54_ ( 
        .D(n52001), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n174) );
  AND2x2_ASAP7_75t_SRAM or1200_cpu_or1200_rf_C164 ( .A(or1200_cpu_rf_rdb), .B(
        n78440), .Y(or1200_cpu_or1200_rf_rf_enb) );
  DFFHQNx3_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_30_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n193), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_30_) );
  DFFHQNx1_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_fract_o_reg_39_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_39_), .CLK(clk_i), 
        .QN(n28192) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_state_reg ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n253), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_state) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_reg_2_ ( 
        .D(n3166), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_reg_4_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n118), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_reg_3_ ( 
        .D(n3165), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_rf_addra_last_reg_3_ ( .D(
        or1200_cpu_or1200_rf_n8), .CLK(clk_i), .QN(
        or1200_cpu_or1200_rf_addra_last_3_) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_reg_25_ ( .D(
        n1588), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_)
         );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_reg_26_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[26]), .CLK(clk_i), 
        .QN(DP_OP_741J1_129_6992_n46) );
  DFFHQNx1_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_reg_2_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n248), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_2_) );
  DFFHQNx3_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_reg_39_ ( 
        .D(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n220), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_39_) );
  ASYNC_DFFHx1_ASAP7_75t_SRAM or1200_immu_top_icpu_vpn_r_reg_13_ ( .D(
        icqmem_adr_qmem[13]), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        n825) );
  DFFHQNx2_ASAP7_75t_SL or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1_reg_2_ ( 
        .D(n1526), .CLK(clk_i), .QN(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]) );
  DFFHQNx2_ASAP7_75t_SRAM or1200_cpu_or1200_fpu_fpu_intfloat_conv_out_reg_23_ ( 
        .D(n78198), .CLK(clk_i), .QN(or1200_cpu_or1200_fpu_result_conv[23]) );
  ASYNC_DFFHx1_ASAP7_75t_SRAM or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_p0_reg_55_ ( 
        .D(n52007), .CLK(clk_i), .RESET(n53192), .SET(rst_i), .QN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_n176) );
  TIELOx1_ASAP7_75t_SL U45068 ( .L(n53192) );
  TIEHIx1_ASAP7_75t_SL U45069 ( .H(n53628) );
  A2O1A1Ixp33_ASAP7_75t_SL U45070 ( .A1(n70077), .A2(n53628), .B(n69823), .C(
        n53628), .Y(n56824) );
  A2O1A1Ixp33_ASAP7_75t_SL U45071 ( .A1(n74839), .A2(n53628), .B(n56809), .C(
        n53628), .Y(n56810) );
  A2O1A1Ixp33_ASAP7_75t_SL U45072 ( .A1(n74745), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_1_), .C(n53628), .Y(
        n56811) );
  A2O1A1Ixp33_ASAP7_75t_SL U45073 ( .A1(n2491), .A2(n53628), .B(n56811), .C(
        n53628), .Y(n56812) );
  A2O1A1Ixp33_ASAP7_75t_SL U45074 ( .A1(n56810), .A2(n53628), .B(n56812), .C(
        n53628), .Y(n56813) );
  A2O1A1Ixp33_ASAP7_75t_SL U45075 ( .A1(n74766), .A2(n53628), .B(n74747), .C(
        n53628), .Y(n56814) );
  A2O1A1Ixp33_ASAP7_75t_SL U45076 ( .A1(n56814), .A2(n53628), .B(n56809), .C(
        n53628), .Y(n56815) );
  A2O1A1Ixp33_ASAP7_75t_SL U45077 ( .A1(n74746), .A2(n53628), .B(n56815), .C(
        n74748), .Y(n56816) );
  A2O1A1Ixp33_ASAP7_75t_SL U45078 ( .A1(n74750), .A2(n53628), .B(n74749), .C(
        n53628), .Y(n56817) );
  O2A1O1Ixp33_ASAP7_75t_SL U45079 ( .A1(n74894), .A2(n76977), .B(n53628), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_in_00), .Y(n56818) );
  A2O1A1Ixp33_ASAP7_75t_SL U45080 ( .A1(n56813), .A2(n53628), .B(n56820), .C(
        n56821), .Y(n3142) );
  O2A1O1Ixp5_ASAP7_75t_SL U45081 ( .A1(n60462), .A2(n61044), .B(n53628), .C(
        n58282), .Y(n56639) );
  A2O1A1Ixp33_ASAP7_75t_SL U45082 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[11]), .A2(
        n53628), .B(n57190), .C(n56808), .Y(n3112) );
  A2O1A1Ixp33_ASAP7_75t_SL U45083 ( .A1(n53628), .A2(n3076), .B(n77567), .C(
        n56633), .Y(n9459) );
  A2O1A1Ixp33_ASAP7_75t_SL U45084 ( .A1(or1200_cpu_or1200_except_n583), .A2(
        n3390), .B(n76579), .C(n53628), .Y(n56806) );
  A2O1A1Ixp33_ASAP7_75t_SL U45085 ( .A1(n59689), .A2(n53628), .B(n3063), .C(
        n56807), .Y(n3064) );
  A2O1A1Ixp33_ASAP7_75t_SL U45086 ( .A1(n57074), .A2(n53628), .B(n3054), .C(
        n56805), .Y(n3055) );
  A2O1A1Ixp33_ASAP7_75t_SL U45087 ( .A1(n59689), .A2(n53628), .B(n3048), .C(
        n56804), .Y(n3049) );
  A2O1A1Ixp33_ASAP7_75t_SL U45088 ( .A1(n63977), .A2(n53628), .B(n63975), .C(
        n53628), .Y(n56802) );
  A2O1A1Ixp33_ASAP7_75t_SL U45089 ( .A1(n59688), .A2(n53628), .B(n3027), .C(
        n56803), .Y(n3028) );
  A2O1A1Ixp33_ASAP7_75t_SL U45090 ( .A1(n59689), .A2(n53628), .B(n3021), .C(
        n56801), .Y(n3022) );
  A2O1A1Ixp33_ASAP7_75t_SL U45091 ( .A1(n59688), .A2(n53628), .B(n3015), .C(
        n56800), .Y(n3016) );
  A2O1A1Ixp33_ASAP7_75t_SL U45092 ( .A1(n53628), .A2(n57074), .B(n3009), .C(
        n55690), .Y(n3010) );
  A2O1A1Ixp33_ASAP7_75t_SL U45093 ( .A1(n76658), .A2(n53628), .B(n76660), .C(
        n53628), .Y(n56798) );
  A2O1A1Ixp33_ASAP7_75t_SL U45094 ( .A1(n76657), .A2(n53628), .B(n76665), .C(
        n77210), .Y(n56799) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45095 ( .A1(n58296), .A2(n77922), .B(n56798), 
        .C(n53628), .D(n56799), .Y(n2967) );
  A2O1A1Ixp33_ASAP7_75t_SL U45096 ( .A1(n75616), .A2(n53628), .B(n2966), .C(
        n56797), .Y(n9326) );
  A2O1A1Ixp33_ASAP7_75t_SL U45097 ( .A1(n2958), .A2(n53628), .B(n57074), .C(
        n56796), .Y(n2959) );
  A2O1A1Ixp33_ASAP7_75t_SL U45098 ( .A1(n53628), .A2(n57074), .B(n2821), .C(
        n56616), .Y(n2822) );
  A2O1A1Ixp33_ASAP7_75t_SL U45099 ( .A1(ex_insn[28]), .A2(n53628), .B(n77567), 
        .C(n56792), .Y(n2811) );
  A2O1A1Ixp33_ASAP7_75t_SL U45100 ( .A1(n53628), .A2(n77246), .B(n2798), .C(
        n56614), .Y(n9334) );
  A2O1A1Ixp33_ASAP7_75t_SL U45101 ( .A1(n53628), .A2(n77399), .B(n56610), .C(
        n58280), .Y(n9471) );
  A2O1A1Ixp33_ASAP7_75t_SL U45102 ( .A1(n53628), .A2(n59689), .B(n2572), .C(
        n56606), .Y(n2573) );
  A2O1A1Ixp33_ASAP7_75t_SL U45103 ( .A1(n53628), .A2(n2514), .B(n57073), .C(
        n54690), .Y(n2515) );
  A2O1A1Ixp33_ASAP7_75t_SL U45104 ( .A1(n53628), .A2(n2496), .B(n57074), .C(
        n56605), .Y(n2497) );
  A2O1A1Ixp33_ASAP7_75t_SL U45105 ( .A1(n69377), .A2(n53628), .B(n70526), .C(
        n56791), .Y(n2454) );
  A2O1A1Ixp33_ASAP7_75t_SL U45106 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_5_), .A2(
        n53628), .B(n56790), .C(n74369), .Y(n2379) );
  A2O1A1Ixp33_ASAP7_75t_SL U45107 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[1]), .A2(n70502), .B(
        n70503), .C(n53628), .Y(n56786) );
  A2O1A1Ixp33_ASAP7_75t_SL U45108 ( .A1(n69750), .A2(n69749), .B(n69754), .C(
        n53628), .Y(n56783) );
  A2O1A1Ixp33_ASAP7_75t_SL U45109 ( .A1(n69752), .A2(n53628), .B(n57081), .C(
        n56784), .Y(n56785) );
  A2O1A1Ixp33_ASAP7_75t_SL U45110 ( .A1(n59621), .A2(n56783), .B(n56785), .C(
        n53628), .Y(n2305) );
  A2O1A1Ixp33_ASAP7_75t_SL U45111 ( .A1(n69911), .A2(n53628), .B(n56777), .C(
        n53628), .Y(n56778) );
  A2O1A1Ixp33_ASAP7_75t_SL U45112 ( .A1(n70502), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[16]), .B(n59621), .C(
        n53628), .Y(n56779) );
  A2O1A1Ixp33_ASAP7_75t_SL U45113 ( .A1(n53628), .A2(n2145), .B(n57073), .C(
        n55222), .Y(n2146) );
  A2O1A1Ixp33_ASAP7_75t_SL U45114 ( .A1(n53628), .A2(n2131), .B(n57073), .C(
        n56574), .Y(n2132) );
  A2O1A1Ixp33_ASAP7_75t_SL U45115 ( .A1(n53628), .A2(n59564), .B(n57073), .C(
        n56091), .Y(n9669) );
  A2O1A1Ixp33_ASAP7_75t_SL U45116 ( .A1(n77246), .A2(n53628), .B(n1983), .C(
        n56776), .Y(n9340) );
  A2O1A1Ixp33_ASAP7_75t_SL U45117 ( .A1(n53628), .A2(n77246), .B(n1978), .C(
        n56573), .Y(n9338) );
  A2O1A1Ixp33_ASAP7_75t_SL U45118 ( .A1(n53628), .A2(n77246), .B(n1961), .C(
        n56572), .Y(n9335) );
  A2O1A1Ixp33_ASAP7_75t_SL U45119 ( .A1(n53628), .A2(n77246), .B(n1945), .C(
        n56571), .Y(n9333) );
  A2O1A1Ixp33_ASAP7_75t_SL U45120 ( .A1(n53628), .A2(n59680), .B(n1824), .C(
        n56567), .Y(or1200_du_N104) );
  A2O1A1Ixp33_ASAP7_75t_SL U45121 ( .A1(n53628), .A2(n77246), .B(n1798), .C(
        n56300), .Y(n9331) );
  A2O1A1Ixp33_ASAP7_75t_SL U45122 ( .A1(n74934), .A2(n53628), .B(n59708), .C(
        n56775), .Y(n9493) );
  A2O1A1Ixp33_ASAP7_75t_SL U45123 ( .A1(n77667), .A2(n53628), .B(n56772), .C(
        n53628), .Y(n56773) );
  A2O1A1Ixp33_ASAP7_75t_SL U45124 ( .A1(n77862), .A2(n77672), .B(n56773), .C(
        n53628), .Y(n1699) );
  A2O1A1Ixp33_ASAP7_75t_SL U45125 ( .A1(n57114), .A2(n53628), .B(n1476), .C(
        n56770), .Y(n9302) );
  A2O1A1Ixp33_ASAP7_75t_SL U45126 ( .A1(n57114), .A2(n53628), .B(n1430), .C(
        n56769), .Y(n9279) );
  A2O1A1Ixp33_ASAP7_75t_SL U45127 ( .A1(n57114), .A2(n53628), .B(n1428), .C(
        n56768), .Y(n9278) );
  A2O1A1Ixp33_ASAP7_75t_SL U45128 ( .A1(n53628), .A2(n74641), .B(n1382), .C(
        n55213), .Y(n9315) );
  A2O1A1Ixp33_ASAP7_75t_SL U45129 ( .A1(n74641), .A2(n53628), .B(n1374), .C(
        n56767), .Y(n9313) );
  A2O1A1Ixp33_ASAP7_75t_SL U45130 ( .A1(n53628), .A2(n74641), .B(n1370), .C(
        n54314), .Y(n9312) );
  A2O1A1Ixp33_ASAP7_75t_SL U45131 ( .A1(n1295), .A2(n53628), .B(n4317), .C(
        n53628), .Y(n56765) );
  A2O1A1Ixp33_ASAP7_75t_SL U45132 ( .A1(n57083), .A2(n53628), .B(n1292), .C(
        n56766), .Y(n1293) );
  A2O1A1Ixp33_ASAP7_75t_SL U45133 ( .A1(n76530), .A2(n53628), .B(n56762), .C(
        n53628), .Y(n56763) );
  A2O1A1Ixp33_ASAP7_75t_SL U45134 ( .A1(n76521), .A2(dbg_dat_i[11]), .B(n56763), .C(n53628), .Y(n56764) );
  A2O1A1Ixp33_ASAP7_75t_SL U45135 ( .A1(n1106), .A2(n53628), .B(n76523), .C(
        n56764), .Y(n9185) );
  A2O1A1Ixp33_ASAP7_75t_SL U45136 ( .A1(n59703), .A2(n53628), .B(n56761), .C(
        n53628), .Y(or1200_immu_top_N34) );
  A2O1A1Ixp33_ASAP7_75t_SL U45137 ( .A1(n59703), .A2(n53628), .B(n56760), .C(
        n53628), .Y(n51954) );
  A2O1A1Ixp33_ASAP7_75t_SL U45138 ( .A1(n59703), .A2(n53628), .B(n56759), .C(
        n53628), .Y(or1200_immu_top_N30) );
  A2O1A1Ixp33_ASAP7_75t_SL U45139 ( .A1(n59703), .A2(n53628), .B(n56758), .C(
        n53628), .Y(or1200_immu_top_N29) );
  A2O1A1Ixp33_ASAP7_75t_SL U45140 ( .A1(n59703), .A2(n53628), .B(n56757), .C(
        n53628), .Y(or1200_immu_top_N26) );
  A2O1A1Ixp33_ASAP7_75t_SL U45141 ( .A1(n59703), .A2(n53628), .B(n56756), .C(
        n53628), .Y(or1200_immu_top_N25) );
  A2O1A1Ixp33_ASAP7_75t_SL U45142 ( .A1(n59703), .A2(n53628), .B(n56755), .C(
        n53628), .Y(or1200_immu_top_N24) );
  A2O1A1Ixp33_ASAP7_75t_SL U45143 ( .A1(n59703), .A2(n53628), .B(n56754), .C(
        n53628), .Y(n51948) );
  O2A1O1Ixp33_ASAP7_75t_SL U45144 ( .A1(n58389), .A2(n68858), .B(n53628), .C(
        n68859), .Y(n56753) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45145 ( .A1(n68856), .A2(n56752), .B(n56753), 
        .C(n53628), .D(n68855), .Y(n51991) );
  A2O1A1Ixp33_ASAP7_75t_SL U45146 ( .A1(n53628), .A2(n65106), .B(n64699), .C(
        n57332), .Y(n56511) );
  A2O1A1Ixp33_ASAP7_75t_SL U45147 ( .A1(or1200_cpu_or1200_mult_mac_n14), .A2(
        n53628), .B(n57105), .C(n56749), .Y(or1200_cpu_or1200_mult_mac_n1502)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45148 ( .A1(n53628), .A2(
        or1200_cpu_or1200_mult_mac_n76), .B(n57105), .C(n56502), .Y(
        or1200_cpu_or1200_mult_mac_n1534) );
  A2O1A1Ixp33_ASAP7_75t_SL U45149 ( .A1(n57105), .A2(n53628), .B(
        or1200_cpu_or1200_mult_mac_n98), .C(n53628), .Y(n56743) );
  A2O1A1Ixp33_ASAP7_75t_SL U45150 ( .A1(n57348), .A2(n56742), .B(n56743), .C(
        n53628), .Y(n56744) );
  A2O1A1Ixp33_ASAP7_75t_SL U45151 ( .A1(n57077), .A2(n53628), .B(
        or1200_cpu_or1200_mult_mac_n100), .C(n56744), .Y(n12970) );
  A2O1A1Ixp33_ASAP7_75t_SL U45152 ( .A1(n53628), .A2(
        or1200_cpu_or1200_mult_mac_n108), .B(n57105), .C(n56499), .Y(
        or1200_cpu_or1200_mult_mac_n1550) );
  A2O1A1Ixp33_ASAP7_75t_SL U45153 ( .A1(n65164), .A2(n53628), .B(n56732), .C(
        n53628), .Y(n56733) );
  A2O1A1Ixp33_ASAP7_75t_SL U45154 ( .A1(n74045), .A2(n53628), .B(n65182), .C(
        n53628), .Y(n56734) );
  A2O1A1Ixp33_ASAP7_75t_SL U45155 ( .A1(or1200_cpu_or1200_mult_mac_n189), .A2(
        n53628), .B(n76889), .C(n56741), .Y(or1200_cpu_or1200_mult_mac_n1569)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45156 ( .A1(n53628), .A2(n69125), .B(n59671), .C(
        n54629), .Y(n54630) );
  A2O1A1Ixp33_ASAP7_75t_SL U45157 ( .A1(n69198), .A2(n53628), .B(n69197), .C(
        n57080), .Y(n56726) );
  A2O1A1Ixp33_ASAP7_75t_SL U45158 ( .A1(n56725), .A2(n53628), .B(n56726), .C(
        n56731), .Y(or1200_cpu_or1200_mult_mac_n1606) );
  A2O1A1Ixp33_ASAP7_75t_SL U45159 ( .A1(n75512), .A2(n53628), .B(n56724), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_N290) );
  A2O1A1Ixp33_ASAP7_75t_SL U45160 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n302), .C(n56485), .Y(
        or1200_cpu_or1200_except_n303) );
  A2O1A1Ixp33_ASAP7_75t_SL U45161 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n305), .C(n56484), .Y(
        or1200_cpu_or1200_except_n306) );
  A2O1A1Ixp33_ASAP7_75t_SL U45162 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n308), .C(n56483), .Y(
        or1200_cpu_or1200_except_n309) );
  A2O1A1Ixp33_ASAP7_75t_SL U45163 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n311), .C(n56482), .Y(
        or1200_cpu_or1200_except_n312) );
  A2O1A1Ixp33_ASAP7_75t_SL U45164 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n314), .C(n56481), .Y(
        or1200_cpu_or1200_except_n315) );
  A2O1A1Ixp33_ASAP7_75t_SL U45165 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n317), .C(n56480), .Y(
        or1200_cpu_or1200_except_n318) );
  A2O1A1Ixp33_ASAP7_75t_SL U45166 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n320), .C(n56479), .Y(
        or1200_cpu_or1200_except_n321) );
  A2O1A1Ixp33_ASAP7_75t_SL U45167 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n323), .C(n56478), .Y(
        or1200_cpu_or1200_except_n324) );
  A2O1A1Ixp33_ASAP7_75t_SL U45168 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n326), .C(n56477), .Y(
        or1200_cpu_or1200_except_n327) );
  A2O1A1Ixp33_ASAP7_75t_SL U45169 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n329), .C(n56476), .Y(
        or1200_cpu_or1200_except_n330) );
  A2O1A1Ixp33_ASAP7_75t_SL U45170 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n332), .C(n56475), .Y(
        or1200_cpu_or1200_except_n333) );
  A2O1A1Ixp33_ASAP7_75t_SL U45171 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n335), .C(n56474), .Y(
        or1200_cpu_or1200_except_n336) );
  A2O1A1Ixp33_ASAP7_75t_SL U45172 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n338), .C(n56473), .Y(
        or1200_cpu_or1200_except_n339) );
  A2O1A1Ixp33_ASAP7_75t_SL U45173 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n341), .C(n56472), .Y(
        or1200_cpu_or1200_except_n342) );
  A2O1A1Ixp33_ASAP7_75t_SL U45174 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n344), .C(n56471), .Y(
        or1200_cpu_or1200_except_n345) );
  A2O1A1Ixp33_ASAP7_75t_SL U45175 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n347), .C(n56470), .Y(
        or1200_cpu_or1200_except_n348) );
  A2O1A1Ixp33_ASAP7_75t_SL U45176 ( .A1(n53628), .A2(n57074), .B(
        or1200_cpu_or1200_except_n350), .C(n56469), .Y(
        or1200_cpu_or1200_except_n351) );
  A2O1A1Ixp33_ASAP7_75t_SL U45177 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n353), .C(n56468), .Y(
        or1200_cpu_or1200_except_n354) );
  A2O1A1Ixp33_ASAP7_75t_SL U45178 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n356), .C(n56722), .Y(
        or1200_cpu_or1200_except_n357) );
  A2O1A1Ixp33_ASAP7_75t_SL U45179 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n359), .C(n56467), .Y(
        or1200_cpu_or1200_except_n360) );
  A2O1A1Ixp33_ASAP7_75t_SL U45180 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n362), .C(n56721), .Y(
        or1200_cpu_or1200_except_n363) );
  A2O1A1Ixp33_ASAP7_75t_SL U45181 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n365), .C(n56466), .Y(
        or1200_cpu_or1200_except_n366) );
  A2O1A1Ixp33_ASAP7_75t_SL U45182 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n368), .C(n56720), .Y(
        or1200_cpu_or1200_except_n369) );
  A2O1A1Ixp33_ASAP7_75t_SL U45183 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n371), .C(n56465), .Y(
        or1200_cpu_or1200_except_n372) );
  A2O1A1Ixp33_ASAP7_75t_SL U45184 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n374), .C(n56719), .Y(
        or1200_cpu_or1200_except_n375) );
  A2O1A1Ixp33_ASAP7_75t_SL U45185 ( .A1(n53628), .A2(n57074), .B(
        or1200_cpu_or1200_except_n377), .C(n56464), .Y(
        or1200_cpu_or1200_except_n378) );
  A2O1A1Ixp33_ASAP7_75t_SL U45186 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n383), .C(n56462), .Y(
        or1200_cpu_or1200_except_n384) );
  A2O1A1Ixp33_ASAP7_75t_SL U45187 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n386), .C(n56461), .Y(
        or1200_cpu_or1200_except_n387) );
  A2O1A1Ixp33_ASAP7_75t_SL U45188 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n389), .C(n56460), .Y(
        or1200_cpu_or1200_except_n390) );
  A2O1A1Ixp33_ASAP7_75t_SL U45189 ( .A1(n74276), .A2(n53628), .B(n56718), .C(
        n74275), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n48) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45190 ( .A1(n72508), .A2(n72504), .B(n53628), 
        .C(n72505), .Y(n56449) );
  A2O1A1Ixp33_ASAP7_75t_SL U45191 ( .A1(n72490), .A2(n72501), .B(n56449), .C(
        n53628), .Y(n56450) );
  A2O1A1Ixp33_ASAP7_75t_SL U45192 ( .A1(n53628), .A2(n72507), .B(n72509), .C(
        n56450), .Y(n56451) );
  A2O1A1Ixp33_ASAP7_75t_SL U45193 ( .A1(n72502), .A2(n56448), .B(n56451), .C(
        n53628), .Y(n56452) );
  A2O1A1Ixp33_ASAP7_75t_SL U45194 ( .A1(n58599), .A2(n72411), .B(n72368), .C(
        n53628), .Y(n56454) );
  A2O1A1Ixp33_ASAP7_75t_SL U45195 ( .A1(n71632), .A2(n53628), .B(n56441), .C(
        n71631), .Y(n56442) );
  A2O1A1Ixp33_ASAP7_75t_SL U45196 ( .A1(n71630), .A2(n53628), .B(n56442), .C(
        n71633), .Y(n56443) );
  A2O1A1Ixp33_ASAP7_75t_SL U45197 ( .A1(n53628), .A2(n71634), .B(n56443), .C(
        n71950), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n136) );
  A2O1A1Ixp33_ASAP7_75t_SL U45198 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_2_), .C(n56436), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n109) );
  A2O1A1Ixp33_ASAP7_75t_SL U45199 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_8_), .C(n56715), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n127) );
  A2O1A1Ixp33_ASAP7_75t_SL U45200 ( .A1(n53320), .A2(n53628), .B(n75942), .C(
        n56714), .Y(n67381) );
  A2O1A1Ixp33_ASAP7_75t_SL U45201 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[15]), .A2(n57217), .B(
        n56711), .C(n53628), .Y(n56712) );
  A2O1A1Ixp33_ASAP7_75t_SL U45202 ( .A1(n70188), .A2(n53628), .B(n56708), .C(
        n70187), .Y(n70195) );
  A2O1A1Ixp33_ASAP7_75t_SL U45203 ( .A1(n70054), .A2(n53628), .B(n78332), .C(
        n53628), .Y(n56702) );
  A2O1A1Ixp33_ASAP7_75t_SL U45204 ( .A1(n70034), .A2(n53628), .B(n78331), .C(
        n53628), .Y(n56703) );
  A2O1A1Ixp33_ASAP7_75t_SL U45205 ( .A1(n78330), .A2(n53628), .B(n70035), .C(
        n53628), .Y(n56704) );
  A2O1A1Ixp33_ASAP7_75t_SL U45206 ( .A1(n56703), .A2(n53628), .B(n56704), .C(
        n53628), .Y(n56705) );
  A2O1A1Ixp33_ASAP7_75t_SL U45207 ( .A1(n56702), .A2(n53628), .B(n56707), .C(
        n53628), .Y(n69904) );
  A2O1A1Ixp33_ASAP7_75t_SL U45208 ( .A1(n61281), .A2(n53628), .B(n77416), .C(
        n53628), .Y(n56701) );
  A2O1A1Ixp33_ASAP7_75t_SL U45209 ( .A1(n65256), .A2(n53628), .B(n65255), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .Y(n56698) );
  A2O1A1Ixp33_ASAP7_75t_SL U45210 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n53628), .B(n70339), .C(n56697), .Y(n70468) );
  A2O1A1Ixp33_ASAP7_75t_SL U45211 ( .A1(n77017), .A2(n53628), .B(n77149), .C(
        n56695), .Y(n78148) );
  A2O1A1Ixp33_ASAP7_75t_SL U45212 ( .A1(n53628), .A2(n69366), .B(n75794), .C(
        n56215), .Y(n78088) );
  A2O1A1Ixp33_ASAP7_75t_SL U45213 ( .A1(n66224), .A2(n53628), .B(n56693), .C(
        n53628), .Y(n75392) );
  A2O1A1Ixp33_ASAP7_75t_SL U45214 ( .A1(n57168), .A2(n53628), .B(n874), .C(
        n53628), .Y(n56692) );
  A2O1A1Ixp33_ASAP7_75t_SL U45215 ( .A1(n56692), .A2(n53628), .B(n63984), .C(
        n53628), .Y(n78261) );
  A2O1A1Ixp33_ASAP7_75t_SL U45216 ( .A1(n57168), .A2(n53628), .B(n1000), .C(
        n53628), .Y(n56691) );
  A2O1A1Ixp33_ASAP7_75t_SL U45217 ( .A1(n56691), .A2(n53628), .B(n75171), .C(
        n53628), .Y(n78262) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45218 ( .A1(n57149), .A2(n75067), .B(n53628), 
        .C(n55530), .Y(n55531) );
  A2O1A1Ixp33_ASAP7_75t_SL U45219 ( .A1(n55533), .A2(n75082), .B(n55534), .C(
        n53628), .Y(n75138) );
  A2O1A1Ixp33_ASAP7_75t_SL U45220 ( .A1(n69303), .A2(n53628), .B(n69302), .C(
        n53628), .Y(n56690) );
  A2O1A1Ixp33_ASAP7_75t_SL U45221 ( .A1(n69305), .A2(n69304), .B(n56690), .C(
        n53628), .Y(n69306) );
  A2O1A1Ixp33_ASAP7_75t_SL U45222 ( .A1(n68757), .A2(n53628), .B(n56688), .C(
        n53628), .Y(n68760) );
  A2O1A1Ixp33_ASAP7_75t_SL U45223 ( .A1(n75989), .A2(n53628), .B(n56686), .C(
        n53628), .Y(n75990) );
  A2O1A1Ixp33_ASAP7_75t_SL U45224 ( .A1(or1200_cpu_or1200_mult_mac_n299), .A2(
        n53628), .B(n56684), .C(n53628), .Y(n63385) );
  A2O1A1Ixp33_ASAP7_75t_SL U45225 ( .A1(n63776), .A2(n53628), .B(n56683), .C(
        n53628), .Y(n63889) );
  A2O1A1Ixp33_ASAP7_75t_SL U45226 ( .A1(n69017), .A2(n53628), .B(n56681), .C(
        n69016), .Y(n69020) );
  A2O1A1Ixp33_ASAP7_75t_SL U45227 ( .A1(or1200_cpu_or1200_mult_mac_n257), .A2(
        n53628), .B(n56680), .C(n53628), .Y(n75133) );
  A2O1A1Ixp33_ASAP7_75t_SL U45228 ( .A1(n59581), .A2(n53628), .B(n77744), .C(
        n53628), .Y(n56678) );
  A2O1A1Ixp33_ASAP7_75t_SL U45229 ( .A1(n59551), .A2(n53628), .B(n77745), .C(
        n53628), .Y(n56679) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45230 ( .A1(n77746), .A2(n78327), .B(n56678), 
        .C(n53628), .D(n56679), .Y(n4240) );
  A2O1A1Ixp33_ASAP7_75t_SL U45231 ( .A1(n77704), .A2(n53628), .B(n59709), .C(
        n56677), .Y(n4302) );
  A2O1A1Ixp33_ASAP7_75t_SL U45232 ( .A1(n57208), .A2(n53628), .B(n71984), .C(
        n53628), .Y(n56671) );
  A2O1A1Ixp33_ASAP7_75t_SL U45233 ( .A1(n56671), .A2(n53628), .B(n56674), .C(
        n53628), .Y(n56675) );
  A2O1A1Ixp33_ASAP7_75t_SL U45234 ( .A1(n71793), .A2(n53628), .B(n56670), .C(
        n53628), .Y(n71791) );
  A2O1A1Ixp33_ASAP7_75t_SL U45235 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_17_), 
        .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_), 
        .C(n53628), .Y(n56669) );
  A2O1A1Ixp33_ASAP7_75t_SL U45236 ( .A1(n70855), .A2(n53628), .B(n70856), .C(
        n53628), .Y(n56668) );
  A2O1A1Ixp33_ASAP7_75t_SL U45237 ( .A1(n53628), .A2(n59562), .B(n65745), .C(
        n55741), .Y(n66119) );
  A2O1A1Ixp33_ASAP7_75t_SL U45238 ( .A1(n66080), .A2(n53628), .B(n65970), .C(
        n53628), .Y(n56666) );
  A2O1A1Ixp33_ASAP7_75t_SL U45239 ( .A1(n65939), .A2(n53628), .B(n65974), .C(
        n53628), .Y(n56667) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45240 ( .A1(n65978), .A2(n66007), .B(n56666), 
        .C(n53628), .D(n56667), .Y(n65991) );
  A2O1A1Ixp33_ASAP7_75t_SL U45241 ( .A1(n53628), .A2(n59630), .B(n73123), .C(
        n56387), .Y(n73322) );
  A2O1A1Ixp33_ASAP7_75t_SL U45242 ( .A1(n73708), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .C(
        n53628), .Y(n56665) );
  A2O1A1Ixp33_ASAP7_75t_SL U45243 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[1]), .B(n56665), .C(
        n53628), .Y(n73739) );
  A2O1A1Ixp33_ASAP7_75t_SL U45244 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_5_), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_4_), .C(n53628), .Y(
        n56664) );
  A2O1A1Ixp33_ASAP7_75t_SL U45245 ( .A1(n2773), .A2(n53628), .B(n56661), .C(
        n53628), .Y(n60277) );
  A2O1A1Ixp33_ASAP7_75t_SL U45246 ( .A1(n75276), .A2(n56378), .B(n56380), .C(
        n53628), .Y(n75280) );
  A2O1A1Ixp33_ASAP7_75t_SL U45247 ( .A1(n69036), .A2(n53628), .B(n69035), .C(
        n69034), .Y(n56658) );
  A2O1A1Ixp33_ASAP7_75t_SL U45248 ( .A1(n56657), .A2(n56658), .B(n69037), .C(
        n53628), .Y(n56659) );
  A2O1A1Ixp33_ASAP7_75t_SL U45249 ( .A1(n69038), .A2(n53628), .B(n56659), .C(
        n53628), .Y(n69040) );
  O2A1O1Ixp5_ASAP7_75t_SL U45250 ( .A1(n71392), .A2(n71391), .B(n53628), .C(
        n56376), .Y(n71397) );
  A2O1A1Ixp33_ASAP7_75t_SL U45251 ( .A1(n69227), .A2(n53628), .B(n69226), .C(
        n53628), .Y(n56656) );
  A2O1A1Ixp33_ASAP7_75t_SL U45252 ( .A1(n69228), .A2(n69227), .B(n56656), .C(
        n53628), .Y(n69230) );
  A2O1A1Ixp33_ASAP7_75t_SL U45253 ( .A1(n73975), .A2(n53628), .B(n73974), .C(
        n53628), .Y(n56654) );
  A2O1A1Ixp33_ASAP7_75t_SL U45254 ( .A1(n73591), .A2(n56365), .B(n73555), .C(
        n53628), .Y(n73551) );
  A2O1A1Ixp33_ASAP7_75t_SL U45255 ( .A1(n59012), .A2(n53628), .B(n64502), .C(
        n56652), .Y(n64541) );
  OAI21xp5_ASAP7_75t_SL U45256 ( .A1(n59283), .A2(n67826), .B(n53628), .Y(
        n56651) );
  A2O1A1Ixp33_ASAP7_75t_SL U45257 ( .A1(n69902), .A2(n53628), .B(n69900), .C(
        n69828), .Y(n56354) );
  A2O1A1Ixp33_ASAP7_75t_SL U45258 ( .A1(n69996), .A2(n69872), .B(n56354), .C(
        n53628), .Y(n56355) );
  A2O1A1Ixp33_ASAP7_75t_SL U45259 ( .A1(n60458), .A2(n53628), .B(n60464), .C(
        n53628), .Y(n56642) );
  A2O1A1Ixp33_ASAP7_75t_SL U45260 ( .A1(n77488), .A2(n53628), .B(n3109), .C(
        n53628), .Y(n56634) );
  A2O1A1Ixp33_ASAP7_75t_SL U45261 ( .A1(n61297), .A2(n53628), .B(n56635), .C(
        n61287), .Y(n56636) );
  A2O1A1Ixp33_ASAP7_75t_SL U45262 ( .A1(n59689), .A2(n53628), .B(n3060), .C(
        n56631), .Y(n3061) );
  A2O1A1Ixp33_ASAP7_75t_SL U45263 ( .A1(n57073), .A2(n53628), .B(n3051), .C(
        n56630), .Y(n3052) );
  A2O1A1Ixp33_ASAP7_75t_SL U45264 ( .A1(n53628), .A2(n59689), .B(n3045), .C(
        n55909), .Y(n3046) );
  A2O1A1Ixp33_ASAP7_75t_SL U45265 ( .A1(n53628), .A2(n57074), .B(n3033), .C(
        n56342), .Y(n3034) );
  A2O1A1Ixp33_ASAP7_75t_SL U45266 ( .A1(n59688), .A2(n53628), .B(n3018), .C(
        n56629), .Y(n3019) );
  A2O1A1Ixp33_ASAP7_75t_SL U45267 ( .A1(n57074), .A2(n53628), .B(n3003), .C(
        n56628), .Y(n3004) );
  A2O1A1Ixp33_ASAP7_75t_SL U45268 ( .A1(n77301), .A2(n53628), .B(n56622), .C(
        n53628), .Y(n51976) );
  A2O1A1Ixp33_ASAP7_75t_SL U45269 ( .A1(n53628), .A2(n57144), .B(n77878), .C(
        n55473), .Y(n2942) );
  A2O1A1Ixp33_ASAP7_75t_SL U45270 ( .A1(n77171), .A2(n53628), .B(n56621), .C(
        n53628), .Y(n52499) );
  A2O1A1Ixp33_ASAP7_75t_SL U45271 ( .A1(n53628), .A2(n57202), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[29]), .C(n56329), 
        .Y(n2869) );
  A2O1A1Ixp33_ASAP7_75t_SL U45272 ( .A1(n53628), .A2(n59627), .B(n72786), .C(
        n56118), .Y(n2838) );
  A2O1A1Ixp33_ASAP7_75t_SL U45273 ( .A1(n53628), .A2(n77246), .B(n2796), .C(
        n56324), .Y(n9330) );
  A2O1A1Ixp33_ASAP7_75t_SL U45274 ( .A1(n2577), .A2(n53628), .B(n77567), .C(
        n56609), .Y(n9494) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45275 ( .A1(n65331), .A2(n55894), .B(n53628), 
        .C(n55895), .Y(n2487) );
  A2O1A1Ixp33_ASAP7_75t_SL U45276 ( .A1(n74677), .A2(n74686), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .C(
        n53628), .Y(n56598) );
  A2O1A1Ixp33_ASAP7_75t_SL U45277 ( .A1(n74706), .A2(n53628), .B(n70544), .C(
        n56601), .Y(n56602) );
  A2O1A1Ixp33_ASAP7_75t_SL U45278 ( .A1(n70553), .A2(n53628), .B(n2448), .C(
        n56603), .Y(n56604) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45279 ( .A1(n70549), .A2(n70550), .B(n56597), 
        .C(n53628), .D(n56604), .Y(n2436) );
  A2O1A1Ixp33_ASAP7_75t_SL U45280 ( .A1(n77301), .A2(n53628), .B(n56595), .C(
        n53628), .Y(n51959) );
  A2O1A1Ixp33_ASAP7_75t_SL U45281 ( .A1(n77301), .A2(n53628), .B(n56594), .C(
        n53628), .Y(n2422) );
  A2O1A1Ixp33_ASAP7_75t_SL U45282 ( .A1(n77301), .A2(n53628), .B(n56593), .C(
        n53628), .Y(n51975) );
  A2O1A1Ixp33_ASAP7_75t_SL U45283 ( .A1(n77301), .A2(n53628), .B(n56592), .C(
        n53628), .Y(n51973) );
  A2O1A1Ixp33_ASAP7_75t_SL U45284 ( .A1(n77301), .A2(n53628), .B(n56591), .C(
        n53628), .Y(n2377) );
  A2O1A1Ixp33_ASAP7_75t_SL U45285 ( .A1(n77301), .A2(n53628), .B(n56590), .C(
        n53628), .Y(n51972) );
  A2O1A1Ixp33_ASAP7_75t_SL U45286 ( .A1(n77301), .A2(n53628), .B(n56589), .C(
        n53628), .Y(n51971) );
  A2O1A1Ixp33_ASAP7_75t_SL U45287 ( .A1(n77301), .A2(n53628), .B(n56588), .C(
        n53628), .Y(n51970) );
  A2O1A1Ixp33_ASAP7_75t_SL U45288 ( .A1(n77301), .A2(n53628), .B(n56587), .C(
        n53628), .Y(n51960) );
  A2O1A1Ixp33_ASAP7_75t_SL U45289 ( .A1(n77301), .A2(n53628), .B(n56586), .C(
        n53628), .Y(n51969) );
  A2O1A1Ixp33_ASAP7_75t_SL U45290 ( .A1(n77301), .A2(n53628), .B(n56585), .C(
        n53628), .Y(n51968) );
  A2O1A1Ixp33_ASAP7_75t_SL U45291 ( .A1(n77301), .A2(n53628), .B(n56584), .C(
        n53628), .Y(n51967) );
  A2O1A1Ixp33_ASAP7_75t_SL U45292 ( .A1(n77301), .A2(n53628), .B(n56583), .C(
        n53628), .Y(n51966) );
  A2O1A1Ixp33_ASAP7_75t_SL U45293 ( .A1(n69721), .A2(n69722), .B(n69729), .C(
        n53628), .Y(n56580) );
  A2O1A1Ixp33_ASAP7_75t_SL U45294 ( .A1(n57081), .A2(n53628), .B(n69724), .C(
        n53628), .Y(n56581) );
  A2O1A1Ixp33_ASAP7_75t_SL U45295 ( .A1(n70504), .A2(n53628), .B(n70422), .C(
        n53628), .Y(n56582) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45296 ( .A1(n56580), .A2(n59621), .B(n56581), 
        .C(n53628), .D(n56582), .Y(n2311) );
  A2O1A1Ixp33_ASAP7_75t_SL U45297 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[6]), .A2(n70502), .B(
        n70510), .C(n53628), .Y(n56575) );
  A2O1A1Ixp33_ASAP7_75t_SL U45298 ( .A1(n77901), .A2(n77212), .B(n56569), .C(
        n53628), .Y(n56570) );
  A2O1A1Ixp33_ASAP7_75t_SL U45299 ( .A1(n1936), .A2(n53628), .B(n77214), .C(
        n56570), .Y(or1200_cpu_to_sr[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL U45300 ( .A1(n53628), .A2(n77246), .B(n57404), .C(
        n56298), .Y(n9328) );
  A2O1A1Ixp33_ASAP7_75t_SL U45301 ( .A1(n53628), .A2(n59680), .B(n1721), .C(
        n56083), .Y(or1200_du_N95) );
  A2O1A1Ixp33_ASAP7_75t_SL U45302 ( .A1(n77614), .A2(n53628), .B(n77645), .C(
        n53628), .Y(n56563) );
  A2O1A1Ixp33_ASAP7_75t_SL U45303 ( .A1(n56563), .A2(n53628), .B(n56566), .C(
        n53628), .Y(n1706) );
  A2O1A1Ixp33_ASAP7_75t_SL U45304 ( .A1(n77301), .A2(n53628), .B(n56562), .C(
        n53628), .Y(n51965) );
  A2O1A1Ixp33_ASAP7_75t_SL U45305 ( .A1(n77301), .A2(n53628), .B(n56561), .C(
        n53628), .Y(n51964) );
  A2O1A1Ixp33_ASAP7_75t_SL U45306 ( .A1(n77301), .A2(n53628), .B(n56560), .C(
        n53628), .Y(n51963) );
  A2O1A1Ixp33_ASAP7_75t_SL U45307 ( .A1(n77301), .A2(n53628), .B(n56559), .C(
        n53628), .Y(n51962) );
  A2O1A1Ixp33_ASAP7_75t_SL U45308 ( .A1(n59629), .A2(n53628), .B(n72700), .C(
        n56558), .Y(n1638) );
  A2O1A1Ixp33_ASAP7_75t_SL U45309 ( .A1(n77301), .A2(n53628), .B(n56557), .C(
        n53628), .Y(n51961) );
  A2O1A1Ixp33_ASAP7_75t_SL U45310 ( .A1(n57190), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_), .B(n56082), .C(
        n53628), .Y(n78374) );
  A2O1A1Ixp33_ASAP7_75t_SL U45311 ( .A1(n57114), .A2(n53628), .B(n1484), .C(
        n56556), .Y(n9306) );
  A2O1A1Ixp33_ASAP7_75t_SL U45312 ( .A1(n57114), .A2(n53628), .B(n1426), .C(
        n56555), .Y(n9277) );
  A2O1A1Ixp33_ASAP7_75t_SL U45313 ( .A1(n74641), .A2(n53628), .B(n1420), .C(
        n56554), .Y(n9325) );
  A2O1A1Ixp33_ASAP7_75t_SL U45314 ( .A1(n56542), .A2(n53628), .B(n76227), .C(
        n53628), .Y(n56543) );
  A2O1A1Ixp33_ASAP7_75t_SL U45315 ( .A1(n56536), .A2(n53628), .B(n63255), .C(
        n53628), .Y(n56537) );
  A2O1A1Ixp33_ASAP7_75t_SL U45316 ( .A1(n74641), .A2(n53628), .B(n1358), .C(
        n56531), .Y(n9309) );
  A2O1A1Ixp33_ASAP7_75t_SL U45317 ( .A1(n1290), .A2(n53628), .B(n4317), .C(
        n53628), .Y(n56520) );
  A2O1A1Ixp33_ASAP7_75t_SL U45318 ( .A1(n57083), .A2(n53628), .B(n1287), .C(
        n56521), .Y(n1288) );
  A2O1A1Ixp33_ASAP7_75t_SL U45319 ( .A1(n59703), .A2(n53628), .B(n56518), .C(
        n53628), .Y(or1200_immu_top_N33) );
  A2O1A1Ixp33_ASAP7_75t_SL U45320 ( .A1(n59703), .A2(n53628), .B(n56517), .C(
        n53628), .Y(n51953) );
  A2O1A1Ixp33_ASAP7_75t_SL U45321 ( .A1(n59703), .A2(n53628), .B(n56516), .C(
        n53628), .Y(n51951) );
  A2O1A1Ixp33_ASAP7_75t_SL U45322 ( .A1(n59703), .A2(n53628), .B(n56515), .C(
        n53628), .Y(n51947) );
  A2O1A1Ixp33_ASAP7_75t_SL U45323 ( .A1(n78264), .A2(n4132), .B(n59703), .C(
        n53628), .Y(n51946) );
  A2O1A1Ixp33_ASAP7_75t_SL U45324 ( .A1(n58863), .A2(n53628), .B(n76633), .C(
        n53628), .Y(n56500) );
  A2O1A1Ixp33_ASAP7_75t_SL U45325 ( .A1(or1200_cpu_or1200_mult_mac_n78), .A2(
        n53628), .B(n57077), .C(n53628), .Y(n56501) );
  A2O1A1Ixp33_ASAP7_75t_SL U45326 ( .A1(n56500), .A2(n53628), .B(n56501), .C(
        n53628), .Y(n56502) );
  A2O1A1Ixp33_ASAP7_75t_SL U45327 ( .A1(n58931), .A2(n53628), .B(n76633), .C(
        n53628), .Y(n56497) );
  A2O1A1Ixp33_ASAP7_75t_SL U45328 ( .A1(or1200_cpu_or1200_mult_mac_n110), .A2(
        n53628), .B(n57077), .C(n53628), .Y(n56498) );
  A2O1A1Ixp33_ASAP7_75t_SL U45329 ( .A1(n56497), .A2(n53628), .B(n56498), .C(
        n53628), .Y(n56499) );
  A2O1A1Ixp33_ASAP7_75t_SL U45330 ( .A1(or1200_cpu_or1200_mult_mac_n185), .A2(
        n53628), .B(n76889), .C(n53628), .Y(n56487) );
  A2O1A1Ixp33_ASAP7_75t_SL U45331 ( .A1(n77875), .A2(n76888), .B(n56487), .C(
        n53628), .Y(n56488) );
  A2O1A1Ixp33_ASAP7_75t_SL U45332 ( .A1(n65129), .A2(n53628), .B(n65100), .C(
        n65131), .Y(n56489) );
  A2O1A1Ixp33_ASAP7_75t_SL U45333 ( .A1(n59671), .A2(n53628), .B(n56489), .C(
        n56491), .Y(n56492) );
  A2O1A1Ixp33_ASAP7_75t_SL U45334 ( .A1(n59672), .A2(n56489), .B(n56491), .C(
        n53628), .Y(n56493) );
  A2O1A1Ixp33_ASAP7_75t_SL U45335 ( .A1(n76906), .A2(n53628), .B(n65126), .C(
        n56493), .Y(n56494) );
  A2O1A1Ixp33_ASAP7_75t_SL U45336 ( .A1(n53628), .A2(n55815), .B(n55818), .C(
        n55829), .Y(n55830) );
  A2O1A1Ixp33_ASAP7_75t_SL U45337 ( .A1(n75652), .A2(n53628), .B(n75135), .C(
        n57080), .Y(n55808) );
  A2O1A1Ixp33_ASAP7_75t_SL U45338 ( .A1(or1200_cpu_or1200_except_n290), .A2(
        n53628), .B(n77439), .C(n56486), .Y(or1200_cpu_or1200_except_n1786) );
  A2O1A1Ixp33_ASAP7_75t_SL U45339 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n380), .C(n56463), .Y(
        or1200_cpu_or1200_except_n381) );
  A2O1A1Ixp33_ASAP7_75t_SL U45340 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_spr_dat_ppc[20]), .C(n56241), .Y(
        or1200_cpu_or1200_except_n453) );
  A2O1A1Ixp33_ASAP7_75t_SL U45341 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_spr_dat_ppc[24]), .C(n56459), .Y(
        or1200_cpu_or1200_except_n465) );
  A2O1A1Ixp33_ASAP7_75t_SL U45342 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_spr_dat_ppc[26]), .C(n56027), .Y(
        or1200_cpu_or1200_except_n471) );
  A2O1A1Ixp33_ASAP7_75t_SL U45343 ( .A1(n76671), .A2(n53628), .B(n57331), .C(
        n56458), .Y(or1200_cpu_or1200_except_n682) );
  A2O1A1Ixp33_ASAP7_75t_SL U45344 ( .A1(n74245), .A2(n53628), .B(n74492), .C(
        n53628), .Y(n56455) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45345 ( .A1(n74246), .A2(n74493), .B(n74276), 
        .C(n53628), .D(n56455), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n50) );
  A2O1A1Ixp33_ASAP7_75t_SL U45346 ( .A1(n28210), .A2(n53628), .B(n70690), .C(
        n53628), .Y(n56434) );
  A2O1A1Ixp33_ASAP7_75t_SL U45347 ( .A1(n53628), .A2(n75925), .B(
        or1200_cpu_or1200_mult_mac_n54), .C(n55997), .Y(n76003) );
  A2O1A1Ixp33_ASAP7_75t_SL U45348 ( .A1(n71537), .A2(n53628), .B(n56428), .C(
        n53628), .Y(n71539) );
  A2O1A1Ixp33_ASAP7_75t_SL U45349 ( .A1(n70122), .A2(n53628), .B(n70121), .C(
        n53628), .Y(n56425) );
  A2O1A1Ixp33_ASAP7_75t_SL U45350 ( .A1(n70103), .A2(n53628), .B(n56422), .C(
        n53628), .Y(n70525) );
  A2O1A1Ixp33_ASAP7_75t_SL U45351 ( .A1(n74667), .A2(n53628), .B(n56419), .C(
        n53628), .Y(n74693) );
  A2O1A1Ixp33_ASAP7_75t_SL U45352 ( .A1(n77147), .A2(n53628), .B(n55988), .C(
        n55989), .Y(n78144) );
  A2O1A1Ixp33_ASAP7_75t_SL U45353 ( .A1(n57168), .A2(n53628), .B(n901), .C(
        n53628), .Y(n56418) );
  A2O1A1Ixp33_ASAP7_75t_SL U45354 ( .A1(n56418), .A2(n53628), .B(n63925), .C(
        n53628), .Y(n78256) );
  A2O1A1Ixp33_ASAP7_75t_SL U45355 ( .A1(n57160), .A2(n53628), .B(n56417), .C(
        n53628), .Y(n64259) );
  A2O1A1Ixp33_ASAP7_75t_SL U45356 ( .A1(n57160), .A2(n53628), .B(n56416), .C(
        n53628), .Y(n75161) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45357 ( .A1(n57321), .A2(n57456), .B(n53628), 
        .C(n59638), .Y(n56414) );
  A2O1A1Ixp33_ASAP7_75t_SL U45358 ( .A1(n69102), .A2(n53628), .B(n56413), .C(
        n53628), .Y(n69099) );
  A2O1A1Ixp33_ASAP7_75t_SL U45359 ( .A1(n75006), .A2(n53628), .B(n75009), .C(
        n53628), .Y(n56410) );
  A2O1A1Ixp33_ASAP7_75t_SL U45360 ( .A1(n75000), .A2(n53628), .B(n68820), .C(
        n56410), .Y(n68823) );
  A2O1A1Ixp33_ASAP7_75t_SL U45361 ( .A1(n68878), .A2(n53628), .B(n56409), .C(
        n53628), .Y(n68861) );
  A2O1A1Ixp33_ASAP7_75t_SL U45362 ( .A1(n69088), .A2(n53628), .B(n56407), .C(
        n53628), .Y(n69072) );
  A2O1A1Ixp33_ASAP7_75t_SL U45363 ( .A1(n69200), .A2(n53628), .B(n56406), .C(
        n53628), .Y(n69198) );
  A2O1A1Ixp33_ASAP7_75t_SL U45364 ( .A1(n59442), .A2(n53628), .B(n77744), .C(
        n53628), .Y(n56403) );
  A2O1A1Ixp33_ASAP7_75t_SL U45365 ( .A1(n59543), .A2(n53628), .B(n77745), .C(
        n53628), .Y(n56404) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45366 ( .A1(n77746), .A2(n77732), .B(n56403), 
        .C(n53628), .D(n56404), .Y(n4254) );
  A2O1A1Ixp33_ASAP7_75t_SL U45367 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_), 
        .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_), 
        .C(n53628), .Y(n56400) );
  A2O1A1Ixp33_ASAP7_75t_SL U45368 ( .A1(n70750), .A2(n53628), .B(n56399), .C(
        n53628), .Y(n70746) );
  A2O1A1Ixp33_ASAP7_75t_SL U45369 ( .A1(n71005), .A2(n53628), .B(n71006), .C(
        n53628), .Y(n56398) );
  A2O1A1Ixp33_ASAP7_75t_SL U45370 ( .A1(n53628), .A2(n65855), .B(n65646), .C(
        n53683), .Y(n66128) );
  A2O1A1Ixp33_ASAP7_75t_SL U45371 ( .A1(n65974), .A2(n53628), .B(n65969), .C(
        n53628), .Y(n56394) );
  A2O1A1Ixp33_ASAP7_75t_SL U45372 ( .A1(n65970), .A2(n53628), .B(n65966), .C(
        n53628), .Y(n56395) );
  A2O1A1Ixp33_ASAP7_75t_SL U45373 ( .A1(n65967), .A2(n66024), .B(n56395), .C(
        n53628), .Y(n56396) );
  A2O1A1Ixp33_ASAP7_75t_SL U45374 ( .A1(n66027), .A2(n53628), .B(n65971), .C(
        n56396), .Y(n56397) );
  A2O1A1Ixp33_ASAP7_75t_SL U45375 ( .A1(n56394), .A2(n53628), .B(n56397), .C(
        n53628), .Y(n65989) );
  O2A1O1Ixp33_ASAP7_75t_SL U45376 ( .A1(n75947), .A2(n58803), .B(n53628), .C(
        n59595), .Y(n56391) );
  A2O1A1Ixp33_ASAP7_75t_SL U45377 ( .A1(n58094), .A2(n53628), .B(n56388), .C(
        n53628), .Y(n68585) );
  A2O1A1Ixp33_ASAP7_75t_SL U45378 ( .A1(n53628), .A2(n59630), .B(n73180), .C(
        n56163), .Y(n73272) );
  A2O1A1Ixp33_ASAP7_75t_SL U45379 ( .A1(n53628), .A2(n59630), .B(n73141), .C(
        n55958), .Y(n73280) );
  A2O1A1Ixp33_ASAP7_75t_SL U45380 ( .A1(n3331), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .C(
        n53628), .Y(n56386) );
  A2O1A1Ixp33_ASAP7_75t_SL U45381 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[2]), .B(n56386), .C(
        n53628), .Y(n73725) );
  A2O1A1Ixp33_ASAP7_75t_SL U45382 ( .A1(n75738), .A2(n53628), .B(
        or1200_cpu_or1200_mult_mac_n347), .C(n53628), .Y(n56384) );
  A2O1A1Ixp33_ASAP7_75t_SL U45383 ( .A1(n75736), .A2(n76429), .B(n56384), .C(
        n53628), .Y(n56385) );
  A2O1A1Ixp33_ASAP7_75t_SL U45384 ( .A1(n72944), .A2(n53628), .B(n56382), .C(
        n53628), .Y(n72967) );
  A2O1A1Ixp33_ASAP7_75t_SL U45385 ( .A1(n75278), .A2(n53628), .B(n75277), .C(
        n53628), .Y(n56378) );
  A2O1A1Ixp33_ASAP7_75t_SL U45386 ( .A1(n75283), .A2(n53628), .B(n56379), .C(
        n53628), .Y(n56380) );
  A2O1A1Ixp33_ASAP7_75t_SL U45387 ( .A1(n71413), .A2(n53628), .B(n56377), .C(
        n53628), .Y(n71251) );
  A2O1A1Ixp33_ASAP7_75t_SL U45388 ( .A1(n57187), .A2(n65823), .B(n56373), .C(
        n53628), .Y(n56374) );
  A2O1A1Ixp33_ASAP7_75t_SL U45389 ( .A1(or1200_cpu_or1200_mult_mac_n98), .A2(
        n53628), .B(n56369), .C(n53628), .Y(n56370) );
  A2O1A1Ixp33_ASAP7_75t_SL U45390 ( .A1(n57121), .A2(n63501), .B(n56370), .C(
        n53628), .Y(n77115) );
  A2O1A1Ixp33_ASAP7_75t_SL U45391 ( .A1(n70103), .A2(n53628), .B(n56368), .C(
        n53628), .Y(n69627) );
  A2O1A1Ixp33_ASAP7_75t_SL U45392 ( .A1(n68602), .A2(n53628), .B(n59670), .C(
        n53628), .Y(n56366) );
  A2O1A1Ixp33_ASAP7_75t_SL U45393 ( .A1(n68603), .A2(n59670), .B(n56366), .C(
        n53628), .Y(n56367) );
  A2O1A1Ixp33_ASAP7_75t_SL U45394 ( .A1(n75076), .A2(n53628), .B(n68604), .C(
        n56367), .Y(n68612) );
  A2O1A1Ixp33_ASAP7_75t_SL U45395 ( .A1(n66988), .A2(n56363), .B(n69138), .C(
        n53628), .Y(n56364) );
  A2O1A1Ixp33_ASAP7_75t_SL U45396 ( .A1(n56364), .A2(n53628), .B(n69137), .C(
        n53628), .Y(n67104) );
  INVx1_ASAP7_75t_SL U45397 ( .A(n59648), .Y(n53226) );
  INVx1_ASAP7_75t_SL U45398 ( .A(n67964), .Y(n53240) );
  A2O1A1Ixp33_ASAP7_75t_SL U45399 ( .A1(n72678), .A2(n53628), .B(n56138), .C(
        n56139), .Y(n27978) );
  A2O1A1Ixp33_ASAP7_75t_SL U45400 ( .A1(n71527), .A2(n53628), .B(n71528), .C(
        n53628), .Y(n56357) );
  A2O1A1Ixp33_ASAP7_75t_SL U45401 ( .A1(n78054), .A2(n59701), .B(n56350), .C(
        n53628), .Y(n56351) );
  A2O1A1Ixp33_ASAP7_75t_SL U45402 ( .A1(n78163), .A2(n53628), .B(n77491), .C(
        n53628), .Y(n56346) );
  A2O1A1Ixp33_ASAP7_75t_SL U45403 ( .A1(n77469), .A2(n56346), .B(n77486), .C(
        n53628), .Y(n56347) );
  A2O1A1Ixp33_ASAP7_75t_SL U45404 ( .A1(n77764), .A2(n53628), .B(n77470), .C(
        n53628), .Y(n56348) );
  A2O1A1Ixp33_ASAP7_75t_SL U45405 ( .A1(n78157), .A2(n53628), .B(n56348), .C(
        n53628), .Y(n56349) );
  A2O1A1Ixp33_ASAP7_75t_SL U45406 ( .A1(n56347), .A2(n53628), .B(n3111), .C(
        n56349), .Y(n9391) );
  A2O1A1Ixp33_ASAP7_75t_SL U45407 ( .A1(n3078), .A2(n53628), .B(n77454), .C(
        n56345), .Y(n9677) );
  A2O1A1Ixp33_ASAP7_75t_SL U45408 ( .A1(n53628), .A2(n59688), .B(n3071), .C(
        n55910), .Y(n3072) );
  A2O1A1Ixp33_ASAP7_75t_SL U45409 ( .A1(n59688), .A2(n53628), .B(n3057), .C(
        n56343), .Y(n3058) );
  A2O1A1Ixp33_ASAP7_75t_SL U45410 ( .A1(n64162), .A2(n53628), .B(n64163), .C(
        n53628), .Y(n56333) );
  A2O1A1Ixp33_ASAP7_75t_SL U45411 ( .A1(n57144), .A2(n53628), .B(n56333), .C(
        n53628), .Y(n56334) );
  A2O1A1Ixp33_ASAP7_75t_SL U45412 ( .A1(n57144), .A2(n53628), .B(n56331), .C(
        n56332), .Y(n2998) );
  A2O1A1Ixp33_ASAP7_75t_SL U45413 ( .A1(n76948), .A2(n74899), .B(n74844), .C(
        n53628), .Y(n56330) );
  A2O1A1Ixp33_ASAP7_75t_SL U45414 ( .A1(n74741), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[29]), .C(n53628), 
        .Y(n56327) );
  A2O1A1Ixp33_ASAP7_75t_SL U45415 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_1_), 
        .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[29]), .C(
        n53628), .Y(n56328) );
  A2O1A1Ixp33_ASAP7_75t_SL U45416 ( .A1(n56327), .A2(n53628), .B(n56328), .C(
        n53628), .Y(n56329) );
  A2O1A1Ixp33_ASAP7_75t_SL U45417 ( .A1(n77301), .A2(n53628), .B(n56326), .C(
        n53628), .Y(n2852) );
  A2O1A1Ixp33_ASAP7_75t_SL U45418 ( .A1(n53628), .A2(n57074), .B(wb_insn[28]), 
        .C(n55678), .Y(n2808) );
  A2O1A1Ixp33_ASAP7_75t_SL U45419 ( .A1(n53628), .A2(n59689), .B(n2804), .C(
        n56117), .Y(n2805) );
  A2O1A1Ixp33_ASAP7_75t_SL U45420 ( .A1(n57190), .A2(n53628), .B(n72884), .C(
        n56325), .Y(n2799) );
  A2O1A1Ixp33_ASAP7_75t_SL U45421 ( .A1(n53628), .A2(n77246), .B(n2785), .C(
        n56116), .Y(n9337) );
  A2O1A1Ixp33_ASAP7_75t_SL U45422 ( .A1(n53447), .A2(n53628), .B(n77346), .C(
        n53628), .Y(n56322) );
  A2O1A1Ixp33_ASAP7_75t_SL U45423 ( .A1(n77345), .A2(n56322), .B(n59156), .C(
        n53628), .Y(n56323) );
  A2O1A1Ixp33_ASAP7_75t_SL U45424 ( .A1(n2614), .A2(n53628), .B(n77567), .C(
        n56321), .Y(n9203) );
  A2O1A1Ixp33_ASAP7_75t_SL U45425 ( .A1(n2532), .A2(n53628), .B(n59688), .C(
        n56320), .Y(n2533) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45426 ( .A1(n65387), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_8_), .B(n65317), .C(
        n53628), .D(n65354), .Y(n56319) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45427 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_8_), .A2(n65357), .B(
        n56319), .C(n53628), .D(n65331), .Y(n2488) );
  A2O1A1Ixp33_ASAP7_75t_SL U45428 ( .A1(n53628), .A2(n2461), .B(n59688), .C(
        n56114), .Y(n2462) );
  A2O1A1Ixp33_ASAP7_75t_SL U45429 ( .A1(n74681), .A2(n53628), .B(n70553), .C(
        n53628), .Y(n56304) );
  A2O1A1Ixp33_ASAP7_75t_SL U45430 ( .A1(n70551), .A2(n53628), .B(n2448), .C(
        n53628), .Y(n56305) );
  A2O1A1Ixp33_ASAP7_75t_SL U45431 ( .A1(n56304), .A2(n53628), .B(n56305), .C(
        n53628), .Y(n56306) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45432 ( .A1(n70538), .A2(n70539), .B(n56308), 
        .C(n53628), .D(n70537), .Y(n56309) );
  A2O1A1Ixp33_ASAP7_75t_SL U45433 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_2_), .A2(
        n53628), .B(n70540), .C(n53628), .Y(n56313) );
  A2O1A1Ixp33_ASAP7_75t_SL U45434 ( .A1(n74674), .A2(n53628), .B(n59633), .C(
        n53628), .Y(n56314) );
  A2O1A1Ixp33_ASAP7_75t_SL U45435 ( .A1(n56313), .A2(n53628), .B(n56314), .C(
        n53628), .Y(n56315) );
  A2O1A1Ixp33_ASAP7_75t_SL U45436 ( .A1(n77301), .A2(n53628), .B(n56303), .C(
        n53628), .Y(n51974) );
  A2O1A1Ixp33_ASAP7_75t_SL U45437 ( .A1(n70530), .A2(n53628), .B(n27525), .C(
        n53628), .Y(n56302) );
  A2O1A1Ixp33_ASAP7_75t_SL U45438 ( .A1(n56302), .A2(n53628), .B(n70503), .C(
        n53628), .Y(n2210) );
  A2O1A1Ixp33_ASAP7_75t_SL U45439 ( .A1(n53628), .A2(n57144), .B(n77902), .C(
        n55445), .Y(n2197) );
  A2O1A1Ixp33_ASAP7_75t_SL U45440 ( .A1(n53628), .A2(n2119), .B(n57073), .C(
        n56092), .Y(n2120) );
  A2O1A1Ixp33_ASAP7_75t_SL U45441 ( .A1(n53628), .A2(n59689), .B(n2023), .C(
        n55439), .Y(n2024) );
  A2O1A1Ixp33_ASAP7_75t_SL U45442 ( .A1(n53628), .A2(n59680), .B(n1976), .C(
        n56090), .Y(or1200_du_N98) );
  A2O1A1Ixp33_ASAP7_75t_SL U45443 ( .A1(n53628), .A2(n77246), .B(n1938), .C(
        n56089), .Y(n9329) );
  A2O1A1Ixp33_ASAP7_75t_SL U45444 ( .A1(n59703), .A2(n53628), .B(n56301), .C(
        n53628), .Y(n9467) );
  A2O1A1Ixp33_ASAP7_75t_SL U45445 ( .A1(n53628), .A2(n77246), .B(n1832), .C(
        n56088), .Y(n9336) );
  A2O1A1Ixp33_ASAP7_75t_SL U45446 ( .A1(n53628), .A2(n59680), .B(n1826), .C(
        n56087), .Y(or1200_du_N103) );
  A2O1A1Ixp33_ASAP7_75t_SL U45447 ( .A1(n53628), .A2(n77246), .B(n1815), .C(
        n56086), .Y(n9332) );
  A2O1A1Ixp33_ASAP7_75t_SL U45448 ( .A1(n59629), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_11_), .C(n56299), .Y(
        n1780) );
  A2O1A1Ixp33_ASAP7_75t_SL U45449 ( .A1(n57083), .A2(n53628), .B(dwb_sel_o[0]), 
        .C(n56297), .Y(n1749) );
  A2O1A1Ixp33_ASAP7_75t_SL U45450 ( .A1(n77590), .A2(n53628), .B(n77645), .C(
        n53628), .Y(n56292) );
  A2O1A1Ixp33_ASAP7_75t_SL U45451 ( .A1(n56292), .A2(n53628), .B(n56295), .C(
        n53628), .Y(n1713) );
  A2O1A1Ixp33_ASAP7_75t_SL U45452 ( .A1(n57190), .A2(n53628), .B(n56291), .C(
        n53628), .Y(n1543) );
  A2O1A1Ixp33_ASAP7_75t_SL U45453 ( .A1(n57114), .A2(n53628), .B(n1474), .C(
        n56289), .Y(n9301) );
  A2O1A1Ixp33_ASAP7_75t_SL U45454 ( .A1(n53628), .A2(n74641), .B(n1400), .C(
        n55018), .Y(n9320) );
  A2O1A1Ixp33_ASAP7_75t_SL U45455 ( .A1(n59703), .A2(n53628), .B(n56283), .C(
        n53628), .Y(or1200_immu_top_N20) );
  A2O1A1Ixp33_ASAP7_75t_SL U45456 ( .A1(n59703), .A2(n53628), .B(n56282), .C(
        n53628), .Y(n51949) );
  A2O1A1Ixp33_ASAP7_75t_SL U45457 ( .A1(n64699), .A2(n53628), .B(n64095), .C(
        n53628), .Y(n56279) );
  A2O1A1Ixp33_ASAP7_75t_SL U45458 ( .A1(n63370), .A2(n53628), .B(n63369), .C(
        n53628), .Y(n56277) );
  A2O1A1Ixp33_ASAP7_75t_SL U45459 ( .A1(or1200_cpu_or1200_mult_mac_n18), .A2(
        n53628), .B(n56274), .C(n53628), .Y(n56275) );
  A2O1A1Ixp33_ASAP7_75t_SL U45460 ( .A1(n76195), .A2(n56273), .B(n56275), .C(
        n53628), .Y(n56276) );
  A2O1A1Ixp33_ASAP7_75t_SL U45461 ( .A1(or1200_cpu_or1200_mult_mac_n20), .A2(
        n53628), .B(n76158), .C(n56276), .Y(or1200_cpu_or1200_mult_mac_n1504)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45462 ( .A1(n53628), .A2(
        or1200_cpu_or1200_mult_mac_n82), .B(n57105), .C(n55840), .Y(
        or1200_cpu_or1200_mult_mac_n1537) );
  A2O1A1Ixp33_ASAP7_75t_SL U45463 ( .A1(or1200_cpu_or1200_mult_mac_n92), .A2(
        n53628), .B(n57077), .C(n53628), .Y(n56269) );
  A2O1A1Ixp33_ASAP7_75t_SL U45464 ( .A1(n53241), .A2(n56268), .B(n56269), .C(
        n53628), .Y(n56270) );
  A2O1A1Ixp33_ASAP7_75t_SL U45465 ( .A1(or1200_cpu_or1200_mult_mac_n90), .A2(
        n53628), .B(n57105), .C(n56270), .Y(or1200_cpu_or1200_mult_mac_n1541)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45466 ( .A1(n53628), .A2(n57105), .B(
        or1200_cpu_or1200_mult_mac_n112), .C(n56060), .Y(
        or1200_cpu_or1200_mult_mac_n1552) );
  A2O1A1Ixp33_ASAP7_75t_SL U45467 ( .A1(n63516), .A2(n53628), .B(n56255), .C(
        n53628), .Y(n56256) );
  A2O1A1Ixp33_ASAP7_75t_SL U45468 ( .A1(n76906), .A2(n53628), .B(n63532), .C(
        n53628), .Y(n56257) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45469 ( .A1(n59672), .A2(n56256), .B(n56257), 
        .C(n53628), .D(n56258), .Y(n56259) );
  A2O1A1Ixp33_ASAP7_75t_SL U45470 ( .A1(n56256), .A2(n53628), .B(n59671), .C(
        n53628), .Y(n56260) );
  A2O1A1Ixp33_ASAP7_75t_SL U45471 ( .A1(n56260), .A2(n53628), .B(n56262), .C(
        n53628), .Y(n56263) );
  A2O1A1Ixp33_ASAP7_75t_SL U45472 ( .A1(n56259), .A2(n53628), .B(n56263), .C(
        n53628), .Y(n56264) );
  A2O1A1Ixp33_ASAP7_75t_SL U45473 ( .A1(or1200_cpu_or1200_mult_mac_n173), .A2(
        n53628), .B(n76889), .C(n53628), .Y(n56265) );
  A2O1A1Ixp33_ASAP7_75t_SL U45474 ( .A1(n56264), .A2(n53628), .B(n56265), .C(
        n53628), .Y(n56266) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45475 ( .A1(n75290), .A2(n54430), .B(n53628), 
        .C(n59671), .Y(n54431) );
  A2O1A1Ixp33_ASAP7_75t_SL U45476 ( .A1(n53628), .A2(n75294), .B(n75293), .C(
        n54432), .Y(n54433) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45477 ( .A1(n75294), .A2(n54434), .B(n53628), 
        .C(n75293), .Y(n54435) );
  A2O1A1Ixp33_ASAP7_75t_SL U45478 ( .A1(n53628), .A2(n54430), .B(n75290), .C(
        n57079), .Y(n54436) );
  A2O1A1Ixp33_ASAP7_75t_SL U45479 ( .A1(n53628), .A2(n54431), .B(n54433), .C(
        n54437), .Y(n54438) );
  A2O1A1Ixp33_ASAP7_75t_SL U45480 ( .A1(n75117), .A2(n53628), .B(n76906), .C(
        n53628), .Y(n56245) );
  A2O1A1Ixp33_ASAP7_75t_SL U45481 ( .A1(n75118), .A2(n53628), .B(n59671), .C(
        n53628), .Y(n56249) );
  A2O1A1Ixp33_ASAP7_75t_SL U45482 ( .A1(n56249), .A2(n53628), .B(n56250), .C(
        n53628), .Y(n56251) );
  A2O1A1Ixp33_ASAP7_75t_SL U45483 ( .A1(n56245), .A2(n53628), .B(n56248), .C(
        n56253), .Y(n56254) );
  A2O1A1Ixp33_ASAP7_75t_SL U45484 ( .A1(n53628), .A2(n77209), .B(
        or1200_cpu_or1200_except_n122), .C(n56036), .Y(
        or1200_cpu_or1200_except_n1735) );
  A2O1A1Ixp33_ASAP7_75t_SL U45485 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n401), .C(n56035), .Y(
        or1200_cpu_or1200_except_n402) );
  A2O1A1Ixp33_ASAP7_75t_SL U45486 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n404), .C(n56034), .Y(
        or1200_cpu_or1200_except_n405) );
  A2O1A1Ixp33_ASAP7_75t_SL U45487 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n407), .C(n56033), .Y(
        or1200_cpu_or1200_except_n408) );
  A2O1A1Ixp33_ASAP7_75t_SL U45488 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n416), .C(n55166), .Y(
        or1200_cpu_or1200_except_n417) );
  A2O1A1Ixp33_ASAP7_75t_SL U45489 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n419), .C(n56032), .Y(
        or1200_cpu_or1200_except_n420) );
  A2O1A1Ixp33_ASAP7_75t_SL U45490 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n422), .C(n55373), .Y(
        or1200_cpu_or1200_except_n423) );
  A2O1A1Ixp33_ASAP7_75t_SL U45491 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n425), .C(n55372), .Y(
        or1200_cpu_or1200_except_n426) );
  A2O1A1Ixp33_ASAP7_75t_SL U45492 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n431), .C(n56031), .Y(
        or1200_cpu_or1200_except_n432) );
  A2O1A1Ixp33_ASAP7_75t_SL U45493 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n434), .C(n56242), .Y(
        or1200_cpu_or1200_except_n435) );
  A2O1A1Ixp33_ASAP7_75t_SL U45494 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n446), .C(n56030), .Y(
        or1200_cpu_or1200_except_n447) );
  A2O1A1Ixp33_ASAP7_75t_SL U45495 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_spr_dat_ppc[19]), .C(n56029), .Y(
        or1200_cpu_or1200_except_n450) );
  A2O1A1Ixp33_ASAP7_75t_SL U45496 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_spr_dat_ppc[21]), .C(n55802), .Y(
        or1200_cpu_or1200_except_n456) );
  A2O1A1Ixp33_ASAP7_75t_SL U45497 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_spr_dat_ppc[22]), .C(n56240), .Y(
        or1200_cpu_or1200_except_n459) );
  A2O1A1Ixp33_ASAP7_75t_SL U45498 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n461), .C(n56028), .Y(
        or1200_cpu_or1200_except_n462) );
  A2O1A1Ixp33_ASAP7_75t_SL U45499 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n467), .C(n56239), .Y(
        or1200_cpu_or1200_except_n468) );
  A2O1A1Ixp33_ASAP7_75t_SL U45500 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_spr_dat_ppc[27]), .C(n55602), .Y(
        or1200_cpu_or1200_except_n474) );
  A2O1A1Ixp33_ASAP7_75t_SL U45501 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_spr_dat_ppc[29]), .C(n56238), .Y(
        or1200_cpu_or1200_except_n480) );
  A2O1A1Ixp33_ASAP7_75t_SL U45502 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n482), .C(n56026), .Y(
        or1200_cpu_or1200_except_n483) );
  A2O1A1Ixp33_ASAP7_75t_SL U45503 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_spr_dat_ppc[31]), .C(n56025), .Y(
        or1200_cpu_or1200_except_n486) );
  A2O1A1Ixp33_ASAP7_75t_SL U45504 ( .A1(n74492), .A2(n53628), .B(n56236), .C(
        n53628), .Y(n56237) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45505 ( .A1(n74493), .A2(n56234), .B(n74276), 
        .C(n53628), .D(n56237), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n54) );
  A2O1A1Ixp33_ASAP7_75t_SL U45506 ( .A1(n70690), .A2(n71353), .B(n59699), .C(
        n53628), .Y(n56230) );
  A2O1A1Ixp33_ASAP7_75t_SL U45507 ( .A1(n56230), .A2(n53628), .B(n56231), .C(
        n53628), .Y(n56232) );
  A2O1A1Ixp33_ASAP7_75t_SL U45508 ( .A1(n56229), .A2(n53628), .B(n56232), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n106) );
  A2O1A1Ixp33_ASAP7_75t_SL U45509 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .A2(
        n53628), .B(n73765), .C(n56226), .Y(n73796) );
  A2O1A1Ixp33_ASAP7_75t_SL U45510 ( .A1(or1200_cpu_or1200_except_n619), .A2(
        n53628), .B(n2630), .C(n53628), .Y(n56225) );
  A2O1A1Ixp33_ASAP7_75t_SL U45511 ( .A1(n56225), .A2(n53628), .B(n63994), .C(
        n53628), .Y(n63975) );
  A2O1A1Ixp33_ASAP7_75t_SL U45512 ( .A1(n70003), .A2(n53628), .B(n56223), .C(
        n53628), .Y(n69987) );
  A2O1A1Ixp33_ASAP7_75t_SL U45513 ( .A1(n53628), .A2(n77148), .B(n55987), .C(
        n53628), .Y(n55988) );
  A2O1A1Ixp33_ASAP7_75t_SL U45514 ( .A1(n57168), .A2(n53628), .B(n919), .C(
        n53628), .Y(n56213) );
  A2O1A1Ixp33_ASAP7_75t_SL U45515 ( .A1(n56213), .A2(n53628), .B(n63920), .C(
        n53628), .Y(n78188) );
  A2O1A1Ixp33_ASAP7_75t_SL U45516 ( .A1(n57160), .A2(n53628), .B(n56212), .C(
        n53628), .Y(n75174) );
  A2O1A1Ixp33_ASAP7_75t_SL U45517 ( .A1(or1200_cpu_or1200_mult_mac_n331), .A2(
        n53628), .B(n56202), .C(n53628), .Y(n65144) );
  A2O1A1Ixp33_ASAP7_75t_SL U45518 ( .A1(n69132), .A2(n53628), .B(n56200), .C(
        n53628), .Y(n69162) );
  A2O1A1Ixp33_ASAP7_75t_SL U45519 ( .A1(or1200_cpu_or1200_mult_mac_n247), .A2(
        n53628), .B(n69258), .C(n53628), .Y(n56198) );
  A2O1A1Ixp33_ASAP7_75t_SL U45520 ( .A1(n69256), .A2(n56197), .B(n56198), .C(
        n53628), .Y(n56199) );
  A2O1A1Ixp33_ASAP7_75t_SL U45521 ( .A1(n59539), .A2(n53628), .B(n77745), .C(
        n53628), .Y(n56193) );
  A2O1A1Ixp33_ASAP7_75t_SL U45522 ( .A1(n59549), .A2(n53628), .B(n77741), .C(
        n53628), .Y(n56194) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45523 ( .A1(n78004), .A2(n77742), .B(n56193), 
        .C(n53628), .D(n56194), .Y(n4246) );
  A2O1A1Ixp33_ASAP7_75t_SL U45524 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_0_), .A2(
        n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_1_), .C(
        n53628), .Y(n56192) );
  A2O1A1Ixp33_ASAP7_75t_SL U45525 ( .A1(n57203), .A2(n53628), .B(n72306), .C(
        n53628), .Y(n56187) );
  A2O1A1Ixp33_ASAP7_75t_SL U45526 ( .A1(n57127), .A2(n53628), .B(n72308), .C(
        n53628), .Y(n56188) );
  A2O1A1Ixp33_ASAP7_75t_SL U45527 ( .A1(n72309), .A2(n53628), .B(n57123), .C(
        n53628), .Y(n56189) );
  A2O1A1Ixp33_ASAP7_75t_SL U45528 ( .A1(n56188), .A2(n53628), .B(n56189), .C(
        n53628), .Y(n56190) );
  A2O1A1Ixp33_ASAP7_75t_SL U45529 ( .A1(n57125), .A2(n53628), .B(n72307), .C(
        n56190), .Y(n56191) );
  A2O1A1Ixp33_ASAP7_75t_SL U45530 ( .A1(n56187), .A2(n53628), .B(n56191), .C(
        n53628), .Y(n72472) );
  A2O1A1Ixp33_ASAP7_75t_SL U45531 ( .A1(n57123), .A2(n53628), .B(n71950), .C(
        n53628), .Y(n56186) );
  A2O1A1Ixp33_ASAP7_75t_SL U45532 ( .A1(n56186), .A2(n53628), .B(n71951), .C(
        n53628), .Y(n72440) );
  A2O1A1Ixp33_ASAP7_75t_SL U45533 ( .A1(n57208), .A2(n53628), .B(n72212), .C(
        n53628), .Y(n56180) );
  A2O1A1Ixp33_ASAP7_75t_SL U45534 ( .A1(n56180), .A2(n53628), .B(n56183), .C(
        n53628), .Y(n56184) );
  A2O1A1Ixp33_ASAP7_75t_SL U45535 ( .A1(n71890), .A2(n53628), .B(n72154), .C(
        n53628), .Y(n56176) );
  A2O1A1Ixp33_ASAP7_75t_SL U45536 ( .A1(n58422), .A2(n53628), .B(n72080), .C(
        n53628), .Y(n56177) );
  A2O1A1Ixp33_ASAP7_75t_SL U45537 ( .A1(n57207), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_33_), 
        .B(n56177), .C(n53628), .Y(n56178) );
  A2O1A1Ixp33_ASAP7_75t_SL U45538 ( .A1(n57208), .A2(n53628), .B(n72132), .C(
        n56178), .Y(n56179) );
  A2O1A1Ixp33_ASAP7_75t_SL U45539 ( .A1(n56176), .A2(n53628), .B(n56179), .C(
        n53628), .Y(n72050) );
  A2O1A1Ixp33_ASAP7_75t_SL U45540 ( .A1(n70799), .A2(n56175), .B(n70800), .C(
        n53628), .Y(n70785) );
  A2O1A1Ixp33_ASAP7_75t_SL U45541 ( .A1(n78402), .A2(n53628), .B(n56172), .C(
        n53628), .Y(n71050) );
  A2O1A1Ixp33_ASAP7_75t_SL U45542 ( .A1(n66181), .A2(n53628), .B(n65630), .C(
        n53628), .Y(n56167) );
  A2O1A1Ixp33_ASAP7_75t_SL U45543 ( .A1(n65646), .A2(n53628), .B(n65635), .C(
        n53628), .Y(n56168) );
  A2O1A1Ixp33_ASAP7_75t_SL U45544 ( .A1(n56167), .A2(n53628), .B(n56168), .C(
        n53628), .Y(n56169) );
  A2O1A1Ixp33_ASAP7_75t_SL U45545 ( .A1(n65970), .A2(n53628), .B(n66075), .C(
        n53628), .Y(n56165) );
  A2O1A1Ixp33_ASAP7_75t_SL U45546 ( .A1(n65965), .A2(n53628), .B(n65974), .C(
        n53628), .Y(n56166) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45547 ( .A1(n65978), .A2(n65964), .B(n56165), 
        .C(n53628), .D(n56166), .Y(n65990) );
  A2O1A1Ixp33_ASAP7_75t_SL U45548 ( .A1(n71746), .A2(n53628), .B(n56164), .C(
        n53628), .Y(n71727) );
  A2O1A1Ixp33_ASAP7_75t_SL U45549 ( .A1(n53628), .A2(n59630), .B(n73129), .C(
        n54052), .Y(n73292) );
  A2O1A1Ixp33_ASAP7_75t_SL U45550 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[2]), .A2(
        n56162), .B(n70133), .C(n53628), .Y(n70132) );
  A2O1A1Ixp33_ASAP7_75t_SL U45551 ( .A1(n77418), .A2(n56160), .B(n77416), .C(
        n53628), .Y(n77417) );
  A2O1A1Ixp33_ASAP7_75t_SL U45552 ( .A1(n61560), .A2(n53628), .B(n61559), .C(
        n61399), .Y(n56159) );
  A2O1A1Ixp33_ASAP7_75t_SL U45553 ( .A1(n69138), .A2(n53628), .B(n53500), .C(
        n53628), .Y(n56153) );
  O2A1O1Ixp33_ASAP7_75t_SL U45554 ( .A1(n69137), .A2(n69142), .B(n53628), .C(
        n56153), .Y(n56154) );
  A2O1A1Ixp33_ASAP7_75t_SL U45555 ( .A1(n56154), .A2(n53628), .B(n56155), .C(
        n53628), .Y(n56156) );
  A2O1A1Ixp33_ASAP7_75t_SL U45556 ( .A1(n63892), .A2(n53628), .B(n63891), .C(
        n56152), .Y(n65081) );
  A2O1A1Ixp33_ASAP7_75t_SL U45557 ( .A1(or1200_cpu_or1200_mult_mac_n261), .A2(
        n53628), .B(n56151), .C(n53628), .Y(n75653) );
  A2O1A1Ixp33_ASAP7_75t_SL U45558 ( .A1(n59631), .A2(n53628), .B(n73265), .C(
        n56150), .Y(n73268) );
  A2O1A1Ixp33_ASAP7_75t_SL U45559 ( .A1(n76383), .A2(n53628), .B(n56149), .C(
        n53628), .Y(n76460) );
  A2O1A1Ixp33_ASAP7_75t_SL U45560 ( .A1(n57120), .A2(n64917), .B(n55269), .C(
        n53628), .Y(n61971) );
  A2O1A1Ixp33_ASAP7_75t_SL U45561 ( .A1(n67179), .A2(n53628), .B(n67190), .C(
        n67187), .Y(n55932) );
  A2O1A1Ixp33_ASAP7_75t_SL U45562 ( .A1(n53628), .A2(n67193), .B(n55932), .C(
        n55935), .Y(n67208) );
  A2O1A1Ixp33_ASAP7_75t_SL U45563 ( .A1(n59548), .A2(n53628), .B(n57183), .C(
        n57120), .Y(n56144) );
  A2O1A1Ixp33_ASAP7_75t_SL U45564 ( .A1(n59440), .A2(n53628), .B(n56143), .C(
        n53628), .Y(n66368) );
  A2O1A1Ixp33_ASAP7_75t_SL U45565 ( .A1(n66962), .A2(n53628), .B(n56141), .C(
        n53628), .Y(n56142) );
  A2O1A1Ixp33_ASAP7_75t_SL U45566 ( .A1(n66963), .A2(n59102), .B(n56142), .C(
        n53628), .Y(n68450) );
  OAI21xp5_ASAP7_75t_SL U45567 ( .A1(n68455), .A2(n56140), .B(n53628), .Y(
        n66722) );
  A2O1A1Ixp33_ASAP7_75t_SL U45568 ( .A1(n73833), .A2(n53628), .B(n59704), .C(
        n53628), .Y(n56135) );
  A2O1A1Ixp33_ASAP7_75t_SL U45569 ( .A1(n73652), .A2(n53628), .B(n56134), .C(
        n53628), .Y(n3281) );
  A2O1A1Ixp33_ASAP7_75t_SL U45570 ( .A1(n78382), .A2(n53628), .B(n71539), .C(
        n53628), .Y(n56131) );
  O2A1O1Ixp33_ASAP7_75t_SL U45571 ( .A1(n55924), .A2(n55925), .B(n53628), .C(
        n69798), .Y(n55926) );
  A2O1A1Ixp33_ASAP7_75t_SL U45572 ( .A1(n70030), .A2(n53628), .B(n69878), .C(
        n55926), .Y(n3216) );
  A2O1A1Ixp33_ASAP7_75t_SL U45573 ( .A1(n74934), .A2(n53628), .B(n59554), .C(
        n53628), .Y(n56123) );
  A2O1A1Ixp33_ASAP7_75t_SL U45574 ( .A1(n3141), .A2(n53628), .B(n74916), .C(
        n53628), .Y(n56124) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45575 ( .A1(n74921), .A2(
        or1200_cpu_or1200_fpu_ine_conv), .B(n56123), .C(n53628), .D(n56124), 
        .Y(n56125) );
  A2O1A1Ixp33_ASAP7_75t_SL U45576 ( .A1(n57144), .A2(n53628), .B(n77462), .C(
        n56122), .Y(n3066) );
  A2O1A1Ixp33_ASAP7_75t_SL U45577 ( .A1(n59688), .A2(n53628), .B(n3024), .C(
        n56121), .Y(n3025) );
  A2O1A1Ixp33_ASAP7_75t_SL U45578 ( .A1(n74846), .A2(n74899), .B(n74885), .C(
        n53628), .Y(n56120) );
  A2O1A1Ixp33_ASAP7_75t_SL U45579 ( .A1(n53628), .A2(n57202), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[28]), .C(n55900), 
        .Y(n2864) );
  A2O1A1Ixp33_ASAP7_75t_SL U45580 ( .A1(n53628), .A2(n57074), .B(n2816), .C(
        n55897), .Y(n2817) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45581 ( .A1(n57084), .A2(n55238), .B(n53628), 
        .C(n2773), .Y(n55239) );
  A2O1A1Ixp33_ASAP7_75t_SL U45582 ( .A1(n53628), .A2(n2544), .B(n57074), .C(
        n54511), .Y(n2545) );
  A2O1A1Ixp33_ASAP7_75t_SL U45583 ( .A1(n2542), .A2(n53628), .B(n77567), .C(
        n56115), .Y(n9204) );
  A2O1A1Ixp33_ASAP7_75t_SL U45584 ( .A1(n2865), .A2(n53628), .B(n65322), .C(
        n65308), .Y(n55675) );
  A2O1A1Ixp33_ASAP7_75t_SL U45585 ( .A1(n70534), .A2(n70541), .B(n70469), .C(
        n53628), .Y(n56099) );
  A2O1A1Ixp33_ASAP7_75t_SL U45586 ( .A1(n70471), .A2(n53628), .B(n70536), .C(
        n53628), .Y(n56103) );
  A2O1A1Ixp33_ASAP7_75t_SL U45587 ( .A1(n70387), .A2(n53628), .B(n70466), .C(
        n53628), .Y(n56104) );
  O2A1O1Ixp33_ASAP7_75t_SL U45588 ( .A1(n56103), .A2(n56104), .B(n53628), .C(
        n56106), .Y(n56107) );
  A2O1A1Ixp33_ASAP7_75t_SL U45589 ( .A1(n56099), .A2(n53628), .B(n56102), .C(
        n56107), .Y(n2429) );
  A2O1A1Ixp33_ASAP7_75t_SL U45590 ( .A1(n53628), .A2(n55883), .B(n55885), .C(
        n59621), .Y(n55886) );
  A2O1A1Ixp33_ASAP7_75t_SL U45591 ( .A1(n53628), .A2(n70506), .B(n70422), .C(
        n53628), .Y(n55888) );
  A2O1A1Ixp33_ASAP7_75t_SL U45592 ( .A1(n53628), .A2(n55887), .B(n55888), .C(
        n53628), .Y(n2309) );
  A2O1A1Ixp33_ASAP7_75t_SL U45593 ( .A1(n53628), .A2(n57074), .B(n2076), .C(
        n55878), .Y(n2077) );
  A2O1A1Ixp33_ASAP7_75t_SL U45594 ( .A1(n53628), .A2(n1951), .B(n77214), .C(
        n54471), .Y(or1200_cpu_to_sr[6]) );
  A2O1A1Ixp33_ASAP7_75t_SL U45595 ( .A1(n57083), .A2(n53628), .B(dwb_sel_o[1]), 
        .C(n56085), .Y(n1746) );
  A2O1A1Ixp33_ASAP7_75t_SL U45596 ( .A1(n77672), .A2(n77864), .B(n55871), .C(
        n53628), .Y(n1700) );
  A2O1A1Ixp33_ASAP7_75t_SL U45597 ( .A1(n59626), .A2(n53628), .B(n78376), .C(
        n53628), .Y(n56082) );
  A2O1A1Ixp33_ASAP7_75t_SL U45598 ( .A1(n75616), .A2(n53628), .B(n1510), .C(
        n56081), .Y(n9327) );
  A2O1A1Ixp33_ASAP7_75t_SL U45599 ( .A1(n57114), .A2(n53628), .B(n1482), .C(
        n56080), .Y(n9305) );
  A2O1A1Ixp33_ASAP7_75t_SL U45600 ( .A1(n53628), .A2(n74641), .B(n1388), .C(
        n55652), .Y(n9317) );
  A2O1A1Ixp33_ASAP7_75t_SL U45601 ( .A1(n53628), .A2(n74641), .B(n1384), .C(
        n54816), .Y(n9316) );
  A2O1A1Ixp33_ASAP7_75t_SL U45602 ( .A1(n59703), .A2(n53628), .B(n56073), .C(
        n53628), .Y(or1200_immu_top_N27) );
  A2O1A1Ixp33_ASAP7_75t_SL U45603 ( .A1(n59703), .A2(n53628), .B(n56072), .C(
        n53628), .Y(or1200_immu_top_N21) );
  A2O1A1Ixp33_ASAP7_75t_SL U45604 ( .A1(n4106), .A2(n53628), .B(n56069), .C(
        n53628), .Y(n56070) );
  A2O1A1Ixp33_ASAP7_75t_SL U45605 ( .A1(n65232), .A2(n59701), .B(n56070), .C(
        n53628), .Y(n56071) );
  A2O1A1Ixp33_ASAP7_75t_SL U45606 ( .A1(n771), .A2(n53628), .B(n76523), .C(
        n56071), .Y(n9170) );
  A2O1A1Ixp33_ASAP7_75t_SL U45607 ( .A1(n63296), .A2(n53628), .B(n63299), .C(
        n53628), .Y(n56062) );
  A2O1A1Ixp33_ASAP7_75t_SL U45608 ( .A1(n76633), .A2(n53628), .B(n57108), .C(
        n53628), .Y(n56058) );
  A2O1A1Ixp33_ASAP7_75t_SL U45609 ( .A1(n57077), .A2(n53628), .B(
        or1200_cpu_or1200_mult_mac_n114), .C(n53628), .Y(n56059) );
  A2O1A1Ixp33_ASAP7_75t_SL U45610 ( .A1(n56058), .A2(n53628), .B(n56059), .C(
        n53628), .Y(n56060) );
  A2O1A1Ixp33_ASAP7_75t_SL U45611 ( .A1(or1200_cpu_or1200_mult_mac_n143), .A2(
        n53628), .B(n76889), .C(n55399), .Y(or1200_cpu_or1200_mult_mac_n1592)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45612 ( .A1(or1200_cpu_or1200_mult_mac_n183), .A2(
        n53628), .B(n76889), .C(n53628), .Y(n56048) );
  A2O1A1Ixp33_ASAP7_75t_SL U45613 ( .A1(n77877), .A2(n76888), .B(n56048), .C(
        n53628), .Y(n56049) );
  A2O1A1Ixp33_ASAP7_75t_SL U45614 ( .A1(n65074), .A2(n56050), .B(n65094), .C(
        n53628), .Y(n56051) );
  A2O1A1Ixp33_ASAP7_75t_SL U45615 ( .A1(n65129), .A2(n53628), .B(n56052), .C(
        n53628), .Y(n56053) );
  A2O1A1Ixp33_ASAP7_75t_SL U45616 ( .A1(n65100), .A2(n53628), .B(n59671), .C(
        n56053), .Y(n56054) );
  A2O1A1Ixp33_ASAP7_75t_SL U45617 ( .A1(n65100), .A2(n59672), .B(n56053), .C(
        n53628), .Y(n56055) );
  A2O1A1Ixp33_ASAP7_75t_SL U45618 ( .A1(n76906), .A2(n53628), .B(n56051), .C(
        n56055), .Y(n56056) );
  A2O1A1Ixp33_ASAP7_75t_SL U45619 ( .A1(n55820), .A2(n53628), .B(
        or1200_cpu_or1200_mult_mac_n381), .C(n53628), .Y(n55821) );
  A2O1A1Ixp33_ASAP7_75t_SL U45620 ( .A1(n76906), .A2(n53628), .B(n56037), .C(
        n53628), .Y(n56038) );
  A2O1A1Ixp33_ASAP7_75t_SL U45621 ( .A1(n75659), .A2(n53628), .B(n75663), .C(
        n56039), .Y(n56040) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45622 ( .A1(n75141), .A2(n75661), .B(n59671), 
        .C(n53628), .D(n75660), .Y(n56041) );
  O2A1O1Ixp5_ASAP7_75t_SL U45623 ( .A1(n56041), .A2(n75659), .B(n53628), .C(
        n75663), .Y(n56042) );
  A2O1A1Ixp33_ASAP7_75t_SL U45624 ( .A1(n56038), .A2(n53628), .B(n56040), .C(
        n56044), .Y(n56045) );
  A2O1A1Ixp33_ASAP7_75t_SL U45625 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n428), .C(n54625), .Y(
        or1200_cpu_or1200_except_n429) );
  A2O1A1Ixp33_ASAP7_75t_SL U45626 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n440), .C(n55803), .Y(
        or1200_cpu_or1200_except_n441) );
  A2O1A1Ixp33_ASAP7_75t_SL U45627 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_spr_dat_ppc[17]), .C(n55603), .Y(
        or1200_cpu_or1200_except_n444) );
  A2O1A1Ixp33_ASAP7_75t_SL U45628 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n652), .C(n55369), .Y(
        or1200_cpu_or1200_except_n1814) );
  O2A1O1Ixp33_ASAP7_75t_SL U45629 ( .A1(n55790), .A2(n55792), .B(n53628), .C(
        n55793), .Y(n55794) );
  A2O1A1Ixp33_ASAP7_75t_SL U45630 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_23_), 
        .A2(n74493), .B(n55796), .C(n53628), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n45) );
  A2O1A1Ixp33_ASAP7_75t_SL U45631 ( .A1(n72499), .A2(n53628), .B(n72290), .C(
        n53628), .Y(n56008) );
  A2O1A1Ixp33_ASAP7_75t_SL U45632 ( .A1(n57192), .A2(n53628), .B(n72285), .C(
        n53628), .Y(n56009) );
  A2O1A1Ixp33_ASAP7_75t_SL U45633 ( .A1(n56008), .A2(n53628), .B(n56009), .C(
        n53628), .Y(n56010) );
  A2O1A1Ixp33_ASAP7_75t_SL U45634 ( .A1(n57125), .A2(n53628), .B(n72250), .C(
        n53628), .Y(n56012) );
  A2O1A1Ixp33_ASAP7_75t_SL U45635 ( .A1(n72348), .A2(n53628), .B(n57123), .C(
        n53628), .Y(n56013) );
  A2O1A1Ixp33_ASAP7_75t_SL U45636 ( .A1(n56012), .A2(n53628), .B(n56013), .C(
        n53628), .Y(n56014) );
  A2O1A1Ixp33_ASAP7_75t_SL U45637 ( .A1(n72502), .A2(n56016), .B(n56020), .C(
        n53628), .Y(n56021) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45638 ( .A1(n53628), .A2(n56011), .B(n72368), 
        .C(n53628), .D(n56023), .Y(n56024) );
  A2O1A1Ixp33_ASAP7_75t_SL U45639 ( .A1(n71494), .A2(n53628), .B(n56006), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_N2435)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45640 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_3_), .C(n55572), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n112) );
  A2O1A1Ixp33_ASAP7_75t_SL U45641 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_13_), .C(n55340), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n142) );
  A2O1A1Ixp33_ASAP7_75t_SL U45642 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_16_), .C(n56005), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n151) );
  A2O1A1Ixp33_ASAP7_75t_SL U45643 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_28_), .C(n56002), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n187) );
  O2A1O1Ixp5_ASAP7_75t_SL U45644 ( .A1(n58206), .A2(n59465), .B(n53628), .C(
        n55998), .Y(n58460) );
  A2O1A1Ixp33_ASAP7_75t_SL U45645 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .A2(
        n53628), .B(n55995), .C(n53628), .Y(n73686) );
  A2O1A1Ixp33_ASAP7_75t_SL U45646 ( .A1(n74141), .A2(n53628), .B(n55991), .C(
        n53628), .Y(n74181) );
  A2O1A1Ixp33_ASAP7_75t_SL U45647 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_6_), 
        .A2(n53628), .B(or1200_cpu_or1200_fpu_fpu_op_r_5_), .C(n53628), .Y(
        n55990) );
  A2O1A1Ixp33_ASAP7_75t_SL U45648 ( .A1(n77150), .A2(n53628), .B(n77149), .C(
        n53628), .Y(n55987) );
  A2O1A1Ixp33_ASAP7_75t_SL U45649 ( .A1(n57168), .A2(n53628), .B(n839), .C(
        n53628), .Y(n55985) );
  A2O1A1Ixp33_ASAP7_75t_SL U45650 ( .A1(n57160), .A2(n53628), .B(n76570), .C(
        n53628), .Y(n55986) );
  O2A1O1Ixp5_ASAP7_75t_SL U45651 ( .A1(n76568), .A2(n55985), .B(n53628), .C(
        n55986), .Y(n4093) );
  A2O1A1Ixp33_ASAP7_75t_SL U45652 ( .A1(n57168), .A2(n53628), .B(n883), .C(
        n53628), .Y(n55984) );
  A2O1A1Ixp33_ASAP7_75t_SL U45653 ( .A1(n55984), .A2(n53628), .B(n63987), .C(
        n53628), .Y(n78254) );
  A2O1A1Ixp33_ASAP7_75t_SL U45654 ( .A1(n53628), .A2(n57130), .B(n55529), .C(
        n53628), .Y(n59295) );
  A2O1A1Ixp33_ASAP7_75t_SL U45655 ( .A1(n68834), .A2(n53628), .B(n58442), .C(
        n53628), .Y(n55982) );
  A2O1A1Ixp33_ASAP7_75t_SL U45656 ( .A1(n68721), .A2(n53628), .B(n58442), .C(
        n58867), .Y(n55983) );
  A2O1A1Ixp33_ASAP7_75t_SL U45657 ( .A1(n53625), .A2(n55982), .B(n55983), .C(
        n53628), .Y(n68855) );
  A2O1A1Ixp33_ASAP7_75t_SL U45658 ( .A1(n68818), .A2(n53628), .B(n55979), .C(
        n53628), .Y(n68799) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45659 ( .A1(n68987), .A2(n68993), .B(n53628), 
        .C(n55976), .Y(n68950) );
  A2O1A1Ixp33_ASAP7_75t_SL U45660 ( .A1(n77443), .A2(n53628), .B(n77435), .C(
        n53628), .Y(n55973) );
  A2O1A1Ixp33_ASAP7_75t_SL U45661 ( .A1(n55973), .A2(n53628), .B(n77434), .C(
        n53628), .Y(n55974) );
  A2O1A1Ixp33_ASAP7_75t_SL U45662 ( .A1(n77437), .A2(n53628), .B(n55974), .C(
        n53628), .Y(n77439) );
  A2O1A1Ixp33_ASAP7_75t_SL U45663 ( .A1(n74235), .A2(n53628), .B(n55972), .C(
        n53628), .Y(n74236) );
  A2O1A1Ixp33_ASAP7_75t_SL U45664 ( .A1(n57208), .A2(n53628), .B(n71993), .C(
        n53628), .Y(n55966) );
  A2O1A1Ixp33_ASAP7_75t_SL U45665 ( .A1(n55966), .A2(n53628), .B(n55969), .C(
        n53628), .Y(n55970) );
  A2O1A1Ixp33_ASAP7_75t_SL U45666 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_31_), .A2(n53628), 
        .B(n55965), .C(n53628), .Y(n71292) );
  A2O1A1Ixp33_ASAP7_75t_SL U45667 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[33]), .A2(n66182), 
        .B(n55515), .C(n53628), .Y(n55516) );
  A2O1A1Ixp33_ASAP7_75t_SL U45668 ( .A1(n65966), .A2(n53628), .B(n65974), .C(
        n53628), .Y(n55962) );
  A2O1A1Ixp33_ASAP7_75t_SL U45669 ( .A1(n65978), .A2(n65967), .B(n55962), .C(
        n53628), .Y(n55963) );
  A2O1A1Ixp33_ASAP7_75t_SL U45670 ( .A1(n65965), .A2(n53628), .B(n65970), .C(
        n55963), .Y(n55964) );
  A2O1A1Ixp33_ASAP7_75t_SL U45671 ( .A1(n65964), .A2(n66024), .B(n55964), .C(
        n53628), .Y(n66043) );
  A2O1A1Ixp33_ASAP7_75t_SL U45672 ( .A1(n65026), .A2(n65027), .B(n65025), .C(
        n53628), .Y(n55960) );
  A2O1A1Ixp33_ASAP7_75t_SL U45673 ( .A1(n55960), .A2(n53628), .B(n55961), .C(
        n53628), .Y(n68262) );
  OAI21xp5_ASAP7_75t_SL U45674 ( .A1(n65029), .A2(n65028), .B(n53628), .Y(
        n55961) );
  A2O1A1Ixp33_ASAP7_75t_SL U45675 ( .A1(n67536), .A2(n53628), .B(n67535), .C(
        n55959), .Y(n67691) );
  A2O1A1Ixp33_ASAP7_75t_SL U45676 ( .A1(n53628), .A2(n59630), .B(n73119), .C(
        n55735), .Y(n73325) );
  A2O1A1Ixp33_ASAP7_75t_SL U45677 ( .A1(n53628), .A2(n70103), .B(n69776), .C(
        n55733), .Y(n69786) );
  A2O1A1Ixp33_ASAP7_75t_SL U45678 ( .A1(n59538), .A2(n53628), .B(n55954), .C(
        n53628), .Y(n61518) );
  A2O1A1Ixp33_ASAP7_75t_SL U45679 ( .A1(n76461), .A2(n53628), .B(n77066), .C(
        n53628), .Y(n55952) );
  A2O1A1Ixp33_ASAP7_75t_SL U45680 ( .A1(or1200_cpu_or1200_mult_mac_n159), .A2(
        n53628), .B(n77057), .C(n53628), .Y(n55953) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45681 ( .A1(n76753), .A2(n63409), .B(n55952), 
        .C(n53628), .D(n55953), .Y(n61354) );
  A2O1A1Ixp33_ASAP7_75t_SL U45682 ( .A1(n75189), .A2(n53628), .B(n75791), .C(
        n53628), .Y(n55950) );
  A2O1A1Ixp33_ASAP7_75t_SL U45683 ( .A1(n75190), .A2(n53628), .B(n55950), .C(
        n53628), .Y(n77175) );
  A2O1A1Ixp33_ASAP7_75t_SL U45684 ( .A1(or1200_cpu_or1200_mult_mac_n239), .A2(
        n53628), .B(n55949), .C(n53628), .Y(n69203) );
  A2O1A1Ixp33_ASAP7_75t_SL U45685 ( .A1(n57203), .A2(n53628), .B(n72079), .C(
        n53628), .Y(n55944) );
  A2O1A1Ixp33_ASAP7_75t_SL U45686 ( .A1(n57127), .A2(n53628), .B(n72141), .C(
        n53628), .Y(n55945) );
  A2O1A1Ixp33_ASAP7_75t_SL U45687 ( .A1(n72080), .A2(n53628), .B(n57123), .C(
        n53628), .Y(n55946) );
  A2O1A1Ixp33_ASAP7_75t_SL U45688 ( .A1(n55945), .A2(n53628), .B(n55946), .C(
        n53628), .Y(n55947) );
  A2O1A1Ixp33_ASAP7_75t_SL U45689 ( .A1(n57125), .A2(n53628), .B(n72132), .C(
        n55947), .Y(n55948) );
  A2O1A1Ixp33_ASAP7_75t_SL U45690 ( .A1(n55944), .A2(n53628), .B(n55948), .C(
        n53628), .Y(n72270) );
  A2O1A1Ixp33_ASAP7_75t_SL U45691 ( .A1(n59526), .A2(n53628), .B(n71377), .C(
        n55280), .Y(n71359) );
  A2O1A1Ixp33_ASAP7_75t_SL U45692 ( .A1(n59631), .A2(n53628), .B(n73264), .C(
        n53628), .Y(n55943) );
  A2O1A1Ixp33_ASAP7_75t_SL U45693 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[2]), .A2(
        n53628), .B(n55941), .C(n53628), .Y(n70133) );
  A2O1A1Ixp33_ASAP7_75t_SL U45694 ( .A1(n73968), .A2(n53628), .B(n55939), .C(
        n53628), .Y(n76434) );
  A2O1A1Ixp33_ASAP7_75t_SL U45695 ( .A1(n67191), .A2(n53628), .B(n55933), .C(
        n53628), .Y(n55934) );
  A2O1A1Ixp33_ASAP7_75t_SL U45696 ( .A1(n59604), .A2(n53628), .B(n59620), .C(
        n55931), .Y(n64380) );
  OAI21xp5_ASAP7_75t_SL U45697 ( .A1(n66829), .A2(n55930), .B(n53628), .Y(
        n58476) );
  A2O1A1Ixp33_ASAP7_75t_SL U45698 ( .A1(n66794), .A2(n66726), .B(n53264), .C(
        n53628), .Y(n66969) );
  A2O1A1Ixp33_ASAP7_75t_SL U45699 ( .A1(n73828), .A2(n53628), .B(n59704), .C(
        n53628), .Y(n55929) );
  A2O1A1Ixp33_ASAP7_75t_SL U45700 ( .A1(n69902), .A2(n53628), .B(n69926), .C(
        n53628), .Y(n55924) );
  A2O1A1Ixp33_ASAP7_75t_SL U45701 ( .A1(n69877), .A2(n53628), .B(n69932), .C(
        n53628), .Y(n55925) );
  A2O1A1Ixp33_ASAP7_75t_SL U45702 ( .A1(n70580), .A2(n53628), .B(n55918), .C(
        n53628), .Y(n55919) );
  A2O1A1Ixp33_ASAP7_75t_SL U45703 ( .A1(n70579), .A2(n53628), .B(n55919), .C(
        n55923), .Y(n51978) );
  A2O1A1Ixp33_ASAP7_75t_SL U45704 ( .A1(n59629), .A2(n53628), .B(n72786), .C(
        n55917), .Y(n3124) );
  A2O1A1Ixp33_ASAP7_75t_SL U45705 ( .A1(n74847), .A2(n77194), .B(n74872), .C(
        n53628), .Y(n55901) );
  A2O1A1Ixp33_ASAP7_75t_SL U45706 ( .A1(n74899), .A2(n55902), .B(n74885), .C(
        n53628), .Y(n55903) );
  A2O1A1Ixp33_ASAP7_75t_SL U45707 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_6_), .A2(n53628), 
        .B(n55901), .C(n55903), .Y(n52489) );
  A2O1A1Ixp33_ASAP7_75t_SL U45708 ( .A1(n74741), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[28]), .C(n53628), 
        .Y(n55898) );
  A2O1A1Ixp33_ASAP7_75t_SL U45709 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_1_), 
        .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[28]), .C(
        n53628), .Y(n55899) );
  A2O1A1Ixp33_ASAP7_75t_SL U45710 ( .A1(n55898), .A2(n53628), .B(n55899), .C(
        n53628), .Y(n55900) );
  A2O1A1Ixp33_ASAP7_75t_SL U45711 ( .A1(n53628), .A2(n77233), .B(n77295), .C(
        n54857), .Y(or1200_du_N107) );
  A2O1A1Ixp33_ASAP7_75t_SL U45712 ( .A1(n53628), .A2(n57144), .B(n77857), .C(
        n55234), .Y(n2559) );
  A2O1A1Ixp33_ASAP7_75t_SL U45713 ( .A1(n65322), .A2(n53628), .B(n55893), .C(
        n53628), .Y(n55894) );
  A2O1A1Ixp33_ASAP7_75t_SL U45714 ( .A1(n65354), .A2(n53628), .B(n65306), .C(
        n53628), .Y(n55895) );
  A2O1A1Ixp33_ASAP7_75t_SL U45715 ( .A1(n53628), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_4_), .B(n69381), .C(
        n55462), .Y(n2452) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45716 ( .A1(n70471), .A2(n70473), .B(n53628), 
        .C(n70472), .Y(n55451) );
  A2O1A1Ixp33_ASAP7_75t_SL U45717 ( .A1(n69726), .A2(n55879), .B(n55882), .C(
        n53628), .Y(n55883) );
  A2O1A1Ixp33_ASAP7_75t_SL U45718 ( .A1(n69727), .A2(n53628), .B(n55884), .C(
        n53628), .Y(n55885) );
  A2O1A1Ixp33_ASAP7_75t_SL U45719 ( .A1(n57081), .A2(n53628), .B(n69731), .C(
        n55886), .Y(n55887) );
  A2O1A1Ixp33_ASAP7_75t_SL U45720 ( .A1(n53628), .A2(n2157), .B(n57073), .C(
        n55666), .Y(n2158) );
  A2O1A1Ixp33_ASAP7_75t_SL U45721 ( .A1(n57074), .A2(n53628), .B(n2056), .C(
        n55877), .Y(n2057) );
  A2O1A1Ixp33_ASAP7_75t_SL U45722 ( .A1(n57144), .A2(n53628), .B(n76628), .C(
        n55875), .Y(n1959) );
  A2O1A1Ixp33_ASAP7_75t_SL U45723 ( .A1(n57190), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .B(n55438), .C(
        n53628), .Y(n1859) );
  A2O1A1Ixp33_ASAP7_75t_SL U45724 ( .A1(n59680), .A2(n53628), .B(n1757), .C(
        n55874), .Y(or1200_du_N97) );
  A2O1A1Ixp33_ASAP7_75t_SL U45725 ( .A1(dwb_sel_o[2]), .A2(n53628), .B(n57083), 
        .C(n55873), .Y(n1743) );
  A2O1A1Ixp33_ASAP7_75t_SL U45726 ( .A1(n77666), .A2(n53628), .B(n55870), .C(
        n53628), .Y(n55871) );
  A2O1A1Ixp33_ASAP7_75t_SL U45727 ( .A1(n59627), .A2(n53628), .B(n72700), .C(
        n55869), .Y(n1632) );
  A2O1A1Ixp33_ASAP7_75t_SL U45728 ( .A1(n53628), .A2(n1492), .B(n54828), .C(
        n54830), .Y(n9672) );
  A2O1A1Ixp33_ASAP7_75t_SL U45729 ( .A1(n57114), .A2(n53628), .B(n1480), .C(
        n55868), .Y(n9304) );
  A2O1A1Ixp33_ASAP7_75t_SL U45730 ( .A1(n53628), .A2(n74641), .B(n1412), .C(
        n54663), .Y(n9323) );
  A2O1A1Ixp33_ASAP7_75t_SL U45731 ( .A1(n53628), .A2(n74641), .B(n1408), .C(
        n55215), .Y(n9322) );
  A2O1A1Ixp33_ASAP7_75t_SL U45732 ( .A1(n74641), .A2(n53628), .B(n1396), .C(
        n55867), .Y(n9319) );
  A2O1A1Ixp33_ASAP7_75t_SL U45733 ( .A1(n57083), .A2(n53628), .B(n1349), .C(
        n55856), .Y(n1350) );
  A2O1A1Ixp33_ASAP7_75t_SL U45734 ( .A1(n75198), .A2(n53628), .B(n76890), .C(
        n55852), .Y(n9247) );
  A2O1A1Ixp33_ASAP7_75t_SL U45735 ( .A1(n55850), .A2(n53628), .B(n76545), .C(
        n53628), .Y(n55851) );
  A2O1A1Ixp33_ASAP7_75t_SL U45736 ( .A1(n63281), .A2(n53628), .B(n63280), .C(
        n63298), .Y(n55411) );
  A2O1A1Ixp33_ASAP7_75t_SL U45737 ( .A1(n53628), .A2(n63279), .B(n55410), .C(
        n55411), .Y(n55412) );
  A2O1A1Ixp33_ASAP7_75t_SL U45738 ( .A1(n76193), .A2(n53628), .B(n55843), .C(
        n53628), .Y(n55844) );
  A2O1A1Ixp33_ASAP7_75t_SL U45739 ( .A1(or1200_cpu_or1200_mult_mac_n2), .A2(
        n53628), .B(n57105), .C(n55845), .Y(or1200_cpu_or1200_mult_mac_n1496)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45740 ( .A1(n58021), .A2(n53628), .B(n76633), .C(
        n53628), .Y(n55838) );
  A2O1A1Ixp33_ASAP7_75t_SL U45741 ( .A1(or1200_cpu_or1200_mult_mac_n84), .A2(
        n53628), .B(n57077), .C(n53628), .Y(n55839) );
  A2O1A1Ixp33_ASAP7_75t_SL U45742 ( .A1(n55838), .A2(n53628), .B(n55839), .C(
        n53628), .Y(n55840) );
  A2O1A1Ixp33_ASAP7_75t_SL U45743 ( .A1(n76897), .A2(n53628), .B(n63770), .C(
        n63889), .Y(n55832) );
  A2O1A1Ixp33_ASAP7_75t_SL U45744 ( .A1(n63775), .A2(n55831), .B(n76906), .C(
        n53628), .Y(n55834) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45745 ( .A1(n63770), .A2(n57079), .B(n55834), 
        .C(n53628), .D(n63889), .Y(n55835) );
  A2O1A1Ixp33_ASAP7_75t_SL U45746 ( .A1(n55833), .A2(n53628), .B(n55835), .C(
        n53628), .Y(n55836) );
  A2O1A1Ixp33_ASAP7_75t_SL U45747 ( .A1(n76888), .A2(n77888), .B(n55836), .C(
        n53628), .Y(n55837) );
  A2O1A1Ixp33_ASAP7_75t_SL U45748 ( .A1(or1200_cpu_or1200_mult_mac_n175), .A2(
        n53628), .B(n76889), .C(n55837), .Y(or1200_cpu_or1200_mult_mac_n1576)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45749 ( .A1(n53628), .A2(n53959), .B(n59671), .C(
        n53960), .Y(n53961) );
  A2O1A1Ixp33_ASAP7_75t_SL U45750 ( .A1(n59672), .A2(n53959), .B(n53960), .C(
        n53628), .Y(n53962) );
  A2O1A1Ixp33_ASAP7_75t_SL U45751 ( .A1(n53628), .A2(n76906), .B(n53958), .C(
        n53962), .Y(n53963) );
  A2O1A1Ixp33_ASAP7_75t_SL U45752 ( .A1(n76906), .A2(n53628), .B(n69162), .C(
        n53628), .Y(n55815) );
  A2O1A1Ixp33_ASAP7_75t_SL U45753 ( .A1(n69213), .A2(n53628), .B(n59671), .C(
        n53628), .Y(n55820) );
  A2O1A1Ixp33_ASAP7_75t_SL U45754 ( .A1(n75141), .A2(n55805), .B(n76897), .C(
        n53628), .Y(n55806) );
  A2O1A1Ixp33_ASAP7_75t_SL U45755 ( .A1(n55807), .A2(n53628), .B(n55808), .C(
        n55809), .Y(n55810) );
  A2O1A1Ixp33_ASAP7_75t_SL U45756 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n413), .C(n55167), .Y(
        or1200_cpu_or1200_except_n414) );
  A2O1A1Ixp33_ASAP7_75t_SL U45757 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n619), .C(n55599), .Y(
        or1200_cpu_or1200_except_n1803) );
  A2O1A1Ixp33_ASAP7_75t_SL U45758 ( .A1(or1200_cpu_or1200_except_n631), .A2(
        n53628), .B(n57093), .C(n55801), .Y(or1200_cpu_or1200_except_n1807) );
  A2O1A1Ixp33_ASAP7_75t_SL U45759 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n643), .C(n53951), .Y(
        or1200_cpu_or1200_except_n1811) );
  A2O1A1Ixp33_ASAP7_75t_SL U45760 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n655), .C(n55163), .Y(
        or1200_cpu_or1200_except_n1815) );
  A2O1A1Ixp33_ASAP7_75t_SL U45761 ( .A1(n53628), .A2(n76671), .B(n2966), .C(
        n55597), .Y(or1200_cpu_or1200_except_n685) );
  A2O1A1Ixp33_ASAP7_75t_SL U45762 ( .A1(n74488), .A2(n53628), .B(n55789), .C(
        n53628), .Y(n55790) );
  A2O1A1Ixp33_ASAP7_75t_SL U45763 ( .A1(n74489), .A2(n53628), .B(n55791), .C(
        n53628), .Y(n55792) );
  A2O1A1Ixp33_ASAP7_75t_SL U45764 ( .A1(n74730), .A2(n53628), .B(n74728), .C(
        n53628), .Y(n55793) );
  A2O1A1Ixp33_ASAP7_75t_SL U45765 ( .A1(n72509), .A2(n53628), .B(n59624), .C(
        n53628), .Y(n55781) );
  A2O1A1Ixp33_ASAP7_75t_SL U45766 ( .A1(n72472), .A2(n53628), .B(n59623), .C(
        n53628), .Y(n55782) );
  A2O1A1Ixp33_ASAP7_75t_SL U45767 ( .A1(n72371), .A2(n53628), .B(n72434), .C(
        n53628), .Y(n55783) );
  O2A1O1Ixp5_ASAP7_75t_SL U45768 ( .A1(n55781), .A2(n55782), .B(n53628), .C(
        n55783), .Y(n55784) );
  A2O1A1Ixp33_ASAP7_75t_SL U45769 ( .A1(n59622), .A2(n53628), .B(n72506), .C(
        n55784), .Y(n55785) );
  A2O1A1Ixp33_ASAP7_75t_SL U45770 ( .A1(n72510), .A2(n55785), .B(n55786), .C(
        n53628), .Y(n55787) );
  A2O1A1Ixp33_ASAP7_75t_SL U45771 ( .A1(n53628), .A2(n70713), .B(n55568), .C(
        n55571), .Y(n55572) );
  A2O1A1Ixp33_ASAP7_75t_SL U45772 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_5_), .C(n54412), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n118) );
  A2O1A1Ixp33_ASAP7_75t_SL U45773 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_10_), .C(n55567), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n133) );
  A2O1A1Ixp33_ASAP7_75t_SL U45774 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_14_), .C(n55562), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n145) );
  A2O1A1Ixp33_ASAP7_75t_SL U45775 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_18_), .C(n54407), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n157) );
  A2O1A1Ixp33_ASAP7_75t_SL U45776 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_26_), .C(n55557), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n181) );
  A2O1A1Ixp33_ASAP7_75t_SL U45777 ( .A1(n67515), .A2(n53628), .B(n58884), .C(
        n67514), .Y(n55780) );
  A2O1A1Ixp33_ASAP7_75t_SL U45778 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[11]), .A2(n59632), .B(
        n55779), .C(n53628), .Y(n73771) );
  A2O1A1Ixp33_ASAP7_75t_SL U45779 ( .A1(n57217), .A2(n73767), .B(n55773), .C(
        n53628), .Y(n55774) );
  A2O1A1Ixp33_ASAP7_75t_SL U45780 ( .A1(n72600), .A2(n53628), .B(n55770), .C(
        n53628), .Y(n71526) );
  A2O1A1Ixp33_ASAP7_75t_SL U45781 ( .A1(n70201), .A2(n53628), .B(n55769), .C(
        n53628), .Y(n70204) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45782 ( .A1(n76861), .A2(n76860), .B(n53628), 
        .C(n76859), .Y(n55767) );
  A2O1A1Ixp33_ASAP7_75t_SL U45783 ( .A1(n76862), .A2(n53628), .B(n55767), .C(
        n53628), .Y(n55768) );
  A2O1A1Ixp33_ASAP7_75t_SL U45784 ( .A1(n75191), .A2(n53628), .B(n55764), .C(
        n53628), .Y(n55765) );
  A2O1A1Ixp33_ASAP7_75t_SL U45785 ( .A1(n57168), .A2(n53628), .B(n892), .C(
        n53628), .Y(n55763) );
  A2O1A1Ixp33_ASAP7_75t_SL U45786 ( .A1(n55763), .A2(n53628), .B(n63930), .C(
        n53628), .Y(n78255) );
  A2O1A1Ixp33_ASAP7_75t_SL U45787 ( .A1(n57160), .A2(n53628), .B(n55762), .C(
        n53628), .Y(n75171) );
  O2A1O1Ixp33_ASAP7_75t_SL U45788 ( .A1(n76151), .A2(n76148), .B(n53628), .C(
        n55760), .Y(n76150) );
  A2O1A1Ixp33_ASAP7_75t_SL U45789 ( .A1(n76040), .A2(n55758), .B(n76041), .C(
        n53628), .Y(n55759) );
  A2O1A1Ixp33_ASAP7_75t_SL U45790 ( .A1(n76042), .A2(n53628), .B(n55759), .C(
        n53628), .Y(n76054) );
  A2O1A1Ixp33_ASAP7_75t_SL U45791 ( .A1(n63399), .A2(n53628), .B(n63326), .C(
        n55757), .Y(n63335) );
  A2O1A1Ixp33_ASAP7_75t_SL U45792 ( .A1(n53453), .A2(n53628), .B(n55754), .C(
        n53628), .Y(n75019) );
  A2O1A1Ixp33_ASAP7_75t_SL U45793 ( .A1(or1200_cpu_or1200_mult_mac_n209), .A2(
        n53628), .B(n55753), .C(n53628), .Y(n68872) );
  A2O1A1Ixp33_ASAP7_75t_SL U45794 ( .A1(n59710), .A2(n53628), .B(n77744), .C(
        n53628), .Y(n55750) );
  A2O1A1Ixp33_ASAP7_75t_SL U45795 ( .A1(n59554), .A2(n53628), .B(n77745), .C(
        n53628), .Y(n55751) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45796 ( .A1(n77746), .A2(n77730), .B(n55750), 
        .C(n53628), .D(n55751), .Y(n4256) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45797 ( .A1(n74237), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_4_), .B(
        n74236), .C(n53628), .D(n55748), .Y(n55749) );
  A2O1A1Ixp33_ASAP7_75t_SL U45798 ( .A1(n71869), .A2(n53628), .B(n58422), .C(
        n53628), .Y(n55746) );
  A2O1A1Ixp33_ASAP7_75t_SL U45799 ( .A1(n71835), .A2(n53628), .B(n57208), .C(
        n53628), .Y(n55747) );
  A2O1A1Ixp33_ASAP7_75t_SL U45800 ( .A1(n55746), .A2(n53628), .B(n55747), .C(
        n53628), .Y(n72390) );
  A2O1A1Ixp33_ASAP7_75t_SL U45801 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_), 
        .A2(n53628), .B(n71601), .C(n53628), .Y(n55745) );
  A2O1A1Ixp33_ASAP7_75t_SL U45802 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .A2(n53628), .B(n71540), .C(n53628), .Y(n55743) );
  A2O1A1Ixp33_ASAP7_75t_SL U45803 ( .A1(n65953), .A2(n53628), .B(n55736), .C(
        n55737), .Y(n55738) );
  A2O1A1Ixp33_ASAP7_75t_SL U45804 ( .A1(n65952), .A2(n66022), .B(n55738), .C(
        n53628), .Y(n55739) );
  A2O1A1Ixp33_ASAP7_75t_SL U45805 ( .A1(n53628), .A2(n59631), .B(n73381), .C(
        n55507), .Y(n73391) );
  A2O1A1Ixp33_ASAP7_75t_SL U45806 ( .A1(n70139), .A2(n53628), .B(n55734), .C(
        n53628), .Y(n70163) );
  A2O1A1Ixp33_ASAP7_75t_SL U45807 ( .A1(n76394), .A2(n53628), .B(n55731), .C(
        n53628), .Y(n76459) );
  A2O1A1Ixp33_ASAP7_75t_SL U45808 ( .A1(n74690), .A2(n53628), .B(n55730), .C(
        n53628), .Y(n74703) );
  A2O1A1Ixp33_ASAP7_75t_SL U45809 ( .A1(n59850), .A2(n53628), .B(n55729), .C(
        n53628), .Y(n77147) );
  A2O1A1Ixp33_ASAP7_75t_SL U45810 ( .A1(n68614), .A2(n68615), .B(n75057), .C(
        n53628), .Y(n68620) );
  A2O1A1Ixp33_ASAP7_75t_SL U45811 ( .A1(n57203), .A2(n53628), .B(n71993), .C(
        n53628), .Y(n55723) );
  A2O1A1Ixp33_ASAP7_75t_SL U45812 ( .A1(n57127), .A2(n53628), .B(n72005), .C(
        n53628), .Y(n55724) );
  A2O1A1Ixp33_ASAP7_75t_SL U45813 ( .A1(n71995), .A2(n53628), .B(n57123), .C(
        n53628), .Y(n55725) );
  A2O1A1Ixp33_ASAP7_75t_SL U45814 ( .A1(n55724), .A2(n53628), .B(n55725), .C(
        n53628), .Y(n55726) );
  A2O1A1Ixp33_ASAP7_75t_SL U45815 ( .A1(n57125), .A2(n53628), .B(n71994), .C(
        n55726), .Y(n55727) );
  A2O1A1Ixp33_ASAP7_75t_SL U45816 ( .A1(n55723), .A2(n53628), .B(n55727), .C(
        n53628), .Y(n72186) );
  A2O1A1Ixp33_ASAP7_75t_SL U45817 ( .A1(n57208), .A2(n53628), .B(n72341), .C(
        n53628), .Y(n55717) );
  A2O1A1Ixp33_ASAP7_75t_SL U45818 ( .A1(n55717), .A2(n53628), .B(n55720), .C(
        n53628), .Y(n55721) );
  A2O1A1Ixp33_ASAP7_75t_SL U45819 ( .A1(n65545), .A2(n53628), .B(n55716), .C(
        n53628), .Y(n65419) );
  A2O1A1Ixp33_ASAP7_75t_SL U45820 ( .A1(n61509), .A2(n53628), .B(n61510), .C(
        n53628), .Y(n55714) );
  A2O1A1Ixp33_ASAP7_75t_SL U45821 ( .A1(n59577), .A2(n53628), .B(n55712), .C(
        n53628), .Y(n62089) );
  A2O1A1Ixp33_ASAP7_75t_SL U45822 ( .A1(n67463), .A2(n53628), .B(n58851), .C(
        n53628), .Y(n55709) );
  OAI21xp5_ASAP7_75t_SL U45823 ( .A1(n67945), .A2(n53565), .B(n53628), .Y(
        n55703) );
  A2O1A1Ixp33_ASAP7_75t_SL U45824 ( .A1(n58658), .A2(n53628), .B(n67241), .C(
        n55704), .Y(n57026) );
  A2O1A1Ixp33_ASAP7_75t_SL U45825 ( .A1(n72675), .A2(n53628), .B(n55481), .C(
        n55482), .Y(n27977) );
  A2O1A1Ixp33_ASAP7_75t_SL U45826 ( .A1(n73658), .A2(n53628), .B(n73655), .C(
        n53628), .Y(n55700) );
  A2O1A1Ixp33_ASAP7_75t_SL U45827 ( .A1(n73661), .A2(n53628), .B(n55700), .C(
        n73660), .Y(n3277) );
  A2O1A1Ixp33_ASAP7_75t_SL U45828 ( .A1(n71522), .A2(n53628), .B(n55695), .C(
        n53628), .Y(n55696) );
  A2O1A1Ixp33_ASAP7_75t_SL U45829 ( .A1(n69873), .A2(n69953), .B(n55693), .C(
        n53628), .Y(n55694) );
  A2O1A1Ixp33_ASAP7_75t_SL U45830 ( .A1(n69902), .A2(n53628), .B(n69956), .C(
        n55694), .Y(n3215) );
  A2O1A1Ixp33_ASAP7_75t_SL U45831 ( .A1(n77415), .A2(n53628), .B(n55691), .C(
        n53628), .Y(dwb_biu_N36) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45832 ( .A1(n77472), .A2(n77475), .B(n53628), 
        .C(n3086), .Y(n55244) );
  A2O1A1Ixp33_ASAP7_75t_SL U45833 ( .A1(n53628), .A2(n59689), .B(n3042), .C(
        n55477), .Y(n3043) );
  A2O1A1Ixp33_ASAP7_75t_SL U45834 ( .A1(n57074), .A2(n53628), .B(n2985), .C(
        n53628), .Y(n55682) );
  A2O1A1Ixp33_ASAP7_75t_SL U45835 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_10_), .A2(n53628), 
        .B(n77171), .C(n53628), .Y(n55680) );
  A2O1A1Ixp33_ASAP7_75t_SL U45836 ( .A1(n74904), .A2(n53628), .B(n74878), .C(
        n55680), .Y(n55681) );
  A2O1A1Ixp33_ASAP7_75t_SL U45837 ( .A1(n2843), .A2(n53628), .B(n57074), .C(
        n55679), .Y(n2844) );
  A2O1A1Ixp33_ASAP7_75t_SL U45838 ( .A1(n74797), .A2(n53628), .B(n55676), .C(
        n53628), .Y(n9565) );
  A2O1A1Ixp33_ASAP7_75t_SL U45839 ( .A1(n65275), .A2(n53628), .B(n55672), .C(
        n65346), .Y(n55673) );
  A2O1A1Ixp33_ASAP7_75t_SL U45840 ( .A1(n65275), .A2(n55672), .B(n55673), .C(
        n53628), .Y(n55674) );
  A2O1A1Ixp33_ASAP7_75t_SL U45841 ( .A1(n55674), .A2(n53628), .B(n55675), .C(
        n53628), .Y(n2482) );
  A2O1A1Ixp33_ASAP7_75t_SL U45842 ( .A1(n70470), .A2(n55455), .B(n70469), .C(
        n53628), .Y(n55456) );
  A2O1A1Ixp33_ASAP7_75t_SL U45843 ( .A1(n70551), .A2(n53628), .B(n74685), .C(
        n53628), .Y(n55461) );
  A2O1A1Ixp33_ASAP7_75t_SL U45844 ( .A1(n53628), .A2(n55460), .B(n55461), .C(
        n53628), .Y(n2412) );
  A2O1A1Ixp33_ASAP7_75t_SL U45845 ( .A1(n53628), .A2(n69735), .B(n69734), .C(
        n69762), .Y(n54835) );
  A2O1A1Ixp33_ASAP7_75t_SL U45846 ( .A1(n53628), .A2(n2107), .B(n57073), .C(
        n55442), .Y(n2108) );
  A2O1A1Ixp33_ASAP7_75t_SL U45847 ( .A1(n53628), .A2(n57074), .B(n2059), .C(
        n54833), .Y(n2060) );
  A2O1A1Ixp33_ASAP7_75t_SL U45848 ( .A1(n59627), .A2(n53628), .B(n73046), .C(
        n55665), .Y(n2017) );
  A2O1A1Ixp33_ASAP7_75t_SL U45849 ( .A1(n77980), .A2(n53628), .B(n77233), .C(
        n53628), .Y(n55663) );
  A2O1A1Ixp33_ASAP7_75t_SL U45850 ( .A1(n77246), .A2(n53628), .B(n1755), .C(
        n55662), .Y(n9339) );
  A2O1A1Ixp33_ASAP7_75t_SL U45851 ( .A1(n74934), .A2(n53628), .B(n59710), .C(
        n53628), .Y(n55658) );
  A2O1A1Ixp33_ASAP7_75t_SL U45852 ( .A1(n1717), .A2(n53628), .B(n55659), .C(
        n53628), .Y(n55660) );
  A2O1A1Ixp33_ASAP7_75t_SL U45853 ( .A1(n55658), .A2(n53628), .B(n55660), .C(
        n53628), .Y(n55661) );
  A2O1A1Ixp33_ASAP7_75t_SL U45854 ( .A1(n77847), .A2(n53628), .B(n77673), .C(
        n53628), .Y(n55657) );
  A2O1A1Ixp33_ASAP7_75t_SL U45855 ( .A1(n57114), .A2(n53628), .B(n1472), .C(
        n55655), .Y(n9300) );
  A2O1A1Ixp33_ASAP7_75t_SL U45856 ( .A1(n53628), .A2(n74641), .B(n1416), .C(
        n55426), .Y(n9324) );
  A2O1A1Ixp33_ASAP7_75t_SL U45857 ( .A1(n77287), .A2(n53628), .B(n76634), .C(
        n53628), .Y(n55653) );
  A2O1A1Ixp33_ASAP7_75t_SL U45858 ( .A1(n4097), .A2(n53628), .B(n55646), .C(
        n53628), .Y(n55647) );
  A2O1A1Ixp33_ASAP7_75t_SL U45859 ( .A1(n75631), .A2(n59701), .B(n55647), .C(
        n53628), .Y(n55648) );
  A2O1A1Ixp33_ASAP7_75t_SL U45860 ( .A1(n75632), .A2(n53628), .B(n77249), .C(
        n55648), .Y(n9166) );
  A2O1A1Ixp33_ASAP7_75t_SL U45861 ( .A1(n63277), .A2(n55403), .B(n63296), .C(
        n53628), .Y(n55404) );
  A2O1A1Ixp33_ASAP7_75t_SL U45862 ( .A1(n68911), .A2(n53628), .B(n55633), .C(
        n69053), .Y(n55634) );
  A2O1A1Ixp33_ASAP7_75t_SL U45863 ( .A1(n69052), .A2(n53628), .B(n55636), .C(
        n53628), .Y(n55637) );
  A2O1A1Ixp33_ASAP7_75t_SL U45864 ( .A1(n76906), .A2(n53628), .B(n55634), .C(
        n55639), .Y(n55640) );
  A2O1A1Ixp33_ASAP7_75t_SL U45865 ( .A1(n69112), .A2(n53628), .B(n69091), .C(
        n69111), .Y(n55623) );
  A2O1A1Ixp33_ASAP7_75t_SL U45866 ( .A1(n69092), .A2(n53628), .B(n76906), .C(
        n53628), .Y(n55625) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45867 ( .A1(n57079), .A2(n55624), .B(n69093), 
        .C(n53628), .D(n55625), .Y(n55626) );
  A2O1A1Ixp33_ASAP7_75t_SL U45868 ( .A1(n69113), .A2(n53628), .B(n76906), .C(
        n53628), .Y(n55628) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45869 ( .A1(n59673), .A2(n77901), .B(n55627), 
        .C(n53628), .D(n55628), .Y(n55629) );
  A2O1A1Ixp33_ASAP7_75t_SL U45870 ( .A1(n74570), .A2(n53628), .B(n55607), .C(
        n74571), .Y(n55608) );
  A2O1A1Ixp33_ASAP7_75t_SL U45871 ( .A1(n76906), .A2(n53628), .B(n55609), .C(
        n53628), .Y(n55613) );
  A2O1A1Ixp33_ASAP7_75t_SL U45872 ( .A1(n55613), .A2(n53628), .B(n55614), .C(
        n53628), .Y(n55615) );
  A2O1A1Ixp33_ASAP7_75t_SL U45873 ( .A1(or1200_cpu_or1200_except_n288), .A2(
        n53628), .B(n77441), .C(n55606), .Y(or1200_cpu_or1200_except_n1785) );
  A2O1A1Ixp33_ASAP7_75t_SL U45874 ( .A1(n53628), .A2(n59688), .B(
        or1200_cpu_or1200_except_n410), .C(n54994), .Y(
        or1200_cpu_or1200_except_n411) );
  A2O1A1Ixp33_ASAP7_75t_SL U45875 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n437), .C(n55604), .Y(
        or1200_cpu_or1200_except_n438) );
  A2O1A1Ixp33_ASAP7_75t_SL U45876 ( .A1(n57074), .A2(n53628), .B(
        or1200_cpu_or1200_except_n476), .C(n55601), .Y(
        or1200_cpu_or1200_except_n477) );
  A2O1A1Ixp33_ASAP7_75t_SL U45877 ( .A1(or1200_cpu_or1200_except_n616), .A2(
        n53628), .B(n57093), .C(n55600), .Y(or1200_cpu_or1200_except_n1802) );
  A2O1A1Ixp33_ASAP7_75t_SL U45878 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n640), .C(n54127), .Y(
        or1200_cpu_or1200_except_n1810) );
  A2O1A1Ixp33_ASAP7_75t_SL U45879 ( .A1(or1200_cpu_or1200_except_n664), .A2(
        n53628), .B(n57093), .C(n55598), .Y(or1200_cpu_or1200_except_n1818) );
  A2O1A1Ixp33_ASAP7_75t_SL U45880 ( .A1(or1200_cpu_or1200_except_n684), .A2(
        n53628), .B(n55595), .C(n53628), .Y(n55596) );
  A2O1A1Ixp33_ASAP7_75t_SL U45881 ( .A1(n74245), .A2(n53628), .B(n74230), .C(
        n53628), .Y(n55592) );
  A2O1A1Ixp33_ASAP7_75t_SL U45882 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .A2(
        n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_2_), 
        .C(n53628), .Y(n55580) );
  A2O1A1Ixp33_ASAP7_75t_SL U45883 ( .A1(n72517), .A2(n72366), .B(n72482), .C(
        n53628), .Y(n55581) );
  A2O1A1Ixp33_ASAP7_75t_SL U45884 ( .A1(n57203), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_), 
        .C(n55581), .Y(n55582) );
  A2O1A1Ixp33_ASAP7_75t_SL U45885 ( .A1(n55580), .A2(n53628), .B(n55582), .C(
        n53628), .Y(n55583) );
  A2O1A1Ixp33_ASAP7_75t_SL U45886 ( .A1(n72489), .A2(n72492), .B(n55583), .C(
        n53628), .Y(n55584) );
  A2O1A1Ixp33_ASAP7_75t_SL U45887 ( .A1(n72507), .A2(n53628), .B(n72436), .C(
        n55584), .Y(n55585) );
  A2O1A1Ixp33_ASAP7_75t_SL U45888 ( .A1(n72488), .A2(n53628), .B(n72503), .C(
        n72500), .Y(n55586) );
  A2O1A1Ixp33_ASAP7_75t_SL U45889 ( .A1(n55585), .A2(n53628), .B(n55586), .C(
        n53628), .Y(n55587) );
  A2O1A1Ixp33_ASAP7_75t_SL U45890 ( .A1(n72499), .A2(n53628), .B(n72396), .C(
        n55591), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n59) );
  A2O1A1Ixp33_ASAP7_75t_SL U45891 ( .A1(n72132), .A2(n72154), .B(n71565), .C(
        n53628), .Y(n55575) );
  A2O1A1Ixp33_ASAP7_75t_SL U45892 ( .A1(n71628), .A2(n53628), .B(n71541), .C(
        n55576), .Y(n55577) );
  A2O1A1Ixp33_ASAP7_75t_SL U45893 ( .A1(n55574), .A2(n53628), .B(n55577), .C(
        n53628), .Y(n55578) );
  A2O1A1Ixp33_ASAP7_75t_SL U45894 ( .A1(n59699), .A2(n53628), .B(n70714), .C(
        n53628), .Y(n55568) );
  A2O1A1Ixp33_ASAP7_75t_SL U45895 ( .A1(n70805), .A2(n70794), .B(n55563), .C(
        n53628), .Y(n55564) );
  A2O1A1Ixp33_ASAP7_75t_SL U45896 ( .A1(n59698), .A2(n53628), .B(n55565), .C(
        n53628), .Y(n55566) );
  A2O1A1Ixp33_ASAP7_75t_SL U45897 ( .A1(n70859), .A2(n53628), .B(n70858), .C(
        n53628), .Y(n55559) );
  A2O1A1Ixp33_ASAP7_75t_SL U45898 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_22_), .C(n53937), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n169) );
  A2O1A1Ixp33_ASAP7_75t_SL U45899 ( .A1(n59698), .A2(n53628), .B(n55553), .C(
        n53628), .Y(n55554) );
  A2O1A1Ixp33_ASAP7_75t_SL U45900 ( .A1(n71083), .A2(n53628), .B(n71081), .C(
        n53628), .Y(n55555) );
  A2O1A1Ixp33_ASAP7_75t_SL U45901 ( .A1(n59697), .A2(n53628), .B(n70650), .C(
        n53628), .Y(n55552) );
  A2O1A1Ixp33_ASAP7_75t_SL U45902 ( .A1(n55552), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_start_i), .C(n53628), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n253) );
  A2O1A1Ixp33_ASAP7_75t_SL U45903 ( .A1(n59632), .A2(n73695), .B(n55136), .C(
        n53628), .Y(n73781) );
  A2O1A1Ixp33_ASAP7_75t_SL U45904 ( .A1(n74460), .A2(n53628), .B(n55551), .C(
        n53628), .Y(n74462) );
  A2O1A1Ixp33_ASAP7_75t_SL U45905 ( .A1(n62044), .A2(n53628), .B(n55543), .C(
        n53628), .Y(n55544) );
  A2O1A1Ixp33_ASAP7_75t_SL U45906 ( .A1(n55544), .A2(n53628), .B(n55548), .C(
        n53628), .Y(n62066) );
  A2O1A1Ixp33_ASAP7_75t_SL U45907 ( .A1(n76991), .A2(n53628), .B(n55542), .C(
        n53628), .Y(n77206) );
  A2O1A1Ixp33_ASAP7_75t_SL U45908 ( .A1(n62477), .A2(n53628), .B(n57312), .C(
        n55541), .Y(n77890) );
  A2O1A1Ixp33_ASAP7_75t_SL U45909 ( .A1(n62477), .A2(n53628), .B(n57068), .C(
        n55540), .Y(n77871) );
  A2O1A1Ixp33_ASAP7_75t_SL U45910 ( .A1(n62477), .A2(n53628), .B(n59578), .C(
        n55538), .Y(n77875) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45911 ( .A1(n58451), .A2(n55537), .B(n76580), 
        .C(n53628), .D(n76581), .Y(n4092) );
  A2O1A1Ixp33_ASAP7_75t_SL U45912 ( .A1(n57160), .A2(n53628), .B(n55536), .C(
        n53628), .Y(n63925) );
  A2O1A1Ixp33_ASAP7_75t_SL U45913 ( .A1(n57168), .A2(n53628), .B(n1027), .C(
        n53628), .Y(n55535) );
  A2O1A1Ixp33_ASAP7_75t_SL U45914 ( .A1(n55535), .A2(n53628), .B(n77383), .C(
        n53628), .Y(n78183) );
  A2O1A1Ixp33_ASAP7_75t_SL U45915 ( .A1(n75082), .A2(n53628), .B(n75079), .C(
        n53628), .Y(n55534) );
  A2O1A1Ixp33_ASAP7_75t_SL U45916 ( .A1(n63782), .A2(n53628), .B(n55528), .C(
        n53628), .Y(n63430) );
  A2O1A1Ixp33_ASAP7_75t_SL U45917 ( .A1(n64172), .A2(n53628), .B(n55527), .C(
        n53628), .Y(n63786) );
  A2O1A1Ixp33_ASAP7_75t_SL U45918 ( .A1(n68782), .A2(n53628), .B(n55526), .C(
        n53628), .Y(n68768) );
  A2O1A1Ixp33_ASAP7_75t_SL U45919 ( .A1(n57123), .A2(n53628), .B(n72318), .C(
        n53628), .Y(n55521) );
  A2O1A1Ixp33_ASAP7_75t_SL U45920 ( .A1(n57203), .A2(n53628), .B(n72317), .C(
        n53628), .Y(n55522) );
  A2O1A1Ixp33_ASAP7_75t_SL U45921 ( .A1(n57125), .A2(n53628), .B(n72310), .C(
        n53628), .Y(n55523) );
  O2A1O1Ixp5_ASAP7_75t_SL U45922 ( .A1(n55521), .A2(n55522), .B(n53628), .C(
        n55523), .Y(n55524) );
  A2O1A1Ixp33_ASAP7_75t_SL U45923 ( .A1(n57127), .A2(n53628), .B(n72311), .C(
        n55524), .Y(n72464) );
  A2O1A1Ixp33_ASAP7_75t_SL U45924 ( .A1(n71899), .A2(n72163), .B(n57207), .C(
        n53628), .Y(n55518) );
  A2O1A1Ixp33_ASAP7_75t_SL U45925 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_), 
        .A2(n53628), .B(n57208), .C(n55518), .Y(n55519) );
  A2O1A1Ixp33_ASAP7_75t_SL U45926 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_), 
        .A2(n53628), .B(n71890), .C(n53628), .Y(n55520) );
  A2O1A1Ixp33_ASAP7_75t_SL U45927 ( .A1(n53628), .A2(n65743), .B(n65646), .C(
        n53628), .Y(n55514) );
  A2O1A1Ixp33_ASAP7_75t_SL U45928 ( .A1(n65859), .A2(n53628), .B(n65653), .C(
        n53628), .Y(n55515) );
  A2O1A1Ixp33_ASAP7_75t_SL U45929 ( .A1(n65711), .A2(n53628), .B(n66181), .C(
        n55516), .Y(n55517) );
  A2O1A1Ixp33_ASAP7_75t_SL U45930 ( .A1(n55514), .A2(n53628), .B(n55517), .C(
        n53628), .Y(n66101) );
  A2O1A1Ixp33_ASAP7_75t_SL U45931 ( .A1(n66022), .A2(n65958), .B(n55511), .C(
        n53628), .Y(n55512) );
  O2A1O1Ixp33_ASAP7_75t_SL U45932 ( .A1(n57201), .A2(n63177), .B(n53628), .C(
        n55508), .Y(n63180) );
  A2O1A1Ixp33_ASAP7_75t_SL U45933 ( .A1(n61418), .A2(n76753), .B(n55504), .C(
        n53628), .Y(n61423) );
  A2O1A1Ixp33_ASAP7_75t_SL U45934 ( .A1(or1200_cpu_or1200_except_n498), .A2(
        n61651), .B(n62263), .C(n53628), .Y(n54226) );
  A2O1A1Ixp33_ASAP7_75t_SL U45935 ( .A1(n62464), .A2(n53628), .B(n55502), .C(
        n55503), .Y(n76299) );
  A2O1A1Ixp33_ASAP7_75t_SL U45936 ( .A1(n63886), .A2(n55500), .B(n64747), .C(
        n53628), .Y(n65105) );
  A2O1A1Ixp33_ASAP7_75t_SL U45937 ( .A1(or1200_cpu_or1200_mult_mac_n259), .A2(
        n53628), .B(n55498), .C(n53628), .Y(n75651) );
  A2O1A1Ixp33_ASAP7_75t_SL U45938 ( .A1(n71380), .A2(n55496), .B(n71385), .C(
        n53628), .Y(n71400) );
  A2O1A1Ixp33_ASAP7_75t_SL U45939 ( .A1(n53628), .A2(n78339), .B(n57190), .C(
        n54548), .Y(n72937) );
  A2O1A1Ixp33_ASAP7_75t_SL U45940 ( .A1(n77090), .A2(
        or1200_cpu_or1200_fpu_result_conv[23]), .B(n55493), .C(n53628), .Y(
        n55494) );
  A2O1A1Ixp33_ASAP7_75t_SL U45941 ( .A1(or1200_cpu_or1200_mult_mac_n187), .A2(
        n53628), .B(n75723), .C(n55494), .Y(n75578) );
  A2O1A1Ixp33_ASAP7_75t_SL U45942 ( .A1(n57685), .A2(n53628), .B(n55491), .C(
        n57684), .Y(n59247) );
  A2O1A1Ixp33_ASAP7_75t_SL U45943 ( .A1(n57218), .A2(n53628), .B(n57120), .C(
        n53628), .Y(n55490) );
  A2O1A1Ixp33_ASAP7_75t_SL U45944 ( .A1(n53628), .A2(n59549), .B(n61979), .C(
        n57120), .Y(n55270) );
  A2O1A1Ixp33_ASAP7_75t_SL U45945 ( .A1(n67077), .A2(n53628), .B(n55483), .C(
        n53628), .Y(n55484) );
  A2O1A1Ixp33_ASAP7_75t_SL U45946 ( .A1(n67078), .A2(n59447), .B(n55484), .C(
        n53628), .Y(n67132) );
  A2O1A1Ixp33_ASAP7_75t_SL U45947 ( .A1(n53628), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[6]), .B(n73563), 
        .C(n54713), .Y(n3274) );
  A2O1A1Ixp33_ASAP7_75t_SL U45948 ( .A1(n53628), .A2(n69902), .B(n70001), .C(
        n55249), .Y(n3213) );
  A2O1A1Ixp33_ASAP7_75t_SL U45949 ( .A1(n53628), .A2(n70582), .B(n70574), .C(
        n53628), .Y(n54864) );
  A2O1A1Ixp33_ASAP7_75t_SL U45950 ( .A1(n70575), .A2(n53628), .B(n70579), .C(
        n53628), .Y(n54869) );
  A2O1A1Ixp33_ASAP7_75t_SL U45951 ( .A1(n53628), .A2(n54869), .B(n54864), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[3]), .Y(
        n54870) );
  A2O1A1Ixp33_ASAP7_75t_SL U45952 ( .A1(n53628), .A2(n57144), .B(n55058), .C(
        n55059), .Y(n3001) );
  A2O1A1Ixp33_ASAP7_75t_SL U45953 ( .A1(n2941), .A2(n53628), .B(n55471), .C(
        n53628), .Y(n55472) );
  A2O1A1Ixp33_ASAP7_75t_SL U45954 ( .A1(n77194), .A2(n77193), .B(n77196), .C(
        n53628), .Y(n55240) );
  A2O1A1Ixp33_ASAP7_75t_SL U45955 ( .A1(n53628), .A2(n57074), .B(n2666), .C(
        n55236), .Y(n2667) );
  A2O1A1Ixp33_ASAP7_75t_SL U45956 ( .A1(n70540), .A2(n53628), .B(n74674), .C(
        n53628), .Y(n55447) );
  A2O1A1Ixp33_ASAP7_75t_SL U45957 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_6_), .A2(
        n53628), .B(n59633), .C(n53628), .Y(n55448) );
  A2O1A1Ixp33_ASAP7_75t_SL U45958 ( .A1(n55447), .A2(n53628), .B(n55448), .C(
        n53628), .Y(n55449) );
  A2O1A1Ixp33_ASAP7_75t_SL U45959 ( .A1(n70541), .A2(n55450), .B(n55451), .C(
        n53628), .Y(n55452) );
  A2O1A1Ixp33_ASAP7_75t_SL U45960 ( .A1(n2196), .A2(n53628), .B(n55443), .C(
        n53628), .Y(n55444) );
  A2O1A1Ixp33_ASAP7_75t_SL U45961 ( .A1(n2073), .A2(n53628), .B(n59689), .C(
        n55441), .Y(n2074) );
  A2O1A1Ixp33_ASAP7_75t_SL U45962 ( .A1(n53628), .A2(n59627), .B(n72779), .C(
        n55219), .Y(n1952) );
  A2O1A1Ixp33_ASAP7_75t_SL U45963 ( .A1(n59626), .A2(n53628), .B(n78372), .C(
        n53628), .Y(n55438) );
  A2O1A1Ixp33_ASAP7_75t_SL U45964 ( .A1(n59680), .A2(n53628), .B(n1807), .C(
        n53628), .Y(n55435) );
  A2O1A1Ixp33_ASAP7_75t_SL U45965 ( .A1(n59680), .A2(n77968), .B(n55435), .C(
        n53628), .Y(n55436) );
  A2O1A1Ixp33_ASAP7_75t_SL U45966 ( .A1(n77847), .A2(n53628), .B(n77583), .C(
        n55433), .Y(n55434) );
  A2O1A1Ixp33_ASAP7_75t_SL U45967 ( .A1(n77584), .A2(n77675), .B(n55434), .C(
        n53628), .Y(n1715) );
  A2O1A1Ixp33_ASAP7_75t_SL U45968 ( .A1(n57114), .A2(n53628), .B(n1470), .C(
        n55432), .Y(n9299) );
  A2O1A1Ixp33_ASAP7_75t_SL U45969 ( .A1(n53628), .A2(n74641), .B(n1404), .C(
        n55214), .Y(n9321) );
  A2O1A1Ixp33_ASAP7_75t_SL U45970 ( .A1(n53628), .A2(n74641), .B(n1378), .C(
        n55012), .Y(n9314) );
  A2O1A1Ixp33_ASAP7_75t_SL U45971 ( .A1(n77287), .A2(n53628), .B(n77140), .C(
        n53628), .Y(n55419) );
  A2O1A1Ixp33_ASAP7_75t_SL U45972 ( .A1(n1121), .A2(n53628), .B(n76892), .C(
        n53628), .Y(n55417) );
  A2O1A1Ixp33_ASAP7_75t_SL U45973 ( .A1(n59703), .A2(n53628), .B(n55416), .C(
        n53628), .Y(n51950) );
  A2O1A1Ixp33_ASAP7_75t_SL U45974 ( .A1(n4132), .A2(n53628), .B(n55413), .C(
        n53628), .Y(n55414) );
  A2O1A1Ixp33_ASAP7_75t_SL U45975 ( .A1(n63969), .A2(n59701), .B(n55414), .C(
        n53628), .Y(n55415) );
  A2O1A1Ixp33_ASAP7_75t_SL U45976 ( .A1(n823), .A2(n53628), .B(n76523), .C(
        n55415), .Y(n9183) );
  A2O1A1Ixp33_ASAP7_75t_SL U45977 ( .A1(n63278), .A2(n53628), .B(n57486), .C(
        n53628), .Y(n55405) );
  A2O1A1Ixp33_ASAP7_75t_SL U45978 ( .A1(n59656), .A2(n53628), .B(n67227), .C(
        n53628), .Y(n55406) );
  A2O1A1Ixp33_ASAP7_75t_SL U45979 ( .A1(n63274), .A2(n53628), .B(n55393), .C(
        n59674), .Y(n55394) );
  A2O1A1Ixp33_ASAP7_75t_SL U45980 ( .A1(n63274), .A2(n55393), .B(n55394), .C(
        n53628), .Y(n55395) );
  A2O1A1Ixp33_ASAP7_75t_SL U45981 ( .A1(n63275), .A2(n53628), .B(n55393), .C(
        n53628), .Y(n55396) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U45982 ( .A1(n63275), .A2(n55393), .B(n76897), 
        .C(n53628), .D(n55396), .Y(n55397) );
  A2O1A1Ixp33_ASAP7_75t_SL U45983 ( .A1(n77585), .A2(n53628), .B(n65182), .C(
        n53628), .Y(n55398) );
  O2A1O1Ixp33_ASAP7_75t_SL U45984 ( .A1(n55395), .A2(n55397), .B(n53628), .C(
        n55398), .Y(n55399) );
  A2O1A1Ixp33_ASAP7_75t_SL U45985 ( .A1(or1200_cpu_or1200_mult_mac_n203), .A2(
        n53628), .B(n76889), .C(n53628), .Y(n55383) );
  A2O1A1Ixp33_ASAP7_75t_SL U45986 ( .A1(n77854), .A2(n76888), .B(n55383), .C(
        n53628), .Y(n55384) );
  A2O1A1Ixp33_ASAP7_75t_SL U45987 ( .A1(n76887), .A2(n53628), .B(n59671), .C(
        n55388), .Y(n55389) );
  A2O1A1Ixp33_ASAP7_75t_SL U45988 ( .A1(n76887), .A2(n57079), .B(n55388), .C(
        n53628), .Y(n55390) );
  A2O1A1Ixp33_ASAP7_75t_SL U45989 ( .A1(n76906), .A2(n53628), .B(n55386), .C(
        n55390), .Y(n55391) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U45990 ( .A1(n76897), .A2(n69021), .B(n53628), 
        .C(n55184), .Y(n55185) );
  A2O1A1Ixp33_ASAP7_75t_SL U45991 ( .A1(n69021), .A2(n57079), .B(n55183), .C(
        n53628), .Y(n55188) );
  A2O1A1Ixp33_ASAP7_75t_SL U45992 ( .A1(n57080), .A2(n69020), .B(n55182), .C(
        n53628), .Y(n55189) );
  A2O1A1Ixp33_ASAP7_75t_SL U45993 ( .A1(or1200_cpu_or1200_mult_mac_n223), .A2(
        n53628), .B(n76909), .C(n55191), .Y(or1200_cpu_or1200_mult_mac_n1615)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U45994 ( .A1(n76906), .A2(n53628), .B(n74116), .C(
        n74115), .Y(n54798) );
  A2O1A1Ixp33_ASAP7_75t_SL U45995 ( .A1(n57080), .A2(n74116), .B(n74115), .C(
        n53628), .Y(n54799) );
  A2O1A1Ixp33_ASAP7_75t_SL U45996 ( .A1(n53628), .A2(n74117), .B(n59671), .C(
        n54799), .Y(n54800) );
  A2O1A1Ixp33_ASAP7_75t_SL U45997 ( .A1(n69313), .A2(n53628), .B(n59671), .C(
        n55378), .Y(n55379) );
  A2O1A1Ixp33_ASAP7_75t_SL U45998 ( .A1(n69313), .A2(n59672), .B(n55378), .C(
        n53628), .Y(n55380) );
  A2O1A1Ixp33_ASAP7_75t_SL U45999 ( .A1(n76906), .A2(n53628), .B(n69310), .C(
        n55380), .Y(n55381) );
  A2O1A1Ixp33_ASAP7_75t_SL U46000 ( .A1(or1200_cpu_or1200_except_n592), .A2(
        n53628), .B(n57072), .C(n55371), .Y(or1200_cpu_or1200_except_n1794) );
  A2O1A1Ixp33_ASAP7_75t_SL U46001 ( .A1(or1200_cpu_or1200_except_n625), .A2(
        n53628), .B(n57093), .C(n55370), .Y(or1200_cpu_or1200_except_n1805) );
  A2O1A1Ixp33_ASAP7_75t_SL U46002 ( .A1(or1200_cpu_or1200_except_n658), .A2(
        n53628), .B(n57093), .C(n55368), .Y(or1200_cpu_or1200_except_n1816) );
  A2O1A1Ixp33_ASAP7_75t_SL U46003 ( .A1(n2966), .A2(n1510), .B(n58037), .C(
        n53628), .Y(n55355) );
  A2O1A1Ixp33_ASAP7_75t_SL U46004 ( .A1(n76674), .A2(n76673), .B(n76672), .C(
        n53628), .Y(n55356) );
  A2O1A1Ixp33_ASAP7_75t_SL U46005 ( .A1(or1200_cpu_or1200_except_n552), .A2(
        n53628), .B(n55354), .C(n55367), .Y(or1200_cpu_or1200_except_n553) );
  A2O1A1Ixp33_ASAP7_75t_SL U46006 ( .A1(n894), .A2(n53628), .B(n53428), .C(
        n53628), .Y(n55352) );
  A2O1A1Ixp33_ASAP7_75t_SL U46007 ( .A1(n64011), .A2(n57090), .B(n55352), .C(
        n53628), .Y(n55353) );
  A2O1A1Ixp33_ASAP7_75t_SL U46008 ( .A1(n901), .A2(n53628), .B(n77276), .C(
        n55353), .Y(or1200_cpu_or1200_except_n629) );
  A2O1A1Ixp33_ASAP7_75t_SL U46009 ( .A1(n57123), .A2(n53628), .B(n72360), .C(
        n53628), .Y(n55341) );
  A2O1A1Ixp33_ASAP7_75t_SL U46010 ( .A1(n57125), .A2(n53628), .B(n72348), .C(
        n53628), .Y(n55342) );
  A2O1A1Ixp33_ASAP7_75t_SL U46011 ( .A1(n55341), .A2(n53628), .B(n55342), .C(
        n53628), .Y(n55343) );
  A2O1A1Ixp33_ASAP7_75t_SL U46012 ( .A1(n72507), .A2(n53628), .B(n72479), .C(
        n55346), .Y(n55347) );
  A2O1A1Ixp33_ASAP7_75t_SL U46013 ( .A1(n72508), .A2(n53628), .B(n72481), .C(
        n72500), .Y(n55348) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46014 ( .A1(n72490), .A2(n72480), .B(n55347), 
        .C(n53628), .D(n55348), .Y(n55349) );
  A2O1A1Ixp33_ASAP7_75t_SL U46015 ( .A1(n57192), .A2(n53628), .B(n72383), .C(
        n72469), .Y(n55350) );
  A2O1A1Ixp33_ASAP7_75t_SL U46016 ( .A1(n72499), .A2(n53628), .B(n72389), .C(
        n55351), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n61) );
  A2O1A1Ixp33_ASAP7_75t_SL U46017 ( .A1(n53628), .A2(n70716), .B(n59697), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_4_), .Y(n54972) );
  A2O1A1Ixp33_ASAP7_75t_SL U46018 ( .A1(n53628), .A2(n57211), .B(n28213), .C(
        n54974), .Y(n54975) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46019 ( .A1(n70797), .A2(n70783), .B(n53628), 
        .C(n59699), .Y(n54966) );
  A2O1A1Ixp33_ASAP7_75t_SL U46020 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_9_), .C(n54970), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n130) );
  A2O1A1Ixp33_ASAP7_75t_SL U46021 ( .A1(n70842), .A2(n70849), .B(n55336), .C(
        n53628), .Y(n55337) );
  A2O1A1Ixp33_ASAP7_75t_SL U46022 ( .A1(n55338), .A2(n53628), .B(n59699), .C(
        n53628), .Y(n55339) );
  A2O1A1Ixp33_ASAP7_75t_SL U46023 ( .A1(n66147), .A2(n53628), .B(n66104), .C(
        n53628), .Y(n55324) );
  A2O1A1Ixp33_ASAP7_75t_SL U46024 ( .A1(n66105), .A2(n53628), .B(n66106), .C(
        n53628), .Y(n55325) );
  A2O1A1Ixp33_ASAP7_75t_SL U46025 ( .A1(n66122), .A2(n53628), .B(n66102), .C(
        n53628), .Y(n55326) );
  A2O1A1Ixp33_ASAP7_75t_SL U46026 ( .A1(n66103), .A2(n53628), .B(n66153), .C(
        n53628), .Y(n55327) );
  A2O1A1Ixp33_ASAP7_75t_SL U46027 ( .A1(n55326), .A2(n53628), .B(n55327), .C(
        n53628), .Y(n55328) );
  A2O1A1Ixp33_ASAP7_75t_SL U46028 ( .A1(n66109), .A2(n53628), .B(n66160), .C(
        n53628), .Y(n55329) );
  A2O1A1Ixp33_ASAP7_75t_SL U46029 ( .A1(n66158), .A2(n53628), .B(n66107), .C(
        n53628), .Y(n55330) );
  A2O1A1Ixp33_ASAP7_75t_SL U46030 ( .A1(n66108), .A2(n53628), .B(n66156), .C(
        n53628), .Y(n55331) );
  O2A1O1Ixp5_ASAP7_75t_SL U46031 ( .A1(n55329), .A2(n55330), .B(n53628), .C(
        n55331), .Y(n55332) );
  O2A1O1Ixp5_ASAP7_75t_SL U46032 ( .A1(n55324), .A2(n55325), .B(n53628), .C(
        n55333), .Y(n55334) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46033 ( .A1(n66112), .A2(n55334), .B(n66111), 
        .C(n53628), .D(n55335), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n7) );
  A2O1A1Ixp33_ASAP7_75t_SL U46034 ( .A1(n71528), .A2(n53628), .B(n71527), .C(
        n53628), .Y(n55323) );
  A2O1A1Ixp33_ASAP7_75t_SL U46035 ( .A1(n71526), .A2(n53628), .B(n55323), .C(
        n53628), .Y(n71530) );
  A2O1A1Ixp33_ASAP7_75t_SL U46036 ( .A1(n66184), .A2(n53628), .B(n66185), .C(
        n53628), .Y(n55322) );
  A2O1A1Ixp33_ASAP7_75t_SL U46037 ( .A1(n55322), .A2(n53628), .B(n66186), .C(
        n53628), .Y(n74089) );
  A2O1A1Ixp33_ASAP7_75t_SL U46038 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[2]), 
        .A2(n73890), .B(n73869), .C(n53628), .Y(n74103) );
  A2O1A1Ixp33_ASAP7_75t_SL U46039 ( .A1(n74808), .A2(n53628), .B(n55318), .C(
        n53628), .Y(n74813) );
  A2O1A1Ixp33_ASAP7_75t_SL U46040 ( .A1(n57160), .A2(n53628), .B(n55314), .C(
        n53628), .Y(n63930) );
  A2O1A1Ixp33_ASAP7_75t_SL U46041 ( .A1(n57168), .A2(n53628), .B(n1018), .C(
        n53628), .Y(n55313) );
  A2O1A1Ixp33_ASAP7_75t_SL U46042 ( .A1(n55313), .A2(n53628), .B(n75631), .C(
        n53628), .Y(n78185) );
  A2O1A1Ixp33_ASAP7_75t_SL U46043 ( .A1(n65169), .A2(n65168), .B(n55310), .C(
        n53628), .Y(n65149) );
  A2O1A1Ixp33_ASAP7_75t_SL U46044 ( .A1(or1200_cpu_or1200_mult_mac_n211), .A2(
        n53628), .B(n55309), .C(n53628), .Y(n68873) );
  A2O1A1Ixp33_ASAP7_75t_SL U46045 ( .A1(n53628), .A2(n71869), .B(n57208), .C(
        n54743), .Y(n72285) );
  A2O1A1Ixp33_ASAP7_75t_SL U46046 ( .A1(n57203), .A2(n53628), .B(n72212), .C(
        n53628), .Y(n55304) );
  A2O1A1Ixp33_ASAP7_75t_SL U46047 ( .A1(n57123), .A2(n53628), .B(n72219), .C(
        n53628), .Y(n55305) );
  A2O1A1Ixp33_ASAP7_75t_SL U46048 ( .A1(n57125), .A2(n53628), .B(n72234), .C(
        n53628), .Y(n55306) );
  A2O1A1Ixp33_ASAP7_75t_SL U46049 ( .A1(n55305), .A2(n53628), .B(n55306), .C(
        n53628), .Y(n55307) );
  A2O1A1Ixp33_ASAP7_75t_SL U46050 ( .A1(n57127), .A2(n53628), .B(n72253), .C(
        n55307), .Y(n55308) );
  A2O1A1Ixp33_ASAP7_75t_SL U46051 ( .A1(n55304), .A2(n53628), .B(n55308), .C(
        n53628), .Y(n72371) );
  A2O1A1Ixp33_ASAP7_75t_SL U46052 ( .A1(n71899), .A2(n53628), .B(n71898), .C(
        n54246), .Y(n72120) );
  A2O1A1Ixp33_ASAP7_75t_SL U46053 ( .A1(n72308), .A2(n53628), .B(n57208), .C(
        n53628), .Y(n55298) );
  A2O1A1Ixp33_ASAP7_75t_SL U46054 ( .A1(n55298), .A2(n53628), .B(n55301), .C(
        n53628), .Y(n55302) );
  A2O1A1Ixp33_ASAP7_75t_SL U46055 ( .A1(n55295), .A2(n53628), .B(n55296), .C(
        n53628), .Y(n55297) );
  A2O1A1Ixp33_ASAP7_75t_SL U46056 ( .A1(or1200_cpu_or1200_mult_mac_n102), .A2(
        n53628), .B(n61826), .C(n55289), .Y(n61833) );
  A2O1A1Ixp33_ASAP7_75t_SL U46057 ( .A1(n61639), .A2(n53628), .B(n55287), .C(
        n53628), .Y(n55288) );
  A2O1A1Ixp33_ASAP7_75t_SL U46058 ( .A1(n64840), .A2(n55286), .B(n55288), .C(
        n53628), .Y(n61355) );
  A2O1A1Ixp33_ASAP7_75t_SL U46059 ( .A1(n59871), .A2(n53628), .B(n55285), .C(
        n53628), .Y(n75192) );
  A2O1A1Ixp33_ASAP7_75t_SL U46060 ( .A1(n77251), .A2(n53628), .B(n55284), .C(
        n53628), .Y(n76825) );
  A2O1A1Ixp33_ASAP7_75t_SL U46061 ( .A1(n75036), .A2(n53628), .B(n75038), .C(
        n53628), .Y(n55283) );
  A2O1A1Ixp33_ASAP7_75t_SL U46062 ( .A1(n71357), .A2(n53628), .B(n55278), .C(
        n53628), .Y(n55279) );
  A2O1A1Ixp33_ASAP7_75t_SL U46063 ( .A1(n58582), .A2(n53628), .B(n65783), .C(
        n55277), .Y(n65954) );
  A2O1A1Ixp33_ASAP7_75t_SL U46064 ( .A1(n74599), .A2(n53628), .B(n55275), .C(
        n53628), .Y(n76462) );
  A2O1A1Ixp33_ASAP7_75t_SL U46065 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[21]), .A2(
        n53628), .B(n55274), .C(n53628), .Y(n73085) );
  A2O1A1Ixp33_ASAP7_75t_SL U46066 ( .A1(n57190), .A2(n53628), .B(n78431), .C(
        n55273), .Y(n72902) );
  A2O1A1Ixp33_ASAP7_75t_SL U46067 ( .A1(n57057), .A2(n57141), .B(n64090), .C(
        n53628), .Y(n55272) );
  A2O1A1Ixp33_ASAP7_75t_SL U46068 ( .A1(n57212), .A2(n53628), .B(n1571), .C(
        n53628), .Y(n55271) );
  A2O1A1Ixp33_ASAP7_75t_SL U46069 ( .A1(n55271), .A2(n53628), .B(n74018), .C(
        n53628), .Y(n76338) );
  A2O1A1Ixp33_ASAP7_75t_SL U46070 ( .A1(n57120), .A2(n53628), .B(n77732), .C(
        n53628), .Y(n55269) );
  A2O1A1Ixp33_ASAP7_75t_SL U46071 ( .A1(n59662), .A2(n53628), .B(n57405), .C(
        n53628), .Y(n55260) );
  A2O1A1Ixp33_ASAP7_75t_SL U46072 ( .A1(n57277), .A2(n59662), .B(n55260), .C(
        n53628), .Y(n55261) );
  A2O1A1Ixp33_ASAP7_75t_SL U46073 ( .A1(n66568), .A2(n55259), .B(n55261), .C(
        n53628), .Y(n68596) );
  A2O1A1Ixp33_ASAP7_75t_SL U46074 ( .A1(n53628), .A2(n59602), .B(n75927), .C(
        n54539), .Y(n63214) );
  A2O1A1Ixp33_ASAP7_75t_SL U46075 ( .A1(n58851), .A2(n53628), .B(n66796), .C(
        n55257), .Y(n55258) );
  A2O1A1Ixp33_ASAP7_75t_SL U46076 ( .A1(n66797), .A2(n53628), .B(n55256), .C(
        n55258), .Y(n68466) );
  A2O1A1Ixp33_ASAP7_75t_SL U46077 ( .A1(n53628), .A2(n72673), .B(n72675), .C(
        n72674), .Y(n55071) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46078 ( .A1(n73474), .A2(n73475), .B(n53628), 
        .C(n73476), .Y(n55254) );
  A2O1A1Ixp33_ASAP7_75t_SL U46079 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[4]), .A2(n53628), .B(
        n59704), .C(n53628), .Y(n55251) );
  A2O1A1Ixp33_ASAP7_75t_SL U46080 ( .A1(n73829), .A2(n53628), .B(n55251), .C(
        n53628), .Y(n55252) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46081 ( .A1(n73656), .A2(n73657), .B(n53628), 
        .C(n73659), .Y(n55066) );
  A2O1A1Ixp33_ASAP7_75t_SL U46082 ( .A1(n53628), .A2(n73661), .B(n55067), .C(
        n73660), .Y(n3276) );
  A2O1A1Ixp33_ASAP7_75t_SL U46083 ( .A1(n77767), .A2(n53628), .B(n55244), .C(
        n53628), .Y(n55245) );
  A2O1A1Ixp33_ASAP7_75t_SL U46084 ( .A1(n59689), .A2(n53628), .B(n3036), .C(
        n54711), .Y(n3037) );
  O2A1O1Ixp33_ASAP7_75t_SL U46085 ( .A1(n75541), .A2(n75543), .B(n53628), .C(
        n55056), .Y(n55057) );
  A2O1A1Ixp33_ASAP7_75t_SL U46086 ( .A1(n53628), .A2(n77142), .B(n3418), .C(
        n55050), .Y(or1200_cpu_to_sr[3]) );
  A2O1A1Ixp33_ASAP7_75t_SL U46087 ( .A1(n53628), .A2(n57074), .B(n2791), .C(
        n54856), .Y(n2792) );
  A2O1A1Ixp33_ASAP7_75t_SL U46088 ( .A1(iwb_ack_i), .A2(n53628), .B(n55237), 
        .C(n53628), .Y(n55238) );
  A2O1A1Ixp33_ASAP7_75t_SL U46089 ( .A1(n2558), .A2(n53628), .B(n55232), .C(
        n53628), .Y(n55233) );
  A2O1A1Ixp33_ASAP7_75t_SL U46090 ( .A1(n70531), .A2(n53628), .B(n55230), .C(
        n53628), .Y(n55231) );
  A2O1A1Ixp33_ASAP7_75t_SL U46091 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[0]), .A2(n55229), .B(
        n55231), .C(n53628), .Y(n2449) );
  A2O1A1Ixp33_ASAP7_75t_SL U46092 ( .A1(n74662), .A2(n53628), .B(n70553), .C(
        n53628), .Y(n55223) );
  A2O1A1Ixp33_ASAP7_75t_SL U46093 ( .A1(n2440), .A2(n53628), .B(n70551), .C(
        n53628), .Y(n55224) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46094 ( .A1(n70468), .A2(n70302), .B(n55223), 
        .C(n53628), .D(n55224), .Y(n2400) );
  A2O1A1Ixp33_ASAP7_75t_SL U46095 ( .A1(n2039), .A2(n53628), .B(n57073), .C(
        n55221), .Y(n2040) );
  A2O1A1Ixp33_ASAP7_75t_SL U46096 ( .A1(n53628), .A2(n57144), .B(n77905), .C(
        n55027), .Y(n1805) );
  A2O1A1Ixp33_ASAP7_75t_SL U46097 ( .A1(n53628), .A2(n74934), .B(n59442), .C(
        n54328), .Y(n9492) );
  A2O1A1Ixp33_ASAP7_75t_SL U46098 ( .A1(n77649), .A2(n53628), .B(n55217), .C(
        n53628), .Y(n55218) );
  A2O1A1Ixp33_ASAP7_75t_SL U46099 ( .A1(n77890), .A2(n77672), .B(n55218), .C(
        n53628), .Y(n1684) );
  A2O1A1Ixp33_ASAP7_75t_SL U46100 ( .A1(n57114), .A2(n53628), .B(n1486), .C(
        n55216), .Y(n9307) );
  A2O1A1Ixp33_ASAP7_75t_SL U46101 ( .A1(n4124), .A2(n53628), .B(n55204), .C(
        n53628), .Y(n55205) );
  A2O1A1Ixp33_ASAP7_75t_SL U46102 ( .A1(n63925), .A2(n59701), .B(n55205), .C(
        n53628), .Y(n55206) );
  A2O1A1Ixp33_ASAP7_75t_SL U46103 ( .A1(n807), .A2(n53628), .B(n76523), .C(
        n55206), .Y(n9179) );
  A2O1A1Ixp33_ASAP7_75t_SL U46104 ( .A1(n63363), .A2(n53628), .B(n55007), .C(
        n55008), .Y(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N11) );
  A2O1A1Ixp33_ASAP7_75t_SL U46105 ( .A1(n63509), .A2(n63508), .B(n63517), .C(
        n53628), .Y(n53970) );
  A2O1A1Ixp33_ASAP7_75t_SL U46106 ( .A1(n53628), .A2(n76897), .B(n53975), .C(
        n53976), .Y(n53977) );
  A2O1A1Ixp33_ASAP7_75t_SL U46107 ( .A1(n53628), .A2(
        or1200_cpu_or1200_mult_mac_n171), .B(n76889), .C(n53978), .Y(
        or1200_cpu_or1200_mult_mac_n1578) );
  A2O1A1Ixp33_ASAP7_75t_SL U46108 ( .A1(n68877), .A2(n53628), .B(n68872), .C(
        n53628), .Y(n55194) );
  A2O1A1Ixp33_ASAP7_75t_SL U46109 ( .A1(n76906), .A2(n53628), .B(n68861), .C(
        n55198), .Y(n55199) );
  A2O1A1Ixp33_ASAP7_75t_SL U46110 ( .A1(n69057), .A2(n53628), .B(n55181), .C(
        n53628), .Y(n55182) );
  A2O1A1Ixp33_ASAP7_75t_SL U46111 ( .A1(n69021), .A2(n53628), .B(n55183), .C(
        n53628), .Y(n55184) );
  A2O1A1Ixp33_ASAP7_75t_SL U46112 ( .A1(n59673), .A2(n77992), .B(n55185), .C(
        n53628), .Y(n55186) );
  A2O1A1Ixp33_ASAP7_75t_SL U46113 ( .A1(n55187), .A2(n53628), .B(n55190), .C(
        n53628), .Y(n55191) );
  A2O1A1Ixp33_ASAP7_75t_SL U46114 ( .A1(n75128), .A2(n53628), .B(n75117), .C(
        n53628), .Y(n55170) );
  O2A1O1Ixp33_ASAP7_75t_SL U46115 ( .A1(n55170), .A2(n75133), .B(n53628), .C(
        n76906), .Y(n55171) );
  A2O1A1Ixp33_ASAP7_75t_SL U46116 ( .A1(n75121), .A2(n53628), .B(n75118), .C(
        n75119), .Y(n55173) );
  A2O1A1Ixp33_ASAP7_75t_SL U46117 ( .A1(n59671), .A2(n53628), .B(n55173), .C(
        n53628), .Y(n55176) );
  A2O1A1Ixp33_ASAP7_75t_SL U46118 ( .A1(n55176), .A2(n53628), .B(n55172), .C(
        n53628), .Y(n55177) );
  A2O1A1Ixp33_ASAP7_75t_SL U46119 ( .A1(n55170), .A2(n53628), .B(n75133), .C(
        n57080), .Y(n55178) );
  A2O1A1Ixp33_ASAP7_75t_SL U46120 ( .A1(n55171), .A2(n53628), .B(n55175), .C(
        n55179), .Y(n55180) );
  A2O1A1Ixp33_ASAP7_75t_SL U46121 ( .A1(or1200_cpu_or1200_except_n628), .A2(
        n53628), .B(n57072), .C(n55165), .Y(or1200_cpu_or1200_except_n1806) );
  A2O1A1Ixp33_ASAP7_75t_SL U46122 ( .A1(or1200_cpu_or1200_except_n634), .A2(
        n53628), .B(n57072), .C(n55164), .Y(or1200_cpu_or1200_except_n1808) );
  A2O1A1Ixp33_ASAP7_75t_SL U46123 ( .A1(n858), .A2(n53628), .B(n53428), .C(
        n53628), .Y(n55161) );
  A2O1A1Ixp33_ASAP7_75t_SL U46124 ( .A1(n63960), .A2(n57090), .B(n55161), .C(
        n53628), .Y(n55162) );
  A2O1A1Ixp33_ASAP7_75t_SL U46125 ( .A1(n865), .A2(n53628), .B(n77276), .C(
        n55162), .Y(or1200_cpu_or1200_except_n617) );
  A2O1A1Ixp33_ASAP7_75t_SL U46126 ( .A1(n76671), .A2(n53628), .B(n57404), .C(
        n55160), .Y(or1200_cpu_or1200_except_n691) );
  A2O1A1Ixp33_ASAP7_75t_SL U46127 ( .A1(n74252), .A2(n55157), .B(n74276), .C(
        n53628), .Y(n55158) );
  A2O1A1Ixp33_ASAP7_75t_SL U46128 ( .A1(n74252), .A2(n53628), .B(n55157), .C(
        n55158), .Y(n55159) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46129 ( .A1(n72503), .A2(n72505), .B(n53628), 
        .C(n72504), .Y(n54980) );
  A2O1A1Ixp33_ASAP7_75t_SL U46130 ( .A1(n72502), .A2(n72501), .B(n54980), .C(
        n53628), .Y(n54981) );
  A2O1A1Ixp33_ASAP7_75t_SL U46131 ( .A1(n53628), .A2(n54978), .B(n54984), .C(
        n72515), .Y(n54985) );
  A2O1A1Ixp33_ASAP7_75t_SL U46132 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .A2(
        n72513), .B(n54985), .C(n53628), .Y(n54986) );
  A2O1A1Ixp33_ASAP7_75t_SL U46133 ( .A1(n53628), .A2(n70784), .B(n70775), .C(
        n53628), .Y(n54967) );
  A2O1A1Ixp33_ASAP7_75t_SL U46134 ( .A1(n70797), .A2(n53628), .B(n70783), .C(
        n53628), .Y(n54968) );
  A2O1A1Ixp33_ASAP7_75t_SL U46135 ( .A1(n53628), .A2(n59699), .B(n54968), .C(
        n54967), .Y(n54969) );
  A2O1A1Ixp33_ASAP7_75t_SL U46136 ( .A1(n53628), .A2(n54966), .B(n54967), .C(
        n54969), .Y(n54970) );
  A2O1A1Ixp33_ASAP7_75t_SL U46137 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_15_), .C(n54965), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n148) );
  A2O1A1Ixp33_ASAP7_75t_SL U46138 ( .A1(n66160), .A2(n53628), .B(n66099), .C(
        n53628), .Y(n55142) );
  A2O1A1Ixp33_ASAP7_75t_SL U46139 ( .A1(n66156), .A2(n53628), .B(n66100), .C(
        n53628), .Y(n55143) );
  A2O1A1Ixp33_ASAP7_75t_SL U46140 ( .A1(n66105), .A2(n53628), .B(n66098), .C(
        n53628), .Y(n55146) );
  A2O1A1Ixp33_ASAP7_75t_SL U46141 ( .A1(n66095), .A2(n53628), .B(n66096), .C(
        n53628), .Y(n55149) );
  A2O1A1Ixp33_ASAP7_75t_SL U46142 ( .A1(n66094), .A2(n55148), .B(n55149), .C(
        n53628), .Y(n55150) );
  A2O1A1Ixp33_ASAP7_75t_SL U46143 ( .A1(n66093), .A2(n53628), .B(n55147), .C(
        n55150), .Y(n55151) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46144 ( .A1(n66101), .A2(n55145), .B(n55146), 
        .C(n53628), .D(n55151), .Y(n55152) );
  A2O1A1Ixp33_ASAP7_75t_SL U46145 ( .A1(n66158), .A2(n53628), .B(n55144), .C(
        n55152), .Y(n55153) );
  O2A1O1Ixp5_ASAP7_75t_SL U46146 ( .A1(n55142), .A2(n55143), .B(n53628), .C(
        n55153), .Y(n55154) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46147 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_5_), .A2(n66138), 
        .B(n53628), .C(n66166), .Y(n55155) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46148 ( .A1(n55154), .A2(n66112), .B(n55155), 
        .C(n53628), .D(n55156), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n8) );
  A2O1A1Ixp33_ASAP7_75t_SL U46149 ( .A1(n57217), .A2(n73688), .B(n55139), .C(
        n53628), .Y(n55140) );
  A2O1A1Ixp33_ASAP7_75t_SL U46150 ( .A1(n71533), .A2(n53628), .B(n55132), .C(
        n53628), .Y(n71532) );
  A2O1A1Ixp33_ASAP7_75t_SL U46151 ( .A1(n74706), .A2(n53628), .B(n70382), .C(
        n55131), .Y(n70490) );
  A2O1A1Ixp33_ASAP7_75t_SL U46152 ( .A1(n77759), .A2(n53628), .B(n77758), .C(
        n53628), .Y(n55130) );
  A2O1A1Ixp33_ASAP7_75t_SL U46153 ( .A1(or1200_cpu_or1200_fpu_fpu_arith_done), 
        .A2(n55127), .B(n55129), .C(n53628), .Y(n74756) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46154 ( .A1(n75298), .A2(n74981), .B(n53628), 
        .C(n74982), .Y(n55125) );
  A2O1A1Ixp33_ASAP7_75t_SL U46155 ( .A1(n75429), .A2(n54596), .B(n54598), .C(
        n53628), .Y(n78117) );
  A2O1A1Ixp33_ASAP7_75t_SL U46156 ( .A1(n75190), .A2(n53628), .B(n75189), .C(
        n53628), .Y(n55123) );
  A2O1A1Ixp33_ASAP7_75t_SL U46157 ( .A1(n55123), .A2(n53628), .B(n75791), .C(
        n53628), .Y(n55124) );
  A2O1A1Ixp33_ASAP7_75t_SL U46158 ( .A1(n57168), .A2(n53628), .B(n910), .C(
        n53628), .Y(n55122) );
  A2O1A1Ixp33_ASAP7_75t_SL U46159 ( .A1(n55122), .A2(n53628), .B(n74961), .C(
        n53628), .Y(n78257) );
  A2O1A1Ixp33_ASAP7_75t_SL U46160 ( .A1(n63313), .A2(n53628), .B(n55118), .C(
        n63310), .Y(n63293) );
  A2O1A1Ixp33_ASAP7_75t_SL U46161 ( .A1(n65099), .A2(n65098), .B(n55115), .C(
        n53628), .Y(n65074) );
  A2O1A1Ixp33_ASAP7_75t_SL U46162 ( .A1(n77452), .A2(n53628), .B(n55111), .C(
        n53628), .Y(n77437) );
  A2O1A1Ixp33_ASAP7_75t_SL U46163 ( .A1(n59550), .A2(n53628), .B(n77741), .C(
        n53628), .Y(n55107) );
  A2O1A1Ixp33_ASAP7_75t_SL U46164 ( .A1(n59552), .A2(n53628), .B(n77745), .C(
        n53628), .Y(n55108) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46165 ( .A1(n78003), .A2(n77742), .B(n55107), 
        .C(n53628), .D(n55108), .Y(n4242) );
  A2O1A1Ixp33_ASAP7_75t_SL U46166 ( .A1(n53628), .A2(n71800), .B(n71679), .C(
        n54919), .Y(n54920) );
  A2O1A1Ixp33_ASAP7_75t_SL U46167 ( .A1(n57203), .A2(n53628), .B(n72234), .C(
        n53628), .Y(n55102) );
  A2O1A1Ixp33_ASAP7_75t_SL U46168 ( .A1(n57127), .A2(n53628), .B(n72309), .C(
        n53628), .Y(n55103) );
  A2O1A1Ixp33_ASAP7_75t_SL U46169 ( .A1(n72253), .A2(n53628), .B(n57123), .C(
        n53628), .Y(n55104) );
  A2O1A1Ixp33_ASAP7_75t_SL U46170 ( .A1(n55103), .A2(n53628), .B(n55104), .C(
        n53628), .Y(n55105) );
  A2O1A1Ixp33_ASAP7_75t_SL U46171 ( .A1(n57125), .A2(n53628), .B(n72306), .C(
        n55105), .Y(n55106) );
  A2O1A1Ixp33_ASAP7_75t_SL U46172 ( .A1(n55102), .A2(n53628), .B(n55106), .C(
        n53628), .Y(n72465) );
  A2O1A1Ixp33_ASAP7_75t_SL U46173 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .A2(n58611), .B(n54908), .C(n53628), .Y(n54909) );
  A2O1A1Ixp33_ASAP7_75t_SL U46174 ( .A1(n72154), .A2(n53628), .B(n57208), .C(
        n53628), .Y(n55096) );
  A2O1A1Ixp33_ASAP7_75t_SL U46175 ( .A1(n55096), .A2(n53628), .B(n55099), .C(
        n53628), .Y(n55100) );
  A2O1A1Ixp33_ASAP7_75t_SL U46176 ( .A1(n70990), .A2(n53628), .B(n70991), .C(
        n53628), .Y(n55095) );
  A2O1A1Ixp33_ASAP7_75t_SL U46177 ( .A1(n71792), .A2(n53628), .B(n71727), .C(
        n55094), .Y(n71730) );
  A2O1A1Ixp33_ASAP7_75t_SL U46178 ( .A1(n59626), .A2(n53628), .B(n78433), .C(
        n53628), .Y(n55093) );
  A2O1A1Ixp33_ASAP7_75t_SL U46179 ( .A1(n73047), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[2]), .B(n55093), 
        .C(n53628), .Y(n73027) );
  A2O1A1Ixp33_ASAP7_75t_SL U46180 ( .A1(n72813), .A2(n53628), .B(n55091), .C(
        n53628), .Y(n55092) );
  A2O1A1Ixp33_ASAP7_75t_SL U46181 ( .A1(n72990), .A2(n72814), .B(n55092), .C(
        n53628), .Y(n72851) );
  A2O1A1Ixp33_ASAP7_75t_SL U46182 ( .A1(n75218), .A2(n57191), .B(n55089), .C(
        n53628), .Y(n55090) );
  A2O1A1Ixp33_ASAP7_75t_SL U46183 ( .A1(or1200_cpu_or1200_mult_mac_n345), .A2(
        n53628), .B(n77073), .C(n55090), .Y(n75221) );
  A2O1A1Ixp33_ASAP7_75t_SL U46184 ( .A1(n71080), .A2(n53628), .B(n71083), .C(
        n53628), .Y(n55082) );
  A2O1A1Ixp33_ASAP7_75t_SL U46185 ( .A1(n71081), .A2(n53628), .B(n55082), .C(
        n53628), .Y(n71131) );
  A2O1A1Ixp33_ASAP7_75t_SL U46186 ( .A1(n64757), .A2(n53628), .B(n55081), .C(
        n53628), .Y(n76268) );
  OAI22xp5_ASAP7_75t_SL U46187 ( .A1(n57292), .A2(n75641), .B1(n66480), .B2(
        n75641), .Y(n54720) );
  A2O1A1Ixp33_ASAP7_75t_SL U46188 ( .A1(n66506), .A2(n66507), .B(n54722), .C(
        n53628), .Y(n66512) );
  A2O1A1Ixp33_ASAP7_75t_SL U46189 ( .A1(n64682), .A2(n53628), .B(n64683), .C(
        n64681), .Y(n55079) );
  A2O1A1Ixp33_ASAP7_75t_SL U46190 ( .A1(n64717), .A2(n53628), .B(n55079), .C(
        n55080), .Y(n64707) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46191 ( .A1(n57881), .A2(n77242), .B(n53628), 
        .C(n63130), .Y(n55078) );
  A2O1A1Ixp33_ASAP7_75t_SL U46192 ( .A1(n67974), .A2(n53628), .B(n67628), .C(
        n55076), .Y(n67797) );
  NOR2x1_ASAP7_75t_SL U46193 ( .A(n53588), .B(n57156), .Y(n55075) );
  A2O1A1Ixp33_ASAP7_75t_SL U46194 ( .A1(n72646), .A2(n55073), .B(n55071), .C(
        n53628), .Y(n55074) );
  A2O1A1Ixp33_ASAP7_75t_SL U46195 ( .A1(n73466), .A2(n73467), .B(n73468), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_6_)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46196 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[5]), .A2(n53628), .B(
        n59704), .C(n53628), .Y(n55068) );
  A2O1A1Ixp33_ASAP7_75t_SL U46197 ( .A1(n73829), .A2(n53628), .B(n55068), .C(
        n53628), .Y(n55069) );
  A2O1A1Ixp33_ASAP7_75t_SL U46198 ( .A1(n71512), .A2(n53628), .B(n78329), .C(
        n53628), .Y(n55063) );
  A2O1A1Ixp33_ASAP7_75t_SL U46199 ( .A1(n53628), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[3]), .B(
        n54864), .C(n53628), .Y(n54865) );
  A2O1A1Ixp33_ASAP7_75t_SL U46200 ( .A1(n70575), .A2(n53628), .B(n70579), .C(
        n53628), .Y(n54866) );
  A2O1A1Ixp33_ASAP7_75t_SL U46201 ( .A1(n61319), .A2(n53628), .B(n78067), .C(
        n55062), .Y(n9347) );
  A2O1A1Ixp33_ASAP7_75t_SL U46202 ( .A1(n74899), .A2(n55052), .B(n74885), .C(
        n53628), .Y(n55053) );
  A2O1A1Ixp33_ASAP7_75t_SL U46203 ( .A1(n53628), .A2(n57202), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[27]), .C(n54860), 
        .Y(n2858) );
  A2O1A1Ixp33_ASAP7_75t_SL U46204 ( .A1(n53628), .A2(n57074), .B(n2659), .C(
        n54193), .Y(n2660) );
  A2O1A1Ixp33_ASAP7_75t_SL U46205 ( .A1(n77427), .A2(n53628), .B(n2589), .C(
        n53628), .Y(n55045) );
  A2O1A1Ixp33_ASAP7_75t_SL U46206 ( .A1(n57144), .A2(n53628), .B(n55046), .C(
        n53628), .Y(n9495) );
  A2O1A1Ixp33_ASAP7_75t_SL U46207 ( .A1(n70478), .A2(n53628), .B(n70467), .C(
        n53628), .Y(n55039) );
  A2O1A1Ixp33_ASAP7_75t_SL U46208 ( .A1(n55039), .A2(n59621), .B(n55040), .C(
        n53628), .Y(n2447) );
  A2O1A1Ixp33_ASAP7_75t_SL U46209 ( .A1(n70461), .A2(n53628), .B(n70405), .C(
        n70370), .Y(n55035) );
  A2O1A1Ixp33_ASAP7_75t_SL U46210 ( .A1(n70485), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_11_), .B(
        n55035), .C(n53628), .Y(n55036) );
  A2O1A1Ixp33_ASAP7_75t_SL U46211 ( .A1(n70465), .A2(n53628), .B(n70483), .C(
        n55038), .Y(n2390) );
  A2O1A1Ixp33_ASAP7_75t_SL U46212 ( .A1(n69774), .A2(n69784), .B(n69782), .C(
        n53628), .Y(n55032) );
  A2O1A1Ixp33_ASAP7_75t_SL U46213 ( .A1(n57081), .A2(n53628), .B(n69776), .C(
        n53628), .Y(n55033) );
  A2O1A1Ixp33_ASAP7_75t_SL U46214 ( .A1(n70511), .A2(n53628), .B(n70422), .C(
        n53628), .Y(n55034) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46215 ( .A1(n55032), .A2(n59621), .B(n55033), 
        .C(n53628), .D(n55034), .Y(n2301) );
  A2O1A1Ixp33_ASAP7_75t_SL U46216 ( .A1(n59629), .A2(n53628), .B(n72779), .C(
        n55031), .Y(n1964) );
  A2O1A1Ixp33_ASAP7_75t_SL U46217 ( .A1(n53628), .A2(n1924), .B(n59689), .C(
        n54670), .Y(n1925) );
  A2O1A1Ixp33_ASAP7_75t_SL U46218 ( .A1(n59680), .A2(n53628), .B(n1847), .C(
        n53628), .Y(n55029) );
  A2O1A1Ixp33_ASAP7_75t_SL U46219 ( .A1(n59680), .A2(n77977), .B(n55029), .C(
        n53628), .Y(n55030) );
  A2O1A1Ixp33_ASAP7_75t_SL U46220 ( .A1(n76609), .A2(n53628), .B(n55028), .C(
        n55030), .Y(n18405) );
  A2O1A1Ixp33_ASAP7_75t_SL U46221 ( .A1(n1804), .A2(n53628), .B(n55025), .C(
        n53628), .Y(n55026) );
  A2O1A1Ixp33_ASAP7_75t_SL U46222 ( .A1(n77246), .A2(n53628), .B(n1719), .C(
        n55024), .Y(n9341) );
  A2O1A1Ixp33_ASAP7_75t_SL U46223 ( .A1(n77847), .A2(n53628), .B(n77585), .C(
        n53628), .Y(n55020) );
  A2O1A1Ixp33_ASAP7_75t_SL U46224 ( .A1(n77586), .A2(n53628), .B(n77639), .C(
        n53628), .Y(n55021) );
  O2A1O1Ixp5_ASAP7_75t_SL U46225 ( .A1(n55020), .A2(n55021), .B(n53628), .C(
        n55023), .Y(n1714) );
  A2O1A1Ixp33_ASAP7_75t_SL U46226 ( .A1(n57114), .A2(n53628), .B(n1478), .C(
        n55019), .Y(n9303) );
  A2O1A1Ixp33_ASAP7_75t_SL U46227 ( .A1(n1119), .A2(n1121), .B(n76891), .C(
        n53628), .Y(n54809) );
  A2O1A1Ixp33_ASAP7_75t_SL U46228 ( .A1(n77673), .A2(n53628), .B(n76890), .C(
        n53628), .Y(n54810) );
  A2O1A1Ixp33_ASAP7_75t_SL U46229 ( .A1(n4126), .A2(n53628), .B(n55009), .C(
        n53628), .Y(n55010) );
  A2O1A1Ixp33_ASAP7_75t_SL U46230 ( .A1(n63930), .A2(n59701), .B(n55010), .C(
        n53628), .Y(n55011) );
  A2O1A1Ixp33_ASAP7_75t_SL U46231 ( .A1(n811), .A2(n53628), .B(n76523), .C(
        n55011), .Y(n9180) );
  A2O1A1Ixp33_ASAP7_75t_SL U46232 ( .A1(or1200_cpu_or1200_mult_mac_n145), .A2(
        n53628), .B(n76889), .C(n54651), .Y(or1200_cpu_or1200_mult_mac_n1591)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46233 ( .A1(n69000), .A2(n53432), .B(n68999), .C(
        n53628), .Y(n54997) );
  A2O1A1Ixp33_ASAP7_75t_SL U46234 ( .A1(n54997), .A2(n53628), .B(n68997), .C(
        n53628), .Y(n54998) );
  A2O1A1Ixp33_ASAP7_75t_SL U46235 ( .A1(n54998), .A2(n53628), .B(n54996), .C(
        n53628), .Y(n54999) );
  A2O1A1Ixp33_ASAP7_75t_SL U46236 ( .A1(n69018), .A2(n53628), .B(n55000), .C(
        n59672), .Y(n55001) );
  A2O1A1Ixp33_ASAP7_75t_SL U46237 ( .A1(n54999), .A2(n53628), .B(n55001), .C(
        n55002), .Y(n55003) );
  A2O1A1Ixp33_ASAP7_75t_SL U46238 ( .A1(n75650), .A2(n69002), .B(n55003), .C(
        n53628), .Y(n55004) );
  A2O1A1Ixp33_ASAP7_75t_SL U46239 ( .A1(or1200_cpu_or1200_except_n610), .A2(
        n53628), .B(n57093), .C(n54993), .Y(or1200_cpu_or1200_except_n1800) );
  A2O1A1Ixp33_ASAP7_75t_SL U46240 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n622), .C(n54794), .Y(
        or1200_cpu_or1200_except_n1804) );
  A2O1A1Ixp33_ASAP7_75t_SL U46241 ( .A1(n57093), .A2(n53628), .B(
        or1200_cpu_or1200_except_n649), .C(n54992), .Y(
        or1200_cpu_or1200_except_n1813) );
  A2O1A1Ixp33_ASAP7_75t_SL U46242 ( .A1(or1200_cpu_or1200_except_n661), .A2(
        n53628), .B(n57093), .C(n54991), .Y(or1200_cpu_or1200_except_n1817) );
  A2O1A1Ixp33_ASAP7_75t_SL U46243 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n667), .C(n54793), .Y(
        or1200_cpu_or1200_except_n1819) );
  A2O1A1Ixp33_ASAP7_75t_SL U46244 ( .A1(n1042), .A2(n53628), .B(n54988), .C(
        n53628), .Y(n54989) );
  A2O1A1Ixp33_ASAP7_75t_SL U46245 ( .A1(n77275), .A2(n57090), .B(n54989), .C(
        n53628), .Y(n54990) );
  A2O1A1Ixp33_ASAP7_75t_SL U46246 ( .A1(n1044), .A2(n53628), .B(n77276), .C(
        n54990), .Y(or1200_cpu_or1200_except_n593) );
  A2O1A1Ixp33_ASAP7_75t_SL U46247 ( .A1(n72512), .A2(n72511), .B(n72510), .C(
        n53628), .Y(n54978) );
  A2O1A1Ixp33_ASAP7_75t_SL U46248 ( .A1(n53628), .A2(n72509), .B(n72508), .C(
        n53628), .Y(n54979) );
  A2O1A1Ixp33_ASAP7_75t_SL U46249 ( .A1(n72507), .A2(n53628), .B(n72506), .C(
        n54981), .Y(n54982) );
  A2O1A1Ixp33_ASAP7_75t_SL U46250 ( .A1(n54979), .A2(n53628), .B(n54982), .C(
        n53628), .Y(n54983) );
  A2O1A1Ixp33_ASAP7_75t_SL U46251 ( .A1(n59698), .A2(n53628), .B(n54960), .C(
        n53628), .Y(n54961) );
  A2O1A1Ixp33_ASAP7_75t_SL U46252 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .A2(n53628), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), .C(n53628), 
        .Y(n54956) );
  A2O1A1Ixp33_ASAP7_75t_SL U46253 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .A2(n53628), 
        .B(n54957), .C(n53628), .Y(n54958) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46254 ( .A1(n65662), .A2(n65788), .B(n65661), 
        .C(n53628), .D(n54959), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n62) );
  A2O1A1Ixp33_ASAP7_75t_SL U46255 ( .A1(n57217), .A2(n73687), .B(n54950), .C(
        n53628), .Y(n54951) );
  A2O1A1Ixp33_ASAP7_75t_SL U46256 ( .A1(n57217), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[12]), .B(n54945), .C(
        n53628), .Y(n54946) );
  A2O1A1Ixp33_ASAP7_75t_SL U46257 ( .A1(n70162), .A2(n70163), .B(n70164), .C(
        n53628), .Y(n70179) );
  A2O1A1Ixp33_ASAP7_75t_SL U46258 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_1_), .B(n66184), .C(
        n53628), .Y(n54941) );
  A2O1A1Ixp33_ASAP7_75t_SL U46259 ( .A1(n59562), .A2(n53628), .B(n66180), .C(
        n54941), .Y(n54942) );
  A2O1A1Ixp33_ASAP7_75t_SL U46260 ( .A1(n69911), .A2(n53628), .B(n69910), .C(
        n69909), .Y(n54940) );
  A2O1A1Ixp33_ASAP7_75t_SL U46261 ( .A1(n62477), .A2(n53628), .B(n59548), .C(
        n54939), .Y(n77864) );
  A2O1A1Ixp33_ASAP7_75t_SL U46262 ( .A1(n62477), .A2(n53628), .B(n1571), .C(
        n54938), .Y(n77866) );
  A2O1A1Ixp33_ASAP7_75t_SL U46263 ( .A1(n76695), .A2(n53628), .B(n54936), .C(
        n76639), .Y(n54937) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46264 ( .A1(n76548), .A2(n76550), .B(n53628), 
        .C(n76549), .Y(n54935) );
  A2O1A1Ixp33_ASAP7_75t_SL U46265 ( .A1(n57168), .A2(n53628), .B(n865), .C(
        n53628), .Y(n54931) );
  A2O1A1Ixp33_ASAP7_75t_SL U46266 ( .A1(n54931), .A2(n53628), .B(n63969), .C(
        n53628), .Y(n78264) );
  A2O1A1Ixp33_ASAP7_75t_SL U46267 ( .A1(n57160), .A2(n53628), .B(n54930), .C(
        n53628), .Y(n77383) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46268 ( .A1(n62898), .A2(n57178), .B(n53628), 
        .C(n59435), .Y(n54929) );
  A2O1A1Ixp33_ASAP7_75t_SL U46269 ( .A1(n54929), .A2(n53628), .B(n63281), .C(
        n53628), .Y(n63296) );
  A2O1A1Ixp33_ASAP7_75t_SL U46270 ( .A1(n76088), .A2(n53628), .B(n54927), .C(
        n53628), .Y(n76068) );
  A2O1A1Ixp33_ASAP7_75t_SL U46271 ( .A1(n65084), .A2(n54923), .B(n65081), .C(
        n53628), .Y(n54924) );
  A2O1A1Ixp33_ASAP7_75t_SL U46272 ( .A1(n65076), .A2(n53628), .B(n54924), .C(
        n53628), .Y(n64167) );
  A2O1A1Ixp33_ASAP7_75t_SL U46273 ( .A1(n78150), .A2(n53628), .B(n54921), .C(
        n53628), .Y(n78154) );
  A2O1A1Ixp33_ASAP7_75t_SL U46274 ( .A1(n71676), .A2(n53628), .B(n71677), .C(
        n53628), .Y(n54918) );
  A2O1A1Ixp33_ASAP7_75t_SL U46275 ( .A1(n74098), .A2(n53628), .B(n74097), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_), .Y(
        n54916) );
  A2O1A1Ixp33_ASAP7_75t_SL U46276 ( .A1(n74099), .A2(n53628), .B(n54916), .C(
        n53628), .Y(n74233) );
  A2O1A1Ixp33_ASAP7_75t_SL U46277 ( .A1(n57203), .A2(n53628), .B(n72219), .C(
        n53628), .Y(n54911) );
  A2O1A1Ixp33_ASAP7_75t_SL U46278 ( .A1(n57127), .A2(n53628), .B(n72306), .C(
        n53628), .Y(n54912) );
  A2O1A1Ixp33_ASAP7_75t_SL U46279 ( .A1(n72234), .A2(n53628), .B(n57123), .C(
        n53628), .Y(n54913) );
  A2O1A1Ixp33_ASAP7_75t_SL U46280 ( .A1(n54912), .A2(n53628), .B(n54913), .C(
        n53628), .Y(n54914) );
  A2O1A1Ixp33_ASAP7_75t_SL U46281 ( .A1(n57125), .A2(n53628), .B(n72253), .C(
        n54914), .Y(n54915) );
  A2O1A1Ixp33_ASAP7_75t_SL U46282 ( .A1(n54911), .A2(n53628), .B(n54915), .C(
        n53628), .Y(n72453) );
  A2O1A1Ixp33_ASAP7_75t_SL U46283 ( .A1(n57127), .A2(n53628), .B(n71936), .C(
        n53628), .Y(n54910) );
  A2O1A1Ixp33_ASAP7_75t_SL U46284 ( .A1(n54910), .A2(n53628), .B(n71937), .C(
        n53628), .Y(n72422) );
  A2O1A1Ixp33_ASAP7_75t_SL U46285 ( .A1(n71284), .A2(n53628), .B(n71334), .C(
        n53628), .Y(n54903) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46286 ( .A1(n71194), .A2(n71394), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_35_), .C(n53628), 
        .D(n54903), .Y(n54904) );
  A2O1A1Ixp33_ASAP7_75t_SL U46287 ( .A1(n57187), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .B(n54900), 
        .C(n53628), .Y(n54901) );
  A2O1A1Ixp33_ASAP7_75t_SL U46288 ( .A1(n72999), .A2(n53628), .B(n72711), .C(
        n54897), .Y(n73039) );
  A2O1A1Ixp33_ASAP7_75t_SL U46289 ( .A1(n77066), .A2(n53628), .B(n76463), .C(
        n53628), .Y(n54890) );
  A2O1A1Ixp33_ASAP7_75t_SL U46290 ( .A1(or1200_cpu_or1200_mult_mac_n151), .A2(
        n53628), .B(n77057), .C(n53628), .Y(n54891) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46291 ( .A1(n61633), .A2(n57191), .B(n54890), 
        .C(n53628), .D(n54891), .Y(n54892) );
  A2O1A1Ixp33_ASAP7_75t_SL U46292 ( .A1(or1200_cpu_or1200_mult_mac_n297), .A2(
        n53628), .B(n77073), .C(n54892), .Y(n61634) );
  A2O1A1Ixp33_ASAP7_75t_SL U46293 ( .A1(n76764), .A2(n53628), .B(n62256), .C(
        n53628), .Y(n54887) );
  A2O1A1Ixp33_ASAP7_75t_SL U46294 ( .A1(n61433), .A2(n53628), .B(n61183), .C(
        n62433), .Y(n54888) );
  A2O1A1Ixp33_ASAP7_75t_SL U46295 ( .A1(n59559), .A2(n53628), .B(n75714), .C(
        n54888), .Y(n54889) );
  A2O1A1Ixp33_ASAP7_75t_SL U46296 ( .A1(n54887), .A2(n53628), .B(n54889), .C(
        n53628), .Y(n61196) );
  A2O1A1Ixp33_ASAP7_75t_SL U46297 ( .A1(n75053), .A2(n75052), .B(n75065), .C(
        n53628), .Y(n75071) );
  A2O1A1Ixp33_ASAP7_75t_SL U46298 ( .A1(n75557), .A2(n53628), .B(n65146), .C(
        n65145), .Y(n54883) );
  A2O1A1Ixp33_ASAP7_75t_SL U46299 ( .A1(n65147), .A2(n53628), .B(n54883), .C(
        n53628), .Y(n65174) );
  A2O1A1Ixp33_ASAP7_75t_SL U46300 ( .A1(n69090), .A2(n53628), .B(n69089), .C(
        n53628), .Y(n54881) );
  A2O1A1Ixp33_ASAP7_75t_SL U46301 ( .A1(n67264), .A2(n53628), .B(n67560), .C(
        n53628), .Y(n54879) );
  A2O1A1Ixp33_ASAP7_75t_SL U46302 ( .A1(n53628), .A2(n59668), .B(n59639), .C(
        n54544), .Y(n75038) );
  A2O1A1Ixp33_ASAP7_75t_SL U46303 ( .A1(n71413), .A2(n53628), .B(n78384), .C(
        n53628), .Y(n54878) );
  A2O1A1Ixp33_ASAP7_75t_SL U46304 ( .A1(n54878), .A2(n53628), .B(n71380), .C(
        n53628), .Y(n71385) );
  A2O1A1Ixp33_ASAP7_75t_SL U46305 ( .A1(n59561), .A2(n53628), .B(n54877), .C(
        n53628), .Y(n64188) );
  A2O1A1Ixp33_ASAP7_75t_SL U46306 ( .A1(n58735), .A2(n53628), .B(n64352), .C(
        n54876), .Y(n64432) );
  O2A1O1Ixp33_ASAP7_75t_SL U46307 ( .A1(n64347), .A2(n64349), .B(n53628), .C(
        n64348), .Y(n54875) );
  A2O1A1Ixp33_ASAP7_75t_SL U46308 ( .A1(n53628), .A2(n67974), .B(n63066), .C(
        n54714), .Y(n63157) );
  A2O1A1Ixp33_ASAP7_75t_SL U46309 ( .A1(n53224), .A2(n53223), .B(n57177), .C(
        n53628), .Y(n58116) );
  A2O1A1Ixp33_ASAP7_75t_SL U46310 ( .A1(n73431), .A2(n53628), .B(n73449), .C(
        n53628), .Y(n54874) );
  A2O1A1Ixp33_ASAP7_75t_SL U46311 ( .A1(n3309), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[9]), .C(n73817), .Y(
        n54872) );
  A2O1A1Ixp33_ASAP7_75t_SL U46312 ( .A1(n73831), .A2(n73814), .B(n54872), .C(
        n53628), .Y(n54873) );
  A2O1A1Ixp33_ASAP7_75t_SL U46313 ( .A1(n73816), .A2(n53628), .B(n73815), .C(
        n54873), .Y(n3290) );
  A2O1A1Ixp33_ASAP7_75t_SL U46314 ( .A1(n73661), .A2(n53628), .B(n54871), .C(
        n73660), .Y(n3278) );
  A2O1A1Ixp33_ASAP7_75t_SL U46315 ( .A1(n53628), .A2(n69878), .B(n70085), .C(
        n69828), .Y(n54527) );
  A2O1A1Ixp33_ASAP7_75t_SL U46316 ( .A1(n69873), .A2(n69971), .B(n54527), .C(
        n53628), .Y(n54528) );
  A2O1A1Ixp33_ASAP7_75t_SL U46317 ( .A1(n61995), .A2(n61996), .B(n59500), .C(
        n53628), .Y(n54712) );
  A2O1A1Ixp33_ASAP7_75t_SL U46318 ( .A1(n53628), .A2(n3076), .B(n61997), .C(
        n54712), .Y(n52470) );
  A2O1A1Ixp33_ASAP7_75t_SL U46319 ( .A1(n53628), .A2(n59627), .B(n72691), .C(
        n54517), .Y(n2936) );
  A2O1A1Ixp33_ASAP7_75t_SL U46320 ( .A1(n74741), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[27]), .C(n53628), 
        .Y(n54858) );
  A2O1A1Ixp33_ASAP7_75t_SL U46321 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_1_), 
        .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[27]), .C(
        n53628), .Y(n54859) );
  A2O1A1Ixp33_ASAP7_75t_SL U46322 ( .A1(n54858), .A2(n53628), .B(n54859), .C(
        n53628), .Y(n54860) );
  A2O1A1Ixp33_ASAP7_75t_SL U46323 ( .A1(n53628), .A2(n77142), .B(n2687), .C(
        n54697), .Y(or1200_cpu_to_sr[7]) );
  A2O1A1Ixp33_ASAP7_75t_SL U46324 ( .A1(n53628), .A2(n57074), .B(n2680), .C(
        n54693), .Y(n2681) );
  A2O1A1Ixp33_ASAP7_75t_SL U46325 ( .A1(n2587), .A2(n53628), .B(n77567), .C(
        n54855), .Y(n9196) );
  A2O1A1Ixp33_ASAP7_75t_SL U46326 ( .A1(n65401), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_12_), .B(n54689), .C(
        n53628), .Y(n2477) );
  A2O1A1Ixp33_ASAP7_75t_SL U46327 ( .A1(n70385), .A2(n53628), .B(n54851), .C(
        n53628), .Y(n54852) );
  A2O1A1Ixp33_ASAP7_75t_SL U46328 ( .A1(n27448), .A2(n53628), .B(n54852), .C(
        n53628), .Y(n54853) );
  A2O1A1Ixp33_ASAP7_75t_SL U46329 ( .A1(n70545), .A2(n70465), .B(n54842), .C(
        n53628), .Y(n2384) );
  A2O1A1Ixp33_ASAP7_75t_SL U46330 ( .A1(n58553), .A2(n53628), .B(n54835), .C(
        n53628), .Y(n54836) );
  A2O1A1Ixp33_ASAP7_75t_SL U46331 ( .A1(n54836), .A2(n53628), .B(n54839), .C(
        n53628), .Y(n2307) );
  A2O1A1Ixp33_ASAP7_75t_SL U46332 ( .A1(n57144), .A2(n53628), .B(n76654), .C(
        n54834), .Y(n2194) );
  A2O1A1Ixp33_ASAP7_75t_SL U46333 ( .A1(dwb_sel_o[3]), .A2(n53628), .B(n57083), 
        .C(n54832), .Y(n1740) );
  A2O1A1Ixp33_ASAP7_75t_SL U46334 ( .A1(n53628), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[16]), .B(n57190), .C(n54465), .Y(n1687) );
  A2O1A1Ixp33_ASAP7_75t_SL U46335 ( .A1(n77672), .A2(n77885), .B(n54327), .C(
        n53628), .Y(n1652) );
  A2O1A1Ixp33_ASAP7_75t_SL U46336 ( .A1(n57114), .A2(n53628), .B(n1468), .C(
        n54827), .Y(n9298) );
  A2O1A1Ixp33_ASAP7_75t_SL U46337 ( .A1(n1345), .A2(n53628), .B(n77487), .C(
        n53628), .Y(n54814) );
  A2O1A1Ixp33_ASAP7_75t_SL U46338 ( .A1(n4122), .A2(n53628), .B(n54806), .C(
        n53628), .Y(n54807) );
  A2O1A1Ixp33_ASAP7_75t_SL U46339 ( .A1(n74961), .A2(n59701), .B(n54807), .C(
        n53628), .Y(n54808) );
  A2O1A1Ixp33_ASAP7_75t_SL U46340 ( .A1(n803), .A2(n53628), .B(n76523), .C(
        n54808), .Y(n9178) );
  A2O1A1Ixp33_ASAP7_75t_SL U46341 ( .A1(n63525), .A2(n63440), .B(n63435), .C(
        n53628), .Y(n54446) );
  A2O1A1Ixp33_ASAP7_75t_SL U46342 ( .A1(n53628), .A2(n76897), .B(n54447), .C(
        n54448), .Y(n54449) );
  A2O1A1Ixp33_ASAP7_75t_SL U46343 ( .A1(or1200_cpu_or1200_mult_mac_n161), .A2(
        n53628), .B(n76889), .C(n54450), .Y(or1200_cpu_or1200_mult_mac_n1583)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46344 ( .A1(n68845), .A2(n53628), .B(n68848), .C(
        n53628), .Y(n53959) );
  A2O1A1Ixp33_ASAP7_75t_SL U46345 ( .A1(n68842), .A2(n53628), .B(n68844), .C(
        n53628), .Y(n53960) );
  A2O1A1Ixp33_ASAP7_75t_SL U46346 ( .A1(n53628), .A2(n59689), .B(
        or1200_cpu_or1200_except_n398), .C(n54427), .Y(
        or1200_cpu_or1200_except_n399) );
  A2O1A1Ixp33_ASAP7_75t_SL U46347 ( .A1(n57093), .A2(n53628), .B(
        or1200_cpu_or1200_except_n586), .C(n54795), .Y(
        or1200_cpu_or1200_except_n1792) );
  A2O1A1Ixp33_ASAP7_75t_SL U46348 ( .A1(n867), .A2(n53628), .B(n53428), .C(
        n53628), .Y(n54791) );
  A2O1A1Ixp33_ASAP7_75t_SL U46349 ( .A1(n63972), .A2(n57090), .B(n54791), .C(
        n53628), .Y(n54792) );
  A2O1A1Ixp33_ASAP7_75t_SL U46350 ( .A1(n874), .A2(n53628), .B(n77276), .C(
        n54792), .Y(or1200_cpu_or1200_except_n620) );
  A2O1A1Ixp33_ASAP7_75t_SL U46351 ( .A1(n72494), .A2(n72493), .B(n54615), .C(
        n53628), .Y(n54616) );
  A2O1A1Ixp33_ASAP7_75t_SL U46352 ( .A1(n72499), .A2(n53628), .B(n72498), .C(
        n72515), .Y(n54620) );
  A2O1A1Ixp33_ASAP7_75t_SL U46353 ( .A1(n57192), .A2(n53628), .B(n72487), .C(
        n54621), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n63) );
  A2O1A1Ixp33_ASAP7_75t_SL U46354 ( .A1(n70822), .A2(n53628), .B(n70821), .C(
        n70833), .Y(n54608) );
  A2O1A1Ixp33_ASAP7_75t_SL U46355 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_12_), .C(n54609), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n139) );
  A2O1A1Ixp33_ASAP7_75t_SL U46356 ( .A1(n71399), .A2(n53628), .B(n71407), .C(
        n53628), .Y(n54785) );
  A2O1A1Ixp33_ASAP7_75t_SL U46357 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_46_), .C(n54787), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n241) );
  A2O1A1Ixp33_ASAP7_75t_SL U46358 ( .A1(n65663), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .C(n53628), 
        .Y(n54774) );
  A2O1A1Ixp33_ASAP7_75t_SL U46359 ( .A1(n66122), .A2(n53628), .B(n66099), .C(
        n53628), .Y(n54775) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46360 ( .A1(n65570), .A2(n66097), .B(n54774), 
        .C(n53628), .D(n54775), .Y(n54776) );
  A2O1A1Ixp33_ASAP7_75t_SL U46361 ( .A1(n66147), .A2(n53628), .B(n66100), .C(
        n53628), .Y(n54778) );
  A2O1A1Ixp33_ASAP7_75t_SL U46362 ( .A1(n66153), .A2(n53628), .B(n66098), .C(
        n53628), .Y(n54779) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46363 ( .A1(n66094), .A2(n66116), .B(n54778), 
        .C(n53628), .D(n54779), .Y(n54780) );
  A2O1A1Ixp33_ASAP7_75t_SL U46364 ( .A1(n54777), .A2(n53628), .B(n54782), .C(
        n53628), .Y(n54783) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46365 ( .A1(n66167), .A2(n54783), .B(n54784), 
        .C(n53628), .D(n65577), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n4) );
  A2O1A1Ixp33_ASAP7_75t_SL U46366 ( .A1(n3321), .A2(n57217), .B(n54769), .C(
        n53628), .Y(n54770) );
  A2O1A1Ixp33_ASAP7_75t_SL U46367 ( .A1(n78347), .A2(n53628), .B(n70021), .C(
        n53628), .Y(n54761) );
  A2O1A1Ixp33_ASAP7_75t_SL U46368 ( .A1(n69496), .A2(n53628), .B(n78345), .C(
        n53628), .Y(n54762) );
  A2O1A1Ixp33_ASAP7_75t_SL U46369 ( .A1(n78343), .A2(n53628), .B(n69497), .C(
        n53628), .Y(n54763) );
  A2O1A1Ixp33_ASAP7_75t_SL U46370 ( .A1(n54762), .A2(n53628), .B(n54763), .C(
        n53628), .Y(n54764) );
  A2O1A1Ixp33_ASAP7_75t_SL U46371 ( .A1(n69564), .A2(n53628), .B(n78349), .C(
        n54764), .Y(n54765) );
  A2O1A1Ixp33_ASAP7_75t_SL U46372 ( .A1(n54761), .A2(n53628), .B(n54765), .C(
        n53628), .Y(n69881) );
  A2O1A1Ixp33_ASAP7_75t_SL U46373 ( .A1(n74646), .A2(n70543), .B(n54759), .C(
        n53628), .Y(n54760) );
  A2O1A1Ixp33_ASAP7_75t_SL U46374 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .A2(
        n53628), .B(n70488), .C(n54760), .Y(n70411) );
  A2O1A1Ixp33_ASAP7_75t_SL U46375 ( .A1(n62477), .A2(n53628), .B(n59536), .C(
        n54757), .Y(n77888) );
  A2O1A1Ixp33_ASAP7_75t_SL U46376 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_2_), .A2(
        n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_3_), .C(
        n53628), .Y(n54756) );
  A2O1A1Ixp33_ASAP7_75t_SL U46377 ( .A1(n76994), .A2(n53628), .B(n54753), .C(
        n76612), .Y(n54754) );
  A2O1A1Ixp33_ASAP7_75t_SL U46378 ( .A1(n57168), .A2(n53628), .B(n964), .C(
        n53628), .Y(n54751) );
  A2O1A1Ixp33_ASAP7_75t_SL U46379 ( .A1(n54751), .A2(n53628), .B(n65212), .C(
        n53628), .Y(n78205) );
  A2O1A1Ixp33_ASAP7_75t_SL U46380 ( .A1(n63879), .A2(n53628), .B(n54750), .C(
        n53628), .Y(n63500) );
  A2O1A1Ixp33_ASAP7_75t_SL U46381 ( .A1(n63879), .A2(n53628), .B(n54750), .C(
        n53628), .Y(n53459) );
  A2O1A1Ixp33_ASAP7_75t_SL U46382 ( .A1(n63278), .A2(n53628), .B(n54748), .C(
        n53628), .Y(n54749) );
  A2O1A1Ixp33_ASAP7_75t_SL U46383 ( .A1(n54749), .A2(n53628), .B(n63279), .C(
        n53628), .Y(n63297) );
  A2O1A1Ixp33_ASAP7_75t_SL U46384 ( .A1(n76097), .A2(n53628), .B(n76096), .C(
        n54747), .Y(n76108) );
  A2O1A1Ixp33_ASAP7_75t_SL U46385 ( .A1(n53628), .A2(n76033), .B(n76032), .C(
        n54589), .Y(n76036) );
  A2O1A1Ixp33_ASAP7_75t_SL U46386 ( .A1(n75123), .A2(n53628), .B(n54746), .C(
        n53628), .Y(n75118) );
  A2O1A1Ixp33_ASAP7_75t_SL U46387 ( .A1(n57168), .A2(n53628), .B(n991), .C(
        n53628), .Y(n54744) );
  A2O1A1Ixp33_ASAP7_75t_SL U46388 ( .A1(n54744), .A2(n53628), .B(n75161), .C(
        n53628), .Y(n78204) );
  A2O1A1Ixp33_ASAP7_75t_SL U46389 ( .A1(n53628), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_), 
        .B(n57208), .C(n54579), .Y(n54580) );
  A2O1A1Ixp33_ASAP7_75t_SL U46390 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .A2(n53628), .B(n71890), .C(n53628), .Y(n54736) );
  A2O1A1Ixp33_ASAP7_75t_SL U46391 ( .A1(n58422), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_), 
        .C(n53628), .Y(n54737) );
  A2O1A1Ixp33_ASAP7_75t_SL U46392 ( .A1(n57207), .A2(n72212), .B(n54737), .C(
        n53628), .Y(n54738) );
  A2O1A1Ixp33_ASAP7_75t_SL U46393 ( .A1(n57208), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_), 
        .C(n54738), .Y(n54739) );
  A2O1A1Ixp33_ASAP7_75t_SL U46394 ( .A1(n54736), .A2(n53628), .B(n54739), .C(
        n53628), .Y(n72091) );
  A2O1A1Ixp33_ASAP7_75t_SL U46395 ( .A1(n76768), .A2(n62273), .B(n54735), .C(
        n53628), .Y(n61710) );
  A2O1A1Ixp33_ASAP7_75t_SL U46396 ( .A1(n76801), .A2(n53628), .B(n61626), .C(
        n53628), .Y(n54732) );
  A2O1A1Ixp33_ASAP7_75t_SL U46397 ( .A1(n54732), .A2(n53628), .B(n77117), .C(
        n53628), .Y(n62284) );
  A2O1A1Ixp33_ASAP7_75t_SL U46398 ( .A1(n53628), .A2(n63570), .B(n77093), .C(
        n54555), .Y(n60864) );
  A2O1A1Ixp33_ASAP7_75t_SL U46399 ( .A1(or1200_cpu_or1200_mult_mac_n92), .A2(
        n53628), .B(n61826), .C(n54731), .Y(n63563) );
  A2O1A1Ixp33_ASAP7_75t_SL U46400 ( .A1(n78149), .A2(n53628), .B(n54730), .C(
        n53628), .Y(n77016) );
  A2O1A1Ixp33_ASAP7_75t_SL U46401 ( .A1(n71314), .A2(n53628), .B(n71193), .C(
        n54729), .Y(n71223) );
  A2O1A1Ixp33_ASAP7_75t_SL U46402 ( .A1(n59562), .A2(n53628), .B(n65858), .C(
        n54728), .Y(n65600) );
  A2O1A1Ixp33_ASAP7_75t_SL U46403 ( .A1(n57096), .A2(n53628), .B(n75038), .C(
        n53628), .Y(n54725) );
  A2O1A1Ixp33_ASAP7_75t_SL U46404 ( .A1(n75040), .A2(n59635), .B(n54725), .C(
        n53628), .Y(n54726) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46405 ( .A1(n75063), .A2(n75064), .B(n75039), 
        .C(n53628), .D(n54726), .Y(n54727) );
  A2O1A1Ixp33_ASAP7_75t_SL U46406 ( .A1(n75462), .A2(n75469), .B(n54727), .C(
        n53628), .Y(n59280) );
  OAI21xp5_ASAP7_75t_SL U46407 ( .A1(n57107), .A2(n59455), .B(n54724), .Y(
        n67718) );
  A2O1A1Ixp33_ASAP7_75t_SL U46408 ( .A1(n57696), .A2(n53628), .B(n59502), .C(
        n53628), .Y(n54723) );
  A2O1A1Ixp33_ASAP7_75t_SL U46409 ( .A1(n75901), .A2(n59617), .B(n54723), .C(
        n53628), .Y(n65052) );
  A2O1A1Ixp33_ASAP7_75t_SL U46410 ( .A1(n75848), .A2(n66288), .B(n53455), .C(
        n53628), .Y(n54363) );
  A2O1A1Ixp33_ASAP7_75t_SL U46411 ( .A1(n59705), .A2(n73810), .B(n54531), .C(
        n53628), .Y(n54532) );
  A2O1A1Ixp33_ASAP7_75t_SL U46412 ( .A1(n65227), .A2(n53628), .B(n65219), .C(
        n53628), .Y(n54704) );
  A2O1A1Ixp33_ASAP7_75t_SL U46413 ( .A1(n57144), .A2(n53628), .B(n54706), .C(
        n54707), .Y(n2995) );
  A2O1A1Ixp33_ASAP7_75t_SL U46414 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[22]), .A2(
        n53628), .B(n57190), .C(n54702), .Y(n2946) );
  A2O1A1Ixp33_ASAP7_75t_SL U46415 ( .A1(n74885), .A2(n53628), .B(n54700), .C(
        n53628), .Y(n54701) );
  A2O1A1Ixp33_ASAP7_75t_SL U46416 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_20_), .A2(n53628), 
        .B(n74867), .C(n54701), .Y(n52509) );
  A2O1A1Ixp33_ASAP7_75t_SL U46417 ( .A1(n59629), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_15_), .C(n54699), .Y(
        n2845) );
  A2O1A1Ixp33_ASAP7_75t_SL U46418 ( .A1(n59688), .A2(n53628), .B(n2561), .C(
        n54691), .Y(n2562) );
  A2O1A1Ixp33_ASAP7_75t_SL U46419 ( .A1(n65306), .A2(n53628), .B(n54688), .C(
        n53628), .Y(n54689) );
  A2O1A1Ixp33_ASAP7_75t_SL U46420 ( .A1(n62144), .A2(n53628), .B(n60369), .C(
        n53628), .Y(n54679) );
  A2O1A1Ixp33_ASAP7_75t_SL U46421 ( .A1(n54679), .A2(n53628), .B(n54680), .C(
        n53628), .Y(n54681) );
  A2O1A1Ixp33_ASAP7_75t_SL U46422 ( .A1(n62144), .A2(n53628), .B(n60369), .C(
        n60351), .Y(n54682) );
  A2O1A1Ixp33_ASAP7_75t_SL U46423 ( .A1(n57483), .A2(n53628), .B(n77567), .C(
        n54687), .Y(n2470) );
  A2O1A1Ixp33_ASAP7_75t_SL U46424 ( .A1(n70372), .A2(n53628), .B(n54676), .C(
        n53628), .Y(n54677) );
  A2O1A1Ixp33_ASAP7_75t_SL U46425 ( .A1(n70405), .A2(n53628), .B(n70482), .C(
        n53628), .Y(n54672) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46426 ( .A1(n70545), .A2(n54671), .B(n54672), 
        .C(n53628), .D(n54675), .Y(n2419) );
  A2O1A1Ixp33_ASAP7_75t_SL U46427 ( .A1(n77847), .A2(n53628), .B(n77591), .C(
        n53628), .Y(n54665) );
  A2O1A1Ixp33_ASAP7_75t_SL U46428 ( .A1(n77639), .A2(n53628), .B(n77592), .C(
        n53628), .Y(n54666) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46429 ( .A1(n77675), .A2(n77593), .B(n54665), 
        .C(n53628), .D(n54666), .Y(n1712) );
  A2O1A1Ixp33_ASAP7_75t_SL U46430 ( .A1(n57190), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_), .B(n54150), .C(
        n53628), .Y(n78377) );
  A2O1A1Ixp33_ASAP7_75t_SL U46431 ( .A1(n57114), .A2(n53628), .B(n1466), .C(
        n54664), .Y(n9297) );
  A2O1A1Ixp33_ASAP7_75t_SL U46432 ( .A1(n53628), .A2(n74641), .B(n1392), .C(
        n54459), .Y(n9318) );
  A2O1A1Ixp33_ASAP7_75t_SL U46433 ( .A1(n1345), .A2(n53628), .B(n77489), .C(
        n53628), .Y(n54659) );
  A2O1A1Ixp33_ASAP7_75t_SL U46434 ( .A1(n54659), .A2(n53628), .B(n54660), .C(
        n53628), .Y(n54661) );
  A2O1A1Ixp33_ASAP7_75t_SL U46435 ( .A1(n54658), .A2(n53628), .B(n54661), .C(
        n54662), .Y(n9345) );
  A2O1A1Ixp33_ASAP7_75t_SL U46436 ( .A1(n4120), .A2(n53628), .B(n54655), .C(
        n53628), .Y(n54656) );
  A2O1A1Ixp33_ASAP7_75t_SL U46437 ( .A1(n63920), .A2(n59701), .B(n54656), .C(
        n53628), .Y(n54657) );
  A2O1A1Ixp33_ASAP7_75t_SL U46438 ( .A1(n799), .A2(n53628), .B(n76523), .C(
        n54657), .Y(n9177) );
  A2O1A1Ixp33_ASAP7_75t_SL U46439 ( .A1(n75760), .A2(n53628), .B(n59689), .C(
        n57077), .Y(n54653) );
  A2O1A1Ixp33_ASAP7_75t_SL U46440 ( .A1(n63283), .A2(n53628), .B(n54645), .C(
        n59674), .Y(n54646) );
  A2O1A1Ixp33_ASAP7_75t_SL U46441 ( .A1(n63283), .A2(n54645), .B(n54646), .C(
        n53628), .Y(n54647) );
  A2O1A1Ixp33_ASAP7_75t_SL U46442 ( .A1(n63286), .A2(n53628), .B(n54645), .C(
        n53628), .Y(n54648) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46443 ( .A1(n63286), .A2(n54645), .B(n76897), 
        .C(n53628), .D(n54648), .Y(n54649) );
  A2O1A1Ixp33_ASAP7_75t_SL U46444 ( .A1(n76688), .A2(n53628), .B(n65182), .C(
        n53628), .Y(n54650) );
  O2A1O1Ixp33_ASAP7_75t_SL U46445 ( .A1(n54647), .A2(n54649), .B(n53628), .C(
        n54650), .Y(n54651) );
  A2O1A1Ixp33_ASAP7_75t_SL U46446 ( .A1(n68832), .A2(n57079), .B(n54637), .C(
        n53628), .Y(n54638) );
  A2O1A1Ixp33_ASAP7_75t_SL U46447 ( .A1(n76906), .A2(n53628), .B(n68831), .C(
        n53628), .Y(n54640) );
  A2O1A1Ixp33_ASAP7_75t_SL U46448 ( .A1(n68832), .A2(n53628), .B(n59671), .C(
        n54637), .Y(n54641) );
  A2O1A1Ixp33_ASAP7_75t_SL U46449 ( .A1(n54640), .A2(n53628), .B(n54641), .C(
        n53628), .Y(n54642) );
  A2O1A1Ixp33_ASAP7_75t_SL U46450 ( .A1(n54638), .A2(n54639), .B(n54642), .C(
        n53628), .Y(n54643) );
  A2O1A1Ixp33_ASAP7_75t_SL U46451 ( .A1(n59673), .A2(n77922), .B(n54643), .C(
        n53628), .Y(n54644) );
  A2O1A1Ixp33_ASAP7_75t_SL U46452 ( .A1(or1200_cpu_or1200_mult_mac_n205), .A2(
        n53628), .B(n76909), .C(n54644), .Y(or1200_cpu_or1200_mult_mac_n1624)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46453 ( .A1(n59672), .A2(n69125), .B(n54629), .C(
        n53628), .Y(n54631) );
  A2O1A1Ixp33_ASAP7_75t_SL U46454 ( .A1(or1200_cpu_or1200_except_n595), .A2(
        n53628), .B(n57093), .C(n54624), .Y(or1200_cpu_or1200_except_n1795) );
  A2O1A1Ixp33_ASAP7_75t_SL U46455 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n637), .C(n54276), .Y(
        or1200_cpu_or1200_except_n1809) );
  A2O1A1Ixp33_ASAP7_75t_SL U46456 ( .A1(or1200_cpu_or1200_except_n670), .A2(
        n53628), .B(n57072), .C(n54623), .Y(or1200_cpu_or1200_except_n1820) );
  A2O1A1Ixp33_ASAP7_75t_SL U46457 ( .A1(n74099), .A2(n53628), .B(n74100), .C(
        n74236), .Y(n54622) );
  A2O1A1Ixp33_ASAP7_75t_SL U46458 ( .A1(n54619), .A2(n53628), .B(n54620), .C(
        n53628), .Y(n54621) );
  A2O1A1Ixp33_ASAP7_75t_SL U46459 ( .A1(n71519), .A2(n53628), .B(n54606), .C(
        n53628), .Y(n71517) );
  A2O1A1Ixp33_ASAP7_75t_SL U46460 ( .A1(n74227), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_24_), 
        .C(n53628), .Y(n54603) );
  A2O1A1Ixp33_ASAP7_75t_SL U46461 ( .A1(n54603), .A2(n53628), .B(n74451), .C(
        n53628), .Y(n74453) );
  A2O1A1Ixp33_ASAP7_75t_SL U46462 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[4]), 
        .A2(n53628), .B(n54602), .C(n53628), .Y(n74255) );
  O2A1O1Ixp33_ASAP7_75t_SL U46463 ( .A1(n75802), .A2(n75801), .B(n53628), .C(
        n54601), .Y(n73956) );
  A2O1A1Ixp33_ASAP7_75t_SL U46464 ( .A1(n62477), .A2(n53628), .B(n1868), .C(
        n54600), .Y(n77862) );
  A2O1A1Ixp33_ASAP7_75t_SL U46465 ( .A1(n62477), .A2(n53628), .B(n59549), .C(
        n54599), .Y(n77859) );
  O2A1O1Ixp33_ASAP7_75t_SL U46466 ( .A1(n76205), .A2(n76995), .B(n53628), .C(
        n54252), .Y(n54253) );
  A2O1A1Ixp33_ASAP7_75t_SL U46467 ( .A1(n75424), .A2(n53628), .B(n54595), .C(
        n53628), .Y(n54596) );
  A2O1A1Ixp33_ASAP7_75t_SL U46468 ( .A1(n57160), .A2(n53628), .B(n54593), .C(
        n53628), .Y(n65212) );
  A2O1A1Ixp33_ASAP7_75t_SL U46469 ( .A1(n57160), .A2(n53628), .B(n54592), .C(
        n53628), .Y(n75631) );
  A2O1A1Ixp33_ASAP7_75t_SL U46470 ( .A1(n62906), .A2(n53628), .B(n62907), .C(
        n53628), .Y(n54590) );
  A2O1A1Ixp33_ASAP7_75t_SL U46471 ( .A1(n62908), .A2(n53628), .B(n54590), .C(
        n54591), .Y(n63313) );
  A2O1A1Ixp33_ASAP7_75t_SL U46472 ( .A1(or1200_cpu_or1200_mult_mac_div_cntr_2_), .A2(n53628), .B(or1200_cpu_or1200_mult_mac_div_cntr_3_), .C(n53628), .Y(
        n54588) );
  A2O1A1Ixp33_ASAP7_75t_SL U46473 ( .A1(n69326), .A2(n53628), .B(n54584), .C(
        n53628), .Y(n69310) );
  A2O1A1Ixp33_ASAP7_75t_SL U46474 ( .A1(n77209), .A2(n53628), .B(n54583), .C(
        n53628), .Y(n77442) );
  A2O1A1Ixp33_ASAP7_75t_SL U46475 ( .A1(n72309), .A2(n57207), .B(n54580), .C(
        n53628), .Y(n54581) );
  A2O1A1Ixp33_ASAP7_75t_SL U46476 ( .A1(n57208), .A2(n53628), .B(n72141), .C(
        n53628), .Y(n54573) );
  A2O1A1Ixp33_ASAP7_75t_SL U46477 ( .A1(n54573), .A2(n53628), .B(n54576), .C(
        n53628), .Y(n54577) );
  A2O1A1Ixp33_ASAP7_75t_SL U46478 ( .A1(n71890), .A2(n53628), .B(n71835), .C(
        n53628), .Y(n54569) );
  A2O1A1Ixp33_ASAP7_75t_SL U46479 ( .A1(n72250), .A2(n53628), .B(n58422), .C(
        n53628), .Y(n54570) );
  A2O1A1Ixp33_ASAP7_75t_SL U46480 ( .A1(n57207), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_1_), 
        .B(n54570), .C(n53628), .Y(n54571) );
  A2O1A1Ixp33_ASAP7_75t_SL U46481 ( .A1(n57208), .A2(n53628), .B(n72365), .C(
        n54571), .Y(n54572) );
  A2O1A1Ixp33_ASAP7_75t_SL U46482 ( .A1(n54569), .A2(n53628), .B(n54572), .C(
        n53628), .Y(n72354) );
  A2O1A1Ixp33_ASAP7_75t_SL U46483 ( .A1(n71194), .A2(n53628), .B(n71335), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_35_), .Y(n54566) );
  A2O1A1Ixp33_ASAP7_75t_SL U46484 ( .A1(n71334), .A2(n71315), .B(n54566), .C(
        n53628), .Y(n54567) );
  A2O1A1Ixp33_ASAP7_75t_SL U46485 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]), .A2(n57194), 
        .B(n54564), .C(n53628), .Y(n65971) );
  A2O1A1Ixp33_ASAP7_75t_SL U46486 ( .A1(n59631), .A2(n53628), .B(n73238), .C(
        n53628), .Y(n54560) );
  A2O1A1Ixp33_ASAP7_75t_SL U46487 ( .A1(n53628), .A2(n2345), .B(n70488), .C(
        n54048), .Y(n70398) );
  A2O1A1Ixp33_ASAP7_75t_SL U46488 ( .A1(or1200_cpu_or1200_mult_mac_n96), .A2(
        n53628), .B(n61826), .C(n54551), .Y(n62514) );
  A2O1A1Ixp33_ASAP7_75t_SL U46489 ( .A1(n53431), .A2(n53628), .B(n54550), .C(
        n53628), .Y(n65130) );
  A2O1A1Ixp33_ASAP7_75t_SL U46490 ( .A1(n71950), .A2(n53628), .B(n71460), .C(
        n53628), .Y(n54549) );
  A2O1A1Ixp33_ASAP7_75t_SL U46491 ( .A1(n59544), .A2(n53628), .B(n57120), .C(
        n54546), .Y(n61620) );
  A2O1A1Ixp33_ASAP7_75t_SL U46492 ( .A1(n64971), .A2(n53628), .B(n57037), .C(
        n53628), .Y(n54540) );
  A2O1A1Ixp33_ASAP7_75t_SL U46493 ( .A1(n75032), .A2(n53628), .B(n66466), .C(
        n53628), .Y(n54536) );
  A2O1A1Ixp33_ASAP7_75t_SL U46494 ( .A1(n54536), .A2(n53628), .B(n54538), .C(
        n53628), .Y(n66475) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46495 ( .A1(n73424), .A2(n73425), .B(n53628), 
        .C(n73416), .Y(n54534) );
  A2O1A1Ixp33_ASAP7_75t_SL U46496 ( .A1(n73818), .A2(n53628), .B(n73830), .C(
        n53628), .Y(n54531) );
  A2O1A1Ixp33_ASAP7_75t_SL U46497 ( .A1(n54518), .A2(n53628), .B(n54519), .C(
        n53628), .Y(n54520) );
  A2O1A1Ixp33_ASAP7_75t_SL U46498 ( .A1(n54521), .A2(n53628), .B(n54522), .C(
        n53628), .Y(n54523) );
  A2O1A1Ixp33_ASAP7_75t_SL U46499 ( .A1(n53628), .A2(n59689), .B(n2991), .C(
        n54356), .Y(n2992) );
  A2O1A1Ixp33_ASAP7_75t_SL U46500 ( .A1(n74899), .A2(n54515), .B(n74885), .C(
        n53628), .Y(n54516) );
  A2O1A1Ixp33_ASAP7_75t_SL U46501 ( .A1(n62000), .A2(n60590), .B(n60726), .C(
        n53628), .Y(n54512) );
  A2O1A1Ixp33_ASAP7_75t_SL U46502 ( .A1(n53628), .A2(n57074), .B(n2673), .C(
        n54344), .Y(n2674) );
  A2O1A1Ixp33_ASAP7_75t_SL U46503 ( .A1(n70296), .A2(n54185), .B(n70477), .C(
        n53628), .Y(n54187) );
  A2O1A1Ixp33_ASAP7_75t_SL U46504 ( .A1(n70553), .A2(n53628), .B(n74685), .C(
        n53628), .Y(n54493) );
  A2O1A1Ixp33_ASAP7_75t_SL U46505 ( .A1(n54493), .A2(n53628), .B(n54495), .C(
        n53628), .Y(n54496) );
  A2O1A1Ixp33_ASAP7_75t_SL U46506 ( .A1(n74674), .A2(n53628), .B(n70488), .C(
        n53628), .Y(n54497) );
  A2O1A1Ixp33_ASAP7_75t_SL U46507 ( .A1(n54497), .A2(n53628), .B(n54500), .C(
        n53628), .Y(n54501) );
  A2O1A1Ixp33_ASAP7_75t_SL U46508 ( .A1(n70487), .A2(n53628), .B(n54501), .C(
        n54502), .Y(n54503) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46509 ( .A1(n70490), .A2(n70491), .B(n54496), 
        .C(n53628), .D(n54503), .Y(n54504) );
  A2O1A1Ixp33_ASAP7_75t_SL U46510 ( .A1(n69785), .A2(n53628), .B(n69784), .C(
        n69783), .Y(n54482) );
  A2O1A1Ixp33_ASAP7_75t_SL U46511 ( .A1(n69782), .A2(n53628), .B(n54481), .C(
        n53628), .Y(n54484) );
  A2O1A1Ixp33_ASAP7_75t_SL U46512 ( .A1(n70513), .A2(n53628), .B(n70422), .C(
        n53628), .Y(n54487) );
  A2O1A1Ixp33_ASAP7_75t_SL U46513 ( .A1(n57081), .A2(n53628), .B(n69787), .C(
        n53628), .Y(n54488) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46514 ( .A1(n59621), .A2(n54486), .B(n54487), 
        .C(n53628), .D(n54488), .Y(n2299) );
  A2O1A1Ixp33_ASAP7_75t_SL U46515 ( .A1(n65304), .A2(n53628), .B(n54478), .C(
        n53628), .Y(n54479) );
  A2O1A1Ixp33_ASAP7_75t_SL U46516 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_14_), .A2(n65401), .B(
        n54479), .C(n53628), .Y(n1998) );
  A2O1A1Ixp33_ASAP7_75t_SL U46517 ( .A1(n77847), .A2(n53628), .B(n77594), .C(
        n53628), .Y(n54466) );
  A2O1A1Ixp33_ASAP7_75t_SL U46518 ( .A1(n77639), .A2(n53628), .B(n77595), .C(
        n53628), .Y(n54467) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46519 ( .A1(n77675), .A2(n77596), .B(n54466), 
        .C(n53628), .D(n54467), .Y(n1711) );
  A2O1A1Ixp33_ASAP7_75t_SL U46520 ( .A1(n53628), .A2(n57202), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[23]), .C(n54325), 
        .Y(n1613) );
  A2O1A1Ixp33_ASAP7_75t_SL U46521 ( .A1(n74934), .A2(n53628), .B(n59558), .C(
        n53628), .Y(n54461) );
  A2O1A1Ixp33_ASAP7_75t_SL U46522 ( .A1(n74916), .A2(n53628), .B(n1533), .C(
        n53628), .Y(n54462) );
  A2O1A1Ixp33_ASAP7_75t_SL U46523 ( .A1(n54461), .A2(n53628), .B(n54462), .C(
        n53628), .Y(n54463) );
  A2O1A1Ixp33_ASAP7_75t_SL U46524 ( .A1(n57114), .A2(n53628), .B(n1464), .C(
        n54460), .Y(n9296) );
  A2O1A1Ixp33_ASAP7_75t_SL U46525 ( .A1(n53628), .A2(n77999), .B(n77998), .C(
        n54313), .Y(n9380) );
  A2O1A1Ixp33_ASAP7_75t_SL U46526 ( .A1(n4118), .A2(n53628), .B(n54456), .C(
        n53628), .Y(n54457) );
  A2O1A1Ixp33_ASAP7_75t_SL U46527 ( .A1(n64096), .A2(n59701), .B(n54457), .C(
        n53628), .Y(n54458) );
  A2O1A1Ixp33_ASAP7_75t_SL U46528 ( .A1(n795), .A2(n53628), .B(n76523), .C(
        n54458), .Y(n9176) );
  A2O1A1Ixp33_ASAP7_75t_SL U46529 ( .A1(n63525), .A2(n63440), .B(n63430), .C(
        n53628), .Y(n54439) );
  A2O1A1Ixp33_ASAP7_75t_SL U46530 ( .A1(n54439), .A2(n53628), .B(n76906), .C(
        n53628), .Y(n54440) );
  A2O1A1Ixp33_ASAP7_75t_SL U46531 ( .A1(or1200_cpu_or1200_mult_mac_n307), .A2(
        n53628), .B(n54441), .C(n53628), .Y(n54442) );
  A2O1A1Ixp33_ASAP7_75t_SL U46532 ( .A1(n54442), .A2(n53628), .B(n54444), .C(
        n53628), .Y(n54445) );
  A2O1A1Ixp33_ASAP7_75t_SL U46533 ( .A1(n54445), .A2(n53628), .B(n54446), .C(
        n53628), .Y(n54447) );
  A2O1A1Ixp33_ASAP7_75t_SL U46534 ( .A1(n75291), .A2(n53628), .B(n75292), .C(
        n53628), .Y(n54430) );
  A2O1A1Ixp33_ASAP7_75t_SL U46535 ( .A1(n76906), .A2(n53628), .B(n75295), .C(
        n53628), .Y(n54434) );
  A2O1A1Ixp33_ASAP7_75t_SL U46536 ( .A1(n1011), .A2(n53628), .B(n54988), .C(
        n53628), .Y(n54425) );
  A2O1A1Ixp33_ASAP7_75t_SL U46537 ( .A1(n75640), .A2(n57090), .B(n54425), .C(
        n53628), .Y(n54426) );
  A2O1A1Ixp33_ASAP7_75t_SL U46538 ( .A1(n1018), .A2(n53628), .B(n77276), .C(
        n54426), .Y(or1200_cpu_or1200_except_n668) );
  A2O1A1Ixp33_ASAP7_75t_SL U46539 ( .A1(n57192), .A2(n53628), .B(n72334), .C(
        n53628), .Y(n54415) );
  A2O1A1Ixp33_ASAP7_75t_SL U46540 ( .A1(n72499), .A2(n53628), .B(n72335), .C(
        n53628), .Y(n54416) );
  A2O1A1Ixp33_ASAP7_75t_SL U46541 ( .A1(n72544), .A2(n53628), .B(n72336), .C(
        n53628), .Y(n54417) );
  A2O1A1Ixp33_ASAP7_75t_SL U46542 ( .A1(n72507), .A2(n53628), .B(n72466), .C(
        n54418), .Y(n54419) );
  A2O1A1Ixp33_ASAP7_75t_SL U46543 ( .A1(n72464), .A2(n72492), .B(n54419), .C(
        n53628), .Y(n54420) );
  A2O1A1Ixp33_ASAP7_75t_SL U46544 ( .A1(n54417), .A2(n53628), .B(n54422), .C(
        n53628), .Y(n54423) );
  O2A1O1Ixp33_ASAP7_75t_SL U46545 ( .A1(n54415), .A2(n54416), .B(n53628), .C(
        n54423), .Y(n54424) );
  A2O1A1Ixp33_ASAP7_75t_SL U46546 ( .A1(n71731), .A2(n53628), .B(n71687), .C(
        n71690), .Y(n54413) );
  A2O1A1Ixp33_ASAP7_75t_SL U46547 ( .A1(n73558), .A2(n53628), .B(n54399), .C(
        n53628), .Y(n73656) );
  A2O1A1Ixp33_ASAP7_75t_SL U46548 ( .A1(n62477), .A2(n53628), .B(n59711), .C(
        n54397), .Y(n77922) );
  A2O1A1Ixp33_ASAP7_75t_SL U46549 ( .A1(n74137), .A2(n53628), .B(n54392), .C(
        n74140), .Y(n54393) );
  A2O1A1Ixp33_ASAP7_75t_SL U46550 ( .A1(n74137), .A2(n54392), .B(n54393), .C(
        n53628), .Y(n54394) );
  A2O1A1Ixp33_ASAP7_75t_SL U46551 ( .A1(n74139), .A2(n53628), .B(n54394), .C(
        n53628), .Y(n74180) );
  A2O1A1Ixp33_ASAP7_75t_SL U46552 ( .A1(n73887), .A2(n53628), .B(n54391), .C(
        n53628), .Y(n74256) );
  A2O1A1Ixp33_ASAP7_75t_SL U46553 ( .A1(n53628), .A2(n76861), .B(n54251), .C(
        n53628), .Y(n54252) );
  A2O1A1Ixp33_ASAP7_75t_SL U46554 ( .A1(n54254), .A2(n53628), .B(n54255), .C(
        n54256), .Y(n77976) );
  A2O1A1Ixp33_ASAP7_75t_SL U46555 ( .A1(n57168), .A2(n53628), .B(n973), .C(
        n53628), .Y(n54390) );
  A2O1A1Ixp33_ASAP7_75t_SL U46556 ( .A1(n54390), .A2(n53628), .B(n65193), .C(
        n53628), .Y(n78206) );
  A2O1A1Ixp33_ASAP7_75t_SL U46557 ( .A1(n77723), .A2(n53628), .B(n78003), .C(
        n54389), .Y(n4265) );
  A2O1A1Ixp33_ASAP7_75t_SL U46558 ( .A1(n57208), .A2(n53628), .B(n72234), .C(
        n53628), .Y(n54383) );
  A2O1A1Ixp33_ASAP7_75t_SL U46559 ( .A1(n54383), .A2(n53628), .B(n54386), .C(
        n53628), .Y(n54387) );
  A2O1A1Ixp33_ASAP7_75t_SL U46560 ( .A1(n57187), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[34]), .B(n54380), 
        .C(n53628), .Y(n54381) );
  A2O1A1Ixp33_ASAP7_75t_SL U46561 ( .A1(n53628), .A2(n53872), .B(n53873), .C(
        n53628), .Y(n53874) );
  A2O1A1Ixp33_ASAP7_75t_SL U46562 ( .A1(dbg_stall_i), .A2(n53628), .B(n54374), 
        .C(n53628), .Y(n60290) );
  A2O1A1Ixp33_ASAP7_75t_SL U46563 ( .A1(n58818), .A2(n53628), .B(n53452), .C(
        n53628), .Y(n63879) );
  A2O1A1Ixp33_ASAP7_75t_SL U46564 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_), 
        .C(n53628), .Y(n54373) );
  A2O1A1Ixp33_ASAP7_75t_SL U46565 ( .A1(n71018), .A2(n53628), .B(n71335), .C(
        n53628), .Y(n54370) );
  A2O1A1Ixp33_ASAP7_75t_SL U46566 ( .A1(n71362), .A2(n53628), .B(n71019), .C(
        n53628), .Y(n54371) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46567 ( .A1(n71175), .A2(n71263), .B(n54370), 
        .C(n53628), .D(n54371), .Y(n54372) );
  A2O1A1Ixp33_ASAP7_75t_SL U46568 ( .A1(n71146), .A2(n53628), .B(n71284), .C(
        n54372), .Y(n71020) );
  A2O1A1Ixp33_ASAP7_75t_SL U46569 ( .A1(n59562), .A2(n53628), .B(n65613), .C(
        n54369), .Y(n65587) );
  A2O1A1Ixp33_ASAP7_75t_SL U46570 ( .A1(n57190), .A2(n53628), .B(n78345), .C(
        n54368), .Y(n72916) );
  A2O1A1Ixp33_ASAP7_75t_SL U46571 ( .A1(n75467), .A2(n53628), .B(n53275), .C(
        n53628), .Y(n54366) );
  A2O1A1Ixp33_ASAP7_75t_SL U46572 ( .A1(n59616), .A2(n53628), .B(n58431), .C(
        n54365), .Y(n64538) );
  A2O1A1Ixp33_ASAP7_75t_SL U46573 ( .A1(n75848), .A2(n53455), .B(n54363), .C(
        n53628), .Y(n54364) );
  A2O1A1Ixp33_ASAP7_75t_SL U46574 ( .A1(n61979), .A2(n53628), .B(n54364), .C(
        n53628), .Y(n61983) );
  A2O1A1Ixp33_ASAP7_75t_SL U46575 ( .A1(n66578), .A2(n66579), .B(n68616), .C(
        n53628), .Y(n57965) );
  A2O1A1Ixp33_ASAP7_75t_SL U46576 ( .A1(n59142), .A2(n53628), .B(n66482), .C(
        n53628), .Y(n53630) );
  A2O1A1Ixp33_ASAP7_75t_SL U46577 ( .A1(n73415), .A2(n73414), .B(n73438), .C(
        n53628), .Y(n78216) );
  A2O1A1Ixp33_ASAP7_75t_SL U46578 ( .A1(n3309), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[12]), .C(n73817), .Y(
        n54019) );
  A2O1A1Ixp33_ASAP7_75t_SL U46579 ( .A1(n73808), .A2(n73814), .B(n54019), .C(
        n53628), .Y(n54020) );
  A2O1A1Ixp33_ASAP7_75t_SL U46580 ( .A1(n53628), .A2(n73816), .B(n73809), .C(
        n54020), .Y(n3293) );
  A2O1A1Ixp33_ASAP7_75t_SL U46581 ( .A1(n53628), .A2(n69902), .B(n70067), .C(
        n54202), .Y(n3211) );
  A2O1A1Ixp33_ASAP7_75t_SL U46582 ( .A1(n75157), .A2(n53628), .B(n57144), .C(
        n75156), .Y(n54355) );
  A2O1A1Ixp33_ASAP7_75t_SL U46583 ( .A1(n74726), .A2(n53628), .B(n74725), .C(
        n54352), .Y(n54353) );
  A2O1A1Ixp33_ASAP7_75t_SL U46584 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[22]), .A2(
        n74464), .B(n54353), .C(n53628), .Y(n2952) );
  A2O1A1Ixp33_ASAP7_75t_SL U46585 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_0_), .A2(n53628), 
        .B(n74200), .C(n53628), .Y(n54347) );
  A2O1A1Ixp33_ASAP7_75t_SL U46586 ( .A1(n74202), .A2(n53628), .B(n74201), .C(
        n53628), .Y(n54348) );
  A2O1A1Ixp33_ASAP7_75t_SL U46587 ( .A1(n54347), .A2(n53628), .B(n54348), .C(
        n53628), .Y(n54349) );
  A2O1A1Ixp33_ASAP7_75t_SL U46588 ( .A1(n74212), .A2(n53628), .B(n74211), .C(
        n74210), .Y(n54350) );
  A2O1A1Ixp33_ASAP7_75t_SL U46589 ( .A1(n54349), .A2(n53628), .B(n54350), .C(
        n53628), .Y(n78198) );
  A2O1A1Ixp33_ASAP7_75t_SL U46590 ( .A1(n59629), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_12_), .C(n54346), .Y(
        n2832) );
  A2O1A1Ixp33_ASAP7_75t_SL U46591 ( .A1(n53250), .A2(n53628), .B(n54339), .C(
        n53628), .Y(n54340) );
  A2O1A1Ixp33_ASAP7_75t_SL U46592 ( .A1(n62020), .A2(n77566), .B(n54340), .C(
        n53628), .Y(n54341) );
  A2O1A1Ixp33_ASAP7_75t_SL U46593 ( .A1(n53628), .A2(n70303), .B(n70467), .C(
        n53628), .Y(n54185) );
  A2O1A1Ixp33_ASAP7_75t_SL U46594 ( .A1(n62047), .A2(n53628), .B(n62053), .C(
        n53628), .Y(n54337) );
  A2O1A1Ixp33_ASAP7_75t_SL U46595 ( .A1(n53628), .A2(n59629), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_22_), .C(n54012), .Y(
        n2002) );
  A2O1A1Ixp33_ASAP7_75t_SL U46596 ( .A1(n59689), .A2(n53628), .B(n1973), .C(
        n54336), .Y(n1974) );
  A2O1A1Ixp33_ASAP7_75t_SL U46597 ( .A1(n77986), .A2(n77212), .B(n54334), .C(
        n53628), .Y(n54335) );
  A2O1A1Ixp33_ASAP7_75t_SL U46598 ( .A1(n77142), .A2(n53628), .B(n1943), .C(
        n54335), .Y(or1200_cpu_to_sr[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U46599 ( .A1(n53628), .A2(n57144), .B(n77891), .C(
        n53788), .Y(n1693) );
  A2O1A1Ixp33_ASAP7_75t_SL U46600 ( .A1(n77651), .A2(n53628), .B(n54326), .C(
        n53628), .Y(n54327) );
  A2O1A1Ixp33_ASAP7_75t_SL U46601 ( .A1(n74741), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[23]), .C(n53628), 
        .Y(n54323) );
  A2O1A1Ixp33_ASAP7_75t_SL U46602 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_1_), 
        .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[23]), .C(
        n53628), .Y(n54324) );
  A2O1A1Ixp33_ASAP7_75t_SL U46603 ( .A1(n54323), .A2(n53628), .B(n54324), .C(
        n53628), .Y(n54325) );
  A2O1A1Ixp33_ASAP7_75t_SL U46604 ( .A1(n57190), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_), .B(n54149), .C(
        n53628), .Y(n78359) );
  A2O1A1Ixp33_ASAP7_75t_SL U46605 ( .A1(n78363), .A2(n53628), .B(n57190), .C(
        n53628), .Y(n54321) );
  A2O1A1Ixp33_ASAP7_75t_SL U46606 ( .A1(n78362), .A2(n53628), .B(n59629), .C(
        n53628), .Y(n54322) );
  A2O1A1Ixp33_ASAP7_75t_SL U46607 ( .A1(n54321), .A2(n53628), .B(n54322), .C(
        n53628), .Y(n78223) );
  A2O1A1Ixp33_ASAP7_75t_SL U46608 ( .A1(n57114), .A2(n53628), .B(n1462), .C(
        n54320), .Y(n9295) );
  A2O1A1Ixp33_ASAP7_75t_SL U46609 ( .A1(n77997), .A2(n53628), .B(n1185), .C(
        n53628), .Y(n54312) );
  A2O1A1Ixp33_ASAP7_75t_SL U46610 ( .A1(n4116), .A2(n53628), .B(n54309), .C(
        n53628), .Y(n54310) );
  A2O1A1Ixp33_ASAP7_75t_SL U46611 ( .A1(n64258), .A2(n59701), .B(n54310), .C(
        n53628), .Y(n54311) );
  A2O1A1Ixp33_ASAP7_75t_SL U46612 ( .A1(n791), .A2(n53628), .B(n76523), .C(
        n54311), .Y(n9175) );
  O2A1O1Ixp33_ASAP7_75t_SL U46613 ( .A1(n53992), .A2(n76004), .B(n53628), .C(
        or1200_cpu_or1200_mult_mac_n60), .Y(n53993) );
  A2O1A1Ixp33_ASAP7_75t_SL U46614 ( .A1(n53628), .A2(
        or1200_cpu_or1200_mult_mac_n153), .B(n76889), .C(n54142), .Y(
        or1200_cpu_or1200_mult_mac_n1587) );
  A2O1A1Ixp33_ASAP7_75t_SL U46615 ( .A1(n69000), .A2(n54289), .B(n68995), .C(
        n53628), .Y(n54290) );
  A2O1A1Ixp33_ASAP7_75t_SL U46616 ( .A1(n68996), .A2(n53628), .B(n68997), .C(
        n53628), .Y(n54293) );
  A2O1A1Ixp33_ASAP7_75t_SL U46617 ( .A1(n68971), .A2(n53628), .B(n68988), .C(
        n53628), .Y(n54294) );
  A2O1A1Ixp33_ASAP7_75t_SL U46618 ( .A1(n76906), .A2(n53628), .B(n54294), .C(
        n53628), .Y(n54295) );
  A2O1A1Ixp33_ASAP7_75t_SL U46619 ( .A1(n68996), .A2(n53628), .B(n68997), .C(
        n53628), .Y(n54301) );
  A2O1A1Ixp33_ASAP7_75t_SL U46620 ( .A1(n69257), .A2(
        or1200_cpu_or1200_mult_mac_n247), .B(n69258), .C(n53628), .Y(n54280)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46621 ( .A1(n69260), .A2(n53628), .B(n54280), .C(
        n53628), .Y(n54281) );
  A2O1A1Ixp33_ASAP7_75t_SL U46622 ( .A1(n76906), .A2(n53628), .B(n69254), .C(
        n54283), .Y(n54284) );
  A2O1A1Ixp33_ASAP7_75t_SL U46623 ( .A1(n69254), .A2(n57080), .B(n54283), .C(
        n53628), .Y(n54285) );
  A2O1A1Ixp33_ASAP7_75t_SL U46624 ( .A1(n54281), .A2(n53628), .B(n59671), .C(
        n54285), .Y(n54286) );
  A2O1A1Ixp33_ASAP7_75t_SL U46625 ( .A1(n53628), .A2(
        or1200_cpu_or1200_except_n583), .B(n57093), .C(n54130), .Y(
        or1200_cpu_or1200_except_n1791) );
  A2O1A1Ixp33_ASAP7_75t_SL U46626 ( .A1(or1200_cpu_or1200_except_n604), .A2(
        n53628), .B(n57072), .C(n54277), .Y(or1200_cpu_or1200_except_n1798) );
  A2O1A1Ixp33_ASAP7_75t_SL U46627 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n613), .C(n54128), .Y(
        or1200_cpu_or1200_except_n1801) );
  A2O1A1Ixp33_ASAP7_75t_SL U46628 ( .A1(n72477), .A2(n53628), .B(n72478), .C(
        n53628), .Y(n54268) );
  A2O1A1Ixp33_ASAP7_75t_SL U46629 ( .A1(n72510), .A2(n53628), .B(n54268), .C(
        n53628), .Y(n54269) );
  A2O1A1Ixp33_ASAP7_75t_SL U46630 ( .A1(n72479), .A2(n53628), .B(n72508), .C(
        n72500), .Y(n54270) );
  A2O1A1Ixp33_ASAP7_75t_SL U46631 ( .A1(n72483), .A2(n72494), .B(n54270), .C(
        n53628), .Y(n54271) );
  A2O1A1Ixp33_ASAP7_75t_SL U46632 ( .A1(n72503), .A2(n53628), .B(n72481), .C(
        n54271), .Y(n54272) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46633 ( .A1(n72480), .A2(n54267), .B(n54269), 
        .C(n53628), .D(n54272), .Y(n54273) );
  A2O1A1Ixp33_ASAP7_75t_SL U46634 ( .A1(n72485), .A2(n58599), .B(n54273), .C(
        n53628), .Y(n54274) );
  A2O1A1Ixp33_ASAP7_75t_SL U46635 ( .A1(n53628), .A2(n57211), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_6_), .C(n53729), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n121) );
  A2O1A1Ixp33_ASAP7_75t_SL U46636 ( .A1(n71099), .A2(n53628), .B(n71084), .C(
        n53628), .Y(n54261) );
  A2O1A1Ixp33_ASAP7_75t_SL U46637 ( .A1(n54261), .A2(n53628), .B(n54262), .C(
        n53628), .Y(n54263) );
  A2O1A1Ixp33_ASAP7_75t_SL U46638 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_27_), .A2(n53628), 
        .B(n54263), .C(n54266), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n184) );
  A2O1A1Ixp33_ASAP7_75t_SL U46639 ( .A1(n78380), .A2(n53628), .B(n78381), .C(
        n53628), .Y(n54260) );
  A2O1A1Ixp33_ASAP7_75t_SL U46640 ( .A1(n54260), .A2(n53628), .B(n71530), .C(
        n53628), .Y(n71535) );
  A2O1A1Ixp33_ASAP7_75t_SL U46641 ( .A1(n76813), .A2(n53628), .B(n54259), .C(
        n53628), .Y(n76840) );
  A2O1A1Ixp33_ASAP7_75t_SL U46642 ( .A1(n73887), .A2(n73886), .B(n74256), .C(
        n53628), .Y(n54258) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46643 ( .A1(n73886), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[4]), .B(
        n54258), .C(n53628), .D(n74257), .Y(n74240) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46644 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n70412), .B(n53628), .C(n70411), .Y(n53890) );
  A2O1A1Ixp33_ASAP7_75t_SL U46645 ( .A1(n62477), .A2(n53628), .B(n59442), .C(
        n54257), .Y(n77920) );
  A2O1A1Ixp33_ASAP7_75t_SL U46646 ( .A1(n76206), .A2(n53628), .B(n54253), .C(
        n53628), .Y(n54254) );
  A2O1A1Ixp33_ASAP7_75t_SL U46647 ( .A1(n76550), .A2(n53628), .B(n76549), .C(
        n53628), .Y(n54081) );
  O2A1O1Ixp33_ASAP7_75t_SL U46648 ( .A1(n76548), .A2(n54081), .B(n53628), .C(
        n54084), .Y(n54085) );
  A2O1A1Ixp33_ASAP7_75t_SL U46649 ( .A1(n57168), .A2(n53628), .B(n982), .C(
        n53628), .Y(n54248) );
  A2O1A1Ixp33_ASAP7_75t_SL U46650 ( .A1(n54248), .A2(n53628), .B(n65232), .C(
        n53628), .Y(n78207) );
  A2O1A1Ixp33_ASAP7_75t_SL U46651 ( .A1(n57168), .A2(n53628), .B(n1009), .C(
        n53628), .Y(n54247) );
  A2O1A1Ixp33_ASAP7_75t_SL U46652 ( .A1(n54247), .A2(n53628), .B(n75174), .C(
        n53628), .Y(n78208) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46653 ( .A1(n71690), .A2(n71741), .B(n53628), 
        .C(n71719), .Y(n54072) );
  A2O1A1Ixp33_ASAP7_75t_SL U46654 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[35]), .A2(n66146), 
        .B(n54237), .C(n53628), .Y(n54238) );
  A2O1A1Ixp33_ASAP7_75t_SL U46655 ( .A1(n65670), .A2(n53628), .B(n65582), .C(
        n54238), .Y(n66106) );
  A2O1A1Ixp33_ASAP7_75t_SL U46656 ( .A1(n59627), .A2(n53628), .B(n78429), .C(
        n54235), .Y(n72992) );
  A2O1A1Ixp33_ASAP7_75t_SL U46657 ( .A1(n59632), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[7]), .B(n54232), .C(
        n53628), .Y(n54233) );
  A2O1A1Ixp33_ASAP7_75t_SL U46658 ( .A1(n63573), .A2(n53628), .B(n63572), .C(
        n53628), .Y(n54224) );
  A2O1A1Ixp33_ASAP7_75t_SL U46659 ( .A1(n59572), .A2(n53628), .B(n63571), .C(
        n54224), .Y(n54225) );
  A2O1A1Ixp33_ASAP7_75t_SL U46660 ( .A1(n63574), .A2(n53628), .B(n54225), .C(
        n53628), .Y(n75713) );
  A2O1A1Ixp33_ASAP7_75t_SL U46661 ( .A1(n53628), .A2(n76089), .B(n76088), .C(
        n53854), .Y(n76096) );
  A2O1A1Ixp33_ASAP7_75t_SL U46662 ( .A1(n65142), .A2(n53628), .B(n54220), .C(
        n53628), .Y(n65168) );
  A2O1A1Ixp33_ASAP7_75t_SL U46663 ( .A1(n59564), .A2(n53628), .B(n60978), .C(
        n53628), .Y(n54217) );
  A2O1A1Ixp33_ASAP7_75t_SL U46664 ( .A1(n75927), .A2(n53628), .B(n59594), .C(
        n53628), .Y(n54212) );
  A2O1A1Ixp33_ASAP7_75t_SL U46665 ( .A1(n57097), .A2(n53628), .B(n62965), .C(
        n54213), .Y(n63002) );
  A2O1A1Ixp33_ASAP7_75t_SL U46666 ( .A1(n71355), .A2(n53628), .B(n58301), .C(
        n54211), .Y(n71377) );
  A2O1A1Ixp33_ASAP7_75t_SL U46667 ( .A1(n57362), .A2(n53628), .B(n54209), .C(
        n54210), .Y(n63055) );
  A2O1A1Ixp33_ASAP7_75t_SL U46668 ( .A1(n62088), .A2(n53628), .B(n54207), .C(
        n53628), .Y(n54208) );
  A2O1A1Ixp33_ASAP7_75t_SL U46669 ( .A1(n62073), .A2(n53628), .B(n64146), .C(
        n54208), .Y(n61957) );
  OAI21xp5_ASAP7_75t_SL U46670 ( .A1(n66651), .A2(n54206), .B(n53628), .Y(
        n53264) );
  A2O1A1Ixp33_ASAP7_75t_SL U46671 ( .A1(n3309), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]), .C(n73817), .Y(
        n54203) );
  A2O1A1Ixp33_ASAP7_75t_SL U46672 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .A2(
        n73826), .B(n54203), .C(n53628), .Y(n54204) );
  A2O1A1Ixp33_ASAP7_75t_SL U46673 ( .A1(n57074), .A2(n53628), .B(n2988), .C(
        n54197), .Y(n2989) );
  A2O1A1Ixp33_ASAP7_75t_SL U46674 ( .A1(n74196), .A2(n53628), .B(n74139), .C(
        n53628), .Y(n54196) );
  A2O1A1Ixp33_ASAP7_75t_SL U46675 ( .A1(n54196), .A2(n74140), .B(n74217), .C(
        n53628), .Y(n78197) );
  A2O1A1Ixp33_ASAP7_75t_SL U46676 ( .A1(n59629), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_8_), .C(n54195), .Y(
        n2827) );
  A2O1A1Ixp33_ASAP7_75t_SL U46677 ( .A1(n59629), .A2(n53628), .B(n72842), .C(
        n54194), .Y(n2786) );
  A2O1A1Ixp33_ASAP7_75t_SL U46678 ( .A1(n62000), .A2(n62561), .B(n62072), .C(
        n53628), .Y(n54190) );
  A2O1A1Ixp33_ASAP7_75t_SL U46679 ( .A1(n54169), .A2(n53628), .B(n69801), .C(
        n59621), .Y(n54170) );
  A2O1A1Ixp33_ASAP7_75t_SL U46680 ( .A1(n62054), .A2(n62053), .B(n62056), .C(
        n53628), .Y(n54013) );
  A2O1A1Ixp33_ASAP7_75t_SL U46681 ( .A1(n76990), .A2(n53628), .B(n76693), .C(
        n1828), .Y(n54164) );
  A2O1A1Ixp33_ASAP7_75t_SL U46682 ( .A1(n77847), .A2(n53628), .B(n77597), .C(
        n53628), .Y(n54158) );
  A2O1A1Ixp33_ASAP7_75t_SL U46683 ( .A1(n77639), .A2(n53628), .B(n77598), .C(
        n53628), .Y(n54159) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46684 ( .A1(n77675), .A2(n77599), .B(n54158), 
        .C(n53628), .D(n54159), .Y(n1710) );
  A2O1A1Ixp33_ASAP7_75t_SL U46685 ( .A1(n77214), .A2(n53628), .B(n76237), .C(
        n53628), .Y(n54154) );
  A2O1A1Ixp33_ASAP7_75t_SL U46686 ( .A1(n54154), .A2(n53628), .B(n54157), .C(
        n53628), .Y(n78187) );
  A2O1A1Ixp33_ASAP7_75t_SL U46687 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_1_), 
        .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[24]), .C(
        n53628), .Y(n54151) );
  A2O1A1Ixp33_ASAP7_75t_SL U46688 ( .A1(n74741), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[24]), .C(n53628), 
        .Y(n54152) );
  A2O1A1Ixp33_ASAP7_75t_SL U46689 ( .A1(n54151), .A2(n53628), .B(n54152), .C(
        n53628), .Y(n54153) );
  A2O1A1Ixp33_ASAP7_75t_SL U46690 ( .A1(n57202), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[24]), .C(n54153), 
        .Y(n1611) );
  A2O1A1Ixp33_ASAP7_75t_SL U46691 ( .A1(n59626), .A2(n53628), .B(n78379), .C(
        n53628), .Y(n54150) );
  A2O1A1Ixp33_ASAP7_75t_SL U46692 ( .A1(n57190), .A2(n53628), .B(n78361), .C(
        n53628), .Y(n54149) );
  A2O1A1Ixp33_ASAP7_75t_SL U46693 ( .A1(n57114), .A2(n53628), .B(n1460), .C(
        n54148), .Y(n9294) );
  A2O1A1Ixp33_ASAP7_75t_SL U46694 ( .A1(n77287), .A2(n53628), .B(n76855), .C(
        n53628), .Y(n54146) );
  A2O1A1Ixp33_ASAP7_75t_SL U46695 ( .A1(n4114), .A2(n53628), .B(n54143), .C(
        n53628), .Y(n54144) );
  A2O1A1Ixp33_ASAP7_75t_SL U46696 ( .A1(n64259), .A2(n59701), .B(n54144), .C(
        n53628), .Y(n54145) );
  A2O1A1Ixp33_ASAP7_75t_SL U46697 ( .A1(n787), .A2(n53628), .B(n76523), .C(
        n54145), .Y(n9174) );
  A2O1A1Ixp33_ASAP7_75t_SL U46698 ( .A1(n53628), .A2(n68787), .B(n77600), .C(
        n53628), .Y(n54131) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46699 ( .A1(n63385), .A2(n63352), .B(n53628), 
        .C(n63394), .Y(n54135) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46700 ( .A1(n63352), .A2(n54134), .B(n76897), 
        .C(n53628), .D(n54135), .Y(n54136) );
  A2O1A1Ixp33_ASAP7_75t_SL U46701 ( .A1(n63385), .A2(n53628), .B(n63394), .C(
        n53628), .Y(n54137) );
  A2O1A1Ixp33_ASAP7_75t_SL U46702 ( .A1(n63350), .A2(n53628), .B(n54137), .C(
        n53628), .Y(n54138) );
  A2O1A1Ixp33_ASAP7_75t_SL U46703 ( .A1(n54138), .A2(n53628), .B(n54140), .C(
        n53628), .Y(n54141) );
  O2A1O1Ixp33_ASAP7_75t_SL U46704 ( .A1(n54131), .A2(n54136), .B(n53628), .C(
        n54141), .Y(n54142) );
  A2O1A1Ixp33_ASAP7_75t_SL U46705 ( .A1(n53628), .A2(n57093), .B(
        or1200_cpu_or1200_except_n589), .C(n53953), .Y(
        or1200_cpu_or1200_except_n1793) );
  A2O1A1Ixp33_ASAP7_75t_SL U46706 ( .A1(or1200_cpu_or1200_except_n598), .A2(
        n53628), .B(n57072), .C(n54129), .Y(or1200_cpu_or1200_except_n1796) );
  A2O1A1Ixp33_ASAP7_75t_SL U46707 ( .A1(n72508), .A2(n53628), .B(n72506), .C(
        n53628), .Y(n54117) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46708 ( .A1(n72505), .A2(n72482), .B(n53628), 
        .C(n72504), .Y(n54119) );
  A2O1A1Ixp33_ASAP7_75t_SL U46709 ( .A1(n72494), .A2(n54118), .B(n54119), .C(
        n53628), .Y(n54120) );
  A2O1A1Ixp33_ASAP7_75t_SL U46710 ( .A1(n72509), .A2(n53628), .B(n72503), .C(
        n54120), .Y(n54121) );
  A2O1A1Ixp33_ASAP7_75t_SL U46711 ( .A1(n54117), .A2(n53628), .B(n54121), .C(
        n53628), .Y(n54122) );
  A2O1A1Ixp33_ASAP7_75t_SL U46712 ( .A1(n72471), .A2(n53628), .B(n54124), .C(
        n53628), .Y(n54125) );
  A2O1A1Ixp33_ASAP7_75t_SL U46713 ( .A1(n72476), .A2(n53628), .B(n72475), .C(
        n53628), .Y(n54126) );
  A2O1A1Ixp33_ASAP7_75t_SL U46714 ( .A1(n54123), .A2(n53628), .B(n54125), .C(
        n54126), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n66) );
  A2O1A1Ixp33_ASAP7_75t_SL U46715 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), 
        .A2(n53628), .B(n71563), .C(n53628), .Y(n54105) );
  A2O1A1Ixp33_ASAP7_75t_SL U46716 ( .A1(n71480), .A2(n53628), .B(n71628), .C(
        n53628), .Y(n54106) );
  A2O1A1Ixp33_ASAP7_75t_SL U46717 ( .A1(n71468), .A2(n53628), .B(n54107), .C(
        n54108), .Y(n54109) );
  A2O1A1Ixp33_ASAP7_75t_SL U46718 ( .A1(n71568), .A2(n54106), .B(n54109), .C(
        n53628), .Y(n54110) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46719 ( .A1(n71491), .A2(n54105), .B(n71482), 
        .C(n53628), .D(n54112), .Y(n54113) );
  A2O1A1Ixp33_ASAP7_75t_SL U46720 ( .A1(n72079), .A2(n72054), .B(n71484), .C(
        n53628), .Y(n54114) );
  A2O1A1Ixp33_ASAP7_75t_SL U46721 ( .A1(n71488), .A2(n53628), .B(n54116), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n128) );
  A2O1A1Ixp33_ASAP7_75t_SL U46722 ( .A1(n53628), .A2(n70753), .B(n53725), .C(
        n53728), .Y(n53729) );
  A2O1A1Ixp33_ASAP7_75t_SL U46723 ( .A1(n71155), .A2(n53628), .B(n71292), .C(
        n53628), .Y(n54097) );
  A2O1A1Ixp33_ASAP7_75t_SL U46724 ( .A1(n71137), .A2(n54098), .B(n54099), .C(
        n53628), .Y(n54100) );
  A2O1A1Ixp33_ASAP7_75t_SL U46725 ( .A1(n54100), .A2(n53628), .B(n59698), .C(
        n53628), .Y(n54101) );
  A2O1A1Ixp33_ASAP7_75t_SL U46726 ( .A1(n54097), .A2(n53628), .B(n54101), .C(
        n54103), .Y(n54104) );
  A2O1A1Ixp33_ASAP7_75t_SL U46727 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_31_), .A2(n53628), 
        .B(n57211), .C(n54104), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n196) );
  A2O1A1Ixp33_ASAP7_75t_SL U46728 ( .A1(n2569), .A2(n53628), .B(n77749), .C(
        n3423), .Y(n54093) );
  A2O1A1Ixp33_ASAP7_75t_SL U46729 ( .A1(n62477), .A2(n53628), .B(n59550), .C(
        n54092), .Y(n77856) );
  A2O1A1Ixp33_ASAP7_75t_SL U46730 ( .A1(n62477), .A2(n53628), .B(n1626), .C(
        n54091), .Y(n77880) );
  A2O1A1Ixp33_ASAP7_75t_SL U46731 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[6]), 
        .A2(n53628), .B(n73882), .C(n53628), .Y(n54087) );
  A2O1A1Ixp33_ASAP7_75t_SL U46732 ( .A1(n73885), .A2(n53628), .B(n54087), .C(
        n53628), .Y(n54088) );
  A2O1A1Ixp33_ASAP7_75t_SL U46733 ( .A1(n73891), .A2(n53628), .B(n54088), .C(
        n53628), .Y(n54089) );
  A2O1A1Ixp33_ASAP7_75t_SL U46734 ( .A1(n62477), .A2(n53628), .B(n59582), .C(
        n54086), .Y(n77854) );
  A2O1A1Ixp33_ASAP7_75t_SL U46735 ( .A1(n57160), .A2(n53628), .B(n54080), .C(
        n53628), .Y(n65232) );
  A2O1A1Ixp33_ASAP7_75t_SL U46736 ( .A1(n68996), .A2(n53628), .B(n68995), .C(
        n53628), .Y(n54077) );
  A2O1A1Ixp33_ASAP7_75t_SL U46737 ( .A1(n69213), .A2(n53628), .B(n54075), .C(
        n69212), .Y(n75291) );
  A2O1A1Ixp33_ASAP7_75t_SL U46738 ( .A1(n59580), .A2(n53628), .B(n77745), .C(
        n53628), .Y(n54073) );
  A2O1A1Ixp33_ASAP7_75t_SL U46739 ( .A1(n59548), .A2(n53628), .B(n77741), .C(
        n53628), .Y(n54074) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46740 ( .A1(n57214), .A2(n77742), .B(n54073), 
        .C(n53628), .D(n54074), .Y(n4250) );
  A2O1A1Ixp33_ASAP7_75t_SL U46741 ( .A1(n71890), .A2(n53628), .B(n72005), .C(
        n53628), .Y(n54067) );
  A2O1A1Ixp33_ASAP7_75t_SL U46742 ( .A1(n71993), .A2(n53628), .B(n58422), .C(
        n53628), .Y(n54068) );
  A2O1A1Ixp33_ASAP7_75t_SL U46743 ( .A1(n57207), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .B(n54068), .C(n53628), .Y(n54069) );
  A2O1A1Ixp33_ASAP7_75t_SL U46744 ( .A1(n57208), .A2(n53628), .B(n71995), .C(
        n54069), .Y(n54070) );
  A2O1A1Ixp33_ASAP7_75t_SL U46745 ( .A1(n54067), .A2(n53628), .B(n54070), .C(
        n53628), .Y(n71946) );
  A2O1A1Ixp33_ASAP7_75t_SL U46746 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .A2(n66146), 
        .B(n54064), .C(n53628), .Y(n54065) );
  A2O1A1Ixp33_ASAP7_75t_SL U46747 ( .A1(n65616), .A2(n53628), .B(n65670), .C(
        n54065), .Y(n66159) );
  A2O1A1Ixp33_ASAP7_75t_SL U46748 ( .A1(n66155), .A2(n53628), .B(n54062), .C(
        n53628), .Y(n66112) );
  A2O1A1Ixp33_ASAP7_75t_SL U46749 ( .A1(n58419), .A2(n53628), .B(n65859), .C(
        n53628), .Y(n54059) );
  A2O1A1Ixp33_ASAP7_75t_SL U46750 ( .A1(n57187), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[31]), .B(n54059), 
        .C(n53628), .Y(n54060) );
  A2O1A1Ixp33_ASAP7_75t_SL U46751 ( .A1(n58582), .A2(n53628), .B(n65858), .C(
        n54060), .Y(n54061) );
  A2O1A1Ixp33_ASAP7_75t_SL U46752 ( .A1(n57188), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .B(n54061), 
        .C(n53628), .Y(n66000) );
  A2O1A1Ixp33_ASAP7_75t_SL U46753 ( .A1(n57187), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]), .B(n54056), 
        .C(n53628), .Y(n54057) );
  A2O1A1Ixp33_ASAP7_75t_SL U46754 ( .A1(n65466), .A2(n53628), .B(n54053), .C(
        n53628), .Y(n65661) );
  A2O1A1Ixp33_ASAP7_75t_SL U46755 ( .A1(n70120), .A2(n53628), .B(n54051), .C(
        n53628), .Y(n70122) );
  A2O1A1Ixp33_ASAP7_75t_SL U46756 ( .A1(n61882), .A2(n53628), .B(n61884), .C(
        n53628), .Y(n54049) );
  A2O1A1Ixp33_ASAP7_75t_SL U46757 ( .A1(n63571), .A2(n53628), .B(n59533), .C(
        n54049), .Y(n54050) );
  A2O1A1Ixp33_ASAP7_75t_SL U46758 ( .A1(n62107), .A2(n53628), .B(n54050), .C(
        n53628), .Y(n77100) );
  A2O1A1Ixp33_ASAP7_75t_SL U46759 ( .A1(n75605), .A2(n64754), .B(n75882), .C(
        n53628), .Y(n54043) );
  A2O1A1Ixp33_ASAP7_75t_SL U46760 ( .A1(n57075), .A2(n53628), .B(n59308), .C(
        n53628), .Y(n54042) );
  A2O1A1Ixp33_ASAP7_75t_SL U46761 ( .A1(n54041), .A2(n53628), .B(n54042), .C(
        n53628), .Y(n62857) );
  A2O1A1Ixp33_ASAP7_75t_SL U46762 ( .A1(n54041), .A2(n53628), .B(n54042), .C(
        n53628), .Y(n53458) );
  A2O1A1Ixp33_ASAP7_75t_SL U46763 ( .A1(n76125), .A2(n76126), .B(n54040), .C(
        n53628), .Y(n76144) );
  A2O1A1Ixp33_ASAP7_75t_SL U46764 ( .A1(n57187), .A2(n65824), .B(n54037), .C(
        n53628), .Y(n54038) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46765 ( .A1(n75043), .A2(n75076), .B(n53628), 
        .C(n54034), .Y(n75039) );
  A2O1A1Ixp33_ASAP7_75t_SL U46766 ( .A1(n66425), .A2(n53628), .B(n66488), .C(
        n53628), .Y(n54030) );
  A2O1A1Ixp33_ASAP7_75t_SL U46767 ( .A1(n66486), .A2(n66488), .B(n66492), .C(
        n53628), .Y(n54031) );
  A2O1A1Ixp33_ASAP7_75t_SL U46768 ( .A1(n54030), .A2(n53628), .B(n54031), .C(
        n53628), .Y(n66445) );
  A2O1A1Ixp33_ASAP7_75t_SL U46769 ( .A1(n59578), .A2(n53628), .B(n53232), .C(
        n57120), .Y(n54028) );
  A2O1A1Ixp33_ASAP7_75t_SL U46770 ( .A1(n53595), .A2(n53628), .B(n54026), .C(
        n54027), .Y(n66950) );
  A2O1A1Ixp33_ASAP7_75t_SL U46771 ( .A1(n59653), .A2(n53628), .B(n67712), .C(
        n54021), .Y(n67061) );
  O2A1O1Ixp33_ASAP7_75t_SL U46772 ( .A1(n73440), .A2(n73439), .B(n53628), .C(
        n73438), .Y(n53823) );
  A2O1A1Ixp33_ASAP7_75t_SL U46773 ( .A1(n73438), .A2(n53628), .B(n73439), .C(
        n73440), .Y(n53825) );
  O2A1O1Ixp33_ASAP7_75t_SL U46774 ( .A1(n69973), .A2(n69972), .B(n53628), .C(
        n69878), .Y(n53816) );
  A2O1A1Ixp33_ASAP7_75t_SL U46775 ( .A1(n57073), .A2(n53628), .B(wb_insn[16]), 
        .C(n54018), .Y(n2651) );
  A2O1A1Ixp33_ASAP7_75t_SL U46776 ( .A1(n53628), .A2(n57144), .B(n77860), .C(
        n53810), .Y(n2556) );
  A2O1A1Ixp33_ASAP7_75t_SL U46777 ( .A1(n53628), .A2(n74797), .B(n69343), .C(
        n53807), .Y(n2493) );
  A2O1A1Ixp33_ASAP7_75t_SL U46778 ( .A1(n59521), .A2(n53805), .B(n70477), .C(
        n53628), .Y(n53806) );
  A2O1A1Ixp33_ASAP7_75t_SL U46779 ( .A1(n53628), .A2(n59688), .B(n2042), .C(
        n53797), .Y(n2043) );
  A2O1A1Ixp33_ASAP7_75t_SL U46780 ( .A1(n53628), .A2(n59629), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_), .C(n53796), .Y(
        n2012) );
  A2O1A1Ixp33_ASAP7_75t_SL U46781 ( .A1(n77847), .A2(n53628), .B(n77600), .C(
        n53628), .Y(n54006) );
  A2O1A1Ixp33_ASAP7_75t_SL U46782 ( .A1(n77601), .A2(n53628), .B(n77639), .C(
        n53628), .Y(n54007) );
  A2O1A1Ixp33_ASAP7_75t_SL U46783 ( .A1(n77602), .A2(n53628), .B(n77645), .C(
        n53628), .Y(n54008) );
  O2A1O1Ixp5_ASAP7_75t_SL U46784 ( .A1(n54006), .A2(n54007), .B(n53628), .C(
        n54008), .Y(n1709) );
  A2O1A1Ixp33_ASAP7_75t_SL U46785 ( .A1(n78370), .A2(n53628), .B(n59626), .C(
        n53628), .Y(n54005) );
  A2O1A1Ixp33_ASAP7_75t_SL U46786 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_), .A2(n57190), .B(
        n54005), .C(n53628), .Y(n1558) );
  A2O1A1Ixp33_ASAP7_75t_SL U46787 ( .A1(n57114), .A2(n53628), .B(n1458), .C(
        n54004), .Y(n9293) );
  A2O1A1Ixp33_ASAP7_75t_SL U46788 ( .A1(n74641), .A2(n53628), .B(n1366), .C(
        n53998), .Y(n9311) );
  A2O1A1Ixp33_ASAP7_75t_SL U46789 ( .A1(n4112), .A2(n53628), .B(n53995), .C(
        n53628), .Y(n53996) );
  A2O1A1Ixp33_ASAP7_75t_SL U46790 ( .A1(n65191), .A2(n59701), .B(n53996), .C(
        n53628), .Y(n53997) );
  A2O1A1Ixp33_ASAP7_75t_SL U46791 ( .A1(n783), .A2(n53628), .B(n76523), .C(
        n53997), .Y(n9173) );
  A2O1A1Ixp33_ASAP7_75t_SL U46792 ( .A1(n75990), .A2(n53628), .B(n53991), .C(
        n53628), .Y(n53992) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46793 ( .A1(
        or1200_cpu_or1200_mult_mac_mac_op_r2_0_), .A2(
        or1200_cpu_or1200_mult_mac_mac_op_r2_1_), .B(n53628), .C(
        or1200_cpu_or1200_mult_mac_mac_op_r2_2_), .Y(n53986) );
  A2O1A1Ixp33_ASAP7_75t_SL U46794 ( .A1(n53987), .A2(n53628), .B(n53988), .C(
        n53628), .Y(n53989) );
  A2O1A1Ixp33_ASAP7_75t_SL U46795 ( .A1(or1200_cpu_or1200_mult_mac_n139), .A2(
        n53985), .B(n53989), .C(n53628), .Y(or1200_cpu_or1200_mult_mac_N503)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46796 ( .A1(n63270), .A2(
        or1200_cpu_or1200_mult_mac_n287), .B(n63274), .C(n53628), .Y(n53979)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46797 ( .A1(n53979), .A2(n53628), .B(n53980), .C(
        n53628), .Y(n53981) );
  A2O1A1Ixp33_ASAP7_75t_SL U46798 ( .A1(or1200_cpu_or1200_mult_mac_n141), .A2(
        n53628), .B(n76889), .C(n53628), .Y(n53982) );
  A2O1A1Ixp33_ASAP7_75t_SL U46799 ( .A1(n53981), .A2(n53628), .B(n53982), .C(
        n53628), .Y(n53983) );
  A2O1A1Ixp33_ASAP7_75t_SL U46800 ( .A1(n63507), .A2(n53628), .B(n53965), .C(
        n53628), .Y(n53966) );
  A2O1A1Ixp33_ASAP7_75t_SL U46801 ( .A1(n63517), .A2(n53628), .B(n53966), .C(
        n53628), .Y(n53967) );
  A2O1A1Ixp33_ASAP7_75t_SL U46802 ( .A1(n63513), .A2(n53628), .B(n53967), .C(
        n53628), .Y(n53968) );
  A2O1A1Ixp33_ASAP7_75t_SL U46803 ( .A1(n63510), .A2(n53628), .B(n53973), .C(
        n53628), .Y(n53974) );
  A2O1A1Ixp33_ASAP7_75t_SL U46804 ( .A1(n59674), .A2(n53972), .B(n53977), .C(
        n53628), .Y(n53978) );
  A2O1A1Ixp33_ASAP7_75t_SL U46805 ( .A1(n57072), .A2(n53628), .B(
        or1200_cpu_or1200_except_n607), .C(n53952), .Y(
        or1200_cpu_or1200_except_n1799) );
  A2O1A1Ixp33_ASAP7_75t_SL U46806 ( .A1(n72328), .A2(n53628), .B(n72327), .C(
        n53628), .Y(n53945) );
  A2O1A1Ixp33_ASAP7_75t_SL U46807 ( .A1(n72417), .A2(n72491), .B(n53941), .C(
        n53628), .Y(n53942) );
  A2O1A1Ixp33_ASAP7_75t_SL U46808 ( .A1(n72432), .A2(n53628), .B(n53939), .C(
        n53940), .Y(n53941) );
  A2O1A1Ixp33_ASAP7_75t_SL U46809 ( .A1(n71797), .A2(n53628), .B(n53938), .C(
        n71796), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n110) );
  A2O1A1Ixp33_ASAP7_75t_SL U46810 ( .A1(n53628), .A2(n59699), .B(n70746), .C(
        n53628), .Y(n53725) );
  A2O1A1Ixp33_ASAP7_75t_SL U46811 ( .A1(n66147), .A2(n53628), .B(n66148), .C(
        n53628), .Y(n53914) );
  A2O1A1Ixp33_ASAP7_75t_SL U46812 ( .A1(n66153), .A2(n53628), .B(n66154), .C(
        n53628), .Y(n53915) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46813 ( .A1(n66149), .A2(n66162), .B(n53914), 
        .C(n53628), .D(n53915), .Y(n53916) );
  A2O1A1Ixp33_ASAP7_75t_SL U46814 ( .A1(n66150), .A2(n53628), .B(n53913), .C(
        n53916), .Y(n53917) );
  A2O1A1Ixp33_ASAP7_75t_SL U46815 ( .A1(n66156), .A2(n53628), .B(n66157), .C(
        n53628), .Y(n53918) );
  A2O1A1Ixp33_ASAP7_75t_SL U46816 ( .A1(n66160), .A2(n53628), .B(n66161), .C(
        n53628), .Y(n53919) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46817 ( .A1(n66162), .A2(n66163), .B(n53918), 
        .C(n53628), .D(n53919), .Y(n53920) );
  A2O1A1Ixp33_ASAP7_75t_SL U46818 ( .A1(n66158), .A2(n53628), .B(n66159), .C(
        n53920), .Y(n53921) );
  A2O1A1Ixp33_ASAP7_75t_SL U46819 ( .A1(n66145), .A2(n53628), .B(n66144), .C(
        n53628), .Y(n53922) );
  A2O1A1Ixp33_ASAP7_75t_SL U46820 ( .A1(n53922), .A2(n53628), .B(n66155), .C(
        n53628), .Y(n53923) );
  A2O1A1Ixp33_ASAP7_75t_SL U46821 ( .A1(n53923), .A2(n53628), .B(n53926), .C(
        n66167), .Y(n53927) );
  O2A1O1Ixp5_ASAP7_75t_SL U46822 ( .A1(n53917), .A2(n53921), .B(n53628), .C(
        n53927), .Y(n53928) );
  A2O1A1Ixp33_ASAP7_75t_SL U46823 ( .A1(n53928), .A2(n53628), .B(n53929), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n6) );
  A2O1A1Ixp33_ASAP7_75t_SL U46824 ( .A1(n61297), .A2(n53628), .B(n77488), .C(
        n53628), .Y(n53911) );
  A2O1A1Ixp33_ASAP7_75t_SL U46825 ( .A1(n75765), .A2(n57160), .B(n77208), .C(
        n53628), .Y(n53907) );
  A2O1A1Ixp33_ASAP7_75t_SL U46826 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_9_), .A2(n53628), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_10_), .C(
        n53628), .Y(n53891) );
  A2O1A1Ixp33_ASAP7_75t_SL U46827 ( .A1(n76950), .A2(n53891), .B(n76949), .C(
        n53628), .Y(n53892) );
  A2O1A1Ixp33_ASAP7_75t_SL U46828 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_6_), .A2(n53628), 
        .B(n76948), .C(n53628), .Y(n53893) );
  A2O1A1Ixp33_ASAP7_75t_SL U46829 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_5_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_6_), .B(n53893), 
        .C(n53628), .Y(n53894) );
  A2O1A1Ixp33_ASAP7_75t_SL U46830 ( .A1(n76945), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_22_), .C(n53628), 
        .Y(n53895) );
  A2O1A1Ixp33_ASAP7_75t_SL U46831 ( .A1(n76946), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_3_), .C(n53628), 
        .Y(n53896) );
  A2O1A1Ixp33_ASAP7_75t_SL U46832 ( .A1(n53895), .A2(n53628), .B(n53896), .C(
        n53628), .Y(n53897) );
  A2O1A1Ixp33_ASAP7_75t_SL U46833 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_11_), .A2(n53628), 
        .B(n53900), .C(n76974), .Y(n53901) );
  A2O1A1Ixp33_ASAP7_75t_SL U46834 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_16_), .A2(n53628), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_18_), .C(
        n76947), .Y(n53905) );
  O2A1O1Ixp33_ASAP7_75t_SL U46835 ( .A1(n53892), .A2(n53894), .B(n53628), .C(
        n53906), .Y(n76951) );
  A2O1A1Ixp33_ASAP7_75t_SL U46836 ( .A1(or1200_cpu_or1200_mult_mac_n229), .A2(
        or1200_cpu_or1200_mult_mac_n375), .B(n69106), .C(n53628), .Y(n53887)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46837 ( .A1(n69107), .A2(n53628), .B(n69108), .C(
        n53887), .Y(n53888) );
  A2O1A1Ixp33_ASAP7_75t_SL U46838 ( .A1(n69361), .A2(n53628), .B(n53886), .C(
        n53628), .Y(n78100) );
  A2O1A1Ixp33_ASAP7_75t_SL U46839 ( .A1(n71873), .A2(n53628), .B(n72285), .C(
        n53628), .Y(n53884) );
  A2O1A1Ixp33_ASAP7_75t_SL U46840 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .A2(
        n53628), .B(n72061), .C(n53628), .Y(n53885) );
  A2O1A1Ixp33_ASAP7_75t_SL U46841 ( .A1(n53884), .A2(n53628), .B(n53885), .C(
        n53628), .Y(n72334) );
  A2O1A1Ixp33_ASAP7_75t_SL U46842 ( .A1(n72141), .A2(n53628), .B(n71890), .C(
        n53628), .Y(n53880) );
  A2O1A1Ixp33_ASAP7_75t_SL U46843 ( .A1(n58422), .A2(n53628), .B(n72079), .C(
        n53628), .Y(n53881) );
  A2O1A1Ixp33_ASAP7_75t_SL U46844 ( .A1(n57207), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_), 
        .B(n53881), .C(n53628), .Y(n53882) );
  A2O1A1Ixp33_ASAP7_75t_SL U46845 ( .A1(n57208), .A2(n53628), .B(n72080), .C(
        n53882), .Y(n53883) );
  A2O1A1Ixp33_ASAP7_75t_SL U46846 ( .A1(n53880), .A2(n53628), .B(n53883), .C(
        n53628), .Y(n72025) );
  A2O1A1Ixp33_ASAP7_75t_SL U46847 ( .A1(n72738), .A2(n53628), .B(n73010), .C(
        n53628), .Y(n53872) );
  A2O1A1Ixp33_ASAP7_75t_SL U46848 ( .A1(n72901), .A2(n53628), .B(n72859), .C(
        n53628), .Y(n53873) );
  A2O1A1Ixp33_ASAP7_75t_SL U46849 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[8]), .A2(n57217), .B(
        n53868), .C(n53628), .Y(n53869) );
  A2O1A1Ixp33_ASAP7_75t_SL U46850 ( .A1(n75415), .A2(n53628), .B(n75414), .C(
        n53628), .Y(n53862) );
  A2O1A1Ixp33_ASAP7_75t_SL U46851 ( .A1(n64265), .A2(n53628), .B(n64264), .C(
        n53862), .Y(n65203) );
  A2O1A1Ixp33_ASAP7_75t_SL U46852 ( .A1(or1200_cpu_or1200_mult_mac_n86), .A2(
        n53628), .B(n61826), .C(n53861), .Y(n64316) );
  A2O1A1Ixp33_ASAP7_75t_SL U46853 ( .A1(n63584), .A2(n53628), .B(n75734), .C(
        n53628), .Y(n53856) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46854 ( .A1(n74603), .A2(n59709), .B(n53856), 
        .C(n53628), .D(n53859), .Y(n63585) );
  A2O1A1Ixp33_ASAP7_75t_SL U46855 ( .A1(n57208), .A2(n53628), .B(n72311), .C(
        n53628), .Y(n53848) );
  A2O1A1Ixp33_ASAP7_75t_SL U46856 ( .A1(n53848), .A2(n53628), .B(n53851), .C(
        n53628), .Y(n53852) );
  A2O1A1Ixp33_ASAP7_75t_SL U46857 ( .A1(n62308), .A2(n53628), .B(n53847), .C(
        n53628), .Y(n76278) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46858 ( .A1(n75081), .A2(n75083), .B(n53628), 
        .C(n53846), .Y(n75084) );
  A2O1A1Ixp33_ASAP7_75t_SL U46859 ( .A1(n57178), .A2(n53628), .B(n58701), .C(
        n53628), .Y(n53843) );
  INVx1_ASAP7_75t_SL U46860 ( .A(n76028), .Y(n53256) );
  A2O1A1Ixp33_ASAP7_75t_SL U46861 ( .A1(n59142), .A2(n53628), .B(n53833), .C(
        n53628), .Y(n53834) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46862 ( .A1(n64567), .A2(n53832), .B(n53834), 
        .C(n53628), .D(n66385), .Y(n53835) );
  A2O1A1Ixp33_ASAP7_75t_SL U46863 ( .A1(n53205), .A2(n66372), .B(n53836), .C(
        n53628), .Y(n53837) );
  A2O1A1Ixp33_ASAP7_75t_SL U46864 ( .A1(n66429), .A2(n53831), .B(n53837), .C(
        n53628), .Y(n66438) );
  A2O1A1Ixp33_ASAP7_75t_SL U46865 ( .A1(n57097), .A2(n53628), .B(n63156), .C(
        n53628), .Y(n53830) );
  A2O1A1Ixp33_ASAP7_75t_SL U46866 ( .A1(n59637), .A2(n53628), .B(n67569), .C(
        n53827), .Y(n66666) );
  A2O1A1Ixp33_ASAP7_75t_SL U46867 ( .A1(n57871), .A2(n53628), .B(n58254), .C(
        n53826), .Y(n67932) );
  A2O1A1Ixp33_ASAP7_75t_SL U46868 ( .A1(n73835), .A2(n53628), .B(n73818), .C(
        n53628), .Y(n53820) );
  A2O1A1Ixp33_ASAP7_75t_SL U46869 ( .A1(n3327), .A2(n59705), .B(n53820), .C(
        n53628), .Y(n53821) );
  A2O1A1Ixp33_ASAP7_75t_SL U46870 ( .A1(n69877), .A2(n53628), .B(n70085), .C(
        n53628), .Y(n53817) );
  A2O1A1Ixp33_ASAP7_75t_SL U46871 ( .A1(n53816), .A2(n53628), .B(n53817), .C(
        n53628), .Y(n53818) );
  A2O1A1Ixp33_ASAP7_75t_SL U46872 ( .A1(n57074), .A2(n53628), .B(n2646), .C(
        n53815), .Y(n2647) );
  A2O1A1Ixp33_ASAP7_75t_SL U46873 ( .A1(n2555), .A2(n53628), .B(n53808), .C(
        n53628), .Y(n53809) );
  A2O1A1Ixp33_ASAP7_75t_SL U46874 ( .A1(n62061), .A2(n53798), .B(n62060), .C(
        n53628), .Y(n53799) );
  A2O1A1Ixp33_ASAP7_75t_SL U46875 ( .A1(n65399), .A2(n53628), .B(n53794), .C(
        n53628), .Y(n53795) );
  A2O1A1Ixp33_ASAP7_75t_SL U46876 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_3_), .A2(n65401), .B(
        n53795), .C(n53628), .Y(n1969) );
  A2O1A1Ixp33_ASAP7_75t_SL U46877 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[5]), .A2(n53628), .B(n57190), .C(n53793), .Y(n1833) );
  A2O1A1Ixp33_ASAP7_75t_SL U46878 ( .A1(n77609), .A2(n53628), .B(n77645), .C(
        n53628), .Y(n53789) );
  A2O1A1Ixp33_ASAP7_75t_SL U46879 ( .A1(n53789), .A2(n53628), .B(n53792), .C(
        n53628), .Y(n1708) );
  A2O1A1Ixp33_ASAP7_75t_SL U46880 ( .A1(n1692), .A2(n53628), .B(n53786), .C(
        n53628), .Y(n53787) );
  A2O1A1Ixp33_ASAP7_75t_SL U46881 ( .A1(n57114), .A2(n53628), .B(n1456), .C(
        n53785), .Y(n9292) );
  A2O1A1Ixp33_ASAP7_75t_SL U46882 ( .A1(n74641), .A2(n53628), .B(n1362), .C(
        n53784), .Y(n9310) );
  A2O1A1Ixp33_ASAP7_75t_SL U46883 ( .A1(n77287), .A2(n53628), .B(n74972), .C(
        n53628), .Y(n53782) );
  A2O1A1Ixp33_ASAP7_75t_SL U46884 ( .A1(n4110), .A2(n53628), .B(n53779), .C(
        n53628), .Y(n53780) );
  A2O1A1Ixp33_ASAP7_75t_SL U46885 ( .A1(n65212), .A2(n59701), .B(n53780), .C(
        n53628), .Y(n53781) );
  A2O1A1Ixp33_ASAP7_75t_SL U46886 ( .A1(n65213), .A2(n53628), .B(n76839), .C(
        n53781), .Y(n9172) );
  A2O1A1Ixp33_ASAP7_75t_SL U46887 ( .A1(n68787), .A2(n53628), .B(n77594), .C(
        n53628), .Y(n53772) );
  A2O1A1Ixp33_ASAP7_75t_SL U46888 ( .A1(or1200_cpu_or1200_mult_mac_n149), .A2(
        n53628), .B(n76889), .C(n53778), .Y(or1200_cpu_or1200_mult_mac_n1589)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46889 ( .A1(n68877), .A2(n53628), .B(n68861), .C(
        n53628), .Y(n53760) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U46890 ( .A1(n76906), .A2(n53760), .B(n53628), 
        .C(n68872), .Y(n53761) );
  A2O1A1Ixp33_ASAP7_75t_SL U46891 ( .A1(n68873), .A2(n53628), .B(n53762), .C(
        n53628), .Y(n53763) );
  A2O1A1Ixp33_ASAP7_75t_SL U46892 ( .A1(n68863), .A2(n68881), .B(n68882), .C(
        n53628), .Y(n53764) );
  A2O1A1Ixp33_ASAP7_75t_SL U46893 ( .A1(n59671), .A2(n53628), .B(n53764), .C(
        n53628), .Y(n53767) );
  A2O1A1Ixp33_ASAP7_75t_SL U46894 ( .A1(n53767), .A2(n53628), .B(n53763), .C(
        n53628), .Y(n53768) );
  A2O1A1Ixp33_ASAP7_75t_SL U46895 ( .A1(n53760), .A2(n53628), .B(n68872), .C(
        n57080), .Y(n53769) );
  A2O1A1Ixp33_ASAP7_75t_SL U46896 ( .A1(n53761), .A2(n53628), .B(n53766), .C(
        n53770), .Y(n53771) );
  A2O1A1Ixp33_ASAP7_75t_SL U46897 ( .A1(n69057), .A2(n53628), .B(n69020), .C(
        n69060), .Y(n53748) );
  A2O1A1Ixp33_ASAP7_75t_SL U46898 ( .A1(n76906), .A2(n53628), .B(n53748), .C(
        n53628), .Y(n53749) );
  A2O1A1Ixp33_ASAP7_75t_SL U46899 ( .A1(n69072), .A2(n53628), .B(n59671), .C(
        n53628), .Y(n53753) );
  A2O1A1Ixp33_ASAP7_75t_SL U46900 ( .A1(n53753), .A2(n53628), .B(n53750), .C(
        n53628), .Y(n53754) );
  A2O1A1Ixp33_ASAP7_75t_SL U46901 ( .A1(n53749), .A2(n53628), .B(n53752), .C(
        n53756), .Y(n53757) );
  A2O1A1Ixp33_ASAP7_75t_SL U46902 ( .A1(n77615), .A2(n53628), .B(n76661), .C(
        n53628), .Y(n53742) );
  A2O1A1Ixp33_ASAP7_75t_SL U46903 ( .A1(or1200_cpu_or1200_except_n262), .A2(
        n53628), .B(n76507), .C(n53628), .Y(n53743) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U46904 ( .A1(n77220), .A2(n75531), .B(n53742), 
        .C(n53628), .D(n53743), .Y(n53744) );
  A2O1A1Ixp33_ASAP7_75t_SL U46905 ( .A1(n57093), .A2(n53628), .B(
        or1200_cpu_or1200_except_n646), .C(n53741), .Y(
        or1200_cpu_or1200_except_n1812) );
  A2O1A1Ixp33_ASAP7_75t_SL U46906 ( .A1(n72510), .A2(n53628), .B(n72468), .C(
        n53628), .Y(n53730) );
  A2O1A1Ixp33_ASAP7_75t_SL U46907 ( .A1(n72466), .A2(n53628), .B(n72508), .C(
        n53628), .Y(n53731) );
  A2O1A1Ixp33_ASAP7_75t_SL U46908 ( .A1(n72464), .A2(n72490), .B(n53731), .C(
        n53628), .Y(n53732) );
  A2O1A1Ixp33_ASAP7_75t_SL U46909 ( .A1(n72507), .A2(n53628), .B(n72465), .C(
        n53732), .Y(n53733) );
  A2O1A1Ixp33_ASAP7_75t_SL U46910 ( .A1(n72502), .A2(n72463), .B(n53733), .C(
        n53628), .Y(n53734) );
  A2O1A1Ixp33_ASAP7_75t_SL U46911 ( .A1(n53730), .A2(n53628), .B(n53735), .C(
        n53628), .Y(n53736) );
  A2O1A1Ixp33_ASAP7_75t_SL U46912 ( .A1(n72499), .A2(n53628), .B(n72470), .C(
        n72469), .Y(n53737) );
  A2O1A1Ixp33_ASAP7_75t_SL U46913 ( .A1(n53736), .A2(n53628), .B(n53737), .C(
        n53628), .Y(n53738) );
  A2O1A1Ixp33_ASAP7_75t_SL U46914 ( .A1(n57192), .A2(n53628), .B(n72467), .C(
        n53738), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n68) );
  A2O1A1Ixp33_ASAP7_75t_SL U46915 ( .A1(n57211), .A2(n53628), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_33_), .C(n53724), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n202) );
  A2O1A1Ixp33_ASAP7_75t_SL U46916 ( .A1(n65989), .A2(n53628), .B(n53718), .C(
        n53628), .Y(n53719) );
  A2O1A1Ixp33_ASAP7_75t_SL U46917 ( .A1(n66086), .A2(n66067), .B(n53719), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n11) );
  A2O1A1Ixp33_ASAP7_75t_SL U46918 ( .A1(n70576), .A2(n53715), .B(n70236), .C(
        n53628), .Y(n53716) );
  A2O1A1Ixp33_ASAP7_75t_SL U46919 ( .A1(n70576), .A2(n53628), .B(n53715), .C(
        n53716), .Y(n53717) );
  A2O1A1Ixp33_ASAP7_75t_SL U46920 ( .A1(n78429), .A2(n53628), .B(n70078), .C(
        n53628), .Y(n53714) );
  A2O1A1Ixp33_ASAP7_75t_SL U46921 ( .A1(n76557), .A2(n53628), .B(n76558), .C(
        n53713), .Y(n77408) );
  A2O1A1Ixp33_ASAP7_75t_SL U46922 ( .A1(n1347), .A2(n53628), .B(n77412), .C(
        n57083), .Y(n53709) );
  A2O1A1Ixp33_ASAP7_75t_SL U46923 ( .A1(n57083), .A2(n53628), .B(n59713), .C(
        n53628), .Y(n53710) );
  A2O1A1Ixp33_ASAP7_75t_SL U46924 ( .A1(n64265), .A2(n53628), .B(n65207), .C(
        n53708), .Y(n75419) );
  A2O1A1Ixp33_ASAP7_75t_SL U46925 ( .A1(n53702), .A2(n53628), .B(n53703), .C(
        n53628), .Y(n53704) );
  A2O1A1Ixp33_ASAP7_75t_SL U46926 ( .A1(n53705), .A2(n53628), .B(n53706), .C(
        n53628), .Y(n53707) );
  A2O1A1Ixp33_ASAP7_75t_SL U46927 ( .A1(n77194), .A2(n53700), .B(n74872), .C(
        n53628), .Y(n77197) );
  A2O1A1Ixp33_ASAP7_75t_SL U46928 ( .A1(n74656), .A2(n74686), .B(n53697), .C(
        n53628), .Y(n53698) );
  A2O1A1Ixp33_ASAP7_75t_SL U46929 ( .A1(n70540), .A2(n53628), .B(n74660), .C(
        n53698), .Y(n70473) );
  A2O1A1Ixp33_ASAP7_75t_SL U46930 ( .A1(n77161), .A2(n53628), .B(n53695), .C(
        n53628), .Y(n77201) );
  A2O1A1Ixp33_ASAP7_75t_SL U46931 ( .A1(n75760), .A2(n53628), .B(n53694), .C(
        n53628), .Y(n76631) );
  A2O1A1Ixp33_ASAP7_75t_SL U46932 ( .A1(n69170), .A2(n53628), .B(n53693), .C(
        n53628), .Y(n69194) );
  A2O1A1Ixp33_ASAP7_75t_SL U46933 ( .A1(n74117), .A2(n53628), .B(n53692), .C(
        n53628), .Y(n69260) );
  A2O1A1Ixp33_ASAP7_75t_SL U46934 ( .A1(n53628), .A2(n53690), .B(n75660), .C(
        n53628), .Y(n53691) );
  A2O1A1Ixp33_ASAP7_75t_SL U46935 ( .A1(n59622), .A2(n53628), .B(n72228), .C(
        n53628), .Y(n53684) );
  A2O1A1Ixp33_ASAP7_75t_SL U46936 ( .A1(n72298), .A2(n53628), .B(n59623), .C(
        n53628), .Y(n53685) );
  A2O1A1Ixp33_ASAP7_75t_SL U46937 ( .A1(n59624), .A2(n53628), .B(n72226), .C(
        n53628), .Y(n53686) );
  O2A1O1Ixp5_ASAP7_75t_SL U46938 ( .A1(n53684), .A2(n53685), .B(n53628), .C(
        n53686), .Y(n72484) );
  A2O1A1Ixp33_ASAP7_75t_SL U46939 ( .A1(n71698), .A2(n71678), .B(n71679), .C(
        n53628), .Y(n71801) );
  A2O1A1Ixp33_ASAP7_75t_SL U46940 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[34]), .A2(n57193), 
        .B(n53677), .C(n53628), .Y(n53678) );
  A2O1A1Ixp33_ASAP7_75t_SL U46941 ( .A1(n78373), .A2(n53628), .B(n59626), .C(
        n53628), .Y(n53674) );
  A2O1A1Ixp33_ASAP7_75t_SL U46942 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_), .A2(n57190), .B(n53674), 
        .C(n53628), .Y(n72635) );
  A2O1A1Ixp33_ASAP7_75t_SL U46943 ( .A1(n59630), .A2(n53628), .B(n73133), .C(
        n53672), .Y(n73297) );
  A2O1A1Ixp33_ASAP7_75t_SL U46944 ( .A1(n74103), .A2(n53628), .B(n53671), .C(
        n53628), .Y(n73881) );
  A2O1A1Ixp33_ASAP7_75t_SL U46945 ( .A1(n61434), .A2(n53628), .B(n53666), .C(
        n53628), .Y(n53667) );
  A2O1A1Ixp33_ASAP7_75t_SL U46946 ( .A1(n61648), .A2(n53628), .B(n53660), .C(
        n53628), .Y(n53661) );
  A2O1A1Ixp33_ASAP7_75t_SL U46947 ( .A1(n76859), .A2(n53628), .B(n76861), .C(
        n53628), .Y(n53656) );
  A2O1A1Ixp33_ASAP7_75t_SL U46948 ( .A1(n53656), .A2(n53628), .B(n53657), .C(
        n53628), .Y(n76862) );
  A2O1A1Ixp33_ASAP7_75t_SL U46949 ( .A1(n64114), .A2(n53628), .B(n53655), .C(
        n53628), .Y(n75424) );
  A2O1A1Ixp33_ASAP7_75t_SL U46950 ( .A1(n1095), .A2(n53628), .B(n61268), .C(
        n53628), .Y(n53654) );
  A2O1A1Ixp33_ASAP7_75t_SL U46951 ( .A1(n63542), .A2(n53652), .B(n53653), .C(
        n53628), .Y(n63893) );
  A2O1A1Ixp33_ASAP7_75t_SL U46952 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_), 
        .A2(n53628), .B(n57208), .C(n53628), .Y(n53646) );
  A2O1A1Ixp33_ASAP7_75t_SL U46953 ( .A1(n53646), .A2(n53628), .B(n53649), .C(
        n53628), .Y(n53650) );
  A2O1A1Ixp33_ASAP7_75t_SL U46954 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_1_), .A2(
        n53628), .B(n71655), .C(n53628), .Y(n53645) );
  A2O1A1Ixp33_ASAP7_75t_SL U46955 ( .A1(n71670), .A2(n53628), .B(n53645), .C(
        n53628), .Y(n71648) );
  A2O1A1Ixp33_ASAP7_75t_SL U46956 ( .A1(n71569), .A2(n53628), .B(n53644), .C(
        n53628), .Y(n71556) );
  A2O1A1Ixp33_ASAP7_75t_SL U46957 ( .A1(n71316), .A2(n53628), .B(n53639), .C(
        n53628), .Y(n53640) );
  A2O1A1Ixp33_ASAP7_75t_SL U46958 ( .A1(n71262), .A2(n53628), .B(n71335), .C(
        n53628), .Y(n53641) );
  A2O1A1Ixp33_ASAP7_75t_SL U46959 ( .A1(n71315), .A2(n71376), .B(n53641), .C(
        n53628), .Y(n53642) );
  A2O1A1Ixp33_ASAP7_75t_SL U46960 ( .A1(n71318), .A2(n53628), .B(n71362), .C(
        n53642), .Y(n53643) );
  A2O1A1Ixp33_ASAP7_75t_SL U46961 ( .A1(n53640), .A2(n53628), .B(n53643), .C(
        n53628), .Y(n71264) );
  A2O1A1Ixp33_ASAP7_75t_SL U46962 ( .A1(n59560), .A2(n53628), .B(n53638), .C(
        n59541), .Y(n60934) );
  A2O1A1Ixp33_ASAP7_75t_SL U46963 ( .A1(n75076), .A2(n53628), .B(n75077), .C(
        n75075), .Y(n53637) );
  A2O1A1Ixp33_ASAP7_75t_SL U46964 ( .A1(n67227), .A2(n53628), .B(n57720), .C(
        n53628), .Y(n53633) );
  A2O1A1Ixp33_ASAP7_75t_SL U46965 ( .A1(n57494), .A2(n59440), .B(n53631), .C(
        n53628), .Y(n66574) );
  A2O1A1Ixp33_ASAP7_75t_SL U46966 ( .A1(n59598), .A2(n53628), .B(n75962), .C(
        n53628), .Y(n53629) );
  A2O1A1Ixp33_ASAP7_75t_SL U46967 ( .A1(n76176), .A2(n59599), .B(n53629), .C(
        n53628), .Y(n66994) );
  A2O1A1Ixp33_ASAP7_75t_SL U46968 ( .A1(n56634), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56635) );
  A2O1A1Ixp33_ASAP7_75t_SL U46969 ( .A1(n56541), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56542) );
  A2O1A1Ixp33_ASAP7_75t_SL U46970 ( .A1(n56535), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56536) );
  A2O1A1Ixp33_ASAP7_75t_SL U46971 ( .A1(n55849), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55850) );
  A2O1A1Ixp33_ASAP7_75t_SL U46972 ( .A1(n56437), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56438) );
  A2O1A1Ixp33_ASAP7_75t_SL U46973 ( .A1(n56219), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56220) );
  A2O1A1Ixp33_ASAP7_75t_SL U46974 ( .A1(n55820), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55823) );
  A2O1A1Ixp33_ASAP7_75t_SL U46975 ( .A1(n75139), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55807) );
  A2O1A1Ixp33_ASAP7_75t_SL U46976 ( .A1(n55452), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55453) );
  A2O1A1Ixp33_ASAP7_75t_SL U46977 ( .A1(n53628), .A2(n55453), .B(n53192), .C(
        n53628), .Y(n55454) );
  A2O1A1Ixp33_ASAP7_75t_SL U46978 ( .A1(n55400), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55401) );
  A2O1A1Ixp33_ASAP7_75t_SL U46979 ( .A1(n55186), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55187) );
  A2O1A1Ixp33_ASAP7_75t_SL U46980 ( .A1(n53968), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n53969) );
  A2O1A1Ixp33_ASAP7_75t_SL U46981 ( .A1(n54312), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54313) );
  A2O1A1Ixp33_ASAP7_75t_SL U46982 ( .A1(n54301), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54302) );
  A2O1A1Ixp33_ASAP7_75t_SL U46983 ( .A1(n73484), .A2(n56650), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_0_)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U46984 ( .A1(n73464), .A2(n56646), .B(n53192), .C(
        n53628), .Y(n56647) );
  A2O1A1Ixp33_ASAP7_75t_SL U46985 ( .A1(n56648), .A2(n73459), .B(n53192), .C(
        n56647), .Y(n56649) );
  A2O1A1Ixp33_ASAP7_75t_SL U46986 ( .A1(n70234), .A2(n70593), .B(n53192), .C(
        n70587), .Y(n54358) );
  A2O1A1Ixp33_ASAP7_75t_SL U46987 ( .A1(n70235), .A2(n54357), .B(n53192), .C(
        n54358), .Y(n3163) );
  A2O1A1Ixp33_ASAP7_75t_SL U46988 ( .A1(n56816), .A2(n56819), .B(n53192), .C(
        n53628), .Y(n56820) );
  A2O1A1Ixp33_ASAP7_75t_SL U46989 ( .A1(n2491), .A2(n74892), .B(n53192), .C(
        n53628), .Y(n56821) );
  A2O1A1Ixp33_ASAP7_75t_SL U46990 ( .A1(n56638), .A2(n56640), .B(n53192), .C(
        n53628), .Y(n56641) );
  A2O1A1Ixp33_ASAP7_75t_SL U46991 ( .A1(n60470), .A2(n60469), .B(n53192), .C(
        n53628), .Y(n56643) );
  A2O1A1Ixp33_ASAP7_75t_SL U46992 ( .A1(n59628), .A2(n72817), .B(n53192), .C(
        n72818), .Y(n56808) );
  A2O1A1Ixp33_ASAP7_75t_SL U46993 ( .A1(n61288), .A2(n56637), .B(n53192), .C(
        n53628), .Y(n9384) );
  A2O1A1Ixp33_ASAP7_75t_SL U46994 ( .A1(n61315), .A2(n56632), .B(n53192), .C(
        n53628), .Y(n56633) );
  A2O1A1Ixp33_ASAP7_75t_SL U46995 ( .A1(n59689), .A2(n56806), .B(n53192), .C(
        n53628), .Y(n56807) );
  A2O1A1Ixp33_ASAP7_75t_SL U46996 ( .A1(n75616), .A2(n77873), .B(n53192), .C(
        n53628), .Y(n56797) );
  A2O1A1Ixp33_ASAP7_75t_SL U46997 ( .A1(n77855), .A2(n57073), .B(n53192), .C(
        n53628), .Y(n56796) );
  A2O1A1Ixp33_ASAP7_75t_SL U46998 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[22]), .B(n53192), 
        .C(n53628), .Y(n56623) );
  A2O1A1Ixp33_ASAP7_75t_SL U46999 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[22]), .A2(n56624), 
        .B(n53192), .C(n53628), .Y(n56625) );
  A2O1A1Ixp33_ASAP7_75t_SL U47000 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[22]), .B(
        n53192), .C(n53628), .Y(n56626) );
  A2O1A1Ixp33_ASAP7_75t_SL U47001 ( .A1(n56623), .A2(n56625), .B(n53192), .C(
        n56626), .Y(or1200_cpu_or1200_fpu_fpu_arith_N105) );
  A2O1A1Ixp33_ASAP7_75t_SL U47002 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[31]), .B(n53192), 
        .C(n53628), .Y(n56793) );
  A2O1A1Ixp33_ASAP7_75t_SL U47003 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[31]), .B(
        n53192), .C(n53628), .Y(n56794) );
  A2O1A1Ixp33_ASAP7_75t_SL U47004 ( .A1(n74817), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[31]), .B(n53192), 
        .C(n53628), .Y(n56795) );
  A2O1A1Ixp33_ASAP7_75t_SL U47005 ( .A1(n56793), .A2(n56794), .B(n53192), .C(
        n56795), .Y(or1200_cpu_or1200_fpu_fpu_arith_N114) );
  A2O1A1Ixp33_ASAP7_75t_SL U47006 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[15]), .B(n53192), 
        .C(n53628), .Y(n56617) );
  A2O1A1Ixp33_ASAP7_75t_SL U47007 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[15]), .A2(n56618), 
        .B(n53192), .C(n53628), .Y(n56619) );
  A2O1A1Ixp33_ASAP7_75t_SL U47008 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[15]), .B(
        n53192), .C(n53628), .Y(n56620) );
  A2O1A1Ixp33_ASAP7_75t_SL U47009 ( .A1(n56617), .A2(n56619), .B(n53192), .C(
        n56620), .Y(or1200_cpu_or1200_fpu_fpu_arith_N98) );
  A2O1A1Ixp33_ASAP7_75t_SL U47010 ( .A1(n59691), .A2(n56615), .B(n53192), .C(
        n53628), .Y(n56616) );
  A2O1A1Ixp33_ASAP7_75t_SL U47011 ( .A1(n77983), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56614) );
  A2O1A1Ixp33_ASAP7_75t_SL U47012 ( .A1(n76990), .A2(n56611), .B(n53192), .C(
        n53628), .Y(n56612) );
  A2O1A1Ixp33_ASAP7_75t_SL U47013 ( .A1(n59680), .A2(n77974), .B(n53192), .C(
        n53628), .Y(n56613) );
  A2O1A1Ixp33_ASAP7_75t_SL U47014 ( .A1(n77338), .A2(n77400), .B(n53192), .C(
        n53628), .Y(n56610) );
  A2O1A1Ixp33_ASAP7_75t_SL U47015 ( .A1(n77930), .A2(n59691), .B(n53192), .C(
        n53628), .Y(n56606) );
  A2O1A1Ixp33_ASAP7_75t_SL U47016 ( .A1(n69337), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n54690) );
  A2O1A1Ixp33_ASAP7_75t_SL U47017 ( .A1(n69343), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56605) );
  A2O1A1Ixp33_ASAP7_75t_SL U47018 ( .A1(n69377), .A2(n70529), .B(n53192), .C(
        n53628), .Y(n56791) );
  A2O1A1Ixp33_ASAP7_75t_SL U47019 ( .A1(n56786), .A2(n56787), .B(n53192), .C(
        n53628), .Y(n56788) );
  A2O1A1Ixp33_ASAP7_75t_SL U47020 ( .A1(n70372), .A2(n70509), .B(n53192), .C(
        n53628), .Y(n56784) );
  A2O1A1Ixp33_ASAP7_75t_SL U47021 ( .A1(n56779), .A2(n56780), .B(n53192), .C(
        n53628), .Y(n56781) );
  A2O1A1Ixp33_ASAP7_75t_SL U47022 ( .A1(n74796), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n55222) );
  A2O1A1Ixp33_ASAP7_75t_SL U47023 ( .A1(n76809), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56574) );
  A2O1A1Ixp33_ASAP7_75t_SL U47024 ( .A1(n69336), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56091) );
  A2O1A1Ixp33_ASAP7_75t_SL U47025 ( .A1(n77246), .A2(n77920), .B(n53192), .C(
        n53628), .Y(n56776) );
  A2O1A1Ixp33_ASAP7_75t_SL U47026 ( .A1(n77916), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56573) );
  A2O1A1Ixp33_ASAP7_75t_SL U47027 ( .A1(n77980), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56572) );
  A2O1A1Ixp33_ASAP7_75t_SL U47028 ( .A1(n77986), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56571) );
  A2O1A1Ixp33_ASAP7_75t_SL U47029 ( .A1(n77992), .A2(n59680), .B(n53192), .C(
        n53628), .Y(n56567) );
  A2O1A1Ixp33_ASAP7_75t_SL U47030 ( .A1(n77968), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56300) );
  A2O1A1Ixp33_ASAP7_75t_SL U47031 ( .A1(n74934), .A2(n56774), .B(n53192), .C(
        n53628), .Y(n56775) );
  A2O1A1Ixp33_ASAP7_75t_SL U47032 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_ine_o), .A2(n55656), .B(n53192), .C(
        n53628), .Y(n1531) );
  A2O1A1Ixp33_ASAP7_75t_SL U47033 ( .A1(n59578), .A2(n56771), .B(n53192), .C(
        n53628), .Y(n1506) );
  A2O1A1Ixp33_ASAP7_75t_SL U47034 ( .A1(n57114), .A2(n77977), .B(n53192), .C(
        n53628), .Y(n56770) );
  A2O1A1Ixp33_ASAP7_75t_SL U47035 ( .A1(n57114), .A2(n77859), .B(n53192), .C(
        n53628), .Y(n56769) );
  A2O1A1Ixp33_ASAP7_75t_SL U47036 ( .A1(n57114), .A2(n77856), .B(n53192), .C(
        n53628), .Y(n56768) );
  A2O1A1Ixp33_ASAP7_75t_SL U47037 ( .A1(n77901), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n55213) );
  A2O1A1Ixp33_ASAP7_75t_SL U47038 ( .A1(n74641), .A2(n77896), .B(n53192), .C(
        n53628), .Y(n56767) );
  A2O1A1Ixp33_ASAP7_75t_SL U47039 ( .A1(n77893), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n54314) );
  A2O1A1Ixp33_ASAP7_75t_SL U47040 ( .A1(n76235), .A2(n77287), .B(n53192), .C(
        n53628), .Y(n56538) );
  A2O1A1Ixp33_ASAP7_75t_SL U47041 ( .A1(n1364), .A2(n56539), .B(n53192), .C(
        n53628), .Y(n56540) );
  A2O1A1Ixp33_ASAP7_75t_SL U47042 ( .A1(n56538), .A2(n56540), .B(n53192), .C(
        n53628), .Y(n56541) );
  A2O1A1Ixp33_ASAP7_75t_SL U47043 ( .A1(n53192), .A2(n53628), .B(n56543), .C(
        n53628), .Y(or1200_pic_N63) );
  A2O1A1Ixp33_ASAP7_75t_SL U47044 ( .A1(n75302), .A2(n77287), .B(n53192), .C(
        n53628), .Y(n56532) );
  A2O1A1Ixp33_ASAP7_75t_SL U47045 ( .A1(n1360), .A2(n56533), .B(n53192), .C(
        n53628), .Y(n56534) );
  A2O1A1Ixp33_ASAP7_75t_SL U47046 ( .A1(n56532), .A2(n56534), .B(n53192), .C(
        n53628), .Y(n56535) );
  A2O1A1Ixp33_ASAP7_75t_SL U47047 ( .A1(n53192), .A2(n53628), .B(n56537), .C(
        n53628), .Y(or1200_pic_N64) );
  A2O1A1Ixp33_ASAP7_75t_SL U47048 ( .A1(n56528), .A2(n56530), .B(n53192), .C(
        n53628), .Y(n9348) );
  A2O1A1Ixp33_ASAP7_75t_SL U47049 ( .A1(n56525), .A2(n56527), .B(n53192), .C(
        n53628), .Y(n9351) );
  A2O1A1Ixp33_ASAP7_75t_SL U47050 ( .A1(n56522), .A2(n56524), .B(n53192), .C(
        n53628), .Y(n9349) );
  A2O1A1Ixp33_ASAP7_75t_SL U47051 ( .A1(n77615), .A2(n77287), .B(n53192), .C(
        n53628), .Y(n55846) );
  A2O1A1Ixp33_ASAP7_75t_SL U47052 ( .A1(n1115), .A2(n55847), .B(n53192), .C(
        n53628), .Y(n55848) );
  A2O1A1Ixp33_ASAP7_75t_SL U47053 ( .A1(n55846), .A2(n55848), .B(n53192), .C(
        n53628), .Y(n55849) );
  A2O1A1Ixp33_ASAP7_75t_SL U47054 ( .A1(n53192), .A2(n53628), .B(n55851), .C(
        n53628), .Y(or1200_pic_N58) );
  A2O1A1Ixp33_ASAP7_75t_SL U47055 ( .A1(n56750), .A2(n56751), .B(n53192), .C(
        n53628), .Y(n56752) );
  A2O1A1Ixp33_ASAP7_75t_SL U47056 ( .A1(n64095), .A2(n56512), .B(n53192), .C(
        n53628), .Y(n56513) );
  A2O1A1Ixp33_ASAP7_75t_SL U47057 ( .A1(n76224), .A2(n76226), .B(n53192), .C(
        n53628), .Y(n56509) );
  A2O1A1Ixp33_ASAP7_75t_SL U47058 ( .A1(n56508), .A2(n57245), .B(n53192), .C(
        n56509), .Y(n56510) );
  A2O1A1Ixp33_ASAP7_75t_SL U47059 ( .A1(n76631), .A2(n56496), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1106) );
  A2O1A1Ixp33_ASAP7_75t_SL U47060 ( .A1(n65161), .A2(n56735), .B(n53192), .C(
        n53628), .Y(n56736) );
  A2O1A1Ixp33_ASAP7_75t_SL U47061 ( .A1(n69126), .A2(n75650), .B(n53192), .C(
        n53628), .Y(n54626) );
  A2O1A1Ixp33_ASAP7_75t_SL U47062 ( .A1(n69168), .A2(n54628), .B(n53192), .C(
        n53628), .Y(n54629) );
  A2O1A1Ixp33_ASAP7_75t_SL U47063 ( .A1(n54631), .A2(n54632), .B(n53192), .C(
        n53628), .Y(n54633) );
  A2O1A1Ixp33_ASAP7_75t_SL U47064 ( .A1(n59673), .A2(n77899), .B(n53192), .C(
        n53628), .Y(n54635) );
  A2O1A1Ixp33_ASAP7_75t_SL U47065 ( .A1(n54626), .A2(n54634), .B(n53192), .C(
        n54635), .Y(or1200_cpu_or1200_mult_mac_n1611) );
  A2O1A1Ixp33_ASAP7_75t_SL U47066 ( .A1(n75650), .A2(n69188), .B(n53192), .C(
        n53628), .Y(n56727) );
  A2O1A1Ixp33_ASAP7_75t_SL U47067 ( .A1(n77885), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n56728) );
  A2O1A1Ixp33_ASAP7_75t_SL U47068 ( .A1(n56727), .A2(n56728), .B(n53192), .C(
        n53628), .Y(n56729) );
  A2O1A1Ixp33_ASAP7_75t_SL U47069 ( .A1(n62011), .A2(
        or1200_cpu_or1200_mult_mac_n285), .B(n53192), .C(n62025), .Y(n56724)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U47070 ( .A1(n65402), .A2(n56723), .B(n53192), .C(
        n53628), .Y(n1598) );
  A2O1A1Ixp33_ASAP7_75t_SL U47071 ( .A1(n76680), .A2(n59688), .B(n53192), .C(
        n53628), .Y(n56485) );
  A2O1A1Ixp33_ASAP7_75t_SL U47072 ( .A1(n76858), .A2(n59689), .B(n53192), .C(
        n53628), .Y(n56484) );
  A2O1A1Ixp33_ASAP7_75t_SL U47073 ( .A1(n76997), .A2(n57074), .B(n53192), .C(
        n53628), .Y(n56483) );
  A2O1A1Ixp33_ASAP7_75t_SL U47074 ( .A1(n76210), .A2(n59689), .B(n53192), .C(
        n53628), .Y(n56482) );
  A2O1A1Ixp33_ASAP7_75t_SL U47075 ( .A1(n76617), .A2(n59694), .B(n53192), .C(
        n53628), .Y(n56481) );
  A2O1A1Ixp33_ASAP7_75t_SL U47076 ( .A1(n76700), .A2(n59690), .B(n53192), .C(
        n53628), .Y(n56480) );
  A2O1A1Ixp33_ASAP7_75t_SL U47077 ( .A1(n76643), .A2(n59690), .B(n53192), .C(
        n53628), .Y(n56479) );
  A2O1A1Ixp33_ASAP7_75t_SL U47078 ( .A1(n76249), .A2(n59688), .B(n53192), .C(
        n53628), .Y(n56478) );
  A2O1A1Ixp33_ASAP7_75t_SL U47079 ( .A1(n75780), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56477) );
  A2O1A1Ixp33_ASAP7_75t_SL U47080 ( .A1(n76551), .A2(n59689), .B(n53192), .C(
        n53628), .Y(n56476) );
  A2O1A1Ixp33_ASAP7_75t_SL U47081 ( .A1(n77291), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56475) );
  A2O1A1Ixp33_ASAP7_75t_SL U47082 ( .A1(n77224), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56474) );
  A2O1A1Ixp33_ASAP7_75t_SL U47083 ( .A1(n77018), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56473) );
  A2O1A1Ixp33_ASAP7_75t_SL U47084 ( .A1(n77151), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56472) );
  A2O1A1Ixp33_ASAP7_75t_SL U47085 ( .A1(n76230), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56471) );
  A2O1A1Ixp33_ASAP7_75t_SL U47086 ( .A1(n75301), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56470) );
  A2O1A1Ixp33_ASAP7_75t_SL U47087 ( .A1(n74983), .A2(n59689), .B(n53192), .C(
        n53628), .Y(n56469) );
  A2O1A1Ixp33_ASAP7_75t_SL U47088 ( .A1(n74576), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56468) );
  A2O1A1Ixp33_ASAP7_75t_SL U47089 ( .A1(n59693), .A2(n74126), .B(n53192), .C(
        n53628), .Y(n56722) );
  A2O1A1Ixp33_ASAP7_75t_SL U47090 ( .A1(n75430), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56467) );
  A2O1A1Ixp33_ASAP7_75t_SL U47091 ( .A1(n59693), .A2(n75446), .B(n53192), .C(
        n53628), .Y(n56721) );
  A2O1A1Ixp33_ASAP7_75t_SL U47092 ( .A1(n75619), .A2(n59689), .B(n53192), .C(
        n53628), .Y(n56466) );
  A2O1A1Ixp33_ASAP7_75t_SL U47093 ( .A1(n59693), .A2(n74044), .B(n53192), .C(
        n53628), .Y(n56720) );
  A2O1A1Ixp33_ASAP7_75t_SL U47094 ( .A1(n74083), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56465) );
  A2O1A1Ixp33_ASAP7_75t_SL U47095 ( .A1(n59693), .A2(n69367), .B(n53192), .C(
        n53628), .Y(n56719) );
  A2O1A1Ixp33_ASAP7_75t_SL U47096 ( .A1(n75795), .A2(n59689), .B(n53192), .C(
        n53628), .Y(n56464) );
  A2O1A1Ixp33_ASAP7_75t_SL U47097 ( .A1(n75197), .A2(n59688), .B(n53192), .C(
        n53628), .Y(n56462) );
  A2O1A1Ixp33_ASAP7_75t_SL U47098 ( .A1(n75674), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56461) );
  A2O1A1Ixp33_ASAP7_75t_SL U47099 ( .A1(n76922), .A2(n59690), .B(n53192), .C(
        n53628), .Y(n56460) );
  A2O1A1Ixp33_ASAP7_75t_SL U47100 ( .A1(n56445), .A2(n56446), .B(n53192), .C(
        n53628), .Y(n56447) );
  A2O1A1Ixp33_ASAP7_75t_SL U47101 ( .A1(n56444), .A2(n56447), .B(n53192), .C(
        n53628), .Y(n56448) );
  A2O1A1Ixp33_ASAP7_75t_SL U47102 ( .A1(n71627), .A2(n72163), .B(n53192), .C(
        n53628), .Y(n56437) );
  A2O1A1Ixp33_ASAP7_75t_SL U47103 ( .A1(n71628), .A2(n56440), .B(n53192), .C(
        n53628), .Y(n56441) );
  A2O1A1Ixp33_ASAP7_75t_SL U47104 ( .A1(n71186), .A2(n78421), .B(n53192), .C(
        n53628), .Y(n56716) );
  A2O1A1Ixp33_ASAP7_75t_SL U47105 ( .A1(n59611), .A2(n67736), .B(n53192), .C(
        n53628), .Y(n56714) );
  A2O1A1Ixp33_ASAP7_75t_SL U47106 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[12]), .A2(n59632), .B(
        n53192), .C(n53628), .Y(n56709) );
  A2O1A1Ixp33_ASAP7_75t_SL U47107 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]), .A2(n57204), .B(
        n53192), .C(n53628), .Y(n56710) );
  A2O1A1Ixp33_ASAP7_75t_SL U47108 ( .A1(n56709), .A2(n56710), .B(n53192), .C(
        n53628), .Y(n56711) );
  A2O1A1Ixp33_ASAP7_75t_SL U47109 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[14]), .A2(n57205), .B(
        n53192), .C(n53628), .Y(n56713) );
  A2O1A1Ixp33_ASAP7_75t_SL U47110 ( .A1(n56712), .A2(n56713), .B(n53192), .C(
        n53628), .Y(n73765) );
  A2O1A1Ixp33_ASAP7_75t_SL U47111 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[4]), .A2(n70038), .B(n53192), .C(n53628), .Y(n56706) );
  A2O1A1Ixp33_ASAP7_75t_SL U47112 ( .A1(n56705), .A2(n56706), .B(n53192), .C(
        n53628), .Y(n56707) );
  A2O1A1Ixp33_ASAP7_75t_SL U47113 ( .A1(n3376), .A2(n56701), .B(n53192), .C(
        n53628), .Y(n61282) );
  A2O1A1Ixp33_ASAP7_75t_SL U47114 ( .A1(n62004), .A2(n62003), .B(n53192), .C(
        n56700), .Y(n62005) );
  A2O1A1Ixp33_ASAP7_75t_SL U47115 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n70301), .B(n53192), .C(n53628), .Y(n56697) );
  A2O1A1Ixp33_ASAP7_75t_SL U47116 ( .A1(n69783), .A2(n56224), .B(n53192), .C(
        n53628), .Y(n69774) );
  A2O1A1Ixp33_ASAP7_75t_SL U47117 ( .A1(n69835), .A2(n55321), .B(n53192), .C(
        n53628), .Y(n69818) );
  A2O1A1Ixp33_ASAP7_75t_SL U47118 ( .A1(n70005), .A2(n56696), .B(n53192), .C(
        n53628), .Y(n70013) );
  A2O1A1Ixp33_ASAP7_75t_SL U47119 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_4_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_3_), .B(n53192), .C(n53628), 
        .Y(n56219) );
  A2O1A1Ixp33_ASAP7_75t_SL U47120 ( .A1(n62059), .A2(n56222), .B(n53192), .C(
        n53628), .Y(n62063) );
  A2O1A1Ixp33_ASAP7_75t_SL U47121 ( .A1(n77017), .A2(n77015), .B(n53192), .C(
        n56694), .Y(n56695) );
  A2O1A1Ixp33_ASAP7_75t_SL U47122 ( .A1(n75194), .A2(n56214), .B(n53192), .C(
        n53628), .Y(n56215) );
  A2O1A1Ixp33_ASAP7_75t_SL U47123 ( .A1(n75395), .A2(n75398), .B(n53192), .C(
        n53628), .Y(n56693) );
  A2O1A1Ixp33_ASAP7_75t_SL U47124 ( .A1(n74111), .A2(n56689), .B(n53192), .C(
        n53628), .Y(n58546) );
  A2O1A1Ixp33_ASAP7_75t_SL U47125 ( .A1(n74993), .A2(n55761), .B(n53192), .C(
        n53628), .Y(n75789) );
  A2O1A1Ixp33_ASAP7_75t_SL U47126 ( .A1(n76109), .A2(n56204), .B(n53192), .C(
        n53628), .Y(n76099) );
  A2O1A1Ixp33_ASAP7_75t_SL U47127 ( .A1(n76014), .A2(n56687), .B(n53192), .C(
        n53628), .Y(n76018) );
  A2O1A1Ixp33_ASAP7_75t_SL U47128 ( .A1(n63301), .A2(n56685), .B(n53192), .C(
        n53628), .Y(n63283) );
  A2O1A1Ixp33_ASAP7_75t_SL U47129 ( .A1(n63542), .A2(n56411), .B(n53192), .C(
        n53628), .Y(n63468) );
  A2O1A1Ixp33_ASAP7_75t_SL U47130 ( .A1(n65091), .A2(n55755), .B(n53192), .C(
        n53628), .Y(n65073) );
  A2O1A1Ixp33_ASAP7_75t_SL U47131 ( .A1(or1200_cpu_or1200_mult_mac_n339), .A2(
        n56682), .B(n53192), .C(n53628), .Y(n68790) );
  A2O1A1Ixp33_ASAP7_75t_SL U47132 ( .A1(n68986), .A2(n56408), .B(n53192), .C(
        n53628), .Y(n68951) );
  A2O1A1Ixp33_ASAP7_75t_SL U47133 ( .A1(n77704), .A2(n57500), .B(n53192), .C(
        n53628), .Y(n56677) );
  A2O1A1Ixp33_ASAP7_75t_SL U47134 ( .A1(n72564), .A2(n72576), .B(n53192), .C(
        n53628), .Y(n56401) );
  A2O1A1Ixp33_ASAP7_75t_SL U47135 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_0_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39), .B(n53192), .C(n53628), .Y(n56402) );
  A2O1A1Ixp33_ASAP7_75t_SL U47136 ( .A1(n74493), .A2(n56401), .B(n53192), .C(
        n56402), .Y(n74100) );
  A2O1A1Ixp33_ASAP7_75t_SL U47137 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n56672) );
  A2O1A1Ixp33_ASAP7_75t_SL U47138 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n56673) );
  A2O1A1Ixp33_ASAP7_75t_SL U47139 ( .A1(n56672), .A2(n56673), .B(n53192), .C(
        n53628), .Y(n56674) );
  A2O1A1Ixp33_ASAP7_75t_SL U47140 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n56676) );
  A2O1A1Ixp33_ASAP7_75t_SL U47141 ( .A1(n56675), .A2(n56676), .B(n53192), .C(
        n53628), .Y(n71913) );
  A2O1A1Ixp33_ASAP7_75t_SL U47142 ( .A1(n71790), .A2(n71728), .B(n53192), .C(
        n53628), .Y(n56670) );
  A2O1A1Ixp33_ASAP7_75t_SL U47143 ( .A1(n71505), .A2(n56669), .B(n53192), .C(
        n53628), .Y(n71480) );
  A2O1A1Ixp33_ASAP7_75t_SL U47144 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_38_), .A2(n55742), 
        .B(n53192), .C(n53628), .Y(n71255) );
  A2O1A1Ixp33_ASAP7_75t_SL U47145 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[38]), .A2(n59562), 
        .B(n53192), .C(n53628), .Y(n55741) );
  A2O1A1Ixp33_ASAP7_75t_SL U47146 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[20]), .A2(
        n59631), .B(n53192), .C(n53628), .Y(n56387) );
  A2O1A1Ixp33_ASAP7_75t_SL U47147 ( .A1(n69394), .A2(n56664), .B(n53192), .C(
        n53628), .Y(n69426) );
  A2O1A1Ixp33_ASAP7_75t_SL U47148 ( .A1(n62682), .A2(n64217), .B(n53192), .C(
        n53628), .Y(n56663) );
  A2O1A1Ixp33_ASAP7_75t_SL U47149 ( .A1(n75358), .A2(n56663), .B(n53192), .C(
        n53628), .Y(n74626) );
  A2O1A1Ixp33_ASAP7_75t_SL U47150 ( .A1(n2141), .A2(n76772), .B(n53192), .C(
        n53628), .Y(n56662) );
  A2O1A1Ixp33_ASAP7_75t_SL U47151 ( .A1(n64230), .A2(n56662), .B(n53192), .C(
        n53628), .Y(n62445) );
  A2O1A1Ixp33_ASAP7_75t_SL U47152 ( .A1(n77696), .A2(n75847), .B(n53192), .C(
        n53628), .Y(n56660) );
  A2O1A1Ixp33_ASAP7_75t_SL U47153 ( .A1(n69036), .A2(n69035), .B(n53192), .C(
        n53628), .Y(n56657) );
  A2O1A1Ixp33_ASAP7_75t_SL U47154 ( .A1(n57414), .A2(n56655), .B(n53192), .C(
        n53628), .Y(n57675) );
  A2O1A1Ixp33_ASAP7_75t_SL U47155 ( .A1(n74008), .A2(n55940), .B(n53192), .C(
        n53628), .Y(n76396) );
  A2O1A1Ixp33_ASAP7_75t_SL U47156 ( .A1(n57394), .A2(n57108), .B(n53192), .C(
        n53628), .Y(n56146) );
  A2O1A1Ixp33_ASAP7_75t_SL U47157 ( .A1(n60782), .A2(n60783), .B(n53192), .C(
        n53628), .Y(n56653) );
  A2O1A1Ixp33_ASAP7_75t_SL U47158 ( .A1(n59570), .A2(n56653), .B(n53192), .C(
        n53628), .Y(n61955) );
  A2O1A1Ixp33_ASAP7_75t_SL U47159 ( .A1(n73661), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56644) );
  A2O1A1Ixp33_ASAP7_75t_SL U47160 ( .A1(n73580), .A2(n56644), .B(n53192), .C(
        n53628), .Y(n56645) );
  A2O1A1Ixp33_ASAP7_75t_SL U47161 ( .A1(n73660), .A2(n56645), .B(n53192), .C(
        n53628), .Y(n3280) );
  A2O1A1Ixp33_ASAP7_75t_SL U47162 ( .A1(n61040), .A2(n60447), .B(n53192), .C(
        n53628), .Y(n56638) );
  A2O1A1Ixp33_ASAP7_75t_SL U47163 ( .A1(n56639), .A2(n60446), .B(n53192), .C(
        n53628), .Y(n56640) );
  A2O1A1Ixp33_ASAP7_75t_SL U47164 ( .A1(n53628), .A2(n56636), .B(n53192), .C(
        n53628), .Y(n56637) );
  A2O1A1Ixp33_ASAP7_75t_SL U47165 ( .A1(n57144), .A2(n64013), .B(n53192), .C(
        n53628), .Y(n56337) );
  A2O1A1Ixp33_ASAP7_75t_SL U47166 ( .A1(n59694), .A2(n56627), .B(n53192), .C(
        n53628), .Y(n56628) );
  A2O1A1Ixp33_ASAP7_75t_SL U47167 ( .A1(n53192), .A2(n53628), .B(n55472), .C(
        n53628), .Y(n55473) );
  A2O1A1Ixp33_ASAP7_75t_SL U47168 ( .A1(n78341), .A2(n73047), .B(n53192), .C(
        n53628), .Y(n56118) );
  A2O1A1Ixp33_ASAP7_75t_SL U47169 ( .A1(n77971), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56324) );
  A2O1A1Ixp33_ASAP7_75t_SL U47170 ( .A1(n61158), .A2(n56607), .B(n53192), .C(
        n56608), .Y(n56609) );
  A2O1A1Ixp33_ASAP7_75t_SL U47171 ( .A1(n70546), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .B(
        n53192), .C(n53628), .Y(n56596) );
  A2O1A1Ixp33_ASAP7_75t_SL U47172 ( .A1(n74685), .A2(n70542), .B(n53192), .C(
        n53628), .Y(n56599) );
  A2O1A1Ixp33_ASAP7_75t_SL U47173 ( .A1(n70543), .A2(n74681), .B(n53192), .C(
        n53628), .Y(n56600) );
  A2O1A1Ixp33_ASAP7_75t_SL U47174 ( .A1(n56598), .A2(n56599), .B(n53192), .C(
        n56600), .Y(n56601) );
  A2O1A1Ixp33_ASAP7_75t_SL U47175 ( .A1(n70545), .A2(n56602), .B(n53192), .C(
        n53628), .Y(n56603) );
  A2O1A1Ixp33_ASAP7_75t_SL U47176 ( .A1(n56575), .A2(n56576), .B(n53192), .C(
        n53628), .Y(n56577) );
  A2O1A1Ixp33_ASAP7_75t_SL U47177 ( .A1(n56577), .A2(n56579), .B(n53192), .C(
        n53628), .Y(n2303) );
  A2O1A1Ixp33_ASAP7_75t_SL U47178 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_5_), .A2(n56097), .B(n53192), 
        .C(n53628), .Y(n56098) );
  A2O1A1Ixp33_ASAP7_75t_SL U47179 ( .A1(n75533), .A2(n57198), .B(n53192), .C(
        n53628), .Y(n56568) );
  A2O1A1Ixp33_ASAP7_75t_SL U47180 ( .A1(n77899), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56298) );
  A2O1A1Ixp33_ASAP7_75t_SL U47181 ( .A1(n77922), .A2(n59680), .B(n53192), .C(
        n53628), .Y(n56083) );
  A2O1A1Ixp33_ASAP7_75t_SL U47182 ( .A1(n77613), .A2(n77644), .B(n53192), .C(
        n53628), .Y(n56564) );
  A2O1A1Ixp33_ASAP7_75t_SL U47183 ( .A1(n77968), .A2(n77672), .B(n53192), .C(
        n53628), .Y(n56565) );
  A2O1A1Ixp33_ASAP7_75t_SL U47184 ( .A1(n56564), .A2(n56565), .B(n53192), .C(
        n53628), .Y(n56566) );
  A2O1A1Ixp33_ASAP7_75t_SL U47185 ( .A1(n59629), .A2(n78356), .B(n53192), .C(
        n53628), .Y(n56558) );
  A2O1A1Ixp33_ASAP7_75t_SL U47186 ( .A1(n57114), .A2(n77920), .B(n53192), .C(
        n53628), .Y(n56556) );
  A2O1A1Ixp33_ASAP7_75t_SL U47187 ( .A1(n57114), .A2(n77854), .B(n53192), .C(
        n53628), .Y(n56555) );
  A2O1A1Ixp33_ASAP7_75t_SL U47188 ( .A1(n74641), .A2(n77918), .B(n53192), .C(
        n53628), .Y(n56554) );
  A2O1A1Ixp33_ASAP7_75t_SL U47189 ( .A1(n1406), .A2(n56549), .B(n53192), .C(
        n53628), .Y(n56550) );
  A2O1A1Ixp33_ASAP7_75t_SL U47190 ( .A1(n77287), .A2(n77597), .B(n53192), .C(
        n53628), .Y(n56551) );
  A2O1A1Ixp33_ASAP7_75t_SL U47191 ( .A1(n56550), .A2(n56551), .B(n53192), .C(
        n53628), .Y(n56552) );
  A2O1A1Ixp33_ASAP7_75t_SL U47192 ( .A1(n56552), .A2(n56553), .B(n53192), .C(
        n53628), .Y(or1200_pic_N52) );
  A2O1A1Ixp33_ASAP7_75t_SL U47193 ( .A1(n1372), .A2(n56544), .B(n53192), .C(
        n53628), .Y(n56545) );
  A2O1A1Ixp33_ASAP7_75t_SL U47194 ( .A1(n77287), .A2(n77019), .B(n53192), .C(
        n53628), .Y(n56546) );
  A2O1A1Ixp33_ASAP7_75t_SL U47195 ( .A1(n56545), .A2(n56546), .B(n53192), .C(
        n53628), .Y(n56547) );
  A2O1A1Ixp33_ASAP7_75t_SL U47196 ( .A1(n56547), .A2(n56548), .B(n53192), .C(
        n53628), .Y(or1200_pic_N61) );
  A2O1A1Ixp33_ASAP7_75t_SL U47197 ( .A1(n74641), .A2(n77885), .B(n53192), .C(
        n53628), .Y(n56531) );
  A2O1A1Ixp33_ASAP7_75t_SL U47198 ( .A1(n57142), .A2(n77972), .B(n53192), .C(
        n53628), .Y(n56528) );
  A2O1A1Ixp33_ASAP7_75t_SL U47199 ( .A1(n77973), .A2(n56529), .B(n53192), .C(
        n53628), .Y(n56530) );
  A2O1A1Ixp33_ASAP7_75t_SL U47200 ( .A1(n57142), .A2(n77989), .B(n53192), .C(
        n53628), .Y(n56525) );
  A2O1A1Ixp33_ASAP7_75t_SL U47201 ( .A1(n77987), .A2(n56526), .B(n53192), .C(
        n53628), .Y(n56527) );
  A2O1A1Ixp33_ASAP7_75t_SL U47202 ( .A1(n57142), .A2(n77969), .B(n53192), .C(
        n53628), .Y(n56522) );
  A2O1A1Ixp33_ASAP7_75t_SL U47203 ( .A1(n77970), .A2(n56523), .B(n53192), .C(
        n53628), .Y(n56524) );
  A2O1A1Ixp33_ASAP7_75t_SL U47204 ( .A1(n63370), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56504) );
  A2O1A1Ixp33_ASAP7_75t_SL U47205 ( .A1(n63366), .A2(n56504), .B(n53192), .C(
        n53628), .Y(n56505) );
  A2O1A1Ixp33_ASAP7_75t_SL U47206 ( .A1(n56503), .A2(n56505), .B(n53192), .C(
        n53628), .Y(n56506) );
  A2O1A1Ixp33_ASAP7_75t_SL U47207 ( .A1(n63364), .A2(n57044), .B(n53192), .C(
        n56506), .Y(n56507) );
  A2O1A1Ixp33_ASAP7_75t_SL U47208 ( .A1(n56063), .A2(n56064), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N5) );
  A2O1A1Ixp33_ASAP7_75t_SL U47209 ( .A1(n65145), .A2(n56490), .B(n53192), .C(
        n53628), .Y(n56491) );
  A2O1A1Ixp33_ASAP7_75t_SL U47210 ( .A1(n56488), .A2(n56495), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1571) );
  A2O1A1Ixp33_ASAP7_75t_SL U47211 ( .A1(n75650), .A2(n77042), .B(n53192), .C(
        n53628), .Y(n55813) );
  A2O1A1Ixp33_ASAP7_75t_SL U47212 ( .A1(n77893), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n55814) );
  A2O1A1Ixp33_ASAP7_75t_SL U47213 ( .A1(n55827), .A2(n55828), .B(n53192), .C(
        n53628), .Y(n55829) );
  A2O1A1Ixp33_ASAP7_75t_SL U47214 ( .A1(n55813), .A2(n55814), .B(n53192), .C(
        n55830), .Y(or1200_cpu_or1200_mult_mac_n1609) );
  A2O1A1Ixp33_ASAP7_75t_SL U47215 ( .A1(n59673), .A2(n77862), .B(n53192), .C(
        n53628), .Y(n55809) );
  A2O1A1Ixp33_ASAP7_75t_SL U47216 ( .A1(n55811), .A2(n55812), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1596) );
  A2O1A1Ixp33_ASAP7_75t_SL U47217 ( .A1(or1200_cpu_or1200_except_n290), .A2(
        n77438), .B(n53192), .C(n77440), .Y(n56486) );
  A2O1A1Ixp33_ASAP7_75t_SL U47218 ( .A1(n59693), .A2(n77176), .B(n53192), .C(
        n53628), .Y(n56463) );
  A2O1A1Ixp33_ASAP7_75t_SL U47219 ( .A1(n74129), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56241) );
  A2O1A1Ixp33_ASAP7_75t_SL U47220 ( .A1(n59693), .A2(n74047), .B(n53192), .C(
        n53628), .Y(n56459) );
  A2O1A1Ixp33_ASAP7_75t_SL U47221 ( .A1(n69373), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56027) );
  A2O1A1Ixp33_ASAP7_75t_SL U47222 ( .A1(n76671), .A2(n58146), .B(n53192), .C(
        n53628), .Y(n56458) );
  A2O1A1Ixp33_ASAP7_75t_SL U47223 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_25_), .A2(
        n53628), .B(n53192), .C(n53628), .Y(n56456) );
  A2O1A1Ixp33_ASAP7_75t_SL U47224 ( .A1(n74332), .A2(n56456), .B(n53192), .C(
        n53628), .Y(n56457) );
  A2O1A1Ixp33_ASAP7_75t_SL U47225 ( .A1(n74343), .A2(n56457), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n6) );
  A2O1A1Ixp33_ASAP7_75t_SL U47226 ( .A1(n72367), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_1_), 
        .B(n53192), .C(n53628), .Y(n56444) );
  A2O1A1Ixp33_ASAP7_75t_SL U47227 ( .A1(n59527), .A2(n72366), .B(n53192), .C(
        n53628), .Y(n56445) );
  A2O1A1Ixp33_ASAP7_75t_SL U47228 ( .A1(n72365), .A2(n72364), .B(n53192), .C(
        n53628), .Y(n56446) );
  A2O1A1Ixp33_ASAP7_75t_SL U47229 ( .A1(n71629), .A2(n56438), .B(n53192), .C(
        n53628), .Y(n56439) );
  A2O1A1Ixp33_ASAP7_75t_SL U47230 ( .A1(n53628), .A2(n56439), .B(n53192), .C(
        n53628), .Y(n56440) );
  A2O1A1Ixp33_ASAP7_75t_SL U47231 ( .A1(n66082), .A2(n56433), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n32) );
  A2O1A1Ixp33_ASAP7_75t_SL U47232 ( .A1(or1200_cpu_or1200_mult_mac_n30), .A2(
        n55996), .B(n53192), .C(n53628), .Y(n76109) );
  A2O1A1Ixp33_ASAP7_75t_SL U47233 ( .A1(or1200_cpu_or1200_mult_mac_n30), .A2(
        n55996), .B(n53192), .C(n53628), .Y(n53468) );
  A2O1A1Ixp33_ASAP7_75t_SL U47234 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[19]), .A2(n73641), .B(
        n53192), .C(n53628), .Y(n56429) );
  A2O1A1Ixp33_ASAP7_75t_SL U47235 ( .A1(n73642), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[1]), .B(
        n53192), .C(n53628), .Y(n56430) );
  A2O1A1Ixp33_ASAP7_75t_SL U47236 ( .A1(n58400), .A2(n56429), .B(n53192), .C(
        n56430), .Y(n56431) );
  A2O1A1Ixp33_ASAP7_75t_SL U47237 ( .A1(n57204), .A2(n73687), .B(n53192), .C(
        n53628), .Y(n56432) );
  A2O1A1Ixp33_ASAP7_75t_SL U47238 ( .A1(n56425), .A2(n56426), .B(n53192), .C(
        n53628), .Y(n56427) );
  A2O1A1Ixp33_ASAP7_75t_SL U47239 ( .A1(n70138), .A2(n56427), .B(n53192), .C(
        n53628), .Y(n70141) );
  A2O1A1Ixp33_ASAP7_75t_SL U47240 ( .A1(n70138), .A2(n56427), .B(n53192), .C(
        n53628), .Y(n53434) );
  A2O1A1Ixp33_ASAP7_75t_SL U47241 ( .A1(n61281), .A2(n56424), .B(n53192), .C(
        n53628), .Y(n61283) );
  A2O1A1Ixp33_ASAP7_75t_SL U47242 ( .A1(n69963), .A2(n56423), .B(n53192), .C(
        n53628), .Y(n69934) );
  A2O1A1Ixp33_ASAP7_75t_SL U47243 ( .A1(n65338), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56420) );
  A2O1A1Ixp33_ASAP7_75t_SL U47244 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_3_), .A2(n56420), .B(
        n53192), .C(n53628), .Y(n56421) );
  A2O1A1Ixp33_ASAP7_75t_SL U47245 ( .A1(n65394), .A2(n56421), .B(n53192), .C(
        n53628), .Y(n65399) );
  A2O1A1Ixp33_ASAP7_75t_SL U47246 ( .A1(n55988), .A2(n77147), .B(n53192), .C(
        n53628), .Y(n55989) );
  A2O1A1Ixp33_ASAP7_75t_SL U47247 ( .A1(n54249), .A2(n54250), .B(n53192), .C(
        n53628), .Y(n78072) );
  A2O1A1Ixp33_ASAP7_75t_SL U47248 ( .A1(n75471), .A2(n56415), .B(n53192), .C(
        n53628), .Y(n75472) );
  A2O1A1Ixp33_ASAP7_75t_SL U47249 ( .A1(n63342), .A2(n56412), .B(n53192), .C(
        n53628), .Y(n63316) );
  A2O1A1Ixp33_ASAP7_75t_SL U47250 ( .A1(n69252), .A2(n56405), .B(n53192), .C(
        n53628), .Y(n74116) );
  A2O1A1Ixp33_ASAP7_75t_SL U47251 ( .A1(n71452), .A2(n56400), .B(n53192), .C(
        n53628), .Y(n71487) );
  A2O1A1Ixp33_ASAP7_75t_SL U47252 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .A2(n65621), 
        .B(n53192), .C(n53628), .Y(n53680) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47253 ( .A1(n67268), .A2(n75947), .B(n53192), 
        .C(n56827), .D(n56391), .Y(n56392) );
  A2O1A1Ixp33_ASAP7_75t_SL U47254 ( .A1(n65028), .A2(n65029), .B(n53192), .C(
        n53628), .Y(n56389) );
  A2O1A1Ixp33_ASAP7_75t_SL U47255 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[12]), .A2(
        n59630), .B(n53192), .C(n53628), .Y(n56163) );
  A2O1A1Ixp33_ASAP7_75t_SL U47256 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[14]), .A2(
        n59631), .B(n53192), .C(n53628), .Y(n55958) );
  A2O1A1Ixp33_ASAP7_75t_SL U47257 ( .A1(n75737), .A2(n56385), .B(n53192), .C(
        n53628), .Y(n75739) );
  A2O1A1Ixp33_ASAP7_75t_SL U47258 ( .A1(n73970), .A2(n73980), .B(n53192), .C(
        n53628), .Y(n56383) );
  A2O1A1Ixp33_ASAP7_75t_SL U47259 ( .A1(n75390), .A2(n75386), .B(n53192), .C(
        n56381), .Y(n66224) );
  A2O1A1Ixp33_ASAP7_75t_SL U47260 ( .A1(n57194), .A2(n65821), .B(n53192), .C(
        n53628), .Y(n56371) );
  A2O1A1Ixp33_ASAP7_75t_SL U47261 ( .A1(n65822), .A2(n57193), .B(n53192), .C(
        n53628), .Y(n56372) );
  A2O1A1Ixp33_ASAP7_75t_SL U47262 ( .A1(n56371), .A2(n56372), .B(n53192), .C(
        n53628), .Y(n56373) );
  A2O1A1Ixp33_ASAP7_75t_SL U47263 ( .A1(n57188), .A2(n65824), .B(n53192), .C(
        n53628), .Y(n56375) );
  A2O1A1Ixp33_ASAP7_75t_SL U47264 ( .A1(n56374), .A2(n56375), .B(n53192), .C(
        n53628), .Y(n65939) );
  A2O1A1Ixp33_ASAP7_75t_SL U47265 ( .A1(n57736), .A2(n66987), .B(n53192), .C(
        n53628), .Y(n56363) );
  A2O1A1Ixp33_ASAP7_75t_SL U47266 ( .A1(n59648), .A2(n57180), .B(n53192), .C(
        n53628), .Y(n56362) );
  A2O1A1Ixp33_ASAP7_75t_SL U47267 ( .A1(n67964), .A2(n67963), .B(n53192), .C(
        n53628), .Y(n56361) );
  A2O1A1Ixp33_ASAP7_75t_SL U47268 ( .A1(n66374), .A2(n56360), .B(n53192), .C(
        n53628), .Y(n66387) );
  A2O1A1Ixp33_ASAP7_75t_SL U47269 ( .A1(n72677), .A2(n56137), .B(n53192), .C(
        n53628), .Y(n56138) );
  A2O1A1Ixp33_ASAP7_75t_SL U47270 ( .A1(n56138), .A2(n72678), .B(n53192), .C(
        n53628), .Y(n56139) );
  A2O1A1Ixp33_ASAP7_75t_SL U47271 ( .A1(n71526), .A2(n56357), .B(n53192), .C(
        n53628), .Y(n56358) );
  A2O1A1Ixp33_ASAP7_75t_SL U47272 ( .A1(n56356), .A2(n56358), .B(n53192), .C(
        n53628), .Y(n12871) );
  A2O1A1Ixp33_ASAP7_75t_SL U47273 ( .A1(n69877), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56352) );
  A2O1A1Ixp33_ASAP7_75t_SL U47274 ( .A1(n69904), .A2(n56352), .B(n53192), .C(
        n53628), .Y(n56353) );
  A2O1A1Ixp33_ASAP7_75t_SL U47275 ( .A1(n56353), .A2(n56355), .B(n53192), .C(
        n53628), .Y(n3217) );
  A2O1A1Ixp33_ASAP7_75t_SL U47276 ( .A1(n70575), .A2(n70574), .B(n53192), .C(
        n56127), .Y(n56128) );
  A2O1A1Ixp33_ASAP7_75t_SL U47277 ( .A1(n70575), .A2(n70574), .B(n53192), .C(
        n53628), .Y(n56129) );
  A2O1A1Ixp33_ASAP7_75t_SL U47278 ( .A1(n56129), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[1]), .B(
        n53192), .C(n53628), .Y(n56130) );
  A2O1A1Ixp33_ASAP7_75t_SL U47279 ( .A1(n56128), .A2(n56130), .B(n53192), .C(
        n53628), .Y(n3176) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47280 ( .A1(n77370), .A2(n57160), .B(n53192), 
        .C(n77369), .D(n56351), .Y(or1200_immu_top_N3) );
  A2O1A1Ixp33_ASAP7_75t_SL U47281 ( .A1(n77843), .A2(n56344), .B(n53192), .C(
        n53628), .Y(n56345) );
  A2O1A1Ixp33_ASAP7_75t_SL U47282 ( .A1(n77923), .A2(n59691), .B(n53192), .C(
        n53628), .Y(n55910) );
  A2O1A1Ixp33_ASAP7_75t_SL U47283 ( .A1(n59693), .A2(n56339), .B(n53192), .C(
        n53628), .Y(n56340) );
  A2O1A1Ixp33_ASAP7_75t_SL U47284 ( .A1(or1200_cpu_or1200_except_n613), .A2(
        n56340), .B(n53192), .C(n53628), .Y(n56341) );
  A2O1A1Ixp33_ASAP7_75t_SL U47285 ( .A1(n64162), .A2(n64163), .B(n53192), .C(
        n53628), .Y(n56335) );
  A2O1A1Ixp33_ASAP7_75t_SL U47286 ( .A1(n56334), .A2(n56335), .B(n53192), .C(
        n53628), .Y(n56336) );
  A2O1A1Ixp33_ASAP7_75t_SL U47287 ( .A1(n56336), .A2(n56337), .B(n53192), .C(
        n53628), .Y(n3013) );
  A2O1A1Ixp33_ASAP7_75t_SL U47288 ( .A1(n57144), .A2(n65210), .B(n53192), .C(
        n53628), .Y(n56332) );
  A2O1A1Ixp33_ASAP7_75t_SL U47289 ( .A1(n59691), .A2(n55677), .B(n53192), .C(
        n53628), .Y(n55678) );
  A2O1A1Ixp33_ASAP7_75t_SL U47290 ( .A1(n77919), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56117) );
  A2O1A1Ixp33_ASAP7_75t_SL U47291 ( .A1(n59628), .A2(n78433), .B(n53192), .C(
        n53628), .Y(n56325) );
  A2O1A1Ixp33_ASAP7_75t_SL U47292 ( .A1(n77974), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56116) );
  A2O1A1Ixp33_ASAP7_75t_SL U47293 ( .A1(n77505), .A2(n56323), .B(n53192), .C(
        n53628), .Y(n9477) );
  A2O1A1Ixp33_ASAP7_75t_SL U47294 ( .A1(n59691), .A2(n62052), .B(n53192), .C(
        n53628), .Y(n56320) );
  A2O1A1Ixp33_ASAP7_75t_SL U47295 ( .A1(n69335), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56114) );
  A2O1A1Ixp33_ASAP7_75t_SL U47296 ( .A1(n56108), .A2(n56112), .B(n53192), .C(
        n53628), .Y(n56113) );
  A2O1A1Ixp33_ASAP7_75t_SL U47297 ( .A1(n53628), .A2(n56113), .B(n53192), .C(
        n53628), .Y(n2453) );
  A2O1A1Ixp33_ASAP7_75t_SL U47298 ( .A1(n74706), .A2(n70534), .B(n53192), .C(
        n53628), .Y(n56307) );
  A2O1A1Ixp33_ASAP7_75t_SL U47299 ( .A1(n70533), .A2(n70532), .B(n53192), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .Y(
        n56310) );
  A2O1A1Ixp33_ASAP7_75t_SL U47300 ( .A1(n56309), .A2(n56310), .B(n53192), .C(
        n53628), .Y(n56311) );
  A2O1A1Ixp33_ASAP7_75t_SL U47301 ( .A1(n56306), .A2(n56311), .B(n53192), .C(
        n53628), .Y(n56312) );
  A2O1A1Ixp33_ASAP7_75t_SL U47302 ( .A1(n74677), .A2(n70542), .B(n53192), .C(
        n53628), .Y(n56316) );
  A2O1A1Ixp33_ASAP7_75t_SL U47303 ( .A1(n56315), .A2(n56316), .B(n53192), .C(
        n53628), .Y(n56317) );
  A2O1A1Ixp33_ASAP7_75t_SL U47304 ( .A1(n70541), .A2(n56317), .B(n53192), .C(
        n53628), .Y(n56318) );
  A2O1A1Ixp33_ASAP7_75t_SL U47305 ( .A1(n56312), .A2(n56318), .B(n53192), .C(
        n53628), .Y(n2433) );
  A2O1A1Ixp33_ASAP7_75t_SL U47306 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[6]), .B(n53192), 
        .C(n53628), .Y(n55889) );
  A2O1A1Ixp33_ASAP7_75t_SL U47307 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[6]), .A2(n55890), 
        .B(n53192), .C(n53628), .Y(n55891) );
  A2O1A1Ixp33_ASAP7_75t_SL U47308 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[6]), .B(
        n53192), .C(n53628), .Y(n55892) );
  A2O1A1Ixp33_ASAP7_75t_SL U47309 ( .A1(n55889), .A2(n55891), .B(n53192), .C(
        n55892), .Y(or1200_cpu_or1200_fpu_fpu_arith_N89) );
  A2O1A1Ixp33_ASAP7_75t_SL U47310 ( .A1(n53192), .A2(n53628), .B(n55444), .C(
        n53628), .Y(n55445) );
  A2O1A1Ixp33_ASAP7_75t_SL U47311 ( .A1(n63953), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56092) );
  A2O1A1Ixp33_ASAP7_75t_SL U47312 ( .A1(n77924), .A2(n59691), .B(n53192), .C(
        n53628), .Y(n55439) );
  A2O1A1Ixp33_ASAP7_75t_SL U47313 ( .A1(n77916), .A2(n59680), .B(n53192), .C(
        n53628), .Y(n56090) );
  A2O1A1Ixp33_ASAP7_75t_SL U47314 ( .A1(n77901), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56089) );
  A2O1A1Ixp33_ASAP7_75t_SL U47315 ( .A1(n77977), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56088) );
  A2O1A1Ixp33_ASAP7_75t_SL U47316 ( .A1(n77986), .A2(n59680), .B(n53192), .C(
        n53628), .Y(n56087) );
  A2O1A1Ixp33_ASAP7_75t_SL U47317 ( .A1(n77992), .A2(n77246), .B(n53192), .C(
        n53628), .Y(n56086) );
  A2O1A1Ixp33_ASAP7_75t_SL U47318 ( .A1(n59629), .A2(n72818), .B(n53192), .C(
        n72817), .Y(n56299) );
  A2O1A1Ixp33_ASAP7_75t_SL U47319 ( .A1(n3906), .A2(n56296), .B(n53192), .C(
        n53628), .Y(n56297) );
  A2O1A1Ixp33_ASAP7_75t_SL U47320 ( .A1(n77589), .A2(n77644), .B(n53192), .C(
        n53628), .Y(n56293) );
  A2O1A1Ixp33_ASAP7_75t_SL U47321 ( .A1(n77918), .A2(n77672), .B(n53192), .C(
        n53628), .Y(n56294) );
  A2O1A1Ixp33_ASAP7_75t_SL U47322 ( .A1(n56293), .A2(n56294), .B(n53192), .C(
        n53628), .Y(n56295) );
  A2O1A1Ixp33_ASAP7_75t_SL U47323 ( .A1(n76976), .A2(n56290), .B(n53192), .C(
        n53628), .Y(n1516) );
  A2O1A1Ixp33_ASAP7_75t_SL U47324 ( .A1(n57114), .A2(n77980), .B(n53192), .C(
        n53628), .Y(n56289) );
  A2O1A1Ixp33_ASAP7_75t_SL U47325 ( .A1(n1422), .A2(n56284), .B(n53192), .C(
        n53628), .Y(n56285) );
  A2O1A1Ixp33_ASAP7_75t_SL U47326 ( .A1(n77287), .A2(n77585), .B(n53192), .C(
        n53628), .Y(n56286) );
  A2O1A1Ixp33_ASAP7_75t_SL U47327 ( .A1(n56285), .A2(n56286), .B(n53192), .C(
        n53628), .Y(n56287) );
  A2O1A1Ixp33_ASAP7_75t_SL U47328 ( .A1(n56287), .A2(n56288), .B(n53192), .C(
        n53628), .Y(or1200_pic_N48) );
  A2O1A1Ixp33_ASAP7_75t_SL U47329 ( .A1(n77983), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n55018) );
  A2O1A1Ixp33_ASAP7_75t_SL U47330 ( .A1(n56077), .A2(n56079), .B(n53192), .C(
        n53628), .Y(n9354) );
  A2O1A1Ixp33_ASAP7_75t_SL U47331 ( .A1(n55853), .A2(n55855), .B(n53192), .C(
        n53628), .Y(n9350) );
  A2O1A1Ixp33_ASAP7_75t_SL U47332 ( .A1(n75030), .A2(n56074), .B(n53192), .C(
        n53628), .Y(n56075) );
  A2O1A1Ixp33_ASAP7_75t_SL U47333 ( .A1(n77862), .A2(n75649), .B(n53192), .C(
        n53628), .Y(n56076) );
  A2O1A1Ixp33_ASAP7_75t_SL U47334 ( .A1(n63298), .A2(n63297), .B(n53192), .C(
        n53628), .Y(n56061) );
  A2O1A1Ixp33_ASAP7_75t_SL U47335 ( .A1(n63775), .A2(n63778), .B(n53192), .C(
        n53628), .Y(n56258) );
  A2O1A1Ixp33_ASAP7_75t_SL U47336 ( .A1(n63532), .A2(n59674), .B(n53192), .C(
        n53628), .Y(n56261) );
  A2O1A1Ixp33_ASAP7_75t_SL U47337 ( .A1(n56258), .A2(n56261), .B(n53192), .C(
        n53628), .Y(n56262) );
  A2O1A1Ixp33_ASAP7_75t_SL U47338 ( .A1(n75015), .A2(n77890), .B(n53192), .C(
        n53628), .Y(n56267) );
  A2O1A1Ixp33_ASAP7_75t_SL U47339 ( .A1(n56266), .A2(n56267), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1577) );
  A2O1A1Ixp33_ASAP7_75t_SL U47340 ( .A1(n59673), .A2(n77888), .B(n53192), .C(
        n53628), .Y(n54428) );
  A2O1A1Ixp33_ASAP7_75t_SL U47341 ( .A1(n75650), .A2(n75363), .B(n53192), .C(
        n53628), .Y(n54429) );
  A2O1A1Ixp33_ASAP7_75t_SL U47342 ( .A1(n75295), .A2(n57080), .B(n53192), .C(
        n53628), .Y(n54432) );
  A2O1A1Ixp33_ASAP7_75t_SL U47343 ( .A1(n54435), .A2(n54436), .B(n53192), .C(
        n53628), .Y(n54437) );
  A2O1A1Ixp33_ASAP7_75t_SL U47344 ( .A1(n54428), .A2(n54429), .B(n53192), .C(
        n54438), .Y(or1200_cpu_or1200_mult_mac_n1607) );
  A2O1A1Ixp33_ASAP7_75t_SL U47345 ( .A1(n75650), .A2(n75116), .B(n53192), .C(
        n53628), .Y(n56243) );
  A2O1A1Ixp33_ASAP7_75t_SL U47346 ( .A1(n77866), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n56244) );
  A2O1A1Ixp33_ASAP7_75t_SL U47347 ( .A1(n75117), .A2(n57080), .B(n53192), .C(
        n53628), .Y(n56252) );
  A2O1A1Ixp33_ASAP7_75t_SL U47348 ( .A1(n56251), .A2(n56252), .B(n53192), .C(
        n53628), .Y(n56253) );
  A2O1A1Ixp33_ASAP7_75t_SL U47349 ( .A1(n56243), .A2(n56244), .B(n53192), .C(
        n56254), .Y(or1200_cpu_or1200_mult_mac_n1598) );
  A2O1A1Ixp33_ASAP7_75t_SL U47350 ( .A1(n77208), .A2(n77209), .B(n53192), .C(
        n53628), .Y(n56036) );
  A2O1A1Ixp33_ASAP7_75t_SL U47351 ( .A1(n76857), .A2(n59689), .B(n53192), .C(
        n53628), .Y(n56035) );
  A2O1A1Ixp33_ASAP7_75t_SL U47352 ( .A1(n76999), .A2(n59688), .B(n53192), .C(
        n53628), .Y(n56034) );
  A2O1A1Ixp33_ASAP7_75t_SL U47353 ( .A1(n77277), .A2(n57074), .B(n53192), .C(
        n53628), .Y(n56033) );
  A2O1A1Ixp33_ASAP7_75t_SL U47354 ( .A1(n76851), .A2(n59690), .B(n53192), .C(
        n53628), .Y(n55166) );
  A2O1A1Ixp33_ASAP7_75t_SL U47355 ( .A1(n76253), .A2(n59688), .B(n53192), .C(
        n53628), .Y(n56032) );
  A2O1A1Ixp33_ASAP7_75t_SL U47356 ( .A1(n75783), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n55373) );
  A2O1A1Ixp33_ASAP7_75t_SL U47357 ( .A1(n76553), .A2(n59688), .B(n53192), .C(
        n53628), .Y(n55372) );
  A2O1A1Ixp33_ASAP7_75t_SL U47358 ( .A1(n77227), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56031) );
  A2O1A1Ixp33_ASAP7_75t_SL U47359 ( .A1(n59693), .A2(n77021), .B(n53192), .C(
        n53628), .Y(n56242) );
  A2O1A1Ixp33_ASAP7_75t_SL U47360 ( .A1(n74986), .A2(n57074), .B(n53192), .C(
        n53628), .Y(n56030) );
  A2O1A1Ixp33_ASAP7_75t_SL U47361 ( .A1(n74578), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n56029) );
  A2O1A1Ixp33_ASAP7_75t_SL U47362 ( .A1(n75433), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n55802) );
  A2O1A1Ixp33_ASAP7_75t_SL U47363 ( .A1(n59693), .A2(n75449), .B(n53192), .C(
        n53628), .Y(n56240) );
  A2O1A1Ixp33_ASAP7_75t_SL U47364 ( .A1(n75622), .A2(n59693), .B(n53192), .C(
        n53628), .Y(n56028) );
  A2O1A1Ixp33_ASAP7_75t_SL U47365 ( .A1(n59693), .A2(n74081), .B(n53192), .C(
        n53628), .Y(n56239) );
  A2O1A1Ixp33_ASAP7_75t_SL U47366 ( .A1(n75798), .A2(n57074), .B(n53192), .C(
        n53628), .Y(n55602) );
  A2O1A1Ixp33_ASAP7_75t_SL U47367 ( .A1(n59688), .A2(n75200), .B(n53192), .C(
        n53628), .Y(n56238) );
  A2O1A1Ixp33_ASAP7_75t_SL U47368 ( .A1(n75686), .A2(n57074), .B(n53192), .C(
        n53628), .Y(n56026) );
  A2O1A1Ixp33_ASAP7_75t_SL U47369 ( .A1(n76928), .A2(n59690), .B(n53192), .C(
        n53628), .Y(n56025) );
  A2O1A1Ixp33_ASAP7_75t_SL U47370 ( .A1(n56014), .A2(n56015), .B(n53192), .C(
        n53628), .Y(n56016) );
  A2O1A1Ixp33_ASAP7_75t_SL U47371 ( .A1(n72494), .A2(n72464), .B(n53192), .C(
        n53628), .Y(n56017) );
  A2O1A1Ixp33_ASAP7_75t_SL U47372 ( .A1(n72463), .A2(n72492), .B(n53192), .C(
        n53628), .Y(n56018) );
  A2O1A1Ixp33_ASAP7_75t_SL U47373 ( .A1(n72332), .A2(n72333), .B(n53192), .C(
        n72490), .Y(n56019) );
  A2O1A1Ixp33_ASAP7_75t_SL U47374 ( .A1(n56017), .A2(n56018), .B(n53192), .C(
        n56019), .Y(n56020) );
  A2O1A1Ixp33_ASAP7_75t_SL U47375 ( .A1(n56021), .A2(n72500), .B(n53192), .C(
        n53628), .Y(n56022) );
  A2O1A1Ixp33_ASAP7_75t_SL U47376 ( .A1(n53192), .A2(n53628), .B(n56024), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n60) );
  A2O1A1Ixp33_ASAP7_75t_SL U47377 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_1_), .A2(n71413), 
        .B(n53192), .C(n53628), .Y(n56228) );
  A2O1A1Ixp33_ASAP7_75t_SL U47378 ( .A1(n66082), .A2(n56227), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n33) );
  A2O1A1Ixp33_ASAP7_75t_SL U47379 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .A2(
        n73704), .B(n53192), .C(n53628), .Y(n56226) );
  A2O1A1Ixp33_ASAP7_75t_SL U47380 ( .A1(n70196), .A2(n70195), .B(n53192), .C(
        n53628), .Y(n55994) );
  A2O1A1Ixp33_ASAP7_75t_SL U47381 ( .A1(n56220), .A2(n62056), .B(n53192), .C(
        n53628), .Y(n56221) );
  A2O1A1Ixp33_ASAP7_75t_SL U47382 ( .A1(n53628), .A2(n56221), .B(n53192), .C(
        n53628), .Y(n56222) );
  A2O1A1Ixp33_ASAP7_75t_SL U47383 ( .A1(n74703), .A2(n56218), .B(n53192), .C(
        n53628), .Y(n74708) );
  A2O1A1Ixp33_ASAP7_75t_SL U47384 ( .A1(n78138), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56216) );
  A2O1A1Ixp33_ASAP7_75t_SL U47385 ( .A1(n78139), .A2(n56216), .B(n53192), .C(
        n53628), .Y(n56217) );
  A2O1A1Ixp33_ASAP7_75t_SL U47386 ( .A1(n53628), .A2(n56217), .B(n53192), .C(
        n53628), .Y(n78134) );
  A2O1A1Ixp33_ASAP7_75t_SL U47387 ( .A1(n77952), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56210) );
  A2O1A1Ixp33_ASAP7_75t_SL U47388 ( .A1(n78177), .A2(n56210), .B(n53192), .C(
        n53628), .Y(n56211) );
  A2O1A1Ixp33_ASAP7_75t_SL U47389 ( .A1(n53628), .A2(n56211), .B(n53192), .C(
        n53628), .Y(n77962) );
  A2O1A1Ixp33_ASAP7_75t_SL U47390 ( .A1(n75467), .A2(n56206), .B(n53192), .C(
        n53628), .Y(n56207) );
  A2O1A1Ixp33_ASAP7_75t_SL U47391 ( .A1(n75468), .A2(n59638), .B(n53192), .C(
        n57398), .Y(n56208) );
  A2O1A1Ixp33_ASAP7_75t_SL U47392 ( .A1(n56207), .A2(n56208), .B(n53192), .C(
        n53628), .Y(n56209) );
  A2O1A1Ixp33_ASAP7_75t_SL U47393 ( .A1(n75469), .A2(n56209), .B(n53192), .C(
        n53628), .Y(n75471) );
  A2O1A1Ixp33_ASAP7_75t_SL U47394 ( .A1(n69098), .A2(n69094), .B(n53192), .C(
        n53628), .Y(n55529) );
  A2O1A1Ixp33_ASAP7_75t_SL U47395 ( .A1(n63461), .A2(n56203), .B(n53192), .C(
        n53628), .Y(n63415) );
  A2O1A1Ixp33_ASAP7_75t_SL U47396 ( .A1(n68944), .A2(n56201), .B(n53192), .C(
        n53628), .Y(n68911) );
  A2O1A1Ixp33_ASAP7_75t_SL U47397 ( .A1(n69257), .A2(n56199), .B(n53192), .C(
        n53628), .Y(n69283) );
  A2O1A1Ixp33_ASAP7_75t_SL U47398 ( .A1(n76901), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56195) );
  A2O1A1Ixp33_ASAP7_75t_SL U47399 ( .A1(n76900), .A2(n56195), .B(n53192), .C(
        n53628), .Y(n56196) );
  A2O1A1Ixp33_ASAP7_75t_SL U47400 ( .A1(n53628), .A2(n56196), .B(n53192), .C(
        n53628), .Y(n76902) );
  A2O1A1Ixp33_ASAP7_75t_SL U47401 ( .A1(n77430), .A2(
        or1200_cpu_or1200_except_n120), .B(n53192), .C(n54922), .Y(n77447) );
  A2O1A1Ixp33_ASAP7_75t_SL U47402 ( .A1(n56192), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_22_), .B(
        n53192), .C(n53628), .Y(n74297) );
  A2O1A1Ixp33_ASAP7_75t_SL U47403 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n56181) );
  A2O1A1Ixp33_ASAP7_75t_SL U47404 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n56182) );
  A2O1A1Ixp33_ASAP7_75t_SL U47405 ( .A1(n56181), .A2(n56182), .B(n53192), .C(
        n53628), .Y(n56183) );
  A2O1A1Ixp33_ASAP7_75t_SL U47406 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_25_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n56185) );
  A2O1A1Ixp33_ASAP7_75t_SL U47407 ( .A1(n56184), .A2(n56185), .B(n53192), .C(
        n53628), .Y(n72103) );
  A2O1A1Ixp33_ASAP7_75t_SL U47408 ( .A1(n70803), .A2(n70804), .B(n53192), .C(
        n53628), .Y(n56175) );
  A2O1A1Ixp33_ASAP7_75t_SL U47409 ( .A1(n70837), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n56173) );
  A2O1A1Ixp33_ASAP7_75t_SL U47410 ( .A1(n70835), .A2(n56173), .B(n53192), .C(
        n53628), .Y(n56174) );
  A2O1A1Ixp33_ASAP7_75t_SL U47411 ( .A1(n53628), .A2(n56174), .B(n53192), .C(
        n53628), .Y(n70822) );
  A2O1A1Ixp33_ASAP7_75t_SL U47412 ( .A1(n71252), .A2(n71251), .B(n53192), .C(
        n53628), .Y(n56171) );
  A2O1A1Ixp33_ASAP7_75t_SL U47413 ( .A1(n65670), .A2(n65602), .B(n53192), .C(
        n53628), .Y(n56170) );
  A2O1A1Ixp33_ASAP7_75t_SL U47414 ( .A1(n56169), .A2(n56170), .B(n53192), .C(
        n53628), .Y(n66121) );
  A2O1A1Ixp33_ASAP7_75t_SL U47415 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[16]), .A2(
        n59631), .B(n53192), .C(n53628), .Y(n54052) );
  A2O1A1Ixp33_ASAP7_75t_SL U47416 ( .A1(n59561), .A2(n59583), .B(n53192), .C(
        n53628), .Y(n56161) );
  A2O1A1Ixp33_ASAP7_75t_SL U47417 ( .A1(n75246), .A2(n77060), .B(n53192), .C(
        n53628), .Y(n56158) );
  A2O1A1Ixp33_ASAP7_75t_SL U47418 ( .A1(n53658), .A2(n53659), .B(n53192), .C(
        n53628), .Y(n64856) );
  A2O1A1Ixp33_ASAP7_75t_SL U47419 ( .A1(n69141), .A2(n56156), .B(n53192), .C(
        n53628), .Y(n56157) );
  A2O1A1Ixp33_ASAP7_75t_SL U47420 ( .A1(n69143), .A2(n56157), .B(n53192), .C(
        n53628), .Y(n69145) );
  A2O1A1Ixp33_ASAP7_75t_SL U47421 ( .A1(n63889), .A2(n63890), .B(n53192), .C(
        n53628), .Y(n56152) );
  A2O1A1Ixp33_ASAP7_75t_SL U47422 ( .A1(n54881), .A2(n54882), .B(n53192), .C(
        n53628), .Y(n69107) );
  A2O1A1Ixp33_ASAP7_75t_SL U47423 ( .A1(n59631), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[6]), .B(
        n53192), .C(n53628), .Y(n56150) );
  A2O1A1Ixp33_ASAP7_75t_SL U47424 ( .A1(n72929), .A2(n56148), .B(n53192), .C(
        n53628), .Y(n72944) );
  A2O1A1Ixp33_ASAP7_75t_SL U47425 ( .A1(n53192), .A2(n53628), .B(n55934), .C(
        n53628), .Y(n55935) );
  A2O1A1Ixp33_ASAP7_75t_SL U47426 ( .A1(n73472), .A2(n73473), .B(n53192), .C(
        n73477), .Y(n56136) );
  A2O1A1Ixp33_ASAP7_75t_SL U47427 ( .A1(n71520), .A2(n71518), .B(n53192), .C(
        n56132), .Y(n56133) );
  A2O1A1Ixp33_ASAP7_75t_SL U47428 ( .A1(n74920), .A2(or1200_cpu_or1200_fpu_ine), .B(n53192), .C(n53628), .Y(n56126) );
  A2O1A1Ixp33_ASAP7_75t_SL U47429 ( .A1(n56125), .A2(n56126), .B(n53192), .C(
        n53628), .Y(n9485) );
  A2O1A1Ixp33_ASAP7_75t_SL U47430 ( .A1(n61286), .A2(n55911), .B(n53192), .C(
        n53628), .Y(n55912) );
  A2O1A1Ixp33_ASAP7_75t_SL U47431 ( .A1(n61288), .A2(n55916), .B(n53192), .C(
        n53628), .Y(n9378) );
  A2O1A1Ixp33_ASAP7_75t_SL U47432 ( .A1(n59695), .A2(n77770), .B(n53192), .C(
        n53628), .Y(n56122) );
  A2O1A1Ixp33_ASAP7_75t_SL U47433 ( .A1(n76840), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55906) );
  A2O1A1Ixp33_ASAP7_75t_SL U47434 ( .A1(n76841), .A2(n55907), .B(n53192), .C(
        n53628), .Y(n55908) );
  A2O1A1Ixp33_ASAP7_75t_SL U47435 ( .A1(n77194), .A2(n74844), .B(n53192), .C(
        n53628), .Y(n56119) );
  A2O1A1Ixp33_ASAP7_75t_SL U47436 ( .A1(n59691), .A2(n55896), .B(n53192), .C(
        n53628), .Y(n55897) );
  A2O1A1Ixp33_ASAP7_75t_SL U47437 ( .A1(n57073), .A2(n54510), .B(n53192), .C(
        n53628), .Y(n54511) );
  A2O1A1Ixp33_ASAP7_75t_SL U47438 ( .A1(n69378), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_2_), .B(n53192), .C(
        n53628), .Y(n56108) );
  A2O1A1Ixp33_ASAP7_75t_SL U47439 ( .A1(n53628), .A2(n70502), .B(n53192), .C(
        n53628), .Y(n56109) );
  A2O1A1Ixp33_ASAP7_75t_SL U47440 ( .A1(n69379), .A2(n56109), .B(n53192), .C(
        n53628), .Y(n56110) );
  A2O1A1Ixp33_ASAP7_75t_SL U47441 ( .A1(n53628), .A2(n56110), .B(n53192), .C(
        n53628), .Y(n56111) );
  A2O1A1Ixp33_ASAP7_75t_SL U47442 ( .A1(n70478), .A2(n56111), .B(n53192), .C(
        n53628), .Y(n56112) );
  A2O1A1Ixp33_ASAP7_75t_SL U47443 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_9_), .A2(
        n70476), .B(n53192), .C(n53628), .Y(n56100) );
  A2O1A1Ixp33_ASAP7_75t_SL U47444 ( .A1(n70485), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_8_), .B(
        n53192), .C(n53628), .Y(n56101) );
  A2O1A1Ixp33_ASAP7_75t_SL U47445 ( .A1(n56100), .A2(n56101), .B(n53192), .C(
        n53628), .Y(n56102) );
  A2O1A1Ixp33_ASAP7_75t_SL U47446 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n70388), .B(n53192), .C(n53628), .Y(n56105) );
  A2O1A1Ixp33_ASAP7_75t_SL U47447 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[7]), .B(n53192), 
        .C(n53628), .Y(n55667) );
  A2O1A1Ixp33_ASAP7_75t_SL U47448 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[7]), .A2(n55668), 
        .B(n53192), .C(n53628), .Y(n55669) );
  A2O1A1Ixp33_ASAP7_75t_SL U47449 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[7]), .B(
        n53192), .C(n53628), .Y(n55670) );
  A2O1A1Ixp33_ASAP7_75t_SL U47450 ( .A1(n55667), .A2(n55669), .B(n53192), .C(
        n55670), .Y(or1200_cpu_or1200_fpu_fpu_arith_N90) );
  A2O1A1Ixp33_ASAP7_75t_SL U47451 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[0]), .B(n53192), 
        .C(n53628), .Y(n54847) );
  A2O1A1Ixp33_ASAP7_75t_SL U47452 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[0]), .A2(n54848), 
        .B(n53192), .C(n53628), .Y(n54849) );
  A2O1A1Ixp33_ASAP7_75t_SL U47453 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[0]), .B(
        n53192), .C(n53628), .Y(n54850) );
  A2O1A1Ixp33_ASAP7_75t_SL U47454 ( .A1(n54847), .A2(n54849), .B(n53192), .C(
        n54850), .Y(or1200_cpu_or1200_fpu_fpu_arith_N83) );
  A2O1A1Ixp33_ASAP7_75t_SL U47455 ( .A1(n69726), .A2(n55882), .B(n53192), .C(
        n53628), .Y(n55884) );
  A2O1A1Ixp33_ASAP7_75t_SL U47456 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_5_), .A2(n53628), .B(n53192), 
        .C(n53628), .Y(n56095) );
  A2O1A1Ixp33_ASAP7_75t_SL U47457 ( .A1(n62063), .A2(n56095), .B(n53192), .C(
        n53628), .Y(n56096) );
  A2O1A1Ixp33_ASAP7_75t_SL U47458 ( .A1(n62063), .A2(n62057), .B(n53192), .C(
        n53628), .Y(n56097) );
  A2O1A1Ixp33_ASAP7_75t_SL U47459 ( .A1(n56096), .A2(n56098), .B(n53192), .C(
        n53628), .Y(n2207) );
  A2O1A1Ixp33_ASAP7_75t_SL U47460 ( .A1(n57144), .A2(n2199), .B(n53192), .C(
        n53628), .Y(n56093) );
  A2O1A1Ixp33_ASAP7_75t_SL U47461 ( .A1(n77024), .A2(n56093), .B(n53192), .C(
        n53628), .Y(n56094) );
  A2O1A1Ixp33_ASAP7_75t_SL U47462 ( .A1(n53628), .A2(n56094), .B(n53192), .C(
        n53628), .Y(n2200) );
  A2O1A1Ixp33_ASAP7_75t_SL U47463 ( .A1(n77927), .A2(n59691), .B(n53192), .C(
        n53628), .Y(n55878) );
  A2O1A1Ixp33_ASAP7_75t_SL U47464 ( .A1(n57198), .A2(n76623), .B(n53192), .C(
        n53628), .Y(n54468) );
  A2O1A1Ixp33_ASAP7_75t_SL U47465 ( .A1(n3905), .A2(n56084), .B(n53192), .C(
        n53628), .Y(n56085) );
  A2O1A1Ixp33_ASAP7_75t_SL U47466 ( .A1(n75616), .A2(n77875), .B(n53192), .C(
        n53628), .Y(n56081) );
  A2O1A1Ixp33_ASAP7_75t_SL U47467 ( .A1(n57114), .A2(n77918), .B(n53192), .C(
        n53628), .Y(n56080) );
  A2O1A1Ixp33_ASAP7_75t_SL U47468 ( .A1(n77968), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n55652) );
  A2O1A1Ixp33_ASAP7_75t_SL U47469 ( .A1(n77971), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n54816) );
  A2O1A1Ixp33_ASAP7_75t_SL U47470 ( .A1(n57142), .A2(n77978), .B(n53192), .C(
        n53628), .Y(n56077) );
  A2O1A1Ixp33_ASAP7_75t_SL U47471 ( .A1(n77979), .A2(n56078), .B(n53192), .C(
        n53628), .Y(n56079) );
  A2O1A1Ixp33_ASAP7_75t_SL U47472 ( .A1(n63256), .A2(n56065), .B(n53192), .C(
        n53628), .Y(n56066) );
  A2O1A1Ixp33_ASAP7_75t_SL U47473 ( .A1(n63687), .A2(n56067), .B(n53192), .C(
        n53628), .Y(n56068) );
  A2O1A1Ixp33_ASAP7_75t_SL U47474 ( .A1(n56061), .A2(n56062), .B(n53192), .C(
        n53628), .Y(n56063) );
  A2O1A1Ixp33_ASAP7_75t_SL U47475 ( .A1(n56049), .A2(n56057), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1572) );
  A2O1A1Ixp33_ASAP7_75t_SL U47476 ( .A1(n57079), .A2(n69213), .B(n53192), .C(
        n53628), .Y(n55816) );
  A2O1A1Ixp33_ASAP7_75t_SL U47477 ( .A1(n69162), .A2(n57080), .B(n53192), .C(
        n53628), .Y(n55828) );
  A2O1A1Ixp33_ASAP7_75t_SL U47478 ( .A1(n75139), .A2(n75140), .B(n53192), .C(
        n53628), .Y(n56037) );
  A2O1A1Ixp33_ASAP7_75t_SL U47479 ( .A1(n57080), .A2(n56037), .B(n53192), .C(
        n53628), .Y(n56043) );
  A2O1A1Ixp33_ASAP7_75t_SL U47480 ( .A1(n56042), .A2(n56043), .B(n53192), .C(
        n53628), .Y(n56044) );
  A2O1A1Ixp33_ASAP7_75t_SL U47481 ( .A1(n75650), .A2(n75654), .B(n53192), .C(
        n53628), .Y(n56046) );
  A2O1A1Ixp33_ASAP7_75t_SL U47482 ( .A1(n77859), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n56047) );
  A2O1A1Ixp33_ASAP7_75t_SL U47483 ( .A1(n56045), .A2(n56046), .B(n53192), .C(
        n56047), .Y(or1200_cpu_or1200_mult_mac_n1595) );
  A2O1A1Ixp33_ASAP7_75t_SL U47484 ( .A1(n77288), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n54625) );
  A2O1A1Ixp33_ASAP7_75t_SL U47485 ( .A1(n76232), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n55803) );
  A2O1A1Ixp33_ASAP7_75t_SL U47486 ( .A1(n75312), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n55603) );
  A2O1A1Ixp33_ASAP7_75t_SL U47487 ( .A1(n74081), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n55369) );
  A2O1A1Ixp33_ASAP7_75t_SL U47488 ( .A1(n55794), .A2(n55795), .B(n53192), .C(
        n53628), .Y(n55796) );
  A2O1A1Ixp33_ASAP7_75t_SL U47489 ( .A1(n53628), .A2(n56010), .B(n53192), .C(
        n53628), .Y(n56011) );
  A2O1A1Ixp33_ASAP7_75t_SL U47490 ( .A1(n58447), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_), 
        .B(n53192), .C(n53628), .Y(n56015) );
  A2O1A1Ixp33_ASAP7_75t_SL U47491 ( .A1(n71796), .A2(n56007), .B(n53192), .C(
        n53628), .Y(n28105) );
  A2O1A1Ixp33_ASAP7_75t_SL U47492 ( .A1(n70835), .A2(n70833), .B(n53192), .C(
        n53628), .Y(n55336) );
  A2O1A1Ixp33_ASAP7_75t_SL U47493 ( .A1(n53192), .A2(n53628), .B(n55339), .C(
        n53628), .Y(n55340) );
  A2O1A1Ixp33_ASAP7_75t_SL U47494 ( .A1(n66082), .A2(n55999), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n35) );
  A2O1A1Ixp33_ASAP7_75t_SL U47495 ( .A1(n73623), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .B(
        n53192), .C(n53628), .Y(n55995) );
  A2O1A1Ixp33_ASAP7_75t_SL U47496 ( .A1(n70197), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55992) );
  A2O1A1Ixp33_ASAP7_75t_SL U47497 ( .A1(n70194), .A2(n55992), .B(n53192), .C(
        n53628), .Y(n55993) );
  A2O1A1Ixp33_ASAP7_75t_SL U47498 ( .A1(n55993), .A2(n55994), .B(n53192), .C(
        n53628), .Y(n70198) );
  A2O1A1Ixp33_ASAP7_75t_SL U47499 ( .A1(n74681), .A2(n54756), .B(n53192), .C(
        n53628), .Y(n74671) );
  A2O1A1Ixp33_ASAP7_75t_SL U47500 ( .A1(n55990), .A2(n74809), .B(n53192), .C(
        n53628), .Y(n76491) );
  A2O1A1Ixp33_ASAP7_75t_SL U47501 ( .A1(n74574), .A2(n74575), .B(n53192), .C(
        n53628), .Y(n54933) );
  A2O1A1Ixp33_ASAP7_75t_SL U47502 ( .A1(n63346), .A2(n55981), .B(n53192), .C(
        n53628), .Y(n63347) );
  A2O1A1Ixp33_ASAP7_75t_SL U47503 ( .A1(n63454), .A2(n55980), .B(n53192), .C(
        n53628), .Y(n63467) );
  A2O1A1Ixp33_ASAP7_75t_SL U47504 ( .A1(n68832), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55977) );
  A2O1A1Ixp33_ASAP7_75t_SL U47505 ( .A1(n68885), .A2(n55977), .B(n53192), .C(
        n53628), .Y(n55978) );
  A2O1A1Ixp33_ASAP7_75t_SL U47506 ( .A1(n53628), .A2(n55978), .B(n53192), .C(
        n53628), .Y(n68848) );
  A2O1A1Ixp33_ASAP7_75t_SL U47507 ( .A1(or1200_cpu_or1200_mult_mac_n225), .A2(
        n55975), .B(n53192), .C(n53628), .Y(n69061) );
  A2O1A1Ixp33_ASAP7_75t_SL U47508 ( .A1(n54906), .A2(n54907), .B(n53192), .C(
        n53628), .Y(n54908) );
  A2O1A1Ixp33_ASAP7_75t_SL U47509 ( .A1(n54905), .A2(n54909), .B(n53192), .C(
        n53628), .Y(n72125) );
  A2O1A1Ixp33_ASAP7_75t_SL U47510 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n55967) );
  A2O1A1Ixp33_ASAP7_75t_SL U47511 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n55968) );
  A2O1A1Ixp33_ASAP7_75t_SL U47512 ( .A1(n55967), .A2(n55968), .B(n53192), .C(
        n53628), .Y(n55969) );
  A2O1A1Ixp33_ASAP7_75t_SL U47513 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n55971) );
  A2O1A1Ixp33_ASAP7_75t_SL U47514 ( .A1(n55970), .A2(n55971), .B(n53192), .C(
        n53628), .Y(n71927) );
  A2O1A1Ixp33_ASAP7_75t_SL U47515 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[21]), .A2(
        n59631), .B(n53192), .C(n53628), .Y(n55735) );
  A2O1A1Ixp33_ASAP7_75t_SL U47516 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_33_), .A2(n70103), 
        .B(n53192), .C(n53628), .Y(n55733) );
  A2O1A1Ixp33_ASAP7_75t_SL U47517 ( .A1(n75617), .A2(n55951), .B(n53192), .C(
        n53628), .Y(n74042) );
  A2O1A1Ixp33_ASAP7_75t_SL U47518 ( .A1(n71936), .A2(n54373), .B(n53192), .C(
        n53628), .Y(n71550) );
  A2O1A1Ixp33_ASAP7_75t_SL U47519 ( .A1(n53192), .A2(n53628), .B(n55279), .C(
        n53628), .Y(n55280) );
  A2O1A1Ixp33_ASAP7_75t_SL U47520 ( .A1(n73265), .A2(n74502), .B(n53192), .C(
        n53628), .Y(n55942) );
  A2O1A1Ixp33_ASAP7_75t_SL U47521 ( .A1(n72904), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), .B(
        n53192), .C(n53628), .Y(n55937) );
  A2O1A1Ixp33_ASAP7_75t_SL U47522 ( .A1(n72902), .A2(n72993), .B(n53192), .C(
        n53628), .Y(n55938) );
  A2O1A1Ixp33_ASAP7_75t_SL U47523 ( .A1(n55937), .A2(n55938), .B(n53192), .C(
        n53628), .Y(n72758) );
  A2O1A1Ixp33_ASAP7_75t_SL U47524 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[25]), .A2(
        n55936), .B(n53192), .C(n53628), .Y(n73103) );
  A2O1A1Ixp33_ASAP7_75t_SL U47525 ( .A1(n67264), .A2(n59603), .B(n53192), .C(
        n53628), .Y(n55931) );
  A2O1A1Ixp33_ASAP7_75t_SL U47526 ( .A1(n55701), .A2(n55702), .B(n53192), .C(
        n53628), .Y(n12863) );
  A2O1A1Ixp33_ASAP7_75t_SL U47527 ( .A1(n73661), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55927) );
  A2O1A1Ixp33_ASAP7_75t_SL U47528 ( .A1(n73653), .A2(n55927), .B(n53192), .C(
        n53628), .Y(n55928) );
  A2O1A1Ixp33_ASAP7_75t_SL U47529 ( .A1(n73660), .A2(n55928), .B(n53192), .C(
        n53628), .Y(n3279) );
  A2O1A1Ixp33_ASAP7_75t_SL U47530 ( .A1(n53192), .A2(n53628), .B(n55696), .C(
        n53628), .Y(n55697) );
  A2O1A1Ixp33_ASAP7_75t_SL U47531 ( .A1(n71516), .A2(n71517), .B(n53192), .C(
        n55697), .Y(n55698) );
  A2O1A1Ixp33_ASAP7_75t_SL U47532 ( .A1(n71521), .A2(n55696), .B(n53192), .C(
        n53628), .Y(n55699) );
  A2O1A1Ixp33_ASAP7_75t_SL U47533 ( .A1(n55698), .A2(n55699), .B(n53192), .C(
        n53628), .Y(n3271) );
  A2O1A1Ixp33_ASAP7_75t_SL U47534 ( .A1(n70575), .A2(n55920), .B(n53192), .C(
        n53628), .Y(n55921) );
  A2O1A1Ixp33_ASAP7_75t_SL U47535 ( .A1(n70582), .A2(n55921), .B(n53192), .C(
        n53628), .Y(n55922) );
  A2O1A1Ixp33_ASAP7_75t_SL U47536 ( .A1(n59629), .A2(n78340), .B(n53192), .C(
        n53628), .Y(n55917) );
  A2O1A1Ixp33_ASAP7_75t_SL U47537 ( .A1(n53628), .A2(n3109), .B(n53192), .C(
        n53628), .Y(n55913) );
  A2O1A1Ixp33_ASAP7_75t_SL U47538 ( .A1(n77996), .A2(n55913), .B(n53192), .C(
        n53628), .Y(n55914) );
  A2O1A1Ixp33_ASAP7_75t_SL U47539 ( .A1(n3107), .A2(n55914), .B(n53192), .C(
        n53628), .Y(n55915) );
  A2O1A1Ixp33_ASAP7_75t_SL U47540 ( .A1(n55912), .A2(n55915), .B(n53192), .C(
        n53628), .Y(n55916) );
  A2O1A1Ixp33_ASAP7_75t_SL U47541 ( .A1(n59690), .A2(n55906), .B(n53192), .C(
        n53628), .Y(n55907) );
  A2O1A1Ixp33_ASAP7_75t_SL U47542 ( .A1(n57144), .A2(n63968), .B(n53192), .C(
        n53628), .Y(n55905) );
  A2O1A1Ixp33_ASAP7_75t_SL U47543 ( .A1(n75417), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55687) );
  A2O1A1Ixp33_ASAP7_75t_SL U47544 ( .A1(n75416), .A2(n55688), .B(n53192), .C(
        n53628), .Y(n55689) );
  A2O1A1Ixp33_ASAP7_75t_SL U47545 ( .A1(n53192), .A2(n53628), .B(n55233), .C(
        n53628), .Y(n55234) );
  A2O1A1Ixp33_ASAP7_75t_SL U47546 ( .A1(n2450), .A2(n69383), .B(n53192), .C(
        n53628), .Y(n55462) );
  A2O1A1Ixp33_ASAP7_75t_SL U47547 ( .A1(n55446), .A2(n55449), .B(n53192), .C(
        n53628), .Y(n55450) );
  A2O1A1Ixp33_ASAP7_75t_SL U47548 ( .A1(n70475), .A2(n70474), .B(n53192), .C(
        n70491), .Y(n55457) );
  A2O1A1Ixp33_ASAP7_75t_SL U47549 ( .A1(n53628), .A2(n69729), .B(n53192), .C(
        n53628), .Y(n55880) );
  A2O1A1Ixp33_ASAP7_75t_SL U47550 ( .A1(n69728), .A2(n55880), .B(n53192), .C(
        n53628), .Y(n55881) );
  A2O1A1Ixp33_ASAP7_75t_SL U47551 ( .A1(n53628), .A2(n55881), .B(n53192), .C(
        n53628), .Y(n55882) );
  A2O1A1Ixp33_ASAP7_75t_SL U47552 ( .A1(n74793), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n55666) );
  A2O1A1Ixp33_ASAP7_75t_SL U47553 ( .A1(n61124), .A2(n55876), .B(n53192), .C(
        n53628), .Y(n55877) );
  A2O1A1Ixp33_ASAP7_75t_SL U47554 ( .A1(n57144), .A2(n76626), .B(n53192), .C(
        n53628), .Y(n55875) );
  A2O1A1Ixp33_ASAP7_75t_SL U47555 ( .A1(n59680), .A2(n77918), .B(n53192), .C(
        n53628), .Y(n55874) );
  A2O1A1Ixp33_ASAP7_75t_SL U47556 ( .A1(n3904), .A2(n55872), .B(n53192), .C(
        n53628), .Y(n55873) );
  A2O1A1Ixp33_ASAP7_75t_SL U47557 ( .A1(n57190), .A2(n78357), .B(n53192), .C(
        n53628), .Y(n55869) );
  A2O1A1Ixp33_ASAP7_75t_SL U47558 ( .A1(n74756), .A2(n1494), .B(n53192), .C(
        n53628), .Y(n54828) );
  A2O1A1Ixp33_ASAP7_75t_SL U47559 ( .A1(n62070), .A2(n54829), .B(n53192), .C(
        n53628), .Y(n54830) );
  A2O1A1Ixp33_ASAP7_75t_SL U47560 ( .A1(n57114), .A2(n77916), .B(n53192), .C(
        n53628), .Y(n55868) );
  A2O1A1Ixp33_ASAP7_75t_SL U47561 ( .A1(n77974), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n54663) );
  A2O1A1Ixp33_ASAP7_75t_SL U47562 ( .A1(n77977), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n55215) );
  A2O1A1Ixp33_ASAP7_75t_SL U47563 ( .A1(n74641), .A2(n77986), .B(n53192), .C(
        n53628), .Y(n55867) );
  A2O1A1Ixp33_ASAP7_75t_SL U47564 ( .A1(n1390), .A2(n55862), .B(n53192), .C(
        n53628), .Y(n55863) );
  A2O1A1Ixp33_ASAP7_75t_SL U47565 ( .A1(n77287), .A2(n76508), .B(n53192), .C(
        n53628), .Y(n55864) );
  A2O1A1Ixp33_ASAP7_75t_SL U47566 ( .A1(n55863), .A2(n55864), .B(n53192), .C(
        n53628), .Y(n55865) );
  A2O1A1Ixp33_ASAP7_75t_SL U47567 ( .A1(n55865), .A2(n55866), .B(n53192), .C(
        n53628), .Y(or1200_pic_N56) );
  A2O1A1Ixp33_ASAP7_75t_SL U47568 ( .A1(n1386), .A2(n55857), .B(n53192), .C(
        n53628), .Y(n55858) );
  A2O1A1Ixp33_ASAP7_75t_SL U47569 ( .A1(n77287), .A2(n75781), .B(n53192), .C(
        n53628), .Y(n55859) );
  A2O1A1Ixp33_ASAP7_75t_SL U47570 ( .A1(n55858), .A2(n55859), .B(n53192), .C(
        n53628), .Y(n55860) );
  A2O1A1Ixp33_ASAP7_75t_SL U47571 ( .A1(n55860), .A2(n55861), .B(n53192), .C(
        n53628), .Y(or1200_pic_N57) );
  A2O1A1Ixp33_ASAP7_75t_SL U47572 ( .A1(n55649), .A2(n55651), .B(n53192), .C(
        n53628), .Y(n9353) );
  A2O1A1Ixp33_ASAP7_75t_SL U47573 ( .A1(n57142), .A2(n77963), .B(n53192), .C(
        n53628), .Y(n55853) );
  A2O1A1Ixp33_ASAP7_75t_SL U47574 ( .A1(n77964), .A2(n55854), .B(n53192), .C(
        n53628), .Y(n55855) );
  A2O1A1Ixp33_ASAP7_75t_SL U47575 ( .A1(n76224), .A2(n57245), .B(n53192), .C(
        n55642), .Y(n55643) );
  A2O1A1Ixp33_ASAP7_75t_SL U47576 ( .A1(n76224), .A2(n57245), .B(n53192), .C(
        n53628), .Y(n55644) );
  A2O1A1Ixp33_ASAP7_75t_SL U47577 ( .A1(n55644), .A2(n76226), .B(n53192), .C(
        n53628), .Y(n55645) );
  A2O1A1Ixp33_ASAP7_75t_SL U47578 ( .A1(n55643), .A2(n55645), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N14) );
  A2O1A1Ixp33_ASAP7_75t_SL U47579 ( .A1(n53192), .A2(n53628), .B(n55401), .C(
        n53628), .Y(n55402) );
  A2O1A1Ixp33_ASAP7_75t_SL U47580 ( .A1(n55405), .A2(n55406), .B(n53192), .C(
        n53628), .Y(n55407) );
  A2O1A1Ixp33_ASAP7_75t_SL U47581 ( .A1(n63298), .A2(n55404), .B(n53192), .C(
        n55407), .Y(n55408) );
  A2O1A1Ixp33_ASAP7_75t_SL U47582 ( .A1(n55408), .A2(n55412), .B(n53192), .C(
        n53628), .Y(n58577) );
  A2O1A1Ixp33_ASAP7_75t_SL U47583 ( .A1(n55841), .A2(n55842), .B(n53192), .C(
        n53628), .Y(n55843) );
  A2O1A1Ixp33_ASAP7_75t_SL U47584 ( .A1(n63778), .A2(n63532), .B(n53192), .C(
        n53628), .Y(n55831) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47585 ( .A1(n63775), .A2(n59674), .B(n53192), 
        .C(n55831), .D(n55832), .Y(n55833) );
  A2O1A1Ixp33_ASAP7_75t_SL U47586 ( .A1(n59673), .A2(n77920), .B(n53192), .C(
        n53628), .Y(n53954) );
  A2O1A1Ixp33_ASAP7_75t_SL U47587 ( .A1(n75650), .A2(n68846), .B(n53192), .C(
        n53628), .Y(n53955) );
  A2O1A1Ixp33_ASAP7_75t_SL U47588 ( .A1(n53954), .A2(n53955), .B(n53192), .C(
        n53964), .Y(or1200_cpu_or1200_mult_mac_n1623) );
  A2O1A1Ixp33_ASAP7_75t_SL U47589 ( .A1(n55819), .A2(n55821), .B(n53192), .C(
        n53628), .Y(n55822) );
  A2O1A1Ixp33_ASAP7_75t_SL U47590 ( .A1(or1200_cpu_or1200_mult_mac_n381), .A2(
        n55823), .B(n53192), .C(n53628), .Y(n55824) );
  A2O1A1Ixp33_ASAP7_75t_SL U47591 ( .A1(n53628), .A2(n55824), .B(n53192), .C(
        n53628), .Y(n55825) );
  A2O1A1Ixp33_ASAP7_75t_SL U47592 ( .A1(or1200_cpu_or1200_mult_mac_n235), .A2(
        n55825), .B(n53192), .C(n53628), .Y(n55826) );
  A2O1A1Ixp33_ASAP7_75t_SL U47593 ( .A1(n55822), .A2(n55826), .B(n53192), .C(
        n53628), .Y(n55827) );
  A2O1A1Ixp33_ASAP7_75t_SL U47594 ( .A1(n75822), .A2(n75650), .B(n53192), .C(
        n53628), .Y(n55812) );
  A2O1A1Ixp33_ASAP7_75t_SL U47595 ( .A1(n77247), .A2(n77442), .B(n53192), .C(
        n53628), .Y(n55804) );
  A2O1A1Ixp33_ASAP7_75t_SL U47596 ( .A1(n76704), .A2(n59690), .B(n53192), .C(
        n53628), .Y(n55167) );
  A2O1A1Ixp33_ASAP7_75t_SL U47597 ( .A1(n77021), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n55599) );
  A2O1A1Ixp33_ASAP7_75t_SL U47598 ( .A1(n57072), .A2(n74986), .B(n53192), .C(
        n53628), .Y(n55801) );
  A2O1A1Ixp33_ASAP7_75t_SL U47599 ( .A1(n75449), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n53951) );
  A2O1A1Ixp33_ASAP7_75t_SL U47600 ( .A1(n69373), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n55163) );
  A2O1A1Ixp33_ASAP7_75t_SL U47601 ( .A1(n53192), .A2(n53628), .B(n55596), .C(
        n53628), .Y(n55597) );
  A2O1A1Ixp33_ASAP7_75t_SL U47602 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .A2(n71785), .B(n53192), .C(n71709), .Y(n55798) );
  A2O1A1Ixp33_ASAP7_75t_SL U47603 ( .A1(n55797), .A2(n55798), .B(n53192), .C(
        n53628), .Y(n55799) );
  A2O1A1Ixp33_ASAP7_75t_SL U47604 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_0_), .A2(
        n71799), .B(n53192), .C(n71710), .Y(n55800) );
  A2O1A1Ixp33_ASAP7_75t_SL U47605 ( .A1(n55799), .A2(n55800), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n120) );
  A2O1A1Ixp33_ASAP7_75t_SL U47606 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_22_), 
        .A2(n57103), .B(n53192), .C(n53628), .Y(n55795) );
  A2O1A1Ixp33_ASAP7_75t_SL U47607 ( .A1(n72451), .A2(n72326), .B(n53192), .C(
        n55788), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n70) );
  A2O1A1Ixp33_ASAP7_75t_SL U47608 ( .A1(n53192), .A2(n53628), .B(n55566), .C(
        n53628), .Y(n55567) );
  A2O1A1Ixp33_ASAP7_75t_SL U47609 ( .A1(n70842), .A2(n70862), .B(n53192), .C(
        n53628), .Y(n55558) );
  A2O1A1Ixp33_ASAP7_75t_SL U47610 ( .A1(n55559), .A2(n70849), .B(n53192), .C(
        n55558), .Y(n55560) );
  A2O1A1Ixp33_ASAP7_75t_SL U47611 ( .A1(n57211), .A2(n55561), .B(n53192), .C(
        n53628), .Y(n55562) );
  A2O1A1Ixp33_ASAP7_75t_SL U47612 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[12]), .A2(n57204), .B(
        n53192), .C(n53628), .Y(n55776) );
  A2O1A1Ixp33_ASAP7_75t_SL U47613 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]), .A2(n57205), .B(
        n53192), .C(n53628), .Y(n55777) );
  A2O1A1Ixp33_ASAP7_75t_SL U47614 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[14]), .A2(n57217), .B(
        n53192), .C(n53628), .Y(n55778) );
  A2O1A1Ixp33_ASAP7_75t_SL U47615 ( .A1(n55776), .A2(n55777), .B(n53192), .C(
        n55778), .Y(n55779) );
  A2O1A1Ixp33_ASAP7_75t_SL U47616 ( .A1(n73687), .A2(n59632), .B(n53192), .C(
        n53628), .Y(n55771) );
  A2O1A1Ixp33_ASAP7_75t_SL U47617 ( .A1(n73688), .A2(n57204), .B(n53192), .C(
        n53628), .Y(n55772) );
  A2O1A1Ixp33_ASAP7_75t_SL U47618 ( .A1(n55771), .A2(n55772), .B(n53192), .C(
        n53628), .Y(n55773) );
  A2O1A1Ixp33_ASAP7_75t_SL U47619 ( .A1(n73774), .A2(n57205), .B(n53192), .C(
        n53628), .Y(n55775) );
  A2O1A1Ixp33_ASAP7_75t_SL U47620 ( .A1(n55774), .A2(n55775), .B(n53192), .C(
        n53628), .Y(n73754) );
  A2O1A1Ixp33_ASAP7_75t_SL U47621 ( .A1(n75298), .A2(n75299), .B(n53192), .C(
        n53628), .Y(n55317) );
  A2O1A1Ixp33_ASAP7_75t_SL U47622 ( .A1(n54076), .A2(n54077), .B(n53192), .C(
        n53628), .Y(n68999) );
  A2O1A1Ixp33_ASAP7_75t_SL U47623 ( .A1(n2781), .A2(n55752), .B(n53192), .C(
        n53628), .Y(n77831) );
  A2O1A1Ixp33_ASAP7_75t_SL U47624 ( .A1(n74238), .A2(n55749), .B(n53192), .C(
        n53628), .Y(n74274) );
  A2O1A1Ixp33_ASAP7_75t_SL U47625 ( .A1(n55745), .A2(n71501), .B(n53192), .C(
        n53628), .Y(n71604) );
  A2O1A1Ixp33_ASAP7_75t_SL U47626 ( .A1(n66051), .A2(n65954), .B(n53192), .C(
        n53628), .Y(n55737) );
  A2O1A1Ixp33_ASAP7_75t_SL U47627 ( .A1(n65978), .A2(n65951), .B(n53192), .C(
        n53628), .Y(n55740) );
  A2O1A1Ixp33_ASAP7_75t_SL U47628 ( .A1(n55739), .A2(n55740), .B(n53192), .C(
        n53628), .Y(n66059) );
  A2O1A1Ixp33_ASAP7_75t_SL U47629 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[25]), .A2(
        n59631), .B(n53192), .C(n53628), .Y(n55507) );
  A2O1A1Ixp33_ASAP7_75t_SL U47630 ( .A1(n77060), .A2(n55732), .B(n53192), .C(
        n53628), .Y(n62275) );
  A2O1A1Ixp33_ASAP7_75t_SL U47631 ( .A1(n62910), .A2(n62909), .B(n53192), .C(
        n53628), .Y(n55728) );
  A2O1A1Ixp33_ASAP7_75t_SL U47632 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n55718) );
  A2O1A1Ixp33_ASAP7_75t_SL U47633 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n55719) );
  A2O1A1Ixp33_ASAP7_75t_SL U47634 ( .A1(n55718), .A2(n55719), .B(n53192), .C(
        n53628), .Y(n55720) );
  A2O1A1Ixp33_ASAP7_75t_SL U47635 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n55722) );
  A2O1A1Ixp33_ASAP7_75t_SL U47636 ( .A1(n55721), .A2(n55722), .B(n53192), .C(
        n53628), .Y(n72040) );
  A2O1A1Ixp33_ASAP7_75t_SL U47637 ( .A1(n65578), .A2(n65805), .B(n53192), .C(
        n53628), .Y(n55716) );
  A2O1A1Ixp33_ASAP7_75t_SL U47638 ( .A1(n61732), .A2(n55714), .B(n53192), .C(
        n55715), .Y(n76771) );
  A2O1A1Ixp33_ASAP7_75t_SL U47639 ( .A1(n75644), .A2(n57365), .B(n53192), .C(
        n57078), .Y(n55711) );
  A2O1A1Ixp33_ASAP7_75t_SL U47640 ( .A1(n64607), .A2(n64605), .B(n53192), .C(
        n64606), .Y(n55710) );
  A2O1A1Ixp33_ASAP7_75t_SL U47641 ( .A1(n66474), .A2(n55706), .B(n53192), .C(
        n53628), .Y(n55707) );
  A2O1A1Ixp33_ASAP7_75t_SL U47642 ( .A1(n72674), .A2(n55480), .B(n53192), .C(
        n53628), .Y(n55481) );
  A2O1A1Ixp33_ASAP7_75t_SL U47643 ( .A1(n55481), .A2(n72675), .B(n53192), .C(
        n53628), .Y(n55482) );
  A2O1A1Ixp33_ASAP7_75t_SL U47644 ( .A1(n73470), .A2(n53463), .B(n53192), .C(
        n53628), .Y(n55702) );
  A2O1A1Ixp33_ASAP7_75t_SL U47645 ( .A1(n70059), .A2(n69872), .B(n53192), .C(
        n53628), .Y(n55692) );
  A2O1A1Ixp33_ASAP7_75t_SL U47646 ( .A1(n61997), .A2(n55245), .B(n53192), .C(
        n53628), .Y(n9381) );
  A2O1A1Ixp33_ASAP7_75t_SL U47647 ( .A1(n59694), .A2(n55476), .B(n53192), .C(
        n53628), .Y(n55477) );
  A2O1A1Ixp33_ASAP7_75t_SL U47648 ( .A1(n59694), .A2(n55687), .B(n53192), .C(
        n53628), .Y(n55688) );
  A2O1A1Ixp33_ASAP7_75t_SL U47649 ( .A1(n74854), .A2(n77195), .B(n53192), .C(
        n55681), .Y(n52496) );
  A2O1A1Ixp33_ASAP7_75t_SL U47650 ( .A1(n77458), .A2(n57073), .B(n53192), .C(
        n53628), .Y(n55679) );
  A2O1A1Ixp33_ASAP7_75t_SL U47651 ( .A1(n57198), .A2(n77002), .B(n53192), .C(
        n53628), .Y(n55467) );
  A2O1A1Ixp33_ASAP7_75t_SL U47652 ( .A1(n69378), .A2(n55671), .B(n53192), .C(
        n53628), .Y(n9562) );
  A2O1A1Ixp33_ASAP7_75t_SL U47653 ( .A1(n70486), .A2(n70542), .B(n53192), .C(
        n53628), .Y(n55446) );
  A2O1A1Ixp33_ASAP7_75t_SL U47654 ( .A1(n53628), .A2(n70468), .B(n53192), .C(
        n53628), .Y(n55455) );
  A2O1A1Ixp33_ASAP7_75t_SL U47655 ( .A1(n55458), .A2(n55459), .B(n53192), .C(
        n53628), .Y(n55460) );
  A2O1A1Ixp33_ASAP7_75t_SL U47656 ( .A1(n54837), .A2(n54838), .B(n53192), .C(
        n53628), .Y(n54839) );
  A2O1A1Ixp33_ASAP7_75t_SL U47657 ( .A1(n61161), .A2(n59692), .B(n53192), .C(
        n53628), .Y(n55442) );
  A2O1A1Ixp33_ASAP7_75t_SL U47658 ( .A1(n77926), .A2(n59691), .B(n53192), .C(
        n53628), .Y(n54833) );
  A2O1A1Ixp33_ASAP7_75t_SL U47659 ( .A1(n59628), .A2(n78429), .B(n53192), .C(
        n53628), .Y(n55665) );
  A2O1A1Ixp33_ASAP7_75t_SL U47660 ( .A1(n77201), .A2(n76609), .B(n53192), .C(
        n53628), .Y(n55664) );
  A2O1A1Ixp33_ASAP7_75t_SL U47661 ( .A1(n77246), .A2(n77918), .B(n53192), .C(
        n53628), .Y(n55662) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47662 ( .A1(or1200_cpu_except_type_1_), .A2(
        n74933), .B(n53192), .C(n76826), .D(n55661), .Y(n9491) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47663 ( .A1(n77674), .A2(n77676), .B(n53192), 
        .C(n77675), .D(n55657), .Y(n1696) );
  A2O1A1Ixp33_ASAP7_75t_SL U47664 ( .A1(n57114), .A2(n77983), .B(n53192), .C(
        n53628), .Y(n55655) );
  A2O1A1Ixp33_ASAP7_75t_SL U47665 ( .A1(n77916), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n55426) );
  A2O1A1Ixp33_ASAP7_75t_SL U47666 ( .A1(n57142), .A2(n77981), .B(n53192), .C(
        n53628), .Y(n55649) );
  A2O1A1Ixp33_ASAP7_75t_SL U47667 ( .A1(n77982), .A2(n55650), .B(n53192), .C(
        n53628), .Y(n55651) );
  A2O1A1Ixp33_ASAP7_75t_SL U47668 ( .A1(n77856), .A2(n75649), .B(n53192), .C(
        n53628), .Y(n55418) );
  A2O1A1Ixp33_ASAP7_75t_SL U47669 ( .A1(n53192), .A2(n53628), .B(n55402), .C(
        n53628), .Y(n55403) );
  A2O1A1Ixp33_ASAP7_75t_SL U47670 ( .A1(n53628), .A2(n63277), .B(n53192), .C(
        n55403), .Y(n55409) );
  A2O1A1Ixp33_ASAP7_75t_SL U47671 ( .A1(n53628), .A2(n55409), .B(n53192), .C(
        n53628), .Y(n55410) );
  A2O1A1Ixp33_ASAP7_75t_SL U47672 ( .A1(n59656), .A2(n53331), .B(n53192), .C(
        n53628), .Y(n55400) );
  A2O1A1Ixp33_ASAP7_75t_SL U47673 ( .A1(n68932), .A2(n75650), .B(n53192), .C(
        n53628), .Y(n55631) );
  A2O1A1Ixp33_ASAP7_75t_SL U47674 ( .A1(n77977), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n55632) );
  A2O1A1Ixp33_ASAP7_75t_SL U47675 ( .A1(n68931), .A2(n68912), .B(n53192), .C(
        n53628), .Y(n55635) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47676 ( .A1(n68935), .A2(n57079), .B(n53192), 
        .C(n55635), .D(n55637), .Y(n55639) );
  A2O1A1Ixp33_ASAP7_75t_SL U47677 ( .A1(n55631), .A2(n55632), .B(n53192), .C(
        n55641), .Y(or1200_cpu_or1200_mult_mac_n1619) );
  A2O1A1Ixp33_ASAP7_75t_SL U47678 ( .A1(n55622), .A2(n55623), .B(n53192), .C(
        n53628), .Y(n55624) );
  A2O1A1Ixp33_ASAP7_75t_SL U47679 ( .A1(n75650), .A2(n69110), .B(n53192), .C(
        n53628), .Y(n55630) );
  A2O1A1Ixp33_ASAP7_75t_SL U47680 ( .A1(n55629), .A2(n55630), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1612) );
  A2O1A1Ixp33_ASAP7_75t_SL U47681 ( .A1(n74568), .A2(n74569), .B(n53192), .C(
        n53628), .Y(n55609) );
  A2O1A1Ixp33_ASAP7_75t_SL U47682 ( .A1(n55616), .A2(n59672), .B(n53192), .C(
        n53628), .Y(n55617) );
  A2O1A1Ixp33_ASAP7_75t_SL U47683 ( .A1(n55615), .A2(n55617), .B(n53192), .C(
        n53628), .Y(n55618) );
  A2O1A1Ixp33_ASAP7_75t_SL U47684 ( .A1(n75650), .A2(n74573), .B(n53192), .C(
        n53628), .Y(n55620) );
  A2O1A1Ixp33_ASAP7_75t_SL U47685 ( .A1(n77883), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n55621) );
  A2O1A1Ixp33_ASAP7_75t_SL U47686 ( .A1(n55619), .A2(n55620), .B(n53192), .C(
        n55621), .Y(or1200_cpu_or1200_mult_mac_n1605) );
  A2O1A1Ixp33_ASAP7_75t_SL U47687 ( .A1(n77440), .A2(n55605), .B(n53192), .C(
        n53628), .Y(n55606) );
  A2O1A1Ixp33_ASAP7_75t_SL U47688 ( .A1(n76619), .A2(n57074), .B(n53192), .C(
        n53628), .Y(n54994) );
  A2O1A1Ixp33_ASAP7_75t_SL U47689 ( .A1(n59693), .A2(n77153), .B(n53192), .C(
        n53628), .Y(n55604) );
  A2O1A1Ixp33_ASAP7_75t_SL U47690 ( .A1(n59693), .A2(n77179), .B(n53192), .C(
        n53628), .Y(n55601) );
  A2O1A1Ixp33_ASAP7_75t_SL U47691 ( .A1(n57072), .A2(n77227), .B(n53192), .C(
        n53628), .Y(n55600) );
  A2O1A1Ixp33_ASAP7_75t_SL U47692 ( .A1(n75433), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n54127) );
  A2O1A1Ixp33_ASAP7_75t_SL U47693 ( .A1(n57072), .A2(n75200), .B(n53192), .C(
        n53628), .Y(n55598) );
  A2O1A1Ixp33_ASAP7_75t_SL U47694 ( .A1(n74239), .A2(n55593), .B(n53192), .C(
        n53628), .Y(n55594) );
  A2O1A1Ixp33_ASAP7_75t_SL U47695 ( .A1(n74275), .A2(n55594), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n49) );
  A2O1A1Ixp33_ASAP7_75t_SL U47696 ( .A1(n72390), .A2(n55588), .B(n53192), .C(
        n53628), .Y(n55589) );
  A2O1A1Ixp33_ASAP7_75t_SL U47697 ( .A1(n72515), .A2(n72269), .B(n53192), .C(
        n55589), .Y(n55590) );
  A2O1A1Ixp33_ASAP7_75t_SL U47698 ( .A1(n71547), .A2(n55578), .B(n53192), .C(
        n71612), .Y(n55579) );
  A2O1A1Ixp33_ASAP7_75t_SL U47699 ( .A1(n55573), .A2(n55579), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n135) );
  A2O1A1Ixp33_ASAP7_75t_SL U47700 ( .A1(n59699), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55569) );
  A2O1A1Ixp33_ASAP7_75t_SL U47701 ( .A1(n70714), .A2(n55569), .B(n53192), .C(
        n53628), .Y(n55570) );
  A2O1A1Ixp33_ASAP7_75t_SL U47702 ( .A1(n70713), .A2(n55570), .B(n53192), .C(
        n53628), .Y(n55571) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47703 ( .A1(n70805), .A2(n55563), .B(n53192), 
        .C(n70794), .D(n55564), .Y(n55565) );
  A2O1A1Ixp33_ASAP7_75t_SL U47704 ( .A1(n55137), .A2(n55138), .B(n53192), .C(
        n53628), .Y(n55139) );
  A2O1A1Ixp33_ASAP7_75t_SL U47705 ( .A1(n55140), .A2(n55141), .B(n53192), .C(
        n53628), .Y(n73772) );
  A2O1A1Ixp33_ASAP7_75t_SL U47706 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[12]), .A2(n57205), .B(
        n53192), .C(n53628), .Y(n55133) );
  A2O1A1Ixp33_ASAP7_75t_SL U47707 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[11]), .A2(n57204), .B(
        n53192), .C(n53628), .Y(n55134) );
  A2O1A1Ixp33_ASAP7_75t_SL U47708 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]), .A2(n57217), .B(
        n53192), .C(n53628), .Y(n55135) );
  A2O1A1Ixp33_ASAP7_75t_SL U47709 ( .A1(n55133), .A2(n55134), .B(n53192), .C(
        n55135), .Y(n55136) );
  A2O1A1Ixp33_ASAP7_75t_SL U47710 ( .A1(n2765), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55549) );
  A2O1A1Ixp33_ASAP7_75t_SL U47711 ( .A1(n60277), .A2(n55549), .B(n53192), .C(
        n53628), .Y(n55550) );
  A2O1A1Ixp33_ASAP7_75t_SL U47712 ( .A1(n60278), .A2(n55550), .B(n53192), .C(
        n53628), .Y(n60279) );
  A2O1A1Ixp33_ASAP7_75t_SL U47713 ( .A1(n62060), .A2(n62036), .B(n53192), .C(
        n53628), .Y(n55543) );
  A2O1A1Ixp33_ASAP7_75t_SL U47714 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_0_), .A2(n62046), .B(n53192), 
        .C(n53628), .Y(n55545) );
  A2O1A1Ixp33_ASAP7_75t_SL U47715 ( .A1(n62041), .A2(n74817), .B(n53192), .C(
        n53628), .Y(n55546) );
  A2O1A1Ixp33_ASAP7_75t_SL U47716 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_5_), .A2(n62060), .B(n53192), 
        .C(n62054), .Y(n55547) );
  A2O1A1Ixp33_ASAP7_75t_SL U47717 ( .A1(n75763), .A2(n75764), .B(n53192), .C(
        n53628), .Y(n55542) );
  A2O1A1Ixp33_ASAP7_75t_SL U47718 ( .A1(n62477), .A2(dbg_dat_i[16]), .B(n53192), .C(n53628), .Y(n55541) );
  A2O1A1Ixp33_ASAP7_75t_SL U47719 ( .A1(n62477), .A2(dbg_dat_i[24]), .B(n53192), .C(n53628), .Y(n55540) );
  A2O1A1Ixp33_ASAP7_75t_SL U47720 ( .A1(n74646), .A2(n2345), .B(n53192), .C(
        n55539), .Y(n74694) );
  A2O1A1Ixp33_ASAP7_75t_SL U47721 ( .A1(n62477), .A2(dbg_dat_i[22]), .B(n53192), .C(n53628), .Y(n55538) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47722 ( .A1(n78001), .A2(n3082), .B(n53192), .C(
        n1185), .D(n55525), .Y(n78174) );
  A2O1A1Ixp33_ASAP7_75t_SL U47723 ( .A1(n66024), .A2(n65954), .B(n53192), .C(
        n53628), .Y(n55509) );
  A2O1A1Ixp33_ASAP7_75t_SL U47724 ( .A1(n66051), .A2(n65959), .B(n53192), .C(
        n53628), .Y(n55510) );
  A2O1A1Ixp33_ASAP7_75t_SL U47725 ( .A1(n55509), .A2(n55510), .B(n53192), .C(
        n53628), .Y(n55511) );
  A2O1A1Ixp33_ASAP7_75t_SL U47726 ( .A1(n65978), .A2(n65901), .B(n53192), .C(
        n53628), .Y(n55513) );
  A2O1A1Ixp33_ASAP7_75t_SL U47727 ( .A1(n55512), .A2(n55513), .B(n53192), .C(
        n53628), .Y(n65988) );
  A2O1A1Ixp33_ASAP7_75t_SL U47728 ( .A1(n70185), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55505) );
  A2O1A1Ixp33_ASAP7_75t_SL U47729 ( .A1(n70183), .A2(n55505), .B(n53192), .C(
        n53628), .Y(n55506) );
  A2O1A1Ixp33_ASAP7_75t_SL U47730 ( .A1(n70184), .A2(n55506), .B(n53192), .C(
        n53628), .Y(n70194) );
  A2O1A1Ixp33_ASAP7_75t_SL U47731 ( .A1(
        or1200_cpu_or1200_genpc_pcreg_default[6]), .A2(
        or1200_cpu_or1200_genpc_pcreg_default[5]), .B(n53192), .C(n53628), .Y(
        n55284) );
  A2O1A1Ixp33_ASAP7_75t_SL U47732 ( .A1(n74957), .A2(n55501), .B(n53192), .C(
        n53628), .Y(n63939) );
  A2O1A1Ixp33_ASAP7_75t_SL U47733 ( .A1(n64743), .A2(n64749), .B(n53192), .C(
        n53628), .Y(n55499) );
  A2O1A1Ixp33_ASAP7_75t_SL U47734 ( .A1(n64746), .A2(n55499), .B(n53192), .C(
        n53628), .Y(n55500) );
  A2O1A1Ixp33_ASAP7_75t_SL U47735 ( .A1(n71270), .A2(n71271), .B(n53192), .C(
        n55497), .Y(n71206) );
  A2O1A1Ixp33_ASAP7_75t_SL U47736 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[6]), .A2(n73047), .B(n53192), .C(n53628), .Y(n54548) );
  A2O1A1Ixp33_ASAP7_75t_SL U47737 ( .A1(n76350), .A2(n60980), .B(n53192), .C(
        n53628), .Y(n55495) );
  A2O1A1Ixp33_ASAP7_75t_SL U47738 ( .A1(n77091), .A2(
        or1200_cpu_or1200_fpu_result_arith[23]), .B(n53192), .C(n53628), .Y(
        n55492) );
  A2O1A1Ixp33_ASAP7_75t_SL U47739 ( .A1(n59229), .A2(n66964), .B(n53192), .C(
        n53628), .Y(n55488) );
  A2O1A1Ixp33_ASAP7_75t_SL U47740 ( .A1(n57108), .A2(n57244), .B(n53192), .C(
        n53628), .Y(n55485) );
  A2O1A1Ixp33_ASAP7_75t_SL U47741 ( .A1(n73581), .A2(n73562), .B(n53192), .C(
        n53628), .Y(n54713) );
  A2O1A1Ixp33_ASAP7_75t_SL U47742 ( .A1(n69873), .A2(n69996), .B(n53192), .C(
        n53628), .Y(n55246) );
  A2O1A1Ixp33_ASAP7_75t_SL U47743 ( .A1(n54865), .A2(n54867), .B(n53192), .C(
        n53628), .Y(n54868) );
  A2O1A1Ixp33_ASAP7_75t_SL U47744 ( .A1(n54868), .A2(n54870), .B(n53192), .C(
        n53628), .Y(n3174) );
  A2O1A1Ixp33_ASAP7_75t_SL U47745 ( .A1(n77458), .A2(n55241), .B(n53192), .C(
        n53628), .Y(n55242) );
  A2O1A1Ixp33_ASAP7_75t_SL U47746 ( .A1(n77460), .A2(n77459), .B(n53192), .C(
        n53628), .Y(n55243) );
  A2O1A1Ixp33_ASAP7_75t_SL U47747 ( .A1(n53628), .A2(n76517), .B(n53192), .C(
        n53628), .Y(n55474) );
  A2O1A1Ixp33_ASAP7_75t_SL U47748 ( .A1(n76519), .A2(n55474), .B(n53192), .C(
        n53628), .Y(n55475) );
  A2O1A1Ixp33_ASAP7_75t_SL U47749 ( .A1(n76518), .A2(n55475), .B(n53192), .C(
        n53628), .Y(n55476) );
  A2O1A1Ixp33_ASAP7_75t_SL U47750 ( .A1(n57144), .A2(n75544), .B(n53192), .C(
        n53628), .Y(n55059) );
  A2O1A1Ixp33_ASAP7_75t_SL U47751 ( .A1(n77212), .A2(n77974), .B(n53192), .C(
        n53628), .Y(n55468) );
  A2O1A1Ixp33_ASAP7_75t_SL U47752 ( .A1(n55467), .A2(n55468), .B(n53192), .C(
        n53628), .Y(n55469) );
  A2O1A1Ixp33_ASAP7_75t_SL U47753 ( .A1(n53628), .A2(n55469), .B(n53192), .C(
        n53628), .Y(n55470) );
  A2O1A1Ixp33_ASAP7_75t_SL U47754 ( .A1(n59691), .A2(n55235), .B(n53192), .C(
        n53628), .Y(n55236) );
  A2O1A1Ixp33_ASAP7_75t_SL U47755 ( .A1(n55454), .A2(n55456), .B(n53192), .C(
        n55457), .Y(n55458) );
  A2O1A1Ixp33_ASAP7_75t_SL U47756 ( .A1(n70476), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_3_), .B(
        n53192), .C(n53628), .Y(n55459) );
  A2O1A1Ixp33_ASAP7_75t_SL U47757 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[8]), .B(n53192), 
        .C(n53628), .Y(n55225) );
  A2O1A1Ixp33_ASAP7_75t_SL U47758 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[8]), .A2(n55226), 
        .B(n53192), .C(n53628), .Y(n55227) );
  A2O1A1Ixp33_ASAP7_75t_SL U47759 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[8]), .B(
        n53192), .C(n53628), .Y(n55228) );
  A2O1A1Ixp33_ASAP7_75t_SL U47760 ( .A1(n55225), .A2(n55227), .B(n53192), .C(
        n55228), .Y(or1200_cpu_or1200_fpu_fpu_arith_N91) );
  A2O1A1Ixp33_ASAP7_75t_SL U47761 ( .A1(n59693), .A2(n55440), .B(n53192), .C(
        n53628), .Y(n55441) );
  A2O1A1Ixp33_ASAP7_75t_SL U47762 ( .A1(n78339), .A2(n73047), .B(n53192), .C(
        n53628), .Y(n55219) );
  A2O1A1Ixp33_ASAP7_75t_SL U47763 ( .A1(n77201), .A2(n77206), .B(n53192), .C(
        n53628), .Y(n55437) );
  A2O1A1Ixp33_ASAP7_75t_SL U47764 ( .A1(n55436), .A2(n55437), .B(n53192), .C(
        n53628), .Y(or1200_du_N105) );
  A2O1A1Ixp33_ASAP7_75t_SL U47765 ( .A1(n77582), .A2(n77644), .B(n53192), .C(
        n53628), .Y(n55433) );
  A2O1A1Ixp33_ASAP7_75t_SL U47766 ( .A1(n57114), .A2(n77986), .B(n53192), .C(
        n53628), .Y(n55432) );
  A2O1A1Ixp33_ASAP7_75t_SL U47767 ( .A1(n1418), .A2(n55427), .B(n53192), .C(
        n53628), .Y(n55428) );
  A2O1A1Ixp33_ASAP7_75t_SL U47768 ( .A1(n77287), .A2(n76688), .B(n53192), .C(
        n53628), .Y(n55429) );
  A2O1A1Ixp33_ASAP7_75t_SL U47769 ( .A1(n55428), .A2(n55429), .B(n53192), .C(
        n53628), .Y(n55430) );
  A2O1A1Ixp33_ASAP7_75t_SL U47770 ( .A1(n55430), .A2(n55431), .B(n53192), .C(
        n53628), .Y(or1200_pic_N49) );
  A2O1A1Ixp33_ASAP7_75t_SL U47771 ( .A1(n77980), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n55214) );
  A2O1A1Ixp33_ASAP7_75t_SL U47772 ( .A1(n1398), .A2(n55421), .B(n53192), .C(
        n53628), .Y(n55422) );
  A2O1A1Ixp33_ASAP7_75t_SL U47773 ( .A1(n77287), .A2(n77603), .B(n53192), .C(
        n53628), .Y(n55423) );
  A2O1A1Ixp33_ASAP7_75t_SL U47774 ( .A1(n55422), .A2(n55423), .B(n53192), .C(
        n53628), .Y(n55424) );
  A2O1A1Ixp33_ASAP7_75t_SL U47775 ( .A1(n55424), .A2(n55425), .B(n53192), .C(
        n53628), .Y(or1200_pic_N54) );
  A2O1A1Ixp33_ASAP7_75t_SL U47776 ( .A1(n77899), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n55012) );
  A2O1A1Ixp33_ASAP7_75t_SL U47777 ( .A1(n55210), .A2(n55212), .B(n53192), .C(
        n53628), .Y(n9355) );
  A2O1A1Ixp33_ASAP7_75t_SL U47778 ( .A1(n55207), .A2(n55209), .B(n53192), .C(
        n53628), .Y(n9352) );
  A2O1A1Ixp33_ASAP7_75t_SL U47779 ( .A1(or1200_cpu_or1200_mult_mac_div_cntr_2_), .A2(n53628), .B(n53192), .C(n53628), .Y(n55201) );
  A2O1A1Ixp33_ASAP7_75t_SL U47780 ( .A1(n61811), .A2(n55202), .B(n53192), .C(
        n53628), .Y(n55203) );
  A2O1A1Ixp33_ASAP7_75t_SL U47781 ( .A1(n76884), .A2(n55385), .B(n53192), .C(
        n53628), .Y(n55386) );
  A2O1A1Ixp33_ASAP7_75t_SL U47782 ( .A1(n76886), .A2(n55387), .B(n53192), .C(
        n53628), .Y(n55388) );
  A2O1A1Ixp33_ASAP7_75t_SL U47783 ( .A1(n55384), .A2(n55392), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1562) );
  A2O1A1Ixp33_ASAP7_75t_SL U47784 ( .A1(n53192), .A2(n53628), .B(n55182), .C(
        n53628), .Y(n55183) );
  A2O1A1Ixp33_ASAP7_75t_SL U47785 ( .A1(n77880), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n54796) );
  A2O1A1Ixp33_ASAP7_75t_SL U47786 ( .A1(n74114), .A2(n75650), .B(n53192), .C(
        n53628), .Y(n54797) );
  A2O1A1Ixp33_ASAP7_75t_SL U47787 ( .A1(n54796), .A2(n54797), .B(n53192), .C(
        n54801), .Y(or1200_cpu_or1200_mult_mac_n1604) );
  A2O1A1Ixp33_ASAP7_75t_SL U47788 ( .A1(n75650), .A2(n55374), .B(n53192), .C(
        n53628), .Y(n55375) );
  A2O1A1Ixp33_ASAP7_75t_SL U47789 ( .A1(n77871), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n55376) );
  A2O1A1Ixp33_ASAP7_75t_SL U47790 ( .A1(n55375), .A2(n55376), .B(n53192), .C(
        n55382), .Y(or1200_cpu_or1200_mult_mac_n1600) );
  A2O1A1Ixp33_ASAP7_75t_SL U47791 ( .A1(n57093), .A2(n77277), .B(n53192), .C(
        n53628), .Y(n55371) );
  A2O1A1Ixp33_ASAP7_75t_SL U47792 ( .A1(n57072), .A2(n76232), .B(n53192), .C(
        n53628), .Y(n55370) );
  A2O1A1Ixp33_ASAP7_75t_SL U47793 ( .A1(n57072), .A2(n75798), .B(n53192), .C(
        n53628), .Y(n55368) );
  A2O1A1Ixp33_ASAP7_75t_SL U47794 ( .A1(n59690), .A2(n76676), .B(n53192), .C(
        n53628), .Y(n55362) );
  A2O1A1Ixp33_ASAP7_75t_SL U47795 ( .A1(n55361), .A2(n55362), .B(n53192), .C(
        n53628), .Y(n55363) );
  A2O1A1Ixp33_ASAP7_75t_SL U47796 ( .A1(or1200_cpu_or1200_except_n684), .A2(
        or1200_cpu_or1200_except_n687), .B(n53192), .C(n53628), .Y(n55364) );
  A2O1A1Ixp33_ASAP7_75t_SL U47797 ( .A1(n76677), .A2(n55363), .B(n53192), .C(
        n55364), .Y(n55365) );
  A2O1A1Ixp33_ASAP7_75t_SL U47798 ( .A1(n57343), .A2(n55365), .B(n53192), .C(
        n53628), .Y(n55366) );
  A2O1A1Ixp33_ASAP7_75t_SL U47799 ( .A1(n58447), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_), 
        .B(n53192), .C(n53628), .Y(n55344) );
  A2O1A1Ixp33_ASAP7_75t_SL U47800 ( .A1(n55343), .A2(n55344), .B(n53192), .C(
        n53628), .Y(n55345) );
  A2O1A1Ixp33_ASAP7_75t_SL U47801 ( .A1(n72502), .A2(n55345), .B(n53192), .C(
        n53628), .Y(n55346) );
  A2O1A1Ixp33_ASAP7_75t_SL U47802 ( .A1(n54973), .A2(n54975), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n115) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47803 ( .A1(n70842), .A2(n70849), .B(n53192), 
        .C(n55336), .D(n55337), .Y(n55338) );
  A2O1A1Ixp33_ASAP7_75t_SL U47804 ( .A1(n55328), .A2(n55332), .B(n53192), .C(
        n53628), .Y(n55333) );
  A2O1A1Ixp33_ASAP7_75t_SL U47805 ( .A1(n73697), .A2(n57204), .B(n53192), .C(
        n53628), .Y(n54768) );
  A2O1A1Ixp33_ASAP7_75t_SL U47806 ( .A1(n54770), .A2(n54771), .B(n53192), .C(
        n53628), .Y(n73785) );
  A2O1A1Ixp33_ASAP7_75t_SL U47807 ( .A1(n77752), .A2(n77751), .B(n53192), .C(
        n53628), .Y(n55319) );
  A2O1A1Ixp33_ASAP7_75t_SL U47808 ( .A1(n77754), .A2(n77753), .B(n53192), .C(
        n55319), .Y(n55320) );
  A2O1A1Ixp33_ASAP7_75t_SL U47809 ( .A1(n77760), .A2(n55320), .B(n53192), .C(
        n53628), .Y(n3905) );
  A2O1A1Ixp33_ASAP7_75t_SL U47810 ( .A1(n53628), .A2(n75300), .B(n53192), .C(
        n53628), .Y(n55315) );
  A2O1A1Ixp33_ASAP7_75t_SL U47811 ( .A1(n75297), .A2(n55315), .B(n53192), .C(
        n53628), .Y(n55316) );
  A2O1A1Ixp33_ASAP7_75t_SL U47812 ( .A1(n55316), .A2(n55317), .B(n53192), .C(
        n53628), .Y(n78133) );
  A2O1A1Ixp33_ASAP7_75t_SL U47813 ( .A1(n76144), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55311) );
  A2O1A1Ixp33_ASAP7_75t_SL U47814 ( .A1(n76123), .A2(n55311), .B(n53192), .C(
        n53628), .Y(n55312) );
  A2O1A1Ixp33_ASAP7_75t_SL U47815 ( .A1(n53628), .A2(n55312), .B(n53192), .C(
        n53628), .Y(n76137) );
  A2O1A1Ixp33_ASAP7_75t_SL U47816 ( .A1(n65163), .A2(n65162), .B(n53192), .C(
        n53628), .Y(n55310) );
  A2O1A1Ixp33_ASAP7_75t_SL U47817 ( .A1(n57216), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_2_), 
        .B(n53192), .C(n53628), .Y(n54740) );
  A2O1A1Ixp33_ASAP7_75t_SL U47818 ( .A1(n57216), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_32_), 
        .B(n53192), .C(n53628), .Y(n54244) );
  A2O1A1Ixp33_ASAP7_75t_SL U47819 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n55299) );
  A2O1A1Ixp33_ASAP7_75t_SL U47820 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n55300) );
  A2O1A1Ixp33_ASAP7_75t_SL U47821 ( .A1(n55299), .A2(n55300), .B(n53192), .C(
        n53628), .Y(n55301) );
  A2O1A1Ixp33_ASAP7_75t_SL U47822 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n55303) );
  A2O1A1Ixp33_ASAP7_75t_SL U47823 ( .A1(n55302), .A2(n55303), .B(n53192), .C(
        n53628), .Y(n72090) );
  A2O1A1Ixp33_ASAP7_75t_SL U47824 ( .A1(n72054), .A2(n72132), .B(n53192), .C(
        n53628), .Y(n55296) );
  A2O1A1Ixp33_ASAP7_75t_SL U47825 ( .A1(n71485), .A2(n55297), .B(n53192), .C(
        n53628), .Y(n71496) );
  A2O1A1Ixp33_ASAP7_75t_SL U47826 ( .A1(n71072), .A2(n71071), .B(n53192), .C(
        n53628), .Y(n55294) );
  A2O1A1Ixp33_ASAP7_75t_SL U47827 ( .A1(n61672), .A2(n55290), .B(n53192), .C(
        n53628), .Y(n55291) );
  A2O1A1Ixp33_ASAP7_75t_SL U47828 ( .A1(n57121), .A2(n63490), .B(n53192), .C(
        n53628), .Y(n55289) );
  A2O1A1Ixp33_ASAP7_75t_SL U47829 ( .A1(n57321), .A2(n75046), .B(n53192), .C(
        n53628), .Y(n55282) );
  A2O1A1Ixp33_ASAP7_75t_SL U47830 ( .A1(or1200_cpu_or1200_mult_mac_n305), .A2(
        or1200_cpu_or1200_mult_mac_n159), .B(n53192), .C(n53628), .Y(n55281)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U47831 ( .A1(n63433), .A2(n55281), .B(n53192), .C(
        n53628), .Y(n63458) );
  A2O1A1Ixp33_ASAP7_75t_SL U47832 ( .A1(n58418), .A2(n65781), .B(n53192), .C(
        n53628), .Y(n55276) );
  A2O1A1Ixp33_ASAP7_75t_SL U47833 ( .A1(n57190), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[16]), .B(n53192), .C(n53628), .Y(n55273) );
  A2O1A1Ixp33_ASAP7_75t_SL U47834 ( .A1(n59526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_0_), .B(n53192), .C(
        n53473), .Y(n58307) );
  A2O1A1Ixp33_ASAP7_75t_SL U47835 ( .A1(n67882), .A2(n63156), .B(n53192), .C(
        n53628), .Y(n55263) );
  A2O1A1Ixp33_ASAP7_75t_SL U47836 ( .A1(n59604), .A2(n67920), .B(n53192), .C(
        n53628), .Y(n54539) );
  A2O1A1Ixp33_ASAP7_75t_SL U47837 ( .A1(n67564), .A2(n58851), .B(n53192), .C(
        n53628), .Y(n55257) );
  A2O1A1Ixp33_ASAP7_75t_SL U47838 ( .A1(n55252), .A2(n55253), .B(n53192), .C(
        n53628), .Y(n3285) );
  A2O1A1Ixp33_ASAP7_75t_SL U47839 ( .A1(n69872), .A2(n69997), .B(n53192), .C(
        n53628), .Y(n55247) );
  A2O1A1Ixp33_ASAP7_75t_SL U47840 ( .A1(n55246), .A2(n55247), .B(n53192), .C(
        n53628), .Y(n55248) );
  A2O1A1Ixp33_ASAP7_75t_SL U47841 ( .A1(n53628), .A2(n55248), .B(n53192), .C(
        n53628), .Y(n55249) );
  A2O1A1Ixp33_ASAP7_75t_SL U47842 ( .A1(n57198), .A2(n76866), .B(n53192), .C(
        n53628), .Y(n55047) );
  A2O1A1Ixp33_ASAP7_75t_SL U47843 ( .A1(n77915), .A2(n59691), .B(n53192), .C(
        n53628), .Y(n54856) );
  A2O1A1Ixp33_ASAP7_75t_SL U47844 ( .A1(n70529), .A2(n70530), .B(n53192), .C(
        n53628), .Y(n55229) );
  A2O1A1Ixp33_ASAP7_75t_SL U47845 ( .A1(n59692), .A2(n55220), .B(n53192), .C(
        n53628), .Y(n55221) );
  A2O1A1Ixp33_ASAP7_75t_SL U47846 ( .A1(n53192), .A2(n53628), .B(n55026), .C(
        n53628), .Y(n55027) );
  A2O1A1Ixp33_ASAP7_75t_SL U47847 ( .A1(n65237), .A2(n74934), .B(n53192), .C(
        n53628), .Y(n54328) );
  A2O1A1Ixp33_ASAP7_75t_SL U47848 ( .A1(n57114), .A2(n77922), .B(n53192), .C(
        n53628), .Y(n55216) );
  A2O1A1Ixp33_ASAP7_75t_SL U47849 ( .A1(n57142), .A2(n77975), .B(n53192), .C(
        n53628), .Y(n55210) );
  A2O1A1Ixp33_ASAP7_75t_SL U47850 ( .A1(n77976), .A2(n55211), .B(n53192), .C(
        n53628), .Y(n55212) );
  A2O1A1Ixp33_ASAP7_75t_SL U47851 ( .A1(n57142), .A2(n77984), .B(n53192), .C(
        n53628), .Y(n55207) );
  A2O1A1Ixp33_ASAP7_75t_SL U47852 ( .A1(n77985), .A2(n55208), .B(n53192), .C(
        n53628), .Y(n55209) );
  A2O1A1Ixp33_ASAP7_75t_SL U47853 ( .A1(n54811), .A2(n54813), .B(n53192), .C(
        n53628), .Y(n9245) );
  A2O1A1Ixp33_ASAP7_75t_SL U47854 ( .A1(n63447), .A2(n55006), .B(n53192), .C(
        n53628), .Y(n55007) );
  A2O1A1Ixp33_ASAP7_75t_SL U47855 ( .A1(n55007), .A2(n63363), .B(n53192), .C(
        n53628), .Y(n55008) );
  A2O1A1Ixp33_ASAP7_75t_SL U47856 ( .A1(n76631), .A2(n55201), .B(n53192), .C(
        n53628), .Y(n55202) );
  A2O1A1Ixp33_ASAP7_75t_SL U47857 ( .A1(n77893), .A2(n76888), .B(n53192), .C(
        n53628), .Y(n53976) );
  A2O1A1Ixp33_ASAP7_75t_SL U47858 ( .A1(n68849), .A2(n75650), .B(n53192), .C(
        n53628), .Y(n55192) );
  A2O1A1Ixp33_ASAP7_75t_SL U47859 ( .A1(n77918), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n55193) );
  A2O1A1Ixp33_ASAP7_75t_SL U47860 ( .A1(n68863), .A2(n68862), .B(n53192), .C(
        n53628), .Y(n55195) );
  A2O1A1Ixp33_ASAP7_75t_SL U47861 ( .A1(n57079), .A2(n55195), .B(n53192), .C(
        n53628), .Y(n55196) );
  A2O1A1Ixp33_ASAP7_75t_SL U47862 ( .A1(n55194), .A2(n55196), .B(n53192), .C(
        n53628), .Y(n55197) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47863 ( .A1(n68862), .A2(n68863), .B(n53192), 
        .C(n59672), .D(n55194), .Y(n55198) );
  A2O1A1Ixp33_ASAP7_75t_SL U47864 ( .A1(n55192), .A2(n55193), .B(n53192), .C(
        n55200), .Y(or1200_cpu_or1200_mult_mac_n1622) );
  A2O1A1Ixp33_ASAP7_75t_SL U47865 ( .A1(n75650), .A2(n75126), .B(n53192), .C(
        n53628), .Y(n55168) );
  A2O1A1Ixp33_ASAP7_75t_SL U47866 ( .A1(n77864), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n55169) );
  A2O1A1Ixp33_ASAP7_75t_SL U47867 ( .A1(n57079), .A2(n55173), .B(n53192), .C(
        n53628), .Y(n55174) );
  A2O1A1Ixp33_ASAP7_75t_SL U47868 ( .A1(n55172), .A2(n55174), .B(n53192), .C(
        n53628), .Y(n55175) );
  A2O1A1Ixp33_ASAP7_75t_SL U47869 ( .A1(n55177), .A2(n55178), .B(n53192), .C(
        n53628), .Y(n55179) );
  A2O1A1Ixp33_ASAP7_75t_SL U47870 ( .A1(n55168), .A2(n55169), .B(n53192), .C(
        n55180), .Y(or1200_cpu_or1200_mult_mac_n1597) );
  A2O1A1Ixp33_ASAP7_75t_SL U47871 ( .A1(n57093), .A2(n75312), .B(n53192), .C(
        n53628), .Y(n55165) );
  A2O1A1Ixp33_ASAP7_75t_SL U47872 ( .A1(n57093), .A2(n74578), .B(n53192), .C(
        n53628), .Y(n55164) );
  A2O1A1Ixp33_ASAP7_75t_SL U47873 ( .A1(n76671), .A2(n61157), .B(n53192), .C(
        n53628), .Y(n55160) );
  A2O1A1Ixp33_ASAP7_75t_SL U47874 ( .A1(n74275), .A2(n55159), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n51) );
  A2O1A1Ixp33_ASAP7_75t_SL U47875 ( .A1(n54983), .A2(n72500), .B(n53192), .C(
        n53628), .Y(n54984) );
  A2O1A1Ixp33_ASAP7_75t_SL U47876 ( .A1(n54971), .A2(n54972), .B(n53192), .C(
        n53628), .Y(n54973) );
  A2O1A1Ixp33_ASAP7_75t_SL U47877 ( .A1(n70862), .A2(n70875), .B(n53192), .C(
        n53628), .Y(n54962) );
  A2O1A1Ixp33_ASAP7_75t_SL U47878 ( .A1(n71026), .A2(n70873), .B(n53192), .C(
        n53628), .Y(n54963) );
  A2O1A1Ixp33_ASAP7_75t_SL U47879 ( .A1(n3321), .A2(n57204), .B(n53192), .C(
        n53628), .Y(n55137) );
  A2O1A1Ixp33_ASAP7_75t_SL U47880 ( .A1(n73696), .A2(n59632), .B(n53192), .C(
        n53628), .Y(n55138) );
  A2O1A1Ixp33_ASAP7_75t_SL U47881 ( .A1(n73687), .A2(n57205), .B(n53192), .C(
        n53628), .Y(n55141) );
  A2O1A1Ixp33_ASAP7_75t_SL U47882 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_28_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_27_), .B(
        n53192), .C(n53628), .Y(n53702) );
  A2O1A1Ixp33_ASAP7_75t_SL U47883 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_30_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_29_), .B(
        n53192), .C(n53628), .Y(n53703) );
  A2O1A1Ixp33_ASAP7_75t_SL U47884 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_25_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_26_), .B(
        n53192), .C(n53628), .Y(n53705) );
  A2O1A1Ixp33_ASAP7_75t_SL U47885 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_23_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_24_), .B(
        n53192), .C(n53628), .Y(n53706) );
  A2O1A1Ixp33_ASAP7_75t_SL U47886 ( .A1(n53704), .A2(n53707), .B(n53192), .C(
        n53628), .Y(n74460) );
  A2O1A1Ixp33_ASAP7_75t_SL U47887 ( .A1(n74706), .A2(n70431), .B(n53192), .C(
        n53628), .Y(n55131) );
  A2O1A1Ixp33_ASAP7_75t_SL U47888 ( .A1(n55130), .A2(n77760), .B(n53192), .C(
        n53628), .Y(n3903) );
  A2O1A1Ixp33_ASAP7_75t_SL U47889 ( .A1(n74802), .A2(
        or1200_cpu_or1200_fpu_fpu_conv_shr[6]), .B(n53192), .C(n53628), .Y(
        n55128) );
  A2O1A1Ixp33_ASAP7_75t_SL U47890 ( .A1(n76492), .A2(n55128), .B(n53192), .C(
        n53628), .Y(n55129) );
  A2O1A1Ixp33_ASAP7_75t_SL U47891 ( .A1(n75555), .A2(n55126), .B(n53192), .C(
        n53628), .Y(n77656) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47892 ( .A1(n55123), .A2(n75792), .B(n53192), 
        .C(n75794), .D(n55124), .Y(n78084) );
  A2O1A1Ixp33_ASAP7_75t_SL U47893 ( .A1(n63498), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55120) );
  A2O1A1Ixp33_ASAP7_75t_SL U47894 ( .A1(n63500), .A2(n55120), .B(n53192), .C(
        n53628), .Y(n55121) );
  A2O1A1Ixp33_ASAP7_75t_SL U47895 ( .A1(n55119), .A2(n55121), .B(n53192), .C(
        n53628), .Y(n58281) );
  A2O1A1Ixp33_ASAP7_75t_SL U47896 ( .A1(n76137), .A2(n55117), .B(n53192), .C(
        n53628), .Y(n76127) );
  A2O1A1Ixp33_ASAP7_75t_SL U47897 ( .A1(n65093), .A2(n65092), .B(n53192), .C(
        n53628), .Y(n55115) );
  A2O1A1Ixp33_ASAP7_75t_SL U47898 ( .A1(n65148), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55113) );
  A2O1A1Ixp33_ASAP7_75t_SL U47899 ( .A1(n65174), .A2(n55113), .B(n53192), .C(
        n53628), .Y(n55114) );
  A2O1A1Ixp33_ASAP7_75t_SL U47900 ( .A1(n55112), .A2(n55114), .B(n53192), .C(
        n53628), .Y(n65150) );
  A2O1A1Ixp33_ASAP7_75t_SL U47901 ( .A1(n77431), .A2(n55110), .B(n53192), .C(
        n53628), .Y(n55111) );
  A2O1A1Ixp33_ASAP7_75t_SL U47902 ( .A1(n54917), .A2(n54920), .B(n53192), .C(
        n53628), .Y(n71785) );
  A2O1A1Ixp33_ASAP7_75t_SL U47903 ( .A1(n57216), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_), 
        .B(n53192), .C(n53628), .Y(n54905) );
  A2O1A1Ixp33_ASAP7_75t_SL U47904 ( .A1(n71888), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_17_), 
        .B(n53192), .C(n53628), .Y(n54906) );
  A2O1A1Ixp33_ASAP7_75t_SL U47905 ( .A1(n57207), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_), 
        .B(n53192), .C(n53628), .Y(n54907) );
  A2O1A1Ixp33_ASAP7_75t_SL U47906 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n55097) );
  A2O1A1Ixp33_ASAP7_75t_SL U47907 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_33_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n55098) );
  A2O1A1Ixp33_ASAP7_75t_SL U47908 ( .A1(n55097), .A2(n55098), .B(n53192), .C(
        n53628), .Y(n55099) );
  A2O1A1Ixp33_ASAP7_75t_SL U47909 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n55101) );
  A2O1A1Ixp33_ASAP7_75t_SL U47910 ( .A1(n55100), .A2(n55101), .B(n53192), .C(
        n53628), .Y(n72094) );
  A2O1A1Ixp33_ASAP7_75t_SL U47911 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n72812), .B(n53192), .C(n53628), .Y(n55091) );
  A2O1A1Ixp33_ASAP7_75t_SL U47912 ( .A1(n75219), .A2(n75220), .B(n53192), .C(
        n53628), .Y(n55088) );
  A2O1A1Ixp33_ASAP7_75t_SL U47913 ( .A1(n75037), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55086) );
  A2O1A1Ixp33_ASAP7_75t_SL U47914 ( .A1(n75063), .A2(n55086), .B(n53192), .C(
        n53628), .Y(n55087) );
  A2O1A1Ixp33_ASAP7_75t_SL U47915 ( .A1(n55085), .A2(n55087), .B(n53192), .C(
        n53628), .Y(n75462) );
  A2O1A1Ixp33_ASAP7_75t_SL U47916 ( .A1(n63383), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55083) );
  A2O1A1Ixp33_ASAP7_75t_SL U47917 ( .A1(n63375), .A2(n55083), .B(n53192), .C(
        n53628), .Y(n55084) );
  A2O1A1Ixp33_ASAP7_75t_SL U47918 ( .A1(n63382), .A2(n55084), .B(n53192), .C(
        n53628), .Y(n63342) );
  A2O1A1Ixp33_ASAP7_75t_SL U47919 ( .A1(n65052), .A2(n67901), .B(n53192), .C(
        n53628), .Y(n54880) );
  A2O1A1Ixp33_ASAP7_75t_SL U47920 ( .A1(n66348), .A2(n54718), .B(n53192), .C(
        n53628), .Y(n54719) );
  A2O1A1Ixp33_ASAP7_75t_SL U47921 ( .A1(n64682), .A2(n64683), .B(n53192), .C(
        n53628), .Y(n55080) );
  A2O1A1Ixp33_ASAP7_75t_SL U47922 ( .A1(n67432), .A2(n57180), .B(n53192), .C(
        n53628), .Y(n55077) );
  A2O1A1Ixp33_ASAP7_75t_SL U47923 ( .A1(n72648), .A2(n55072), .B(n53192), .C(
        n53628), .Y(n55073) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47924 ( .A1(n72646), .A2(n55071), .B(n53192), 
        .C(n55073), .D(n55074), .Y(n12855) );
  A2O1A1Ixp33_ASAP7_75t_SL U47925 ( .A1(n55069), .A2(n55070), .B(n53192), .C(
        n53628), .Y(n3286) );
  A2O1A1Ixp33_ASAP7_75t_SL U47926 ( .A1(n69766), .A2(n55063), .B(n53192), .C(
        n53628), .Y(n55064) );
  A2O1A1Ixp33_ASAP7_75t_SL U47927 ( .A1(n69739), .A2(n55064), .B(n53192), .C(
        n53628), .Y(n55065) );
  A2O1A1Ixp33_ASAP7_75t_SL U47928 ( .A1(n69977), .A2(n55065), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[1]) );
  A2O1A1Ixp33_ASAP7_75t_SL U47929 ( .A1(n53628), .A2(n54866), .B(n53192), .C(
        n53628), .Y(n54867) );
  A2O1A1Ixp33_ASAP7_75t_SL U47930 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_), .B(n53192), .C(
        n53628), .Y(n54518) );
  A2O1A1Ixp33_ASAP7_75t_SL U47931 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_), .B(n53192), .C(
        n53628), .Y(n54519) );
  A2O1A1Ixp33_ASAP7_75t_SL U47932 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_30_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_), .B(n53192), .C(
        n53628), .Y(n54521) );
  A2O1A1Ixp33_ASAP7_75t_SL U47933 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .B(n53192), .C(
        n53628), .Y(n54522) );
  A2O1A1Ixp33_ASAP7_75t_SL U47934 ( .A1(n54520), .A2(n54523), .B(n53192), .C(
        n53628), .Y(n3143) );
  A2O1A1Ixp33_ASAP7_75t_SL U47935 ( .A1(n76518), .A2(n63761), .B(n53192), .C(
        n63762), .Y(n55060) );
  A2O1A1Ixp33_ASAP7_75t_SL U47936 ( .A1(n57144), .A2(n63763), .B(n53192), .C(
        n53628), .Y(n55061) );
  A2O1A1Ixp33_ASAP7_75t_SL U47937 ( .A1(n75542), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n55054) );
  A2O1A1Ixp33_ASAP7_75t_SL U47938 ( .A1(n75540), .A2(n55054), .B(n53192), .C(
        n53628), .Y(n55055) );
  A2O1A1Ixp33_ASAP7_75t_SL U47939 ( .A1(n53628), .A2(n55055), .B(n53192), .C(
        n53628), .Y(n55056) );
  A2O1A1Ixp33_ASAP7_75t_SL U47940 ( .A1(n77194), .A2(n77196), .B(n53192), .C(
        n53628), .Y(n55051) );
  A2O1A1Ixp33_ASAP7_75t_SL U47941 ( .A1(n77212), .A2(n77916), .B(n53192), .C(
        n53628), .Y(n55048) );
  A2O1A1Ixp33_ASAP7_75t_SL U47942 ( .A1(n55047), .A2(n55048), .B(n53192), .C(
        n53628), .Y(n55049) );
  A2O1A1Ixp33_ASAP7_75t_SL U47943 ( .A1(n53628), .A2(n55049), .B(n53192), .C(
        n53628), .Y(n55050) );
  A2O1A1Ixp33_ASAP7_75t_SL U47944 ( .A1(n59691), .A2(n54192), .B(n53192), .C(
        n53628), .Y(n54193) );
  A2O1A1Ixp33_ASAP7_75t_SL U47945 ( .A1(n77425), .A2(n77426), .B(n53192), .C(
        n55045), .Y(n55046) );
  A2O1A1Ixp33_ASAP7_75t_SL U47946 ( .A1(n65387), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_8_), .B(n53192), .C(
        n53628), .Y(n55041) );
  A2O1A1Ixp33_ASAP7_75t_SL U47947 ( .A1(n65387), .A2(n65400), .B(n53192), .C(
        n53628), .Y(n55043) );
  A2O1A1Ixp33_ASAP7_75t_SL U47948 ( .A1(n55042), .A2(n55043), .B(n53192), .C(
        n53628), .Y(n55044) );
  A2O1A1Ixp33_ASAP7_75t_SL U47949 ( .A1(n70476), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_12_), .B(
        n53192), .C(n53628), .Y(n55037) );
  A2O1A1Ixp33_ASAP7_75t_SL U47950 ( .A1(n55036), .A2(n55037), .B(n53192), .C(
        n53628), .Y(n55038) );
  A2O1A1Ixp33_ASAP7_75t_SL U47951 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[9]), .B(n53192), 
        .C(n53628), .Y(n54843) );
  A2O1A1Ixp33_ASAP7_75t_SL U47952 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[9]), .A2(n54844), 
        .B(n53192), .C(n53628), .Y(n54845) );
  A2O1A1Ixp33_ASAP7_75t_SL U47953 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[9]), .B(
        n53192), .C(n53628), .Y(n54846) );
  A2O1A1Ixp33_ASAP7_75t_SL U47954 ( .A1(n54843), .A2(n54845), .B(n53192), .C(
        n54846), .Y(or1200_cpu_or1200_fpu_fpu_arith_N92) );
  A2O1A1Ixp33_ASAP7_75t_SL U47955 ( .A1(n59629), .A2(n78338), .B(n53192), .C(
        n53628), .Y(n55031) );
  A2O1A1Ixp33_ASAP7_75t_SL U47956 ( .A1(n59688), .A2(n54669), .B(n53192), .C(
        n53628), .Y(n54670) );
  A2O1A1Ixp33_ASAP7_75t_SL U47957 ( .A1(n76539), .A2(n77201), .B(n53192), .C(
        n53628), .Y(n55028) );
  A2O1A1Ixp33_ASAP7_75t_SL U47958 ( .A1(n77246), .A2(n77922), .B(n53192), .C(
        n53628), .Y(n55024) );
  A2O1A1Ixp33_ASAP7_75t_SL U47959 ( .A1(n57114), .A2(n77974), .B(n53192), .C(
        n53628), .Y(n55019) );
  A2O1A1Ixp33_ASAP7_75t_SL U47960 ( .A1(n1380), .A2(n55013), .B(n53192), .C(
        n53628), .Y(n55014) );
  A2O1A1Ixp33_ASAP7_75t_SL U47961 ( .A1(n77287), .A2(n77295), .B(n53192), .C(
        n53628), .Y(n55015) );
  A2O1A1Ixp33_ASAP7_75t_SL U47962 ( .A1(n55014), .A2(n55015), .B(n53192), .C(
        n53628), .Y(n55016) );
  A2O1A1Ixp33_ASAP7_75t_SL U47963 ( .A1(n55016), .A2(n55017), .B(n53192), .C(
        n53628), .Y(or1200_pic_N59) );
  A2O1A1Ixp33_ASAP7_75t_SL U47964 ( .A1(n76892), .A2(n54812), .B(n53192), .C(
        n53628), .Y(n54813) );
  A2O1A1Ixp33_ASAP7_75t_SL U47965 ( .A1(n76631), .A2(n54805), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1103) );
  A2O1A1Ixp33_ASAP7_75t_SL U47966 ( .A1(n69016), .A2(n69059), .B(n53192), .C(
        n53628), .Y(n54996) );
  A2O1A1Ixp33_ASAP7_75t_SL U47967 ( .A1(n76903), .A2(n77986), .B(n53192), .C(
        n53628), .Y(n55002) );
  A2O1A1Ixp33_ASAP7_75t_SL U47968 ( .A1(n57072), .A2(n76553), .B(n53192), .C(
        n53628), .Y(n54993) );
  A2O1A1Ixp33_ASAP7_75t_SL U47969 ( .A1(n77153), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n54794) );
  A2O1A1Ixp33_ASAP7_75t_SL U47970 ( .A1(n57093), .A2(n74047), .B(n53192), .C(
        n53628), .Y(n54992) );
  A2O1A1Ixp33_ASAP7_75t_SL U47971 ( .A1(n57072), .A2(n77179), .B(n53192), .C(
        n53628), .Y(n54991) );
  A2O1A1Ixp33_ASAP7_75t_SL U47972 ( .A1(n75686), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n54793) );
  A2O1A1Ixp33_ASAP7_75t_SL U47973 ( .A1(n72514), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54976) );
  A2O1A1Ixp33_ASAP7_75t_SL U47974 ( .A1(n58599), .A2(n54976), .B(n53192), .C(
        n53628), .Y(n54977) );
  A2O1A1Ixp33_ASAP7_75t_SL U47975 ( .A1(n54977), .A2(n54986), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n62) );
  A2O1A1Ixp33_ASAP7_75t_SL U47976 ( .A1(n65758), .A2(n65831), .B(n53192), .C(
        n54956), .Y(n54957) );
  A2O1A1Ixp33_ASAP7_75t_SL U47977 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[1]), .A2(n57205), .B(
        n53192), .C(n53628), .Y(n54953) );
  A2O1A1Ixp33_ASAP7_75t_SL U47978 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[2]), .A2(n57217), .B(
        n53192), .C(n53628), .Y(n54954) );
  A2O1A1Ixp33_ASAP7_75t_SL U47979 ( .A1(n74733), .A2(n57204), .B(n53192), .C(
        n53628), .Y(n54955) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U47980 ( .A1(n54953), .A2(n54954), .B(n53192), 
        .C(n54955), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .Y(
        n73830) );
  A2O1A1Ixp33_ASAP7_75t_SL U47981 ( .A1(n73697), .A2(n59632), .B(n53192), .C(
        n53628), .Y(n54948) );
  A2O1A1Ixp33_ASAP7_75t_SL U47982 ( .A1(n73696), .A2(n57204), .B(n53192), .C(
        n53628), .Y(n54949) );
  A2O1A1Ixp33_ASAP7_75t_SL U47983 ( .A1(n54948), .A2(n54949), .B(n53192), .C(
        n53628), .Y(n54950) );
  A2O1A1Ixp33_ASAP7_75t_SL U47984 ( .A1(n3321), .A2(n57205), .B(n53192), .C(
        n53628), .Y(n54952) );
  A2O1A1Ixp33_ASAP7_75t_SL U47985 ( .A1(n54951), .A2(n54952), .B(n53192), .C(
        n53628), .Y(n73778) );
  A2O1A1Ixp33_ASAP7_75t_SL U47986 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[9]), .A2(n59632), .B(
        n53192), .C(n53628), .Y(n54943) );
  A2O1A1Ixp33_ASAP7_75t_SL U47987 ( .A1(n73695), .A2(n57204), .B(n53192), .C(
        n53628), .Y(n54944) );
  A2O1A1Ixp33_ASAP7_75t_SL U47988 ( .A1(n54943), .A2(n54944), .B(n53192), .C(
        n53628), .Y(n54945) );
  A2O1A1Ixp33_ASAP7_75t_SL U47989 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[11]), .A2(n57205), .B(
        n53192), .C(n53628), .Y(n54947) );
  A2O1A1Ixp33_ASAP7_75t_SL U47990 ( .A1(n54946), .A2(n54947), .B(n53192), .C(
        n53628), .Y(n73789) );
  A2O1A1Ixp33_ASAP7_75t_SL U47991 ( .A1(n66181), .A2(n54942), .B(n53192), .C(
        n53628), .Y(n74090) );
  A2O1A1Ixp33_ASAP7_75t_SL U47992 ( .A1(n62477), .A2(dbg_dat_i[27]), .B(n53192), .C(n53628), .Y(n54939) );
  A2O1A1Ixp33_ASAP7_75t_SL U47993 ( .A1(n62477), .A2(dbg_dat_i[26]), .B(n53192), .C(n53628), .Y(n54938) );
  A2O1A1Ixp33_ASAP7_75t_SL U47994 ( .A1(n74125), .A2(n54932), .B(n53192), .C(
        n54933), .Y(n54934) );
  A2O1A1Ixp33_ASAP7_75t_SL U47995 ( .A1(n58850), .A2(n59659), .B(n53192), .C(
        n53628), .Y(n54928) );
  A2O1A1Ixp33_ASAP7_75t_SL U47996 ( .A1(n76133), .A2(n54928), .B(n53192), .C(
        n53628), .Y(n76128) );
  A2O1A1Ixp33_ASAP7_75t_SL U47997 ( .A1(n63520), .A2(n63467), .B(n53192), .C(
        n53628), .Y(n54925) );
  A2O1A1Ixp33_ASAP7_75t_SL U47998 ( .A1(n63506), .A2(n54925), .B(n53192), .C(
        n53628), .Y(n54926) );
  A2O1A1Ixp33_ASAP7_75t_SL U47999 ( .A1(n53628), .A2(n54926), .B(n53192), .C(
        n53628), .Y(n63484) );
  A2O1A1Ixp33_ASAP7_75t_SL U48000 ( .A1(n71677), .A2(n71719), .B(n53192), .C(
        n53628), .Y(n54917) );
  A2O1A1Ixp33_ASAP7_75t_SL U48001 ( .A1(n57194), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]), .B(n53192), 
        .C(n53628), .Y(n54898) );
  A2O1A1Ixp33_ASAP7_75t_SL U48002 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .A2(n57193), 
        .B(n53192), .C(n53628), .Y(n54899) );
  A2O1A1Ixp33_ASAP7_75t_SL U48003 ( .A1(n54898), .A2(n54899), .B(n53192), .C(
        n53628), .Y(n54900) );
  A2O1A1Ixp33_ASAP7_75t_SL U48004 ( .A1(n57188), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[18]), .B(n53192), 
        .C(n53628), .Y(n54902) );
  A2O1A1Ixp33_ASAP7_75t_SL U48005 ( .A1(n54901), .A2(n54902), .B(n53192), .C(
        n53628), .Y(n65995) );
  A2O1A1Ixp33_ASAP7_75t_SL U48006 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n72723), .B(n53192), .C(n53628), .Y(n54894) );
  A2O1A1Ixp33_ASAP7_75t_SL U48007 ( .A1(n72758), .A2(n72990), .B(n53192), .C(
        n53628), .Y(n54895) );
  A2O1A1Ixp33_ASAP7_75t_SL U48008 ( .A1(n54894), .A2(n54895), .B(n53192), .C(
        n53628), .Y(n54896) );
  A2O1A1Ixp33_ASAP7_75t_SL U48009 ( .A1(n54893), .A2(n54896), .B(n53192), .C(
        n53628), .Y(n54897) );
  A2O1A1Ixp33_ASAP7_75t_SL U48010 ( .A1(n62497), .A2(n54884), .B(n53192), .C(
        n53628), .Y(n54885) );
  A2O1A1Ixp33_ASAP7_75t_SL U48011 ( .A1(n53456), .A2(n54886), .B(n53192), .C(
        n53628), .Y(n76264) );
  A2O1A1Ixp33_ASAP7_75t_SL U48012 ( .A1(n72946), .A2(n53855), .B(n53192), .C(
        n53628), .Y(n72953) );
  A2O1A1Ixp33_ASAP7_75t_SL U48013 ( .A1(n69088), .A2(n69108), .B(n53192), .C(
        n53628), .Y(n54882) );
  A2O1A1Ixp33_ASAP7_75t_SL U48014 ( .A1(n59564), .A2(n60978), .B(n53192), .C(
        n53628), .Y(n54216) );
  A2O1A1Ixp33_ASAP7_75t_SL U48015 ( .A1(n53192), .A2(n53628), .B(n54217), .C(
        n53628), .Y(n54218) );
  A2O1A1Ixp33_ASAP7_75t_SL U48016 ( .A1(n57436), .A2(n59668), .B(n53192), .C(
        n53628), .Y(n54544) );
  A2O1A1Ixp33_ASAP7_75t_SL U48017 ( .A1(n68086), .A2(n63113), .B(n53192), .C(
        n53628), .Y(n54714) );
  A2O1A1Ixp33_ASAP7_75t_SL U48018 ( .A1(n57144), .A2(n75418), .B(n53192), .C(
        n53628), .Y(n54863) );
  A2O1A1Ixp33_ASAP7_75t_SL U48019 ( .A1(n78367), .A2(n73047), .B(n53192), .C(
        n53628), .Y(n54517) );
  A2O1A1Ixp33_ASAP7_75t_SL U48020 ( .A1(n57198), .A2(n76708), .B(n53192), .C(
        n53628), .Y(n54694) );
  A2O1A1Ixp33_ASAP7_75t_SL U48021 ( .A1(n59691), .A2(n54692), .B(n53192), .C(
        n53628), .Y(n54693) );
  A2O1A1Ixp33_ASAP7_75t_SL U48022 ( .A1(n62072), .A2(n54854), .B(n53192), .C(
        n53628), .Y(n54855) );
  A2O1A1Ixp33_ASAP7_75t_SL U48023 ( .A1(n70476), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .B(
        n53192), .C(n53628), .Y(n54840) );
  A2O1A1Ixp33_ASAP7_75t_SL U48024 ( .A1(n70485), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_19_), .B(
        n53192), .C(n53628), .Y(n54841) );
  A2O1A1Ixp33_ASAP7_75t_SL U48025 ( .A1(n54840), .A2(n54841), .B(n53192), .C(
        n53628), .Y(n54842) );
  A2O1A1Ixp33_ASAP7_75t_SL U48026 ( .A1(n70502), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[4]), .B(n53192), .C(
        n53628), .Y(n54837) );
  A2O1A1Ixp33_ASAP7_75t_SL U48027 ( .A1(n70508), .A2(n70372), .B(n53192), .C(
        n53628), .Y(n54838) );
  A2O1A1Ixp33_ASAP7_75t_SL U48028 ( .A1(n57144), .A2(n76652), .B(n53192), .C(
        n53628), .Y(n54834) );
  A2O1A1Ixp33_ASAP7_75t_SL U48029 ( .A1(n3903), .A2(n54831), .B(n53192), .C(
        n53628), .Y(n54832) );
  A2O1A1Ixp33_ASAP7_75t_SL U48030 ( .A1(n59628), .A2(n72713), .B(n53192), .C(
        n53628), .Y(n54465) );
  A2O1A1Ixp33_ASAP7_75t_SL U48031 ( .A1(n57114), .A2(n77992), .B(n53192), .C(
        n53628), .Y(n54827) );
  A2O1A1Ixp33_ASAP7_75t_SL U48032 ( .A1(n1424), .A2(n54822), .B(n53192), .C(
        n53628), .Y(n54823) );
  A2O1A1Ixp33_ASAP7_75t_SL U48033 ( .A1(n77287), .A2(n77583), .B(n53192), .C(
        n53628), .Y(n54824) );
  A2O1A1Ixp33_ASAP7_75t_SL U48034 ( .A1(n54823), .A2(n54824), .B(n53192), .C(
        n53628), .Y(n54825) );
  A2O1A1Ixp33_ASAP7_75t_SL U48035 ( .A1(n54825), .A2(n54826), .B(n53192), .C(
        n53628), .Y(or1200_pic_N47) );
  A2O1A1Ixp33_ASAP7_75t_SL U48036 ( .A1(n1402), .A2(n54817), .B(n53192), .C(
        n53628), .Y(n54818) );
  A2O1A1Ixp33_ASAP7_75t_SL U48037 ( .A1(n77287), .A2(n77600), .B(n53192), .C(
        n53628), .Y(n54819) );
  A2O1A1Ixp33_ASAP7_75t_SL U48038 ( .A1(n54818), .A2(n54819), .B(n53192), .C(
        n53628), .Y(n54820) );
  A2O1A1Ixp33_ASAP7_75t_SL U48039 ( .A1(n54820), .A2(n54821), .B(n53192), .C(
        n53628), .Y(or1200_pic_N53) );
  A2O1A1Ixp33_ASAP7_75t_SL U48040 ( .A1(n77490), .A2(n77495), .B(n53192), .C(
        n53628), .Y(n54815) );
  A2O1A1Ixp33_ASAP7_75t_SL U48041 ( .A1(n53628), .A2(
        or1200_cpu_or1200_mult_mac_div_cntr_2_), .B(n53192), .C(n53628), .Y(
        n54802) );
  A2O1A1Ixp33_ASAP7_75t_SL U48042 ( .A1(n61811), .A2(n54802), .B(n53192), .C(
        n53628), .Y(n54803) );
  A2O1A1Ixp33_ASAP7_75t_SL U48043 ( .A1(or1200_cpu_or1200_mult_mac_div_cntr_3_), .A2(n54803), .B(n53192), .C(n53628), .Y(n54804) );
  A2O1A1Ixp33_ASAP7_75t_SL U48044 ( .A1(n61812), .A2(n54804), .B(n53192), .C(
        n53628), .Y(n54805) );
  A2O1A1Ixp33_ASAP7_75t_SL U48045 ( .A1(n77968), .A2(n76888), .B(n53192), .C(
        n53628), .Y(n54448) );
  A2O1A1Ixp33_ASAP7_75t_SL U48046 ( .A1(n76681), .A2(n59688), .B(n53192), .C(
        n53628), .Y(n54427) );
  A2O1A1Ixp33_ASAP7_75t_SL U48047 ( .A1(n57093), .A2(n76857), .B(n53192), .C(
        n53628), .Y(n54795) );
  A2O1A1Ixp33_ASAP7_75t_SL U48048 ( .A1(n72490), .A2(n72489), .B(n53192), .C(
        n53628), .Y(n54614) );
  A2O1A1Ixp33_ASAP7_75t_SL U48049 ( .A1(n72492), .A2(n72491), .B(n53192), .C(
        n53628), .Y(n54617) );
  A2O1A1Ixp33_ASAP7_75t_SL U48050 ( .A1(n72500), .A2(n54616), .B(n53192), .C(
        n54617), .Y(n54618) );
  A2O1A1Ixp33_ASAP7_75t_SL U48051 ( .A1(n71794), .A2(n54789), .B(n53192), .C(
        n53628), .Y(n54790) );
  A2O1A1Ixp33_ASAP7_75t_SL U48052 ( .A1(n71796), .A2(n54790), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n108) );
  A2O1A1Ixp33_ASAP7_75t_SL U48053 ( .A1(n54607), .A2(n54608), .B(n53192), .C(
        n53628), .Y(n54609) );
  A2O1A1Ixp33_ASAP7_75t_SL U48054 ( .A1(n66162), .A2(n66101), .B(n53192), .C(
        n53628), .Y(n54781) );
  A2O1A1Ixp33_ASAP7_75t_SL U48055 ( .A1(n54780), .A2(n54781), .B(n53192), .C(
        n53628), .Y(n54782) );
  A2O1A1Ixp33_ASAP7_75t_SL U48056 ( .A1(n73376), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54772) );
  A2O1A1Ixp33_ASAP7_75t_SL U48057 ( .A1(n73377), .A2(n54772), .B(n53192), .C(
        n53628), .Y(n54773) );
  A2O1A1Ixp33_ASAP7_75t_SL U48058 ( .A1(n73378), .A2(n54773), .B(n53192), .C(
        n53628), .Y(n73402) );
  A2O1A1Ixp33_ASAP7_75t_SL U48059 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]), .A2(n53628), .B(
        n53192), .C(n53628), .Y(n54766) );
  A2O1A1Ixp33_ASAP7_75t_SL U48060 ( .A1(n59632), .A2(n54766), .B(n53192), .C(
        n53628), .Y(n54767) );
  A2O1A1Ixp33_ASAP7_75t_SL U48061 ( .A1(n54767), .A2(n54768), .B(n53192), .C(
        n53628), .Y(n54769) );
  A2O1A1Ixp33_ASAP7_75t_SL U48062 ( .A1(n73696), .A2(n57205), .B(n53192), .C(
        n53628), .Y(n54771) );
  A2O1A1Ixp33_ASAP7_75t_SL U48063 ( .A1(n2345), .A2(n74686), .B(n53192), .C(
        n53628), .Y(n54758) );
  A2O1A1Ixp33_ASAP7_75t_SL U48064 ( .A1(n62477), .A2(dbg_dat_i[17]), .B(n53192), .C(n53628), .Y(n54757) );
  A2O1A1Ixp33_ASAP7_75t_SL U48065 ( .A1(n54752), .A2(n54755), .B(n53192), .C(
        n53628), .Y(n77979) );
  A2O1A1Ixp33_ASAP7_75t_SL U48066 ( .A1(n76616), .A2(n54754), .B(n53192), .C(
        n53628), .Y(n54755) );
  A2O1A1Ixp33_ASAP7_75t_SL U48067 ( .A1(n69000), .A2(n68994), .B(n53192), .C(
        n53628), .Y(n54076) );
  A2O1A1Ixp33_ASAP7_75t_SL U48068 ( .A1(n62011), .A2(n54745), .B(n53192), .C(
        n53628), .Y(n62006) );
  A2O1A1Ixp33_ASAP7_75t_SL U48069 ( .A1(n57207), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_0_), 
        .B(n53192), .C(n53628), .Y(n54741) );
  A2O1A1Ixp33_ASAP7_75t_SL U48070 ( .A1(n54740), .A2(n54741), .B(n53192), .C(
        n53628), .Y(n54742) );
  A2O1A1Ixp33_ASAP7_75t_SL U48071 ( .A1(n53628), .A2(n54742), .B(n53192), .C(
        n53628), .Y(n54743) );
  A2O1A1Ixp33_ASAP7_75t_SL U48072 ( .A1(n57216), .A2(n72253), .B(n53192), .C(
        n53628), .Y(n54579) );
  A2O1A1Ixp33_ASAP7_75t_SL U48073 ( .A1(n54581), .A2(n54582), .B(n53192), .C(
        n53628), .Y(n72118) );
  A2O1A1Ixp33_ASAP7_75t_SL U48074 ( .A1(n54376), .A2(n54377), .B(n53192), .C(
        n53628), .Y(n66072) );
  A2O1A1Ixp33_ASAP7_75t_SL U48075 ( .A1(n72803), .A2(n72804), .B(n53192), .C(
        n72990), .Y(n53871) );
  A2O1A1Ixp33_ASAP7_75t_SL U48076 ( .A1(n53871), .A2(n53878), .B(n53192), .C(
        n53628), .Y(n73005) );
  A2O1A1Ixp33_ASAP7_75t_SL U48077 ( .A1(or1200_cpu_or1200_fpu_result_conv[11]), 
        .A2(n77090), .B(n53192), .C(n53628), .Y(n54733) );
  A2O1A1Ixp33_ASAP7_75t_SL U48078 ( .A1(n77091), .A2(
        or1200_cpu_or1200_fpu_result_arith[11]), .B(n53192), .C(n53628), .Y(
        n54734) );
  A2O1A1Ixp33_ASAP7_75t_SL U48079 ( .A1(n54733), .A2(n54734), .B(n53192), .C(
        n53628), .Y(n54735) );
  A2O1A1Ixp33_ASAP7_75t_SL U48080 ( .A1(or1200_cpu_or1200_fpu_result_arith[14]), .A2(n77091), .B(n53192), .C(n53628), .Y(n54552) );
  A2O1A1Ixp33_ASAP7_75t_SL U48081 ( .A1(n57121), .A2(n63891), .B(n53192), .C(
        n53628), .Y(n54731) );
  A2O1A1Ixp33_ASAP7_75t_SL U48082 ( .A1(n71314), .A2(n71329), .B(n53192), .C(
        n53628), .Y(n54729) );
  A2O1A1Ixp33_ASAP7_75t_SL U48083 ( .A1(n59562), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[34]), .B(n53192), 
        .C(n53628), .Y(n54728) );
  A2O1A1Ixp33_ASAP7_75t_SL U48084 ( .A1(n57107), .A2(n67899), .B(n53192), .C(
        n53628), .Y(n54724) );
  A2O1A1Ixp33_ASAP7_75t_SL U48085 ( .A1(n73813), .A2(n73811), .B(n53192), .C(
        n53628), .Y(n54533) );
  A2O1A1Ixp33_ASAP7_75t_SL U48086 ( .A1(n73817), .A2(n54532), .B(n53192), .C(
        n54533), .Y(n3292) );
  A2O1A1Ixp33_ASAP7_75t_SL U48087 ( .A1(n69983), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54529) );
  A2O1A1Ixp33_ASAP7_75t_SL U48088 ( .A1(n54528), .A2(n54530), .B(n53192), .C(
        n53628), .Y(n3214) );
  A2O1A1Ixp33_ASAP7_75t_SL U48089 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[5]), .A2(
        n70589), .B(n53192), .C(n53628), .Y(n54524) );
  A2O1A1Ixp33_ASAP7_75t_SL U48090 ( .A1(n76528), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54708) );
  A2O1A1Ixp33_ASAP7_75t_SL U48091 ( .A1(n59689), .A2(n54708), .B(n53192), .C(
        n53628), .Y(n54709) );
  A2O1A1Ixp33_ASAP7_75t_SL U48092 ( .A1(n76529), .A2(n54709), .B(n53192), .C(
        n53628), .Y(n54710) );
  A2O1A1Ixp33_ASAP7_75t_SL U48093 ( .A1(n57144), .A2(n65220), .B(n53192), .C(
        n53628), .Y(n54707) );
  A2O1A1Ixp33_ASAP7_75t_SL U48094 ( .A1(n72693), .A2(n59628), .B(n53192), .C(
        n53628), .Y(n54702) );
  A2O1A1Ixp33_ASAP7_75t_SL U48095 ( .A1(n59629), .A2(n72719), .B(n53192), .C(
        n54698), .Y(n54699) );
  A2O1A1Ixp33_ASAP7_75t_SL U48096 ( .A1(n77212), .A2(n77983), .B(n53192), .C(
        n53628), .Y(n54695) );
  A2O1A1Ixp33_ASAP7_75t_SL U48097 ( .A1(n54694), .A2(n54695), .B(n53192), .C(
        n53628), .Y(n54696) );
  A2O1A1Ixp33_ASAP7_75t_SL U48098 ( .A1(n53628), .A2(n54696), .B(n53192), .C(
        n53628), .Y(n54697) );
  A2O1A1Ixp33_ASAP7_75t_SL U48099 ( .A1(n59691), .A2(n77921), .B(n53192), .C(
        n53628), .Y(n54691) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U48100 ( .A1(n60491), .A2(n69343), .B(n53192), 
        .C(n61136), .D(n54684), .Y(n54685) );
  A2O1A1Ixp33_ASAP7_75t_SL U48101 ( .A1(n54685), .A2(n54686), .B(n53192), .C(
        n53628), .Y(n54687) );
  A2O1A1Ixp33_ASAP7_75t_SL U48102 ( .A1(n70384), .A2(n70371), .B(n53192), .C(
        n53628), .Y(n54676) );
  A2O1A1Ixp33_ASAP7_75t_SL U48103 ( .A1(n74644), .A2(n70476), .B(n53192), .C(
        n53628), .Y(n54673) );
  A2O1A1Ixp33_ASAP7_75t_SL U48104 ( .A1(n70485), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_), .B(
        n53192), .C(n53628), .Y(n54674) );
  A2O1A1Ixp33_ASAP7_75t_SL U48105 ( .A1(n54673), .A2(n54674), .B(n53192), .C(
        n53628), .Y(n54675) );
  A2O1A1Ixp33_ASAP7_75t_SL U48106 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[1]), .B(n53192), 
        .C(n53628), .Y(n54489) );
  A2O1A1Ixp33_ASAP7_75t_SL U48107 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[1]), .A2(n54490), 
        .B(n53192), .C(n53628), .Y(n54491) );
  A2O1A1Ixp33_ASAP7_75t_SL U48108 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[1]), .B(
        n53192), .C(n53628), .Y(n54492) );
  A2O1A1Ixp33_ASAP7_75t_SL U48109 ( .A1(n54489), .A2(n54491), .B(n53192), .C(
        n54492), .Y(or1200_cpu_or1200_fpu_fpu_arith_N84) );
  A2O1A1Ixp33_ASAP7_75t_SL U48110 ( .A1(n77683), .A2(n77284), .B(n53192), .C(
        n77679), .Y(n54667) );
  A2O1A1Ixp33_ASAP7_75t_SL U48111 ( .A1(n59680), .A2(n77971), .B(n53192), .C(
        n53628), .Y(n54668) );
  A2O1A1Ixp33_ASAP7_75t_SL U48112 ( .A1(n57114), .A2(n77968), .B(n53192), .C(
        n53628), .Y(n54664) );
  A2O1A1Ixp33_ASAP7_75t_SL U48113 ( .A1(n77992), .A2(n74641), .B(n53192), .C(
        n53628), .Y(n54459) );
  A2O1A1Ixp33_ASAP7_75t_SL U48114 ( .A1(n77494), .A2(n77490), .B(n53192), .C(
        n53628), .Y(n54662) );
  A2O1A1Ixp33_ASAP7_75t_SL U48115 ( .A1(n54652), .A2(n54653), .B(n53192), .C(
        n53628), .Y(n54654) );
  A2O1A1Ixp33_ASAP7_75t_SL U48116 ( .A1(n76633), .A2(n54654), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n136) );
  A2O1A1Ixp33_ASAP7_75t_SL U48117 ( .A1(n68885), .A2(n54636), .B(n53192), .C(
        n53628), .Y(n54637) );
  A2O1A1Ixp33_ASAP7_75t_SL U48118 ( .A1(n57080), .A2(n68831), .B(n53192), .C(
        n53628), .Y(n54639) );
  A2O1A1Ixp33_ASAP7_75t_SL U48119 ( .A1(n69130), .A2(n57080), .B(n53192), .C(
        n53628), .Y(n54632) );
  A2O1A1Ixp33_ASAP7_75t_SL U48120 ( .A1(n57072), .A2(n76619), .B(n53192), .C(
        n53628), .Y(n54624) );
  A2O1A1Ixp33_ASAP7_75t_SL U48121 ( .A1(n74129), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n54276) );
  A2O1A1Ixp33_ASAP7_75t_SL U48122 ( .A1(n57093), .A2(n76928), .B(n53192), .C(
        n53628), .Y(n54623) );
  A2O1A1Ixp33_ASAP7_75t_SL U48123 ( .A1(n53628), .A2(n72488), .B(n53192), .C(
        n53628), .Y(n54612) );
  A2O1A1Ixp33_ASAP7_75t_SL U48124 ( .A1(n72502), .A2(n54612), .B(n53192), .C(
        n53628), .Y(n54613) );
  A2O1A1Ixp33_ASAP7_75t_SL U48125 ( .A1(n54613), .A2(n54614), .B(n53192), .C(
        n53628), .Y(n54615) );
  A2O1A1Ixp33_ASAP7_75t_SL U48126 ( .A1(n71797), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54610) );
  A2O1A1Ixp33_ASAP7_75t_SL U48127 ( .A1(n71795), .A2(n54610), .B(n53192), .C(
        n53628), .Y(n54611) );
  A2O1A1Ixp33_ASAP7_75t_SL U48128 ( .A1(n71796), .A2(n54611), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n111) );
  A2O1A1Ixp33_ASAP7_75t_SL U48129 ( .A1(n59698), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54408) );
  A2O1A1Ixp33_ASAP7_75t_SL U48130 ( .A1(n53628), .A2(n54409), .B(n53192), .C(
        n53628), .Y(n54410) );
  A2O1A1Ixp33_ASAP7_75t_SL U48131 ( .A1(n70938), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54403) );
  A2O1A1Ixp33_ASAP7_75t_SL U48132 ( .A1(n53628), .A2(n54404), .B(n53192), .C(
        n53628), .Y(n54405) );
  A2O1A1Ixp33_ASAP7_75t_SL U48133 ( .A1(n74302), .A2(n74303), .B(n53192), .C(
        n54604), .Y(n54605) );
  A2O1A1Ixp33_ASAP7_75t_SL U48134 ( .A1(n62477), .A2(dbg_dat_i[28]), .B(n53192), .C(n53628), .Y(n54600) );
  A2O1A1Ixp33_ASAP7_75t_SL U48135 ( .A1(n62477), .A2(dbg_dat_i[29]), .B(n53192), .C(n53628), .Y(n54599) );
  A2O1A1Ixp33_ASAP7_75t_SL U48136 ( .A1(n76201), .A2(n76200), .B(n53192), .C(
        n53628), .Y(n54251) );
  A2O1A1Ixp33_ASAP7_75t_SL U48137 ( .A1(n76199), .A2(n76612), .B(n53192), .C(
        n53628), .Y(n54255) );
  A2O1A1Ixp33_ASAP7_75t_SL U48138 ( .A1(n75445), .A2(n54595), .B(n53192), .C(
        n53628), .Y(n54597) );
  A2O1A1Ixp33_ASAP7_75t_SL U48139 ( .A1(n53628), .A2(n54597), .B(n53192), .C(
        n53628), .Y(n54598) );
  A2O1A1Ixp33_ASAP7_75t_SL U48140 ( .A1(n77250), .A2(n54594), .B(n53192), .C(
        n53628), .Y(n77272) );
  A2O1A1Ixp33_ASAP7_75t_SL U48141 ( .A1(n62906), .A2(n62907), .B(n53192), .C(
        n53628), .Y(n54591) );
  A2O1A1Ixp33_ASAP7_75t_SL U48142 ( .A1(n61811), .A2(n54588), .B(n53192), .C(
        n53628), .Y(n61812) );
  A2O1A1Ixp33_ASAP7_75t_SL U48143 ( .A1(n63505), .A2(n63484), .B(n53192), .C(
        n53628), .Y(n54586) );
  A2O1A1Ixp33_ASAP7_75t_SL U48144 ( .A1(n63502), .A2(n54586), .B(n53192), .C(
        n53628), .Y(n54587) );
  A2O1A1Ixp33_ASAP7_75t_SL U48145 ( .A1(n53628), .A2(n54587), .B(n53192), .C(
        n53628), .Y(n63509) );
  A2O1A1Ixp33_ASAP7_75t_SL U48146 ( .A1(or1200_cpu_or1200_mult_mac_n233), .A2(
        n54585), .B(n53192), .C(n53628), .Y(n69166) );
  A2O1A1Ixp33_ASAP7_75t_SL U48147 ( .A1(n77431), .A2(n77447), .B(n53192), .C(
        n53628), .Y(n54583) );
  A2O1A1Ixp33_ASAP7_75t_SL U48148 ( .A1(n71888), .A2(n72307), .B(n53192), .C(
        n53628), .Y(n54582) );
  A2O1A1Ixp33_ASAP7_75t_SL U48149 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_32_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n54574) );
  A2O1A1Ixp33_ASAP7_75t_SL U48150 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n54575) );
  A2O1A1Ixp33_ASAP7_75t_SL U48151 ( .A1(n54574), .A2(n54575), .B(n53192), .C(
        n53628), .Y(n54576) );
  A2O1A1Ixp33_ASAP7_75t_SL U48152 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n54578) );
  A2O1A1Ixp33_ASAP7_75t_SL U48153 ( .A1(n54577), .A2(n54578), .B(n53192), .C(
        n53628), .Y(n72069) );
  A2O1A1Ixp33_ASAP7_75t_SL U48154 ( .A1(n71365), .A2(n71223), .B(n53192), .C(
        n53628), .Y(n54568) );
  A2O1A1Ixp33_ASAP7_75t_SL U48155 ( .A1(n54567), .A2(n54568), .B(n53192), .C(
        n53628), .Y(n71203) );
  A2O1A1Ixp33_ASAP7_75t_SL U48156 ( .A1(n66152), .A2(n54565), .B(n53192), .C(
        n53628), .Y(n66095) );
  A2O1A1Ixp33_ASAP7_75t_SL U48157 ( .A1(n53675), .A2(n53676), .B(n53192), .C(
        n53628), .Y(n53677) );
  A2O1A1Ixp33_ASAP7_75t_SL U48158 ( .A1(n53678), .A2(n53679), .B(n53192), .C(
        n53628), .Y(n66013) );
  A2O1A1Ixp33_ASAP7_75t_SL U48159 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .A2(n57193), 
        .B(n53192), .C(n53628), .Y(n54561) );
  A2O1A1Ixp33_ASAP7_75t_SL U48160 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]), .A2(n57188), 
        .B(n53192), .C(n53628), .Y(n54562) );
  A2O1A1Ixp33_ASAP7_75t_SL U48161 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .A2(n57187), 
        .B(n53192), .C(n53628), .Y(n54563) );
  A2O1A1Ixp33_ASAP7_75t_SL U48162 ( .A1(n54561), .A2(n54562), .B(n53192), .C(
        n54563), .Y(n54564) );
  A2O1A1Ixp33_ASAP7_75t_SL U48163 ( .A1(n73239), .A2(n74502), .B(n53192), .C(
        n53628), .Y(n54559) );
  A2O1A1Ixp33_ASAP7_75t_SL U48164 ( .A1(n59632), .A2(n73823), .B(n53192), .C(
        n53628), .Y(n54556) );
  A2O1A1Ixp33_ASAP7_75t_SL U48165 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[7]), .A2(n57204), .B(
        n53192), .C(n53628), .Y(n54557) );
  A2O1A1Ixp33_ASAP7_75t_SL U48166 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[9]), .A2(n57217), .B(
        n53192), .C(n53628), .Y(n54558) );
  A2O1A1Ixp33_ASAP7_75t_SL U48167 ( .A1(n54556), .A2(n54557), .B(n53192), .C(
        n54558), .Y(n73737) );
  A2O1A1Ixp33_ASAP7_75t_SL U48168 ( .A1(n74680), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_12_), .B(
        n53192), .C(n53628), .Y(n54045) );
  A2O1A1Ixp33_ASAP7_75t_SL U48169 ( .A1(or1200_cpu_or1200_fpu_result_conv[14]), 
        .A2(n77090), .B(n53192), .C(n53628), .Y(n54553) );
  A2O1A1Ixp33_ASAP7_75t_SL U48170 ( .A1(n54552), .A2(n54553), .B(n53192), .C(
        n53628), .Y(n54554) );
  A2O1A1Ixp33_ASAP7_75t_SL U48171 ( .A1(n53628), .A2(n54554), .B(n53192), .C(
        n53628), .Y(n54555) );
  A2O1A1Ixp33_ASAP7_75t_SL U48172 ( .A1(n57121), .A2(n63537), .B(n53192), .C(
        n53628), .Y(n54551) );
  A2O1A1Ixp33_ASAP7_75t_SL U48173 ( .A1(n71599), .A2(n54549), .B(n53192), .C(
        n53628), .Y(n71472) );
  A2O1A1Ixp33_ASAP7_75t_SL U48174 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[4]), .A2(
        n54547), .B(n53192), .C(n53628), .Y(n70168) );
  A2O1A1Ixp33_ASAP7_75t_SL U48175 ( .A1(n62614), .A2(n57120), .B(n53192), .C(
        n54545), .Y(n54546) );
  A2O1A1Ixp33_ASAP7_75t_SL U48176 ( .A1(n61911), .A2(n59256), .B(n53192), .C(
        n53628), .Y(n54543) );
  A2O1A1Ixp33_ASAP7_75t_SL U48177 ( .A1(n59563), .A2(n54542), .B(n53192), .C(
        n53628), .Y(n64189) );
  A2O1A1Ixp33_ASAP7_75t_SL U48178 ( .A1(n59518), .A2(n59659), .B(n53192), .C(
        n57425), .Y(n54537) );
  A2O1A1Ixp33_ASAP7_75t_SL U48179 ( .A1(n70081), .A2(n54529), .B(n53192), .C(
        n53628), .Y(n54530) );
  A2O1A1Ixp33_ASAP7_75t_SL U48180 ( .A1(n70594), .A2(n54524), .B(n53192), .C(
        n54525), .Y(n54526) );
  A2O1A1Ixp33_ASAP7_75t_SL U48181 ( .A1(n77194), .A2(n76945), .B(n53192), .C(
        n53628), .Y(n54514) );
  A2O1A1Ixp33_ASAP7_75t_SL U48182 ( .A1(n62001), .A2(n60497), .B(n53192), .C(
        n53628), .Y(n54513) );
  A2O1A1Ixp33_ASAP7_75t_SL U48183 ( .A1(n54512), .A2(n54513), .B(n53192), .C(
        n53628), .Y(n9465) );
  A2O1A1Ixp33_ASAP7_75t_SL U48184 ( .A1(n59691), .A2(n54343), .B(n53192), .C(
        n53628), .Y(n54344) );
  A2O1A1Ixp33_ASAP7_75t_SL U48185 ( .A1(n70485), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_1_), .B(
        n53192), .C(n53628), .Y(n54494) );
  A2O1A1Ixp33_ASAP7_75t_SL U48186 ( .A1(n70537), .A2(n54494), .B(n53192), .C(
        n53628), .Y(n54495) );
  A2O1A1Ixp33_ASAP7_75t_SL U48187 ( .A1(n70543), .A2(n74677), .B(n53192), .C(
        n53628), .Y(n54498) );
  A2O1A1Ixp33_ASAP7_75t_SL U48188 ( .A1(n70486), .A2(n74686), .B(n53192), .C(
        n53628), .Y(n54499) );
  A2O1A1Ixp33_ASAP7_75t_SL U48189 ( .A1(n54498), .A2(n54499), .B(n53192), .C(
        n53628), .Y(n54500) );
  A2O1A1Ixp33_ASAP7_75t_SL U48190 ( .A1(n70539), .A2(n70489), .B(n53192), .C(
        n53628), .Y(n54502) );
  A2O1A1Ixp33_ASAP7_75t_SL U48191 ( .A1(n70482), .A2(n54505), .B(n53192), .C(
        n53628), .Y(n54506) );
  A2O1A1Ixp33_ASAP7_75t_SL U48192 ( .A1(n70483), .A2(n70484), .B(n53192), .C(
        n53628), .Y(n54507) );
  A2O1A1Ixp33_ASAP7_75t_SL U48193 ( .A1(n54506), .A2(n54507), .B(n53192), .C(
        n53628), .Y(n54508) );
  A2O1A1Ixp33_ASAP7_75t_SL U48194 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .A2(
        n54508), .B(n53192), .C(n53628), .Y(n54509) );
  A2O1A1Ixp33_ASAP7_75t_SL U48195 ( .A1(n54504), .A2(n54509), .B(n53192), .C(
        n53628), .Y(n2432) );
  A2O1A1Ixp33_ASAP7_75t_SL U48196 ( .A1(n69781), .A2(n54480), .B(n53192), .C(
        n53628), .Y(n54481) );
  A2O1A1Ixp33_ASAP7_75t_SL U48197 ( .A1(n54481), .A2(n54482), .B(n53192), .C(
        n53628), .Y(n54483) );
  A2O1A1Ixp33_ASAP7_75t_SL U48198 ( .A1(n69783), .A2(n54484), .B(n53192), .C(
        n53628), .Y(n54485) );
  A2O1A1Ixp33_ASAP7_75t_SL U48199 ( .A1(n54483), .A2(n54485), .B(n53192), .C(
        n53628), .Y(n54486) );
  A2O1A1Ixp33_ASAP7_75t_SL U48200 ( .A1(n54338), .A2(n62062), .B(n53192), .C(
        n53628), .Y(n2205) );
  A2O1A1Ixp33_ASAP7_75t_SL U48201 ( .A1(n77200), .A2(n54473), .B(n53192), .C(
        n53628), .Y(n54474) );
  A2O1A1Ixp33_ASAP7_75t_SL U48202 ( .A1(n54472), .A2(n54475), .B(n53192), .C(
        n53628), .Y(n54476) );
  A2O1A1Ixp33_ASAP7_75t_SL U48203 ( .A1(n59680), .A2(n77920), .B(n53192), .C(
        n53628), .Y(n54477) );
  A2O1A1Ixp33_ASAP7_75t_SL U48204 ( .A1(n54476), .A2(n54477), .B(n53192), .C(
        n53628), .Y(or1200_du_N96) );
  A2O1A1Ixp33_ASAP7_75t_SL U48205 ( .A1(n58296), .A2(n77980), .B(n53192), .C(
        n53628), .Y(n54469) );
  A2O1A1Ixp33_ASAP7_75t_SL U48206 ( .A1(n54468), .A2(n54469), .B(n53192), .C(
        n53628), .Y(n54470) );
  A2O1A1Ixp33_ASAP7_75t_SL U48207 ( .A1(n53628), .A2(n54470), .B(n53192), .C(
        n53628), .Y(n54471) );
  A2O1A1Ixp33_ASAP7_75t_SL U48208 ( .A1(or1200_cpu_or1200_fpu_overflow), .A2(
        n74920), .B(n53192), .C(n53628), .Y(n54464) );
  A2O1A1Ixp33_ASAP7_75t_SL U48209 ( .A1(n54463), .A2(n54464), .B(n53192), .C(
        n53628), .Y(n9490) );
  A2O1A1Ixp33_ASAP7_75t_SL U48210 ( .A1(n57114), .A2(n77971), .B(n53192), .C(
        n53628), .Y(n54460) );
  A2O1A1Ixp33_ASAP7_75t_SL U48211 ( .A1(n58600), .A2(n75935), .B(n53192), .C(
        n53628), .Y(n54454) );
  A2O1A1Ixp33_ASAP7_75t_SL U48212 ( .A1(or1200_cpu_or1200_mult_mac_n307), .A2(
        n54441), .B(n53192), .C(n53628), .Y(n54443) );
  A2O1A1Ixp33_ASAP7_75t_SL U48213 ( .A1(n63435), .A2(n54443), .B(n53192), .C(
        n53628), .Y(n54444) );
  A2O1A1Ixp33_ASAP7_75t_SL U48214 ( .A1(n75650), .A2(n76721), .B(n53192), .C(
        n53628), .Y(n54288) );
  A2O1A1Ixp33_ASAP7_75t_SL U48215 ( .A1(n54300), .A2(n54305), .B(n53192), .C(
        n53628), .Y(n54306) );
  A2O1A1Ixp33_ASAP7_75t_SL U48216 ( .A1(n59673), .A2(n77983), .B(n53192), .C(
        n53628), .Y(n54308) );
  A2O1A1Ixp33_ASAP7_75t_SL U48217 ( .A1(n54288), .A2(n54307), .B(n53192), .C(
        n54308), .Y(or1200_cpu_or1200_mult_mac_n1617) );
  A2O1A1Ixp33_ASAP7_75t_SL U48218 ( .A1(n72502), .A2(n72332), .B(n53192), .C(
        n72333), .Y(n54418) );
  A2O1A1Ixp33_ASAP7_75t_SL U48219 ( .A1(n72490), .A2(n72463), .B(n53192), .C(
        n53628), .Y(n54421) );
  A2O1A1Ixp33_ASAP7_75t_SL U48220 ( .A1(n72500), .A2(n54420), .B(n53192), .C(
        n54421), .Y(n54422) );
  A2O1A1Ixp33_ASAP7_75t_SL U48221 ( .A1(n72486), .A2(n54424), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n64) );
  A2O1A1Ixp33_ASAP7_75t_SL U48222 ( .A1(n71785), .A2(n54413), .B(n53192), .C(
        n53628), .Y(n54414) );
  A2O1A1Ixp33_ASAP7_75t_SL U48223 ( .A1(n71796), .A2(n54414), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n109) );
  A2O1A1Ixp33_ASAP7_75t_SL U48224 ( .A1(n70729), .A2(n54408), .B(n53192), .C(
        n53628), .Y(n54409) );
  A2O1A1Ixp33_ASAP7_75t_SL U48225 ( .A1(n53628), .A2(n59699), .B(n53192), .C(
        n53628), .Y(n54400) );
  A2O1A1Ixp33_ASAP7_75t_SL U48226 ( .A1(n70941), .A2(n54400), .B(n53192), .C(
        n53628), .Y(n54401) );
  A2O1A1Ixp33_ASAP7_75t_SL U48227 ( .A1(n53628), .A2(n54401), .B(n53192), .C(
        n53628), .Y(n54402) );
  A2O1A1Ixp33_ASAP7_75t_SL U48228 ( .A1(n70922), .A2(n54403), .B(n53192), .C(
        n53628), .Y(n54404) );
  A2O1A1Ixp33_ASAP7_75t_SL U48229 ( .A1(n73555), .A2(n73556), .B(n53192), .C(
        n53628), .Y(n54399) );
  A2O1A1Ixp33_ASAP7_75t_SL U48230 ( .A1(n76517), .A2(n54398), .B(n53192), .C(
        n53628), .Y(n76518) );
  A2O1A1Ixp33_ASAP7_75t_SL U48231 ( .A1(n62477), .A2(dbg_dat_i[0]), .B(n53192), 
        .C(n53628), .Y(n54397) );
  A2O1A1Ixp33_ASAP7_75t_SL U48232 ( .A1(n74203), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54395) );
  A2O1A1Ixp33_ASAP7_75t_SL U48233 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_sign), .A2(n54395), .B(n53192), 
        .C(n53628), .Y(n54396) );
  A2O1A1Ixp33_ASAP7_75t_SL U48234 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]), .A2(n54396), .B(
        n53192), .C(n53628), .Y(n74212) );
  A2O1A1Ixp33_ASAP7_75t_SL U48235 ( .A1(n54255), .A2(n54254), .B(n53192), .C(
        n53628), .Y(n54256) );
  A2O1A1Ixp33_ASAP7_75t_SL U48236 ( .A1(n77723), .A2(n59578), .B(n53192), .C(
        n53628), .Y(n54389) );
  A2O1A1Ixp33_ASAP7_75t_SL U48237 ( .A1(n57207), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_), 
        .B(n53192), .C(n53628), .Y(n54243) );
  A2O1A1Ixp33_ASAP7_75t_SL U48238 ( .A1(n53628), .A2(n54245), .B(n53192), .C(
        n53628), .Y(n54246) );
  A2O1A1Ixp33_ASAP7_75t_SL U48239 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_24_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n54384) );
  A2O1A1Ixp33_ASAP7_75t_SL U48240 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n54385) );
  A2O1A1Ixp33_ASAP7_75t_SL U48241 ( .A1(n54384), .A2(n54385), .B(n53192), .C(
        n53628), .Y(n54386) );
  A2O1A1Ixp33_ASAP7_75t_SL U48242 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n54388) );
  A2O1A1Ixp33_ASAP7_75t_SL U48243 ( .A1(n54387), .A2(n54388), .B(n53192), .C(
        n53628), .Y(n72065) );
  A2O1A1Ixp33_ASAP7_75t_SL U48244 ( .A1(n57194), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[35]), .B(n53192), 
        .C(n53628), .Y(n54378) );
  A2O1A1Ixp33_ASAP7_75t_SL U48245 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[36]), .A2(n57193), 
        .B(n53192), .C(n53628), .Y(n54379) );
  A2O1A1Ixp33_ASAP7_75t_SL U48246 ( .A1(n54378), .A2(n54379), .B(n53192), .C(
        n53628), .Y(n54380) );
  A2O1A1Ixp33_ASAP7_75t_SL U48247 ( .A1(n57188), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[33]), .B(n53192), 
        .C(n53628), .Y(n54382) );
  A2O1A1Ixp33_ASAP7_75t_SL U48248 ( .A1(n54381), .A2(n54382), .B(n53192), .C(
        n53628), .Y(n65934) );
  A2O1A1Ixp33_ASAP7_75t_SL U48249 ( .A1(n65978), .A2(n66079), .B(n53192), .C(
        n53628), .Y(n54376) );
  A2O1A1Ixp33_ASAP7_75t_SL U48250 ( .A1(n66023), .A2(n66051), .B(n53192), .C(
        n53628), .Y(n54377) );
  A2O1A1Ixp33_ASAP7_75t_SL U48251 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), 
        .A2(n53875), .B(n53192), .C(n53628), .Y(n53876) );
  A2O1A1Ixp33_ASAP7_75t_SL U48252 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n53877), .B(n53192), .C(n53628), .Y(n53878) );
  A2O1A1Ixp33_ASAP7_75t_SL U48253 ( .A1(n78139), .A2(n54375), .B(n53192), .C(
        n53628), .Y(n75297) );
  A2O1A1Ixp33_ASAP7_75t_SL U48254 ( .A1(n65141), .A2(n65143), .B(n53192), .C(
        n53628), .Y(n54220) );
  A2O1A1Ixp33_ASAP7_75t_SL U48255 ( .A1(n59562), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .B(n53192), 
        .C(n53628), .Y(n54369) );
  A2O1A1Ixp33_ASAP7_75t_SL U48256 ( .A1(n57190), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[9]), .B(n53192), 
        .C(n53628), .Y(n54368) );
  A2O1A1Ixp33_ASAP7_75t_SL U48257 ( .A1(n75048), .A2(n75040), .B(n53192), .C(
        n53628), .Y(n54367) );
  A2O1A1Ixp33_ASAP7_75t_SL U48258 ( .A1(n67610), .A2(n58402), .B(n53192), .C(
        n53628), .Y(n54365) );
  A2O1A1Ixp33_ASAP7_75t_SL U48259 ( .A1(n66424), .A2(n59596), .B(n53192), .C(
        n53628), .Y(n54361) );
  A2O1A1Ixp33_ASAP7_75t_SL U48260 ( .A1(n66422), .A2(n54361), .B(n53192), .C(
        n53628), .Y(n54362) );
  A2O1A1Ixp33_ASAP7_75t_SL U48261 ( .A1(n66423), .A2(n54362), .B(n53192), .C(
        n53628), .Y(n66425) );
  A2O1A1Ixp33_ASAP7_75t_SL U48262 ( .A1(n69873), .A2(n70059), .B(n53192), .C(
        n53628), .Y(n54199) );
  A2O1A1Ixp33_ASAP7_75t_SL U48263 ( .A1(n59629), .A2(n72761), .B(n53192), .C(
        n54345), .Y(n54346) );
  A2O1A1Ixp33_ASAP7_75t_SL U48264 ( .A1(n62001), .A2(n62052), .B(n53192), .C(
        n62003), .Y(n54342) );
  A2O1A1Ixp33_ASAP7_75t_SL U48265 ( .A1(n54341), .A2(n54342), .B(n53192), .C(
        n53628), .Y(n9568) );
  A2O1A1Ixp33_ASAP7_75t_SL U48266 ( .A1(n54186), .A2(n54188), .B(n53192), .C(
        n53628), .Y(n54189) );
  A2O1A1Ixp33_ASAP7_75t_SL U48267 ( .A1(n53628), .A2(n54189), .B(n53192), .C(
        n53628), .Y(n2441) );
  A2O1A1Ixp33_ASAP7_75t_SL U48268 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[2]), .B(n53192), 
        .C(n53628), .Y(n54173) );
  A2O1A1Ixp33_ASAP7_75t_SL U48269 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[2]), .A2(n54174), 
        .B(n53192), .C(n53628), .Y(n54175) );
  A2O1A1Ixp33_ASAP7_75t_SL U48270 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[2]), .B(
        n53192), .C(n53628), .Y(n54176) );
  A2O1A1Ixp33_ASAP7_75t_SL U48271 ( .A1(n54173), .A2(n54175), .B(n53192), .C(
        n54176), .Y(or1200_cpu_or1200_fpu_fpu_arith_N85) );
  A2O1A1Ixp33_ASAP7_75t_SL U48272 ( .A1(n70502), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[9]), .B(n53192), .C(
        n53628), .Y(n54171) );
  A2O1A1Ixp33_ASAP7_75t_SL U48273 ( .A1(n72693), .A2(n59629), .B(n53192), .C(
        n53628), .Y(n54012) );
  A2O1A1Ixp33_ASAP7_75t_SL U48274 ( .A1(n59690), .A2(n77917), .B(n53192), .C(
        n53628), .Y(n54336) );
  A2O1A1Ixp33_ASAP7_75t_SL U48275 ( .A1(n76649), .A2(n57198), .B(n53192), .C(
        n53628), .Y(n54333) );
  A2O1A1Ixp33_ASAP7_75t_SL U48276 ( .A1(n53192), .A2(n53628), .B(n53787), .C(
        n53628), .Y(n53788) );
  A2O1A1Ixp33_ASAP7_75t_SL U48277 ( .A1(n57114), .A2(n77901), .B(n53192), .C(
        n53628), .Y(n54320) );
  A2O1A1Ixp33_ASAP7_75t_SL U48278 ( .A1(n1410), .A2(n54315), .B(n53192), .C(
        n53628), .Y(n54316) );
  A2O1A1Ixp33_ASAP7_75t_SL U48279 ( .A1(n77287), .A2(n77594), .B(n53192), .C(
        n53628), .Y(n54317) );
  A2O1A1Ixp33_ASAP7_75t_SL U48280 ( .A1(n54316), .A2(n54317), .B(n53192), .C(
        n53628), .Y(n54318) );
  A2O1A1Ixp33_ASAP7_75t_SL U48281 ( .A1(n54318), .A2(n54319), .B(n53192), .C(
        n53628), .Y(or1200_pic_N51) );
  A2O1A1Ixp33_ASAP7_75t_SL U48282 ( .A1(n75990), .A2(n76195), .B(n53192), .C(
        n53628), .Y(n53990) );
  A2O1A1Ixp33_ASAP7_75t_SL U48283 ( .A1(n75991), .A2(n58600), .B(n53192), .C(
        n53628), .Y(n53994) );
  A2O1A1Ixp33_ASAP7_75t_SL U48284 ( .A1(n53628), .A2(n68970), .B(n53192), .C(
        n53628), .Y(n54289) );
  A2O1A1Ixp33_ASAP7_75t_SL U48285 ( .A1(n53628), .A2(n59671), .B(n53192), .C(
        n53628), .Y(n54291) );
  A2O1A1Ixp33_ASAP7_75t_SL U48286 ( .A1(n54290), .A2(n54291), .B(n53192), .C(
        n53628), .Y(n54292) );
  A2O1A1Ixp33_ASAP7_75t_SL U48287 ( .A1(n53628), .A2(n68986), .B(n53192), .C(
        n54295), .Y(n54296) );
  A2O1A1Ixp33_ASAP7_75t_SL U48288 ( .A1(n54292), .A2(n54293), .B(n53192), .C(
        n54296), .Y(n54297) );
  A2O1A1Ixp33_ASAP7_75t_SL U48289 ( .A1(n53628), .A2(n68969), .B(n53192), .C(
        n53628), .Y(n54298) );
  A2O1A1Ixp33_ASAP7_75t_SL U48290 ( .A1(n68986), .A2(n54298), .B(n53192), .C(
        n53628), .Y(n54299) );
  A2O1A1Ixp33_ASAP7_75t_SL U48291 ( .A1(n57080), .A2(n54299), .B(n53192), .C(
        n53628), .Y(n54300) );
  A2O1A1Ixp33_ASAP7_75t_SL U48292 ( .A1(n54302), .A2(n54303), .B(n53192), .C(
        n53628), .Y(n54304) );
  A2O1A1Ixp33_ASAP7_75t_SL U48293 ( .A1(n53628), .A2(n54304), .B(n53192), .C(
        n53628), .Y(n54305) );
  A2O1A1Ixp33_ASAP7_75t_SL U48294 ( .A1(n54297), .A2(n54306), .B(n53192), .C(
        n53628), .Y(n54307) );
  A2O1A1Ixp33_ASAP7_75t_SL U48295 ( .A1(n69256), .A2(n75650), .B(n53192), .C(
        n53628), .Y(n54278) );
  A2O1A1Ixp33_ASAP7_75t_SL U48296 ( .A1(n77875), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n54279) );
  A2O1A1Ixp33_ASAP7_75t_SL U48297 ( .A1(n69253), .A2(n54282), .B(n53192), .C(
        n53628), .Y(n54283) );
  A2O1A1Ixp33_ASAP7_75t_SL U48298 ( .A1(n54278), .A2(n54279), .B(n53192), .C(
        n54287), .Y(or1200_cpu_or1200_mult_mac_n1602) );
  A2O1A1Ixp33_ASAP7_75t_SL U48299 ( .A1(n76681), .A2(n57072), .B(n53192), .C(
        n53628), .Y(n54130) );
  A2O1A1Ixp33_ASAP7_75t_SL U48300 ( .A1(n57093), .A2(n76253), .B(n53192), .C(
        n53628), .Y(n54277) );
  A2O1A1Ixp33_ASAP7_75t_SL U48301 ( .A1(n77288), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n54128) );
  A2O1A1Ixp33_ASAP7_75t_SL U48302 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .A2(
        n72484), .B(n53192), .C(n53628), .Y(n54275) );
  A2O1A1Ixp33_ASAP7_75t_SL U48303 ( .A1(n72486), .A2(n54274), .B(n53192), .C(
        n54275), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n65) );
  A2O1A1Ixp33_ASAP7_75t_SL U48304 ( .A1(n71099), .A2(n71130), .B(n53192), .C(
        n71098), .Y(n54264) );
  A2O1A1Ixp33_ASAP7_75t_SL U48305 ( .A1(n57211), .A2(n54265), .B(n53192), .C(
        n53628), .Y(n54266) );
  A2O1A1Ixp33_ASAP7_75t_SL U48306 ( .A1(n53192), .A2(n53628), .B(n53890), .C(
        n53628), .Y(n70475) );
  A2O1A1Ixp33_ASAP7_75t_SL U48307 ( .A1(n62477), .A2(dbg_dat_i[1]), .B(n53192), 
        .C(n53628), .Y(n54257) );
  A2O1A1Ixp33_ASAP7_75t_SL U48308 ( .A1(n75672), .A2(n75671), .B(n53192), .C(
        n53628), .Y(n54250) );
  A2O1A1Ixp33_ASAP7_75t_SL U48309 ( .A1(n54072), .A2(n71801), .B(n53192), .C(
        n71795), .Y(n71709) );
  A2O1A1Ixp33_ASAP7_75t_SL U48310 ( .A1(n72596), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_), .B(
        n53192), .C(n54071), .Y(n74253) );
  A2O1A1Ixp33_ASAP7_75t_SL U48311 ( .A1(n54243), .A2(n54244), .B(n53192), .C(
        n53628), .Y(n54245) );
  A2O1A1Ixp33_ASAP7_75t_SL U48312 ( .A1(n72316), .A2(n54241), .B(n53192), .C(
        n53628), .Y(n54242) );
  A2O1A1Ixp33_ASAP7_75t_SL U48313 ( .A1(n71428), .A2(n54242), .B(n53192), .C(
        n53628), .Y(n71506) );
  A2O1A1Ixp33_ASAP7_75t_SL U48314 ( .A1(n71496), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54239) );
  A2O1A1Ixp33_ASAP7_75t_SL U48315 ( .A1(n71471), .A2(n54239), .B(n53192), .C(
        n53628), .Y(n54240) );
  A2O1A1Ixp33_ASAP7_75t_SL U48316 ( .A1(n71472), .A2(n54240), .B(n53192), .C(
        n53628), .Y(n71488) );
  A2O1A1Ixp33_ASAP7_75t_SL U48317 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[36]), .A2(n66182), 
        .B(n53192), .C(n53628), .Y(n54236) );
  A2O1A1Ixp33_ASAP7_75t_SL U48318 ( .A1(n73047), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[0]), .B(n53192), 
        .C(n53628), .Y(n54235) );
  A2O1A1Ixp33_ASAP7_75t_SL U48319 ( .A1(n57205), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[9]), .B(n53192), .C(
        n53628), .Y(n54230) );
  A2O1A1Ixp33_ASAP7_75t_SL U48320 ( .A1(n57217), .A2(n73695), .B(n53192), .C(
        n53628), .Y(n54231) );
  A2O1A1Ixp33_ASAP7_75t_SL U48321 ( .A1(n54230), .A2(n54231), .B(n53192), .C(
        n53628), .Y(n54232) );
  A2O1A1Ixp33_ASAP7_75t_SL U48322 ( .A1(n57204), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[8]), .B(n53192), .C(
        n53628), .Y(n54234) );
  A2O1A1Ixp33_ASAP7_75t_SL U48323 ( .A1(n54233), .A2(n54234), .B(n53192), .C(
        n53628), .Y(n73722) );
  A2O1A1Ixp33_ASAP7_75t_SL U48324 ( .A1(n77082), .A2(n54226), .B(n53192), .C(
        n53628), .Y(n54227) );
  A2O1A1Ixp33_ASAP7_75t_SL U48325 ( .A1(n77091), .A2(
        or1200_cpu_or1200_fpu_result_arith[5]), .B(n53192), .C(n53628), .Y(
        n54228) );
  A2O1A1Ixp33_ASAP7_75t_SL U48326 ( .A1(n54227), .A2(n54228), .B(n53192), .C(
        n53628), .Y(n54229) );
  A2O1A1Ixp33_ASAP7_75t_SL U48327 ( .A1(n53628), .A2(n54229), .B(n53192), .C(
        n53628), .Y(n61654) );
  A2O1A1Ixp33_ASAP7_75t_SL U48328 ( .A1(n75427), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54222) );
  A2O1A1Ixp33_ASAP7_75t_SL U48329 ( .A1(n75425), .A2(n54222), .B(n53192), .C(
        n53628), .Y(n54223) );
  A2O1A1Ixp33_ASAP7_75t_SL U48330 ( .A1(n54221), .A2(n54223), .B(n53192), .C(
        n53628), .Y(n75429) );
  A2O1A1Ixp33_ASAP7_75t_SL U48331 ( .A1(n60979), .A2(n54216), .B(n53192), .C(
        n54218), .Y(n54219) );
  A2O1A1Ixp33_ASAP7_75t_SL U48332 ( .A1(n75644), .A2(n59668), .B(n53192), .C(
        n53628), .Y(n54214) );
  A2O1A1Ixp33_ASAP7_75t_SL U48333 ( .A1(n75032), .A2(n75031), .B(n53192), .C(
        n75077), .Y(n54215) );
  A2O1A1Ixp33_ASAP7_75t_SL U48334 ( .A1(n71356), .A2(n58315), .B(n53192), .C(
        n53628), .Y(n54211) );
  A2O1A1Ixp33_ASAP7_75t_SL U48335 ( .A1(n57900), .A2(n63114), .B(n53192), .C(
        n58481), .Y(n54210) );
  A2O1A1Ixp33_ASAP7_75t_SL U48336 ( .A1(n73807), .A2(n73813), .B(n53192), .C(
        n53628), .Y(n54205) );
  A2O1A1Ixp33_ASAP7_75t_SL U48337 ( .A1(n54204), .A2(n54205), .B(n53192), .C(
        n53628), .Y(n3294) );
  A2O1A1Ixp33_ASAP7_75t_SL U48338 ( .A1(n70061), .A2(n69872), .B(n53192), .C(
        n53628), .Y(n54200) );
  A2O1A1Ixp33_ASAP7_75t_SL U48339 ( .A1(n54199), .A2(n54200), .B(n53192), .C(
        n53628), .Y(n54201) );
  A2O1A1Ixp33_ASAP7_75t_SL U48340 ( .A1(n53628), .A2(n54201), .B(n53192), .C(
        n53628), .Y(n54202) );
  A2O1A1Ixp33_ASAP7_75t_SL U48341 ( .A1(n70597), .A2(n54198), .B(n53192), .C(
        n53628), .Y(n3158) );
  A2O1A1Ixp33_ASAP7_75t_SL U48342 ( .A1(n59629), .A2(n72793), .B(n53192), .C(
        n53628), .Y(n54195) );
  A2O1A1Ixp33_ASAP7_75t_SL U48343 ( .A1(n59629), .A2(n78334), .B(n53192), .C(
        n53628), .Y(n54194) );
  A2O1A1Ixp33_ASAP7_75t_SL U48344 ( .A1(n54190), .A2(n54191), .B(n53192), .C(
        n53628), .Y(n9235) );
  A2O1A1Ixp33_ASAP7_75t_SL U48345 ( .A1(n59621), .A2(n54185), .B(n53192), .C(
        n53628), .Y(n54186) );
  A2O1A1Ixp33_ASAP7_75t_SL U48346 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[18]), .A2(n54187), 
        .B(n53192), .C(n53628), .Y(n54188) );
  A2O1A1Ixp33_ASAP7_75t_SL U48347 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .A2(
        n70484), .B(n53192), .C(n53628), .Y(n54177) );
  A2O1A1Ixp33_ASAP7_75t_SL U48348 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .A2(
        n70482), .B(n53192), .C(n53628), .Y(n54178) );
  A2O1A1Ixp33_ASAP7_75t_SL U48349 ( .A1(n70490), .A2(n70386), .B(n53192), .C(
        n53628), .Y(n54180) );
  A2O1A1Ixp33_ASAP7_75t_SL U48350 ( .A1(n54179), .A2(n54180), .B(n53192), .C(
        n53628), .Y(n54181) );
  A2O1A1Ixp33_ASAP7_75t_SL U48351 ( .A1(n74656), .A2(n70476), .B(n53192), .C(
        n53628), .Y(n54182) );
  A2O1A1Ixp33_ASAP7_75t_SL U48352 ( .A1(n70485), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_9_), .B(
        n53192), .C(n53628), .Y(n54183) );
  A2O1A1Ixp33_ASAP7_75t_SL U48353 ( .A1(n54181), .A2(n54182), .B(n53192), .C(
        n54183), .Y(n54184) );
  A2O1A1Ixp33_ASAP7_75t_SL U48354 ( .A1(n54177), .A2(n54178), .B(n53192), .C(
        n54184), .Y(n2425) );
  A2O1A1Ixp33_ASAP7_75t_SL U48355 ( .A1(n65402), .A2(n54166), .B(n53192), .C(
        n53628), .Y(n2007) );
  A2O1A1Ixp33_ASAP7_75t_SL U48356 ( .A1(n77983), .A2(n59680), .B(n53192), .C(
        n53628), .Y(n54162) );
  A2O1A1Ixp33_ASAP7_75t_SL U48357 ( .A1(n54163), .A2(n54164), .B(n53192), .C(
        n53628), .Y(n54165) );
  A2O1A1Ixp33_ASAP7_75t_SL U48358 ( .A1(n54162), .A2(n54165), .B(n53192), .C(
        n53628), .Y(n58417) );
  A2O1A1Ixp33_ASAP7_75t_SL U48359 ( .A1(n58296), .A2(n76235), .B(n53192), .C(
        n53628), .Y(n54155) );
  A2O1A1Ixp33_ASAP7_75t_SL U48360 ( .A1(or1200_cpu_or1200_except_n252), .A2(
        n57198), .B(n53192), .C(n53628), .Y(n54156) );
  A2O1A1Ixp33_ASAP7_75t_SL U48361 ( .A1(n54155), .A2(n54156), .B(n53192), .C(
        n53628), .Y(n54157) );
  A2O1A1Ixp33_ASAP7_75t_SL U48362 ( .A1(n57114), .A2(n77899), .B(n53192), .C(
        n53628), .Y(n54148) );
  A2O1A1Ixp33_ASAP7_75t_SL U48363 ( .A1(n54132), .A2(n54133), .B(n53192), .C(
        n53628), .Y(n54134) );
  A2O1A1Ixp33_ASAP7_75t_SL U48364 ( .A1(n63350), .A2(n54137), .B(n53192), .C(
        n53628), .Y(n54139) );
  A2O1A1Ixp33_ASAP7_75t_SL U48365 ( .A1(n59674), .A2(n54139), .B(n53192), .C(
        n53628), .Y(n54140) );
  A2O1A1Ixp33_ASAP7_75t_SL U48366 ( .A1(n53628), .A2(n68841), .B(n53192), .C(
        n53628), .Y(n53956) );
  A2O1A1Ixp33_ASAP7_75t_SL U48367 ( .A1(n53628), .A2(n53957), .B(n53192), .C(
        n53628), .Y(n53958) );
  A2O1A1Ixp33_ASAP7_75t_SL U48368 ( .A1(n76999), .A2(n57093), .B(n53192), .C(
        n53628), .Y(n53953) );
  A2O1A1Ixp33_ASAP7_75t_SL U48369 ( .A1(n57093), .A2(n76704), .B(n53192), .C(
        n53628), .Y(n54129) );
  A2O1A1Ixp33_ASAP7_75t_SL U48370 ( .A1(n71469), .A2(n71591), .B(n53192), .C(
        n53628), .Y(n54108) );
  A2O1A1Ixp33_ASAP7_75t_SL U48371 ( .A1(n71470), .A2(n71605), .B(n53192), .C(
        n72212), .Y(n54111) );
  A2O1A1Ixp33_ASAP7_75t_SL U48372 ( .A1(n54110), .A2(n54111), .B(n53192), .C(
        n53628), .Y(n54112) );
  A2O1A1Ixp33_ASAP7_75t_SL U48373 ( .A1(n71485), .A2(n54114), .B(n53192), .C(
        n53628), .Y(n54115) );
  A2O1A1Ixp33_ASAP7_75t_SL U48374 ( .A1(n54113), .A2(n54115), .B(n53192), .C(
        n53628), .Y(n54116) );
  A2O1A1Ixp33_ASAP7_75t_SL U48375 ( .A1(n59698), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n53933) );
  A2O1A1Ixp33_ASAP7_75t_SL U48376 ( .A1(n53628), .A2(n53934), .B(n53192), .C(
        n53628), .Y(n53935) );
  A2O1A1Ixp33_ASAP7_75t_SL U48377 ( .A1(n57211), .A2(n54100), .B(n53192), .C(
        n53628), .Y(n54102) );
  A2O1A1Ixp33_ASAP7_75t_SL U48378 ( .A1(n54097), .A2(n71186), .B(n53192), .C(
        n54102), .Y(n54103) );
  A2O1A1Ixp33_ASAP7_75t_SL U48379 ( .A1(n61996), .A2(n54096), .B(n53192), .C(
        n53628), .Y(n77472) );
  A2O1A1Ixp33_ASAP7_75t_SL U48380 ( .A1(n77754), .A2(n54094), .B(n53192), .C(
        n53628), .Y(n54095) );
  A2O1A1Ixp33_ASAP7_75t_SL U48381 ( .A1(n77760), .A2(n54095), .B(n53192), .C(
        n53628), .Y(n3906) );
  A2O1A1Ixp33_ASAP7_75t_SL U48382 ( .A1(n62477), .A2(dbg_dat_i[30]), .B(n53192), .C(n53628), .Y(n54092) );
  A2O1A1Ixp33_ASAP7_75t_SL U48383 ( .A1(n62477), .A2(dbg_dat_i[20]), .B(n53192), .C(n53628), .Y(n54091) );
  A2O1A1Ixp33_ASAP7_75t_SL U48384 ( .A1(n73893), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[5]), .B(
        n53192), .C(n53628), .Y(n54090) );
  A2O1A1Ixp33_ASAP7_75t_SL U48385 ( .A1(n54089), .A2(n54090), .B(n53192), .C(
        n53628), .Y(n74278) );
  A2O1A1Ixp33_ASAP7_75t_SL U48386 ( .A1(n62477), .A2(dbg_dat_i[31]), .B(n53192), .C(n53628), .Y(n54086) );
  A2O1A1Ixp33_ASAP7_75t_SL U48387 ( .A1(n76546), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n54082) );
  A2O1A1Ixp33_ASAP7_75t_SL U48388 ( .A1(n76547), .A2(n54082), .B(n53192), .C(
        n53628), .Y(n54083) );
  A2O1A1Ixp33_ASAP7_75t_SL U48389 ( .A1(n53628), .A2(n54083), .B(n53192), .C(
        n53628), .Y(n54084) );
  A2O1A1Ixp33_ASAP7_75t_SL U48390 ( .A1(n63534), .A2(n63515), .B(n53192), .C(
        n53628), .Y(n54078) );
  A2O1A1Ixp33_ASAP7_75t_SL U48391 ( .A1(n63539), .A2(n54078), .B(n53192), .C(
        n53628), .Y(n54079) );
  A2O1A1Ixp33_ASAP7_75t_SL U48392 ( .A1(n53628), .A2(n54079), .B(n53192), .C(
        n53628), .Y(n63516) );
  A2O1A1Ixp33_ASAP7_75t_SL U48393 ( .A1(n70793), .A2(n70792), .B(n53192), .C(
        n53628), .Y(n54066) );
  A2O1A1Ixp33_ASAP7_75t_SL U48394 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .A2(n66182), 
        .B(n53192), .C(n53628), .Y(n54063) );
  A2O1A1Ixp33_ASAP7_75t_SL U48395 ( .A1(n57194), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .B(n53192), 
        .C(n53628), .Y(n54054) );
  A2O1A1Ixp33_ASAP7_75t_SL U48396 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]), .A2(n57193), 
        .B(n53192), .C(n53628), .Y(n54055) );
  A2O1A1Ixp33_ASAP7_75t_SL U48397 ( .A1(n54054), .A2(n54055), .B(n53192), .C(
        n53628), .Y(n54056) );
  A2O1A1Ixp33_ASAP7_75t_SL U48398 ( .A1(n57188), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .B(n53192), 
        .C(n53628), .Y(n54058) );
  A2O1A1Ixp33_ASAP7_75t_SL U48399 ( .A1(n54057), .A2(n54058), .B(n53192), .C(
        n53628), .Y(n66016) );
  A2O1A1Ixp33_ASAP7_75t_SL U48400 ( .A1(n74686), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_15_), .B(
        n53192), .C(n53628), .Y(n54046) );
  A2O1A1Ixp33_ASAP7_75t_SL U48401 ( .A1(n54045), .A2(n54046), .B(n53192), .C(
        n53628), .Y(n54047) );
  A2O1A1Ixp33_ASAP7_75t_SL U48402 ( .A1(n53628), .A2(n54047), .B(n53192), .C(
        n53628), .Y(n54048) );
  A2O1A1Ixp33_ASAP7_75t_SL U48403 ( .A1(n54043), .A2(n54044), .B(n53192), .C(
        n53628), .Y(n64806) );
  A2O1A1Ixp33_ASAP7_75t_SL U48404 ( .A1(n57194), .A2(n65823), .B(n53192), .C(
        n53628), .Y(n54035) );
  A2O1A1Ixp33_ASAP7_75t_SL U48405 ( .A1(n65821), .A2(n57193), .B(n53192), .C(
        n53628), .Y(n54036) );
  A2O1A1Ixp33_ASAP7_75t_SL U48406 ( .A1(n54035), .A2(n54036), .B(n53192), .C(
        n53628), .Y(n54037) );
  A2O1A1Ixp33_ASAP7_75t_SL U48407 ( .A1(n57188), .A2(n65784), .B(n53192), .C(
        n53628), .Y(n54039) );
  A2O1A1Ixp33_ASAP7_75t_SL U48408 ( .A1(n54038), .A2(n54039), .B(n53192), .C(
        n53628), .Y(n65928) );
  A2O1A1Ixp33_ASAP7_75t_SL U48409 ( .A1(n70996), .A2(n54033), .B(n53192), .C(
        n53628), .Y(n70778) );
  A2O1A1Ixp33_ASAP7_75t_SL U48410 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[4]), .A2(
        n54032), .B(n53192), .C(n53628), .Y(n70167) );
  A2O1A1Ixp33_ASAP7_75t_SL U48411 ( .A1(n62629), .A2(n57120), .B(n53192), .C(
        n53838), .Y(n53839) );
  A2O1A1Ixp33_ASAP7_75t_SL U48412 ( .A1(n62629), .A2(n57120), .B(n53192), .C(
        n53628), .Y(n53840) );
  A2O1A1Ixp33_ASAP7_75t_SL U48413 ( .A1(n53840), .A2(n59554), .B(n53192), .C(
        n53628), .Y(n53841) );
  A2O1A1Ixp33_ASAP7_75t_SL U48414 ( .A1(n53839), .A2(n53841), .B(n53192), .C(
        n53628), .Y(n60772) );
  A2O1A1Ixp33_ASAP7_75t_SL U48415 ( .A1(n66750), .A2(n67306), .B(n53192), .C(
        n53628), .Y(n54027) );
  A2O1A1Ixp33_ASAP7_75t_SL U48416 ( .A1(n57239), .A2(n54022), .B(n53192), .C(
        n53628), .Y(n54023) );
  A2O1A1Ixp33_ASAP7_75t_SL U48417 ( .A1(n59653), .A2(n59642), .B(n53192), .C(
        n53628), .Y(n54021) );
  A2O1A1Ixp33_ASAP7_75t_SL U48418 ( .A1(n53192), .A2(n53628), .B(n53823), .C(
        n53628), .Y(n53824) );
  A2O1A1Ixp33_ASAP7_75t_SL U48419 ( .A1(n53824), .A2(n53825), .B(n53192), .C(
        n53628), .Y(n78212) );
  A2O1A1Ixp33_ASAP7_75t_SL U48420 ( .A1(n53818), .A2(n53819), .B(n53192), .C(
        n53628), .Y(n3210) );
  A2O1A1Ixp33_ASAP7_75t_SL U48421 ( .A1(n59690), .A2(n54017), .B(n53192), .C(
        n53628), .Y(n54018) );
  A2O1A1Ixp33_ASAP7_75t_SL U48422 ( .A1(n53192), .A2(n53628), .B(n53809), .C(
        n53628), .Y(n53810) );
  A2O1A1Ixp33_ASAP7_75t_SL U48423 ( .A1(n78436), .A2(n74797), .B(n53192), .C(
        n53628), .Y(n53807) );
  A2O1A1Ixp33_ASAP7_75t_SL U48424 ( .A1(n70296), .A2(n70103), .B(n53192), .C(
        n53628), .Y(n53804) );
  A2O1A1Ixp33_ASAP7_75t_SL U48425 ( .A1(n74538), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[10]), .B(n53192), 
        .C(n53628), .Y(n53800) );
  A2O1A1Ixp33_ASAP7_75t_SL U48426 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[10]), .A2(n53801), 
        .B(n53192), .C(n53628), .Y(n53802) );
  A2O1A1Ixp33_ASAP7_75t_SL U48427 ( .A1(n78437), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[10]), .B(
        n53192), .C(n53628), .Y(n53803) );
  A2O1A1Ixp33_ASAP7_75t_SL U48428 ( .A1(n53800), .A2(n53802), .B(n53192), .C(
        n53803), .Y(or1200_cpu_or1200_fpu_fpu_arith_N93) );
  A2O1A1Ixp33_ASAP7_75t_SL U48429 ( .A1(n62059), .A2(n54013), .B(n53192), .C(
        n53628), .Y(n54014) );
  A2O1A1Ixp33_ASAP7_75t_SL U48430 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_2_), .A2(n62064), .B(n53192), 
        .C(n53628), .Y(n54015) );
  A2O1A1Ixp33_ASAP7_75t_SL U48431 ( .A1(n54014), .A2(n54015), .B(n53192), .C(
        n53628), .Y(n54016) );
  A2O1A1Ixp33_ASAP7_75t_SL U48432 ( .A1(n53628), .A2(n54016), .B(n53192), .C(
        n53628), .Y(n2204) );
  A2O1A1Ixp33_ASAP7_75t_SL U48433 ( .A1(n77925), .A2(n59691), .B(n53192), .C(
        n53628), .Y(n53797) );
  A2O1A1Ixp33_ASAP7_75t_SL U48434 ( .A1(n72870), .A2(n59629), .B(n53192), .C(
        n53628), .Y(n53796) );
  A2O1A1Ixp33_ASAP7_75t_SL U48435 ( .A1(n65400), .A2(n65392), .B(n53192), .C(
        n53628), .Y(n54010) );
  A2O1A1Ixp33_ASAP7_75t_SL U48436 ( .A1(n65395), .A2(n54009), .B(n53192), .C(
        n54011), .Y(n1992) );
  A2O1A1Ixp33_ASAP7_75t_SL U48437 ( .A1(n57114), .A2(n77896), .B(n53192), .C(
        n53628), .Y(n54004) );
  A2O1A1Ixp33_ASAP7_75t_SL U48438 ( .A1(n1376), .A2(n53999), .B(n53192), .C(
        n53628), .Y(n54000) );
  A2O1A1Ixp33_ASAP7_75t_SL U48439 ( .A1(n77287), .A2(n77637), .B(n53192), .C(
        n53628), .Y(n54001) );
  A2O1A1Ixp33_ASAP7_75t_SL U48440 ( .A1(n54000), .A2(n54001), .B(n53192), .C(
        n53628), .Y(n54002) );
  A2O1A1Ixp33_ASAP7_75t_SL U48441 ( .A1(n54002), .A2(n54003), .B(n53192), .C(
        n53628), .Y(or1200_pic_N60) );
  A2O1A1Ixp33_ASAP7_75t_SL U48442 ( .A1(n74641), .A2(n77890), .B(n53192), .C(
        n53628), .Y(n53998) );
  A2O1A1Ixp33_ASAP7_75t_SL U48443 ( .A1(or1200_cpu_or1200_mult_mac_n280), .A2(
        n53986), .B(n53192), .C(n62557), .Y(n53987) );
  A2O1A1Ixp33_ASAP7_75t_SL U48444 ( .A1(or1200_cpu_or1200_mult_mac_n282), .A2(
        or1200_cpu_or1200_mult_mac_n278), .B(n53192), .C(n53628), .Y(n53988)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U48445 ( .A1(n75015), .A2(n77922), .B(n53192), .C(
        n53628), .Y(n53984) );
  A2O1A1Ixp33_ASAP7_75t_SL U48446 ( .A1(n53983), .A2(n53984), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_mult_mac_n1625) );
  A2O1A1Ixp33_ASAP7_75t_SL U48447 ( .A1(n63513), .A2(n53970), .B(n53192), .C(
        n53628), .Y(n53971) );
  A2O1A1Ixp33_ASAP7_75t_SL U48448 ( .A1(n53969), .A2(n53971), .B(n53192), .C(
        n53628), .Y(n53972) );
  A2O1A1Ixp33_ASAP7_75t_SL U48449 ( .A1(n68843), .A2(n53956), .B(n53192), .C(
        n53628), .Y(n53957) );
  A2O1A1Ixp33_ASAP7_75t_SL U48450 ( .A1(n57072), .A2(n75783), .B(n53192), .C(
        n53628), .Y(n53952) );
  A2O1A1Ixp33_ASAP7_75t_SL U48451 ( .A1(n74275), .A2(n53950), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n53) );
  A2O1A1Ixp33_ASAP7_75t_SL U48452 ( .A1(n72469), .A2(n53947), .B(n53192), .C(
        n53628), .Y(n53948) );
  A2O1A1Ixp33_ASAP7_75t_SL U48453 ( .A1(n53945), .A2(n53946), .B(n53192), .C(
        n53628), .Y(n53947) );
  A2O1A1Ixp33_ASAP7_75t_SL U48454 ( .A1(n53942), .A2(n53943), .B(n53192), .C(
        n53628), .Y(n53944) );
  A2O1A1Ixp33_ASAP7_75t_SL U48455 ( .A1(n72493), .A2(n72433), .B(n53192), .C(
        n53628), .Y(n53943) );
  A2O1A1Ixp33_ASAP7_75t_SL U48456 ( .A1(n59625), .A2(n72489), .B(n53192), .C(
        n53628), .Y(n53940) );
  A2O1A1O1Ixp25_ASAP7_75t_SL U48457 ( .A1(n71689), .A2(n71690), .B(n53192), 
        .C(n71735), .D(n71688), .Y(n53938) );
  A2O1A1Ixp33_ASAP7_75t_SL U48458 ( .A1(n53628), .A2(n59699), .B(n53192), .C(
        n53628), .Y(n53726) );
  A2O1A1Ixp33_ASAP7_75t_SL U48459 ( .A1(n70753), .A2(n53727), .B(n53192), .C(
        n53628), .Y(n53728) );
  A2O1A1Ixp33_ASAP7_75t_SL U48460 ( .A1(n71030), .A2(n53933), .B(n53192), .C(
        n53628), .Y(n53934) );
  A2O1A1Ixp33_ASAP7_75t_SL U48461 ( .A1(n71114), .A2(n71111), .B(n53192), .C(
        n53628), .Y(n53930) );
  A2O1A1Ixp33_ASAP7_75t_SL U48462 ( .A1(n71112), .A2(n53930), .B(n53192), .C(
        n53628), .Y(n53931) );
  A2O1A1Ixp33_ASAP7_75t_SL U48463 ( .A1(n59699), .A2(n78398), .B(n53192), .C(
        n53628), .Y(n53932) );
  A2O1A1Ixp33_ASAP7_75t_SL U48464 ( .A1(n66152), .A2(n66151), .B(n53192), .C(
        n53628), .Y(n53913) );
  A2O1A1Ixp33_ASAP7_75t_SL U48465 ( .A1(n66146), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[46]), .B(n53192), 
        .C(n53628), .Y(n53924) );
  A2O1A1Ixp33_ASAP7_75t_SL U48466 ( .A1(n66182), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[47]), .B(n53192), 
        .C(n53628), .Y(n53925) );
  A2O1A1Ixp33_ASAP7_75t_SL U48467 ( .A1(n53924), .A2(n53925), .B(n53192), .C(
        n53628), .Y(n53926) );
  A2O1A1Ixp33_ASAP7_75t_SL U48468 ( .A1(n73572), .A2(n53912), .B(n53192), .C(
        n53628), .Y(n73657) );
  A2O1A1Ixp33_ASAP7_75t_SL U48469 ( .A1(n77484), .A2(n53911), .B(n53192), .C(
        n53628), .Y(n61286) );
  A2O1A1Ixp33_ASAP7_75t_SL U48470 ( .A1(n57074), .A2(n53907), .B(n53192), .C(
        n53628), .Y(n76991) );
  A2O1A1Ixp33_ASAP7_75t_SL U48471 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_2_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_1_), .B(n53192), 
        .C(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_4_), .Y(n53898) );
  A2O1A1Ixp33_ASAP7_75t_SL U48472 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_12_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_14_), .B(n53192), 
        .C(n53628), .Y(n53899) );
  A2O1A1Ixp33_ASAP7_75t_SL U48473 ( .A1(n53897), .A2(n53904), .B(n53192), .C(
        n53905), .Y(n53906) );
  A2O1A1Ixp33_ASAP7_75t_SL U48474 ( .A1(n69109), .A2(n69110), .B(n53192), .C(
        n53628), .Y(n53889) );
  A2O1A1Ixp33_ASAP7_75t_SL U48475 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_36_), .A2(n53879), 
        .B(n53192), .C(n53628), .Y(n71236) );
  A2O1A1Ixp33_ASAP7_75t_SL U48476 ( .A1(n53628), .A2(n72723), .B(n53192), .C(
        n53628), .Y(n53875) );
  A2O1A1Ixp33_ASAP7_75t_SL U48477 ( .A1(n53874), .A2(n53876), .B(n53192), .C(
        n53628), .Y(n53877) );
  A2O1A1Ixp33_ASAP7_75t_SL U48478 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[5]), .A2(n59632), .B(
        n53192), .C(n53628), .Y(n53866) );
  A2O1A1Ixp33_ASAP7_75t_SL U48479 ( .A1(n73823), .A2(n57204), .B(n53192), .C(
        n53628), .Y(n53867) );
  A2O1A1Ixp33_ASAP7_75t_SL U48480 ( .A1(n53866), .A2(n53867), .B(n53192), .C(
        n53628), .Y(n53868) );
  A2O1A1Ixp33_ASAP7_75t_SL U48481 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[7]), .A2(n57205), .B(
        n53192), .C(n53628), .Y(n53870) );
  A2O1A1Ixp33_ASAP7_75t_SL U48482 ( .A1(n53869), .A2(n53870), .B(n53192), .C(
        n53628), .Y(n73751) );
  A2O1A1Ixp33_ASAP7_75t_SL U48483 ( .A1(n71513), .A2(n53865), .B(n53192), .C(
        n53628), .Y(n71515) );
  A2O1A1Ixp33_ASAP7_75t_SL U48484 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[6]), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .B(
        n53192), .C(n53628), .Y(n53864) );
  A2O1A1Ixp33_ASAP7_75t_SL U48485 ( .A1(n57121), .A2(n65095), .B(n53192), .C(
        n53628), .Y(n53861) );
  A2O1A1Ixp33_ASAP7_75t_SL U48486 ( .A1(n61525), .A2(n61538), .B(n53192), .C(
        n53860), .Y(n61224) );
  A2O1A1Ixp33_ASAP7_75t_SL U48487 ( .A1(or1200_cpu_or1200_fpu_result_conv[18]), 
        .A2(n77090), .B(n53192), .C(n53628), .Y(n53857) );
  A2O1A1Ixp33_ASAP7_75t_SL U48488 ( .A1(n77091), .A2(
        or1200_cpu_or1200_fpu_result_arith[18]), .B(n53192), .C(n53628), .Y(
        n53858) );
  A2O1A1Ixp33_ASAP7_75t_SL U48489 ( .A1(n53857), .A2(n53858), .B(n53192), .C(
        n53628), .Y(n53859) );
  A2O1A1Ixp33_ASAP7_75t_SL U48490 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_13_), 
        .A2(n57207), .B(n53192), .C(n53628), .Y(n53849) );
  A2O1A1Ixp33_ASAP7_75t_SL U48491 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_), 
        .A2(n57216), .B(n53192), .C(n53628), .Y(n53850) );
  A2O1A1Ixp33_ASAP7_75t_SL U48492 ( .A1(n53849), .A2(n53850), .B(n53192), .C(
        n53628), .Y(n53851) );
  A2O1A1Ixp33_ASAP7_75t_SL U48493 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .A2(n71888), .B(n53192), .C(n53628), .Y(n53853) );
  A2O1A1Ixp33_ASAP7_75t_SL U48494 ( .A1(n53852), .A2(n53853), .B(n53192), .C(
        n53628), .Y(n72041) );
  A2O1A1Ixp33_ASAP7_75t_SL U48495 ( .A1(n68101), .A2(n67343), .B(n53192), .C(
        n53628), .Y(n53842) );
  NAND2xp5_ASAP7_75t_SL U48496 ( .A(n76028), .B(n64897), .Y(n53632) );
  A2O1A1Ixp33_ASAP7_75t_SL U48497 ( .A1(n66387), .A2(n53835), .B(n53192), .C(
        n53628), .Y(n53836) );
  A2O1A1Ixp33_ASAP7_75t_SL U48498 ( .A1(n67264), .A2(n67364), .B(n53192), .C(
        n53628), .Y(n53829) );
  A2O1A1Ixp33_ASAP7_75t_SL U48499 ( .A1(n77722), .A2(n53455), .B(n53192), .C(
        n53628), .Y(n53828) );
  A2O1A1Ixp33_ASAP7_75t_SL U48500 ( .A1(n59637), .A2(n57167), .B(n53192), .C(
        n53628), .Y(n53827) );
  A2O1A1Ixp33_ASAP7_75t_SL U48501 ( .A1(n73813), .A2(n73812), .B(n53192), .C(
        n53628), .Y(n53822) );
  A2O1A1Ixp33_ASAP7_75t_SL U48502 ( .A1(n73817), .A2(n53821), .B(n53192), .C(
        n53822), .Y(n3291) );
  A2O1A1Ixp33_ASAP7_75t_SL U48503 ( .A1(n70081), .A2(n69876), .B(n53192), .C(
        n53628), .Y(n53819) );
  A2O1A1Ixp33_ASAP7_75t_SL U48504 ( .A1(n59691), .A2(n53814), .B(n53192), .C(
        n53628), .Y(n53815) );
  A2O1A1Ixp33_ASAP7_75t_SL U48505 ( .A1(n2607), .A2(n53628), .B(n53192), .C(
        n53628), .Y(n53812) );
  A2O1A1Ixp33_ASAP7_75t_SL U48506 ( .A1(n62000), .A2(n53812), .B(n53192), .C(
        n53628), .Y(n53813) );
  A2O1A1Ixp33_ASAP7_75t_SL U48507 ( .A1(n53811), .A2(n53813), .B(n53192), .C(
        n53628), .Y(n60727) );
  A2O1A1Ixp33_ASAP7_75t_SL U48508 ( .A1(n62062), .A2(n62063), .B(n53192), .C(
        n53799), .Y(n2202) );
  A2O1A1Ixp33_ASAP7_75t_SL U48509 ( .A1(n72829), .A2(n59628), .B(n53192), .C(
        n53628), .Y(n53793) );
  A2O1A1Ixp33_ASAP7_75t_SL U48510 ( .A1(n77608), .A2(n77644), .B(n53192), .C(
        n53628), .Y(n53790) );
  A2O1A1Ixp33_ASAP7_75t_SL U48511 ( .A1(n77986), .A2(n77672), .B(n53192), .C(
        n53628), .Y(n53791) );
  A2O1A1Ixp33_ASAP7_75t_SL U48512 ( .A1(n53790), .A2(n53791), .B(n53192), .C(
        n53628), .Y(n53792) );
  A2O1A1Ixp33_ASAP7_75t_SL U48513 ( .A1(n57114), .A2(n77893), .B(n53192), .C(
        n53628), .Y(n53785) );
  A2O1A1Ixp33_ASAP7_75t_SL U48514 ( .A1(n74641), .A2(n77888), .B(n53192), .C(
        n53628), .Y(n53784) );
  A2O1A1Ixp33_ASAP7_75t_SL U48515 ( .A1(n75650), .A2(n68864), .B(n53192), .C(
        n53628), .Y(n53758) );
  A2O1A1Ixp33_ASAP7_75t_SL U48516 ( .A1(n77916), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n53759) );
  A2O1A1Ixp33_ASAP7_75t_SL U48517 ( .A1(n53764), .A2(n57079), .B(n53192), .C(
        n53628), .Y(n53765) );
  A2O1A1Ixp33_ASAP7_75t_SL U48518 ( .A1(n53763), .A2(n53765), .B(n53192), .C(
        n53628), .Y(n53766) );
  A2O1A1Ixp33_ASAP7_75t_SL U48519 ( .A1(n53768), .A2(n53769), .B(n53192), .C(
        n53628), .Y(n53770) );
  A2O1A1Ixp33_ASAP7_75t_SL U48520 ( .A1(n53758), .A2(n53759), .B(n53192), .C(
        n53771), .Y(or1200_cpu_or1200_mult_mac_n1621) );
  A2O1A1Ixp33_ASAP7_75t_SL U48521 ( .A1(n69024), .A2(n75650), .B(n53192), .C(
        n53628), .Y(n53746) );
  A2O1A1Ixp33_ASAP7_75t_SL U48522 ( .A1(n77968), .A2(n59673), .B(n53192), .C(
        n53628), .Y(n53747) );
  A2O1A1Ixp33_ASAP7_75t_SL U48523 ( .A1(n69061), .A2(n69066), .B(n53192), .C(
        n53628), .Y(n53750) );
  A2O1A1Ixp33_ASAP7_75t_SL U48524 ( .A1(n59672), .A2(n69072), .B(n53192), .C(
        n53628), .Y(n53751) );
  A2O1A1Ixp33_ASAP7_75t_SL U48525 ( .A1(n53750), .A2(n53751), .B(n53192), .C(
        n53628), .Y(n53752) );
  A2O1A1Ixp33_ASAP7_75t_SL U48526 ( .A1(n57080), .A2(n53748), .B(n53192), .C(
        n53628), .Y(n53755) );
  A2O1A1Ixp33_ASAP7_75t_SL U48527 ( .A1(n53754), .A2(n53755), .B(n53192), .C(
        n53628), .Y(n53756) );
  A2O1A1Ixp33_ASAP7_75t_SL U48528 ( .A1(n53746), .A2(n53747), .B(n53192), .C(
        n53757), .Y(or1200_cpu_or1200_mult_mac_n1614) );
  A2O1A1Ixp33_ASAP7_75t_SL U48529 ( .A1(or1200_cpu_to_sr[11]), .A2(n77217), 
        .B(n53192), .C(n53628), .Y(n53745) );
  A2O1A1Ixp33_ASAP7_75t_SL U48530 ( .A1(n53744), .A2(n53745), .B(n53192), .C(
        n53628), .Y(or1200_cpu_or1200_except_n1741) );
  A2O1A1Ixp33_ASAP7_75t_SL U48531 ( .A1(n57093), .A2(n75622), .B(n53192), .C(
        n53628), .Y(n53741) );
  A2O1A1Ixp33_ASAP7_75t_SL U48532 ( .A1(n72500), .A2(n53734), .B(n53192), .C(
        n53628), .Y(n53735) );
  A2O1A1Ixp33_ASAP7_75t_SL U48533 ( .A1(n70746), .A2(n53726), .B(n53192), .C(
        n53628), .Y(n53727) );
  A2O1A1Ixp33_ASAP7_75t_SL U48534 ( .A1(n71205), .A2(n71180), .B(n53192), .C(
        n53628), .Y(n53720) );
  A2O1A1Ixp33_ASAP7_75t_SL U48535 ( .A1(n53722), .A2(n53723), .B(n53192), .C(
        n53628), .Y(n53724) );
  A2O1A1Ixp33_ASAP7_75t_SL U48536 ( .A1(n70242), .A2(n53717), .B(n53192), .C(
        n53628), .Y(n3164) );
  A2O1A1Ixp33_ASAP7_75t_SL U48537 ( .A1(n70109), .A2(n53714), .B(n53192), .C(
        n53628), .Y(n69577) );
  A2O1A1Ixp33_ASAP7_75t_SL U48538 ( .A1(n76557), .A2(n2623), .B(n53192), .C(
        n53628), .Y(n53713) );
  A2O1A1Ixp33_ASAP7_75t_SL U48539 ( .A1(n53710), .A2(n53711), .B(n53192), .C(
        n53628), .Y(n53712) );
  A2O1A1Ixp33_ASAP7_75t_SL U48540 ( .A1(n53709), .A2(n53712), .B(n53192), .C(
        n53628), .Y(n77415) );
  A2O1A1Ixp33_ASAP7_75t_SL U48541 ( .A1(n64330), .A2(n53701), .B(n53192), .C(
        n53628), .Y(n77876) );
  A2O1A1Ixp33_ASAP7_75t_SL U48542 ( .A1(n74240), .A2(n74243), .B(n53192), .C(
        n53699), .Y(n74734) );
  A2O1A1Ixp33_ASAP7_75t_SL U48543 ( .A1(n74680), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_7_), .B(
        n53192), .C(n53628), .Y(n53696) );
  A2O1A1Ixp33_ASAP7_75t_SL U48544 ( .A1(n77233), .A2(n77162), .B(n53192), .C(
        n53628), .Y(n53695) );
  A2O1A1Ixp33_ASAP7_75t_SL U48545 ( .A1(n75661), .A2(n75662), .B(n53192), .C(
        n53628), .Y(n53688) );
  A2O1A1Ixp33_ASAP7_75t_SL U48546 ( .A1(n53688), .A2(n53689), .B(n53192), .C(
        n53628), .Y(n53690) );
  A2O1A1Ixp33_ASAP7_75t_SL U48547 ( .A1(n65670), .A2(n65587), .B(n53192), .C(
        n53628), .Y(n53681) );
  A2O1A1Ixp33_ASAP7_75t_SL U48548 ( .A1(n53680), .A2(n53681), .B(n53192), .C(
        n53628), .Y(n53682) );
  A2O1A1Ixp33_ASAP7_75t_SL U48549 ( .A1(n53628), .A2(n53682), .B(n53192), .C(
        n53628), .Y(n53683) );
  A2O1A1Ixp33_ASAP7_75t_SL U48550 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[33]), .A2(n57194), 
        .B(n53192), .C(n53628), .Y(n53675) );
  A2O1A1Ixp33_ASAP7_75t_SL U48551 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[32]), .A2(n57187), 
        .B(n53192), .C(n53628), .Y(n53676) );
  A2O1A1Ixp33_ASAP7_75t_SL U48552 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[31]), .A2(n57188), 
        .B(n53192), .C(n53628), .Y(n53679) );
  A2O1A1Ixp33_ASAP7_75t_SL U48553 ( .A1(n72642), .A2(n53673), .B(n53192), .C(
        n53628), .Y(n72664) );
  A2O1A1Ixp33_ASAP7_75t_SL U48554 ( .A1(n59631), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[17]), .B(
        n53192), .C(n53628), .Y(n53672) );
  A2O1A1Ixp33_ASAP7_75t_SL U48555 ( .A1(n76627), .A2(n59587), .B(n53192), .C(
        n53628), .Y(n53664) );
  A2O1A1Ixp33_ASAP7_75t_SL U48556 ( .A1(n77278), .A2(n59583), .B(n53192), .C(
        n53628), .Y(n53665) );
  A2O1A1Ixp33_ASAP7_75t_SL U48557 ( .A1(n60849), .A2(n53664), .B(n53192), .C(
        n53665), .Y(n53666) );
  A2O1A1Ixp33_ASAP7_75t_SL U48558 ( .A1(n61646), .A2(n61647), .B(n53192), .C(
        n53628), .Y(n53660) );
  A2O1A1Ixp33_ASAP7_75t_SL U48559 ( .A1(n61650), .A2(n53661), .B(n53192), .C(
        n53628), .Y(n53662) );
  A2O1A1Ixp33_ASAP7_75t_SL U48560 ( .A1(n61649), .A2(n53662), .B(n53192), .C(
        n53628), .Y(n53663) );
  A2O1A1Ixp33_ASAP7_75t_SL U48561 ( .A1(n61861), .A2(n53663), .B(n53192), .C(
        n53628), .Y(n61655) );
  A2O1A1Ixp33_ASAP7_75t_SL U48562 ( .A1(n61827), .A2(n64825), .B(n53192), .C(
        n53628), .Y(n53658) );
  A2O1A1Ixp33_ASAP7_75t_SL U48563 ( .A1(n65159), .A2(n57121), .B(n53192), .C(
        n53628), .Y(n53659) );
  A2O1A1Ixp33_ASAP7_75t_SL U48564 ( .A1(n76822), .A2(n53654), .B(n53192), .C(
        n53628), .Y(n74954) );
  A2O1A1Ixp33_ASAP7_75t_SL U48565 ( .A1(n72346), .A2(n57207), .B(n53192), .C(
        n53628), .Y(n53647) );
  A2O1A1Ixp33_ASAP7_75t_SL U48566 ( .A1(n57216), .A2(n72362), .B(n53192), .C(
        n53628), .Y(n53648) );
  A2O1A1Ixp33_ASAP7_75t_SL U48567 ( .A1(n53647), .A2(n53648), .B(n53192), .C(
        n53628), .Y(n53649) );
  A2O1A1Ixp33_ASAP7_75t_SL U48568 ( .A1(n72263), .A2(n71888), .B(n53192), .C(
        n53628), .Y(n53651) );
  A2O1A1Ixp33_ASAP7_75t_SL U48569 ( .A1(n53650), .A2(n53651), .B(n53192), .C(
        n53628), .Y(n72084) );
  A2O1A1Ixp33_ASAP7_75t_SL U48570 ( .A1(n71568), .A2(n72317), .B(n53192), .C(
        n53628), .Y(n53644) );
  A2O1A1Ixp33_ASAP7_75t_SL U48571 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .A2(n71263), .B(
        n53192), .C(n53628), .Y(n53639) );
  A2O1A1Ixp33_ASAP7_75t_SL U48572 ( .A1(n57067), .A2(n75074), .B(n53192), .C(
        n53628), .Y(n53636) );
  AND2x4_ASAP7_75t_SL U48573 ( .A(n66266), .B(n66269), .Y(n58807) );
  INVx5_ASAP7_75t_SL U48574 ( .A(n58807), .Y(n59637) );
  NAND2x1_ASAP7_75t_SL U48575 ( .A(n66924), .B(n53201), .Y(n66925) );
  NAND2xp5_ASAP7_75t_SRAM U48576 ( .A(n76057), .B(n67951), .Y(n67847) );
  NAND2xp5_ASAP7_75t_SL U48577 ( .A(n67593), .B(n57818), .Y(n57893) );
  BUFx5_ASAP7_75t_SL U48578 ( .A(n68724), .Y(n53193) );
  INVx1_ASAP7_75t_SL U48579 ( .A(n59477), .Y(n58232) );
  NAND2x1_ASAP7_75t_SL U48580 ( .A(n59477), .B(n66798), .Y(n63826) );
  NOR2x1p5_ASAP7_75t_SL U48581 ( .A(n63123), .B(n63081), .Y(n59477) );
  XNOR2x1_ASAP7_75t_SL U48582 ( .A(n59616), .B(n68087), .Y(n68088) );
  NOR2x1p5_ASAP7_75t_SL U48583 ( .A(n68088), .B(n68383), .Y(n68157) );
  NAND2xp5_ASAP7_75t_SL U48584 ( .A(n53194), .B(n63828), .Y(n63829) );
  INVx1_ASAP7_75t_SL U48585 ( .A(n53195), .Y(n53194) );
  NOR2x1_ASAP7_75t_SL U48586 ( .A(n67228), .B(n67739), .Y(n53195) );
  O2A1O1Ixp5_ASAP7_75t_SL U48587 ( .A1(n58861), .A2(n67866), .B(n53196), .C(
        n64360), .Y(n64476) );
  NAND2xp5_ASAP7_75t_SL U48588 ( .A(n58861), .B(n57422), .Y(n53196) );
  OAI21x1_ASAP7_75t_SL U48589 ( .A1(n63210), .A2(n57097), .B(n56845), .Y(
        n63211) );
  INVx3_ASAP7_75t_SL U48590 ( .A(n62649), .Y(n58424) );
  BUFx5_ASAP7_75t_SL U48591 ( .A(n59619), .Y(n53197) );
  INVx2_ASAP7_75t_SL U48592 ( .A(n53198), .Y(n59011) );
  NAND2x1_ASAP7_75t_SL U48593 ( .A(n68693), .B(n75276), .Y(n53198) );
  NAND2x1_ASAP7_75t_SL U48594 ( .A(n75275), .B(n75274), .Y(n75276) );
  BUFx5_ASAP7_75t_SL U48595 ( .A(n68853), .Y(n53199) );
  INVx1_ASAP7_75t_SL U48596 ( .A(n67368), .Y(n58134) );
  NAND2xp5_ASAP7_75t_SL U48597 ( .A(n59637), .B(n75925), .Y(n67287) );
  INVx5_ASAP7_75t_SL U48598 ( .A(n75942), .Y(n75899) );
  NAND2xp5_ASAP7_75t_SL U48599 ( .A(n59451), .B(n58727), .Y(n68901) );
  AOI21xp5_ASAP7_75t_SL U48600 ( .A1(n68740), .A2(n58006), .B(n59056), .Y(
        n59451) );
  AOI22xp5_ASAP7_75t_SL U48601 ( .A1(n67854), .A2(n53362), .B1(n53200), .B2(
        n67853), .Y(n57937) );
  NOR2x1_ASAP7_75t_SL U48602 ( .A(n57176), .B(n66424), .Y(n53200) );
  INVx1_ASAP7_75t_SL U48603 ( .A(n53202), .Y(n53201) );
  NOR2x1_ASAP7_75t_SL U48604 ( .A(n66962), .B(n67871), .Y(n53202) );
  NAND2xp5_ASAP7_75t_SL U48605 ( .A(n59300), .B(n67413), .Y(n66924) );
  BUFx5_ASAP7_75t_SL U48606 ( .A(n67974), .Y(n53203) );
  NOR2x1p5_ASAP7_75t_SL U48607 ( .A(n57411), .B(n67162), .Y(n67181) );
  NAND2x1p5_ASAP7_75t_SL U48608 ( .A(n67182), .B(n67181), .Y(n67180) );
  NOR2x1_ASAP7_75t_SL U48609 ( .A(n66722), .B(n66721), .Y(n68480) );
  NAND2xp5_ASAP7_75t_SL U48610 ( .A(n53204), .B(n57985), .Y(n68229) );
  NAND2xp33_ASAP7_75t_SRAM U48611 ( .A(n58452), .B(n59188), .Y(n53204) );
  OAI22x1_ASAP7_75t_SL U48612 ( .A1(n53595), .A2(n67958), .B1(n57165), .B2(
        n68003), .Y(n58170) );
  INVx2_ASAP7_75t_SL U48613 ( .A(n67823), .Y(n67958) );
  XNOR2x1_ASAP7_75t_SL U48614 ( .A(n57179), .B(n59504), .Y(n67823) );
  INVx3_ASAP7_75t_SL U48615 ( .A(n59352), .Y(n67922) );
  BUFx2_ASAP7_75t_SL U48616 ( .A(n67901), .Y(n57501) );
  BUFx5_ASAP7_75t_SL U48617 ( .A(n58336), .Y(n53205) );
  NAND2x1_ASAP7_75t_SL U48618 ( .A(n67702), .B(n57358), .Y(n57300) );
  BUFx5_ASAP7_75t_SL U48619 ( .A(n69148), .Y(n53206) );
  BUFx5_ASAP7_75t_SL U48620 ( .A(n67839), .Y(n53207) );
  INVx1_ASAP7_75t_SL U48621 ( .A(n53208), .Y(n66746) );
  AOI31xp67_ASAP7_75t_SL U48622 ( .A1(n66741), .A2(n66742), .A3(n66966), .B(
        n66965), .Y(n53208) );
  NAND2x1_ASAP7_75t_SL U48623 ( .A(n53209), .B(n57261), .Y(n58949) );
  NAND2x1_ASAP7_75t_SL U48624 ( .A(n66288), .B(n57347), .Y(n53209) );
  XNOR2xp5_ASAP7_75t_SL U48625 ( .A(n53211), .B(n53210), .Y(n58073) );
  XOR2xp5_ASAP7_75t_SL U48626 ( .A(n67668), .B(n67669), .Y(n53210) );
  INVx1_ASAP7_75t_SL U48627 ( .A(n56833), .Y(n53211) );
  NOR2x1_ASAP7_75t_SL U48628 ( .A(n76028), .B(n67712), .Y(n67716) );
  NOR2x1_ASAP7_75t_SL U48629 ( .A(n59012), .B(n64466), .Y(n64343) );
  NOR2x1p5_ASAP7_75t_SL U48630 ( .A(n64077), .B(n64343), .Y(n64340) );
  INVx4_ASAP7_75t_SL U48631 ( .A(n59588), .Y(n59591) );
  XOR2xp5_ASAP7_75t_SL U48632 ( .A(n53213), .B(n53212), .Y(n68288) );
  XNOR2xp5_ASAP7_75t_SL U48633 ( .A(n68151), .B(n68152), .Y(n53212) );
  INVx1_ASAP7_75t_SL U48634 ( .A(n68150), .Y(n53213) );
  NAND2x1p5_ASAP7_75t_SL U48635 ( .A(n57494), .B(n59431), .Y(n59430) );
  XNOR2x1_ASAP7_75t_SL U48636 ( .A(n53214), .B(n63241), .Y(n63685) );
  XNOR2x2_ASAP7_75t_SL U48637 ( .A(n53215), .B(n63608), .Y(n53214) );
  INVx2_ASAP7_75t_SL U48638 ( .A(n63607), .Y(n53215) );
  XOR2xp5_ASAP7_75t_SL U48639 ( .A(n53217), .B(n53216), .Y(n51999) );
  OAI21xp5_ASAP7_75t_SL U48640 ( .A1(n68690), .A2(n58881), .B(n68689), .Y(
        n53216) );
  INVx1_ASAP7_75t_SL U48641 ( .A(n68691), .Y(n53217) );
  NAND2x1p5_ASAP7_75t_SL U48642 ( .A(n58134), .B(n67833), .Y(n58875) );
  XNOR2x1_ASAP7_75t_SL U48643 ( .A(n57468), .B(n64048), .Y(n63830) );
  NOR2x1p5_ASAP7_75t_SL U48644 ( .A(n53249), .B(n53248), .Y(n57468) );
  INVx3_ASAP7_75t_SL U48645 ( .A(n58696), .Y(n66424) );
  NOR2x2_ASAP7_75t_SL U48646 ( .A(n66411), .B(n59458), .Y(n58696) );
  NOR2x1_ASAP7_75t_SL U48647 ( .A(n68259), .B(n68258), .Y(n68305) );
  XOR2xp5_ASAP7_75t_SL U48648 ( .A(n53218), .B(n53339), .Y(n68258) );
  INVx1_ASAP7_75t_SL U48649 ( .A(n68172), .Y(n53218) );
  NAND2x1_ASAP7_75t_SL U48650 ( .A(n57942), .B(n67464), .Y(n57997) );
  INVx8_ASAP7_75t_SL U48651 ( .A(n59458), .Y(n67586) );
  HB1xp67_ASAP7_75t_SL U48652 ( .A(n59506), .Y(n53219) );
  NAND2xp5_ASAP7_75t_SL U48653 ( .A(n58810), .B(n57802), .Y(n58844) );
  BUFx3_ASAP7_75t_SL U48654 ( .A(n64913), .Y(n58393) );
  XOR2x1_ASAP7_75t_SL U48655 ( .A(n58393), .B(n64871), .Y(n64873) );
  XNOR2xp5_ASAP7_75t_SL U48656 ( .A(n63135), .B(n63136), .Y(n57298) );
  NOR2x1_ASAP7_75t_SL U48657 ( .A(n63091), .B(n63092), .Y(n63136) );
  AOI22x1_ASAP7_75t_SL U48658 ( .A1(n66928), .A2(n57161), .B1(n66788), .B2(
        n67306), .Y(n68462) );
  INVx1_ASAP7_75t_SL U48659 ( .A(n53589), .Y(n67798) );
  OR2x2_ASAP7_75t_SL U48660 ( .A(n53590), .B(n53591), .Y(n53589) );
  NAND2x1p5_ASAP7_75t_SL U48661 ( .A(n58989), .B(n53237), .Y(n68081) );
  NAND2xp5_ASAP7_75t_SL U48662 ( .A(n67809), .B(n68081), .Y(n67630) );
  XNOR2xp5_ASAP7_75t_SL U48663 ( .A(n53220), .B(n58847), .Y(n68056) );
  INVx1_ASAP7_75t_SL U48664 ( .A(n67764), .Y(n53220) );
  OAI21xp5_ASAP7_75t_SL U48665 ( .A1(n53275), .A2(n59297), .B(n59189), .Y(
        n58050) );
  BUFx5_ASAP7_75t_SL U48666 ( .A(n75962), .Y(n53221) );
  INVx2_ASAP7_75t_SL U48667 ( .A(n57206), .Y(n57752) );
  NAND2xp5_ASAP7_75t_SL U48668 ( .A(n67930), .B(n53558), .Y(n59219) );
  XOR2xp5_ASAP7_75t_SL U48669 ( .A(n53222), .B(n67892), .Y(n67930) );
  INVx1_ASAP7_75t_SL U48670 ( .A(n67893), .Y(n53222) );
  XOR2x2_ASAP7_75t_SL U48671 ( .A(n68038), .B(n53509), .Y(n57570) );
  XNOR2x1_ASAP7_75t_SL U48672 ( .A(n57571), .B(n57570), .Y(n68143) );
  INVx1_ASAP7_75t_SL U48673 ( .A(n59614), .Y(n53223) );
  INVx1_ASAP7_75t_SL U48674 ( .A(n57321), .Y(n53224) );
  NOR2xp67_ASAP7_75t_SL U48675 ( .A(n57979), .B(n58324), .Y(n57977) );
  INVx2_ASAP7_75t_SL U48676 ( .A(n53517), .Y(n64507) );
  AND2x4_ASAP7_75t_SL U48677 ( .A(n59709), .B(n64507), .Y(n59412) );
  INVx1_ASAP7_75t_SL U48678 ( .A(n64573), .Y(n64574) );
  OAI21xp5_ASAP7_75t_SL U48679 ( .A1(n59618), .A2(n53225), .B(n56362), .Y(
        n64573) );
  INVx1_ASAP7_75t_SL U48680 ( .A(n53226), .Y(n53225) );
  OAI21x1_ASAP7_75t_SL U48681 ( .A1(n67587), .A2(n67588), .B(n57671), .Y(
        n67590) );
  NOR2x1p5_ASAP7_75t_SL U48682 ( .A(n53326), .B(n53325), .Y(n68150) );
  NOR2x1_ASAP7_75t_SL U48683 ( .A(n64466), .B(n58884), .Y(n53348) );
  XNOR2xp5_ASAP7_75t_SL U48684 ( .A(n64629), .B(n53227), .Y(n64943) );
  XOR2xp5_ASAP7_75t_SL U48685 ( .A(n53228), .B(n64962), .Y(n53227) );
  INVx1_ASAP7_75t_SL U48686 ( .A(n58822), .Y(n53228) );
  XNOR2xp5_ASAP7_75t_SL U48687 ( .A(n68283), .B(n68282), .Y(n57400) );
  MAJIxp5_ASAP7_75t_SL U48688 ( .A(n65001), .B(n65002), .C(n65003), .Y(n68282)
         );
  INVx2_ASAP7_75t_SL U48689 ( .A(n64991), .Y(n64982) );
  NAND2xp67_ASAP7_75t_SL U48690 ( .A(n68242), .B(n68241), .Y(n68250) );
  NAND2x1p5_ASAP7_75t_SL U48691 ( .A(n58077), .B(n67496), .Y(n58075) );
  NOR2x2_ASAP7_75t_SL U48692 ( .A(n57056), .B(n58076), .Y(n67496) );
  NOR2x1p5_ASAP7_75t_SL U48693 ( .A(n63884), .B(n63883), .Y(n64749) );
  INVx2_ASAP7_75t_SL U48694 ( .A(n68592), .Y(n69037) );
  NOR3xp33_ASAP7_75t_SL U48695 ( .A(n54023), .B(n64336), .C(n64340), .Y(n54024) );
  INVx1_ASAP7_75t_SL U48696 ( .A(n66817), .Y(n66818) );
  XNOR2x2_ASAP7_75t_SL U48697 ( .A(n58385), .B(n68197), .Y(n68326) );
  HB1xp67_ASAP7_75t_SL U48698 ( .A(n74787), .Y(n53229) );
  INVx1_ASAP7_75t_SL U48699 ( .A(n67950), .Y(n67953) );
  NAND2xp5_ASAP7_75t_SL U48700 ( .A(n58857), .B(n53270), .Y(n67950) );
  BUFx2_ASAP7_75t_SL U48701 ( .A(n59400), .Y(n53230) );
  BUFx5_ASAP7_75t_SL U48702 ( .A(n67401), .Y(n53231) );
  BUFx5_ASAP7_75t_SL U48703 ( .A(n66451), .Y(n53232) );
  BUFx5_ASAP7_75t_SL U48704 ( .A(n64688), .Y(n53233) );
  O2A1O1Ixp5_ASAP7_75t_SL U48705 ( .A1(n62610), .A2(n57119), .B(n58206), .C(
        n58460), .Y(n59357) );
  NOR2x1_ASAP7_75t_SL U48706 ( .A(n53615), .B(n62609), .Y(n62610) );
  INVx3_ASAP7_75t_SL U48707 ( .A(n53234), .Y(n57551) );
  NOR2x1_ASAP7_75t_SL U48708 ( .A(n62624), .B(n59419), .Y(n53234) );
  NOR2x1_ASAP7_75t_SL U48709 ( .A(n59654), .B(n58860), .Y(n62624) );
  NOR4xp75_ASAP7_75t_SL U48710 ( .A(n64618), .B(n57209), .C(n57424), .D(n66240), .Y(n64620) );
  NAND2x2_ASAP7_75t_SL U48711 ( .A(n58765), .B(n58444), .Y(n62557) );
  BUFx6f_ASAP7_75t_SL U48712 ( .A(n67965), .Y(n57182) );
  XNOR2xp5_ASAP7_75t_SL U48713 ( .A(n57934), .B(n53235), .Y(n66908) );
  XOR2xp5_ASAP7_75t_SL U48714 ( .A(n66811), .B(n53498), .Y(n53235) );
  O2A1O1Ixp5_ASAP7_75t_SL U48715 ( .A1(n58960), .A2(n65036), .B(n68123), .C(
        n53236), .Y(n53340) );
  NOR2x1_ASAP7_75t_SL U48716 ( .A(n59012), .B(n58959), .Y(n53236) );
  NAND3x1_ASAP7_75t_SL U48717 ( .A(n58465), .B(n64442), .C(n64443), .Y(n58778)
         );
  INVx2_ASAP7_75t_SL U48718 ( .A(n59510), .Y(n67955) );
  NOR2x1_ASAP7_75t_SL U48719 ( .A(n67585), .B(n67739), .Y(n67587) );
  BUFx5_ASAP7_75t_SL U48720 ( .A(n67416), .Y(n53237) );
  INVx4_ASAP7_75t_SL U48721 ( .A(n67738), .Y(n59242) );
  AND2x2_ASAP7_75t_SL U48722 ( .A(n66453), .B(n66452), .Y(n67383) );
  XNOR2x1_ASAP7_75t_SL U48723 ( .A(n57660), .B(n67991), .Y(n68234) );
  AOI21xp5_ASAP7_75t_SL U48724 ( .A1(n57067), .A2(n67556), .B(n59096), .Y(
        n67492) );
  OAI22xp5_ASAP7_75t_SL U48725 ( .A1(n59155), .A2(n67966), .B1(n59012), .B2(
        n68024), .Y(n68216) );
  NAND2xp5_ASAP7_75t_SL U48726 ( .A(n53238), .B(n56361), .Y(n68024) );
  NAND2xp5_ASAP7_75t_SL U48727 ( .A(n53240), .B(n53239), .Y(n53238) );
  INVx1_ASAP7_75t_SL U48728 ( .A(n53303), .Y(n53239) );
  BUFx5_ASAP7_75t_SL U48729 ( .A(n66411), .Y(n53241) );
  INVx2_ASAP7_75t_SL U48730 ( .A(n62555), .Y(n58766) );
  XOR2xp5_ASAP7_75t_SL U48731 ( .A(n57055), .B(n68050), .Y(n58736) );
  BUFx5_ASAP7_75t_SL U48732 ( .A(n57410), .Y(n53242) );
  OAI21x1_ASAP7_75t_SL U48733 ( .A1(n67308), .A2(n67307), .B(n63063), .Y(
        n75906) );
  NOR2x1p5_ASAP7_75t_SL U48734 ( .A(n53244), .B(n53243), .Y(n67307) );
  INVx3_ASAP7_75t_SL U48735 ( .A(n57347), .Y(n53243) );
  INVx2_ASAP7_75t_SL U48736 ( .A(n59539), .Y(n53244) );
  NAND3xp33_ASAP7_75t_SL U48737 ( .A(n62569), .B(n75477), .C(n59438), .Y(
        n59108) );
  INVx3_ASAP7_75t_SL U48738 ( .A(n59484), .Y(n58775) );
  NAND2xp5_ASAP7_75t_SL U48739 ( .A(n64448), .B(n53245), .Y(n64686) );
  NAND2xp5_ASAP7_75t_SL U48740 ( .A(n64449), .B(n64688), .Y(n53245) );
  INVx4_ASAP7_75t_SL U48741 ( .A(n59300), .Y(n57076) );
  NAND2xp5_ASAP7_75t_SL U48742 ( .A(n53246), .B(n67263), .Y(n67353) );
  OAI21xp5_ASAP7_75t_SL U48743 ( .A1(n57107), .A2(n58871), .B(n53247), .Y(
        n53246) );
  NAND2xp5_ASAP7_75t_SL U48744 ( .A(n57107), .B(n67511), .Y(n53247) );
  NOR2x1_ASAP7_75t_SL U48745 ( .A(n63824), .B(n67315), .Y(n53248) );
  NOR2x1_ASAP7_75t_SL U48746 ( .A(n68383), .B(n64538), .Y(n53249) );
  NAND2xp5_ASAP7_75t_SL U48747 ( .A(n58241), .B(n58240), .Y(n58239) );
  NOR2x1_ASAP7_75t_SL U48748 ( .A(n57574), .B(n60657), .Y(n57573) );
  AND2x4_ASAP7_75t_SL U48749 ( .A(n57572), .B(n57573), .Y(n59166) );
  NAND2x1_ASAP7_75t_SL U48750 ( .A(n67593), .B(n67594), .Y(n67602) );
  BUFx6f_ASAP7_75t_SL U48751 ( .A(n59519), .Y(n57405) );
  NOR2x1p5_ASAP7_75t_SL U48752 ( .A(n57284), .B(n57405), .Y(n57361) );
  BUFx5_ASAP7_75t_SL U48753 ( .A(n2526), .Y(n53250) );
  BUFx6f_ASAP7_75t_SL U48754 ( .A(n1651), .Y(n59533) );
  NAND2x1_ASAP7_75t_SL U48755 ( .A(n62571), .B(n62568), .Y(n59107) );
  BUFx5_ASAP7_75t_SL U48756 ( .A(n59099), .Y(n53251) );
  NAND2xp5_ASAP7_75t_SL U48757 ( .A(n75098), .B(n75099), .Y(n68646) );
  NOR2x1p5_ASAP7_75t_SL U48758 ( .A(n53252), .B(n64747), .Y(n65113) );
  NOR2x1_ASAP7_75t_SL U48759 ( .A(n63881), .B(n63880), .Y(n64747) );
  INVx2_ASAP7_75t_SL U48760 ( .A(n53253), .Y(n53252) );
  AOI21x1_ASAP7_75t_SL U48761 ( .A1(n64749), .A2(n64750), .B(n64748), .Y(
        n53253) );
  INVx1_ASAP7_75t_SL U48762 ( .A(n65016), .Y(n53512) );
  NAND2xp5_ASAP7_75t_SL U48763 ( .A(n53254), .B(n53632), .Y(n65016) );
  NAND2xp5_ASAP7_75t_SL U48764 ( .A(n53256), .B(n53255), .Y(n53254) );
  INVx1_ASAP7_75t_SL U48765 ( .A(n67739), .Y(n53255) );
  INVx4_ASAP7_75t_SL U48766 ( .A(n53298), .Y(n68124) );
  HB1xp67_ASAP7_75t_SL U48767 ( .A(n64989), .Y(n53257) );
  NAND2x1_ASAP7_75t_SL U48768 ( .A(n68286), .B(n68175), .Y(n68207) );
  NAND2x1_ASAP7_75t_SL U48769 ( .A(n68285), .B(n68284), .Y(n68286) );
  INVx2_ASAP7_75t_SL U48770 ( .A(n62958), .Y(n57259) );
  BUFx5_ASAP7_75t_SL U48771 ( .A(n63120), .Y(n53258) );
  NAND3x1_ASAP7_75t_SL U48772 ( .A(n53260), .B(n57465), .C(n53259), .Y(n57782)
         );
  INVx2_ASAP7_75t_SL U48773 ( .A(n66451), .Y(n53259) );
  INVx2_ASAP7_75t_SL U48774 ( .A(n64482), .Y(n53260) );
  BUFx5_ASAP7_75t_SL U48775 ( .A(n75903), .Y(n53261) );
  XOR2xp5_ASAP7_75t_SL U48776 ( .A(n53262), .B(n68044), .Y(n68052) );
  INVx1_ASAP7_75t_SL U48777 ( .A(n68045), .Y(n53262) );
  NAND2x2_ASAP7_75t_SL U48778 ( .A(n58673), .B(n57176), .Y(n59204) );
  INVx2_ASAP7_75t_SL U48779 ( .A(n59204), .Y(n67854) );
  XNOR2xp5_ASAP7_75t_SL U48780 ( .A(n68076), .B(n58811), .Y(n68077) );
  BUFx5_ASAP7_75t_SL U48781 ( .A(n67978), .Y(n53263) );
  XNOR2x1_ASAP7_75t_SL U48782 ( .A(n64690), .B(n64689), .Y(n64691) );
  OAI22xp5_ASAP7_75t_SL U48783 ( .A1(n58457), .A2(n59369), .B1(n59368), .B2(
        n59365), .Y(n58046) );
  NOR2x1_ASAP7_75t_SL U48784 ( .A(n66638), .B(n66639), .Y(n67408) );
  NAND3xp33_ASAP7_75t_SL U48785 ( .A(n64896), .B(n57111), .C(n59517), .Y(
        n64929) );
  OAI21xp5_ASAP7_75t_SL U48786 ( .A1(n57781), .A2(n59456), .B(n53265), .Y(
        n56986) );
  NAND2xp5_ASAP7_75t_SL U48787 ( .A(n59468), .B(n57781), .Y(n53265) );
  NAND2xp5_ASAP7_75t_SL U48788 ( .A(n53266), .B(n61207), .Y(n61208) );
  NOR2x1_ASAP7_75t_SL U48789 ( .A(n60657), .B(n53267), .Y(n53266) );
  NAND2xp5_ASAP7_75t_SL U48790 ( .A(n53268), .B(n58268), .Y(n53267) );
  NOR2x1_ASAP7_75t_SL U48791 ( .A(n75628), .B(n60945), .Y(n53268) );
  BUFx5_ASAP7_75t_SL U48792 ( .A(n59453), .Y(n53269) );
  NAND2xp5_ASAP7_75t_SL U48793 ( .A(n75904), .B(n64897), .Y(n53270) );
  INVx4_ASAP7_75t_SL U48794 ( .A(n59662), .Y(n53275) );
  BUFx5_ASAP7_75t_SL U48795 ( .A(n67922), .Y(n53271) );
  NOR4xp75_ASAP7_75t_SL U48796 ( .A(n59275), .B(n59271), .C(n59273), .D(n57132), .Y(n57713) );
  OR2x2_ASAP7_75t_SL U48797 ( .A(n59195), .B(n68650), .Y(n59275) );
  NAND2xp5_ASAP7_75t_SL U48798 ( .A(n76091), .B(n57179), .Y(n66787) );
  INVx3_ASAP7_75t_SL U48799 ( .A(n65024), .Y(n64899) );
  XNOR2x1_ASAP7_75t_SL U48800 ( .A(n64899), .B(n64898), .Y(n64900) );
  NOR2x1_ASAP7_75t_SL U48801 ( .A(n53273), .B(n53272), .Y(n67588) );
  INVx1_ASAP7_75t_SL U48802 ( .A(n64897), .Y(n53272) );
  INVx1_ASAP7_75t_SL U48803 ( .A(n67585), .Y(n53273) );
  NAND2x1_ASAP7_75t_SL U48804 ( .A(n59531), .B(n57531), .Y(n64036) );
  NAND2x1_ASAP7_75t_SL U48805 ( .A(n64036), .B(n53230), .Y(n57427) );
  BUFx5_ASAP7_75t_SL U48806 ( .A(n59490), .Y(n53274) );
  NOR2x2_ASAP7_75t_SL U48807 ( .A(n57108), .B(n68079), .Y(n59297) );
  INVx2_ASAP7_75t_SL U48808 ( .A(n67264), .Y(n57701) );
  XNOR2x2_ASAP7_75t_SL U48809 ( .A(n62714), .B(n62715), .Y(n62697) );
  NAND2xp5_ASAP7_75t_SL U48810 ( .A(n53277), .B(n53276), .Y(n61206) );
  INVx1_ASAP7_75t_SL U48811 ( .A(n60945), .Y(n53276) );
  NOR2x1_ASAP7_75t_SL U48812 ( .A(n53278), .B(n75628), .Y(n53277) );
  INVx1_ASAP7_75t_SL U48813 ( .A(n59530), .Y(n53278) );
  OAI21xp5_ASAP7_75t_SL U48814 ( .A1(n58402), .A2(n75925), .B(n53279), .Y(
        n64410) );
  NAND2xp5_ASAP7_75t_SL U48815 ( .A(n67288), .B(n59616), .Y(n53279) );
  BUFx5_ASAP7_75t_SL U48816 ( .A(n57175), .Y(n53280) );
  NAND2x1_ASAP7_75t_SL U48817 ( .A(n64663), .B(n64664), .Y(n64089) );
  NAND2x1_ASAP7_75t_SL U48818 ( .A(n64088), .B(n64087), .Y(n64664) );
  INVx6_ASAP7_75t_SL U48819 ( .A(n75642), .Y(n59644) );
  INVx6_ASAP7_75t_SL U48820 ( .A(n59644), .Y(n59640) );
  AOI22x1_ASAP7_75t_SL U48821 ( .A1(n67821), .A2(n67824), .B1(n67842), .B2(
        n68118), .Y(n68108) );
  INVx2_ASAP7_75t_SL U48822 ( .A(n68108), .Y(n57155) );
  BUFx6f_ASAP7_75t_SL U48823 ( .A(n58775), .Y(n57365) );
  NOR2x2_ASAP7_75t_SL U48824 ( .A(n57365), .B(n59643), .Y(n67532) );
  NOR2x1_ASAP7_75t_SL U48825 ( .A(n75284), .B(n75285), .Y(n75279) );
  NOR2x1_ASAP7_75t_SL U48826 ( .A(n75280), .B(n75279), .Y(n75281) );
  NOR2x1_ASAP7_75t_SL U48827 ( .A(n53282), .B(n53281), .Y(n57023) );
  INVx1_ASAP7_75t_SL U48828 ( .A(n59617), .Y(n53281) );
  NOR3xp33_ASAP7_75t_SL U48829 ( .A(n59660), .B(n57348), .C(n59456), .Y(n53282) );
  NAND3x1_ASAP7_75t_SL U48830 ( .A(n64456), .B(n64453), .C(n64452), .Y(n64581)
         );
  NOR2x1_ASAP7_75t_SL U48831 ( .A(n67939), .B(n67938), .Y(n67796) );
  BUFx5_ASAP7_75t_SL U48832 ( .A(n67629), .Y(n53283) );
  NAND2x1_ASAP7_75t_SL U48833 ( .A(n59445), .B(n53508), .Y(n62563) );
  NOR2x1p5_ASAP7_75t_SL U48834 ( .A(n62563), .B(n62564), .Y(n62566) );
  INVx2_ASAP7_75t_SL U48835 ( .A(n67492), .Y(n59232) );
  OAI22x1_ASAP7_75t_SL U48836 ( .A1(n59612), .A2(n64615), .B1(n64616), .B2(
        n59491), .Y(n64964) );
  XNOR2xp5_ASAP7_75t_SL U48837 ( .A(n53284), .B(n68164), .Y(n65055) );
  INVx1_ASAP7_75t_SL U48838 ( .A(n68163), .Y(n53284) );
  NAND2xp5_ASAP7_75t_SL U48839 ( .A(n53286), .B(n53285), .Y(n68163) );
  INVx1_ASAP7_75t_SL U48840 ( .A(n53603), .Y(n53285) );
  NAND2xp5_ASAP7_75t_SL U48841 ( .A(n64607), .B(n53605), .Y(n53286) );
  AND2x4_ASAP7_75t_SL U48842 ( .A(n53506), .B(n64897), .Y(n67434) );
  XOR2xp5_ASAP7_75t_SL U48843 ( .A(n53287), .B(n58233), .Y(n68505) );
  INVx1_ASAP7_75t_SL U48844 ( .A(n66940), .Y(n53287) );
  BUFx5_ASAP7_75t_SL U48845 ( .A(n59665), .Y(n53288) );
  NAND2xp5_ASAP7_75t_SL U48846 ( .A(n75642), .B(n67444), .Y(n59179) );
  INVx1_ASAP7_75t_SL U48847 ( .A(n68079), .Y(n56390) );
  INVx2_ASAP7_75t_SL U48848 ( .A(n68079), .Y(n57164) );
  BUFx5_ASAP7_75t_SL U48849 ( .A(n59448), .Y(n53289) );
  INVxp33_ASAP7_75t_SRAM U48850 ( .A(n59608), .Y(n53342) );
  BUFx5_ASAP7_75t_SL U48851 ( .A(n62562), .Y(n53290) );
  BUFx5_ASAP7_75t_SL U48852 ( .A(n59458), .Y(n53291) );
  AND2x4_ASAP7_75t_SL U48853 ( .A(n58215), .B(n58214), .Y(n61923) );
  INVx5_ASAP7_75t_SL U48854 ( .A(n61923), .Y(n62614) );
  NAND2xp5_ASAP7_75t_SL U48855 ( .A(n53292), .B(n66710), .Y(n66720) );
  NAND2xp5_ASAP7_75t_SL U48856 ( .A(n53294), .B(n53293), .Y(n53292) );
  INVx1_ASAP7_75t_SL U48857 ( .A(n66711), .Y(n53293) );
  INVx1_ASAP7_75t_SL U48858 ( .A(n59515), .Y(n53294) );
  NAND2xp5_ASAP7_75t_SL U48859 ( .A(n59595), .B(n67610), .Y(n62918) );
  XNOR2xp5_ASAP7_75t_SL U48860 ( .A(n53295), .B(n67202), .Y(n58375) );
  MAJIxp5_ASAP7_75t_SL U48861 ( .A(n56952), .B(n67200), .C(n67201), .Y(n67202)
         );
  INVx1_ASAP7_75t_SL U48862 ( .A(n67203), .Y(n53295) );
  HB1xp67_ASAP7_75t_SL U48863 ( .A(n68743), .Y(n53296) );
  XOR2xp5_ASAP7_75t_SL U48864 ( .A(n53297), .B(n68466), .Y(n68467) );
  INVx1_ASAP7_75t_SL U48865 ( .A(n68465), .Y(n53297) );
  NOR2x1_ASAP7_75t_SL U48866 ( .A(n59089), .B(n58895), .Y(n58894) );
  AND2x2_ASAP7_75t_SL U48867 ( .A(n53533), .B(n62571), .Y(n58765) );
  NAND2x1_ASAP7_75t_SL U48868 ( .A(n59655), .B(n64506), .Y(n64648) );
  BUFx5_ASAP7_75t_SL U48869 ( .A(n66625), .Y(n53298) );
  INVx2_ASAP7_75t_SL U48870 ( .A(n64438), .Y(n64444) );
  INVx4_ASAP7_75t_SL U48871 ( .A(n59352), .Y(n57179) );
  NOR2x2_ASAP7_75t_SL U48872 ( .A(n59292), .B(n53299), .Y(n65072) );
  NOR2x1p5_ASAP7_75t_SL U48873 ( .A(n64621), .B(n64622), .Y(n53299) );
  BUFx5_ASAP7_75t_SL U48874 ( .A(n59591), .Y(n53300) );
  A2O1A1Ixp33_ASAP7_75t_SL U48875 ( .A1(n57171), .A2(n67821), .B(n57826), .C(
        n57828), .Y(n67447) );
  NAND3xp33_ASAP7_75t_SL U48876 ( .A(n53302), .B(n57467), .C(n53301), .Y(
        n57684) );
  INVx1_ASAP7_75t_SL U48877 ( .A(n64472), .Y(n53301) );
  INVx1_ASAP7_75t_SL U48878 ( .A(n57150), .Y(n53302) );
  XNOR2xp5_ASAP7_75t_SL U48879 ( .A(n67501), .B(n67502), .Y(n53555) );
  AOI22xp5_ASAP7_75t_SL U48880 ( .A1(n67411), .A2(n59171), .B1(n67381), .B2(
        n58025), .Y(n67502) );
  NAND2x1_ASAP7_75t_SL U48881 ( .A(or1200_cpu_or1200_except_ex_freeze_prev), 
        .B(n76677), .Y(n62572) );
  NOR2x1_ASAP7_75t_SL U48882 ( .A(n57808), .B(n59529), .Y(n57807) );
  XNOR2xp5_ASAP7_75t_SL U48883 ( .A(n66980), .B(n58320), .Y(n58340) );
  XNOR2xp5_ASAP7_75t_SL U48884 ( .A(n66842), .B(n66709), .Y(n66980) );
  BUFx5_ASAP7_75t_SL U48885 ( .A(n57182), .Y(n53303) );
  NAND3x1_ASAP7_75t_SL U48886 ( .A(n59185), .B(n57326), .C(n53304), .Y(n63174)
         );
  INVx1_ASAP7_75t_SL U48887 ( .A(n59182), .Y(n53304) );
  AOI21xp5_ASAP7_75t_SL U48888 ( .A1(n75103), .A2(n58380), .B(n53305), .Y(
        n51986) );
  INVx1_ASAP7_75t_SL U48889 ( .A(n53306), .Y(n53305) );
  OAI21xp5_ASAP7_75t_SL U48890 ( .A1(n57444), .A2(n75095), .B(n75115), .Y(
        n53306) );
  A2O1A1Ixp33_ASAP7_75t_SL U48891 ( .A1(n57366), .A2(n59660), .B(n64563), .C(
        n64562), .Y(n64564) );
  NAND2xp5_ASAP7_75t_SL U48892 ( .A(n53307), .B(n57375), .Y(n64562) );
  NAND2xp5_ASAP7_75t_SL U48893 ( .A(n53309), .B(n53308), .Y(n53307) );
  INVx1_ASAP7_75t_SL U48894 ( .A(n64490), .Y(n53308) );
  NAND2xp5_ASAP7_75t_SL U48895 ( .A(n59505), .B(n75912), .Y(n53309) );
  BUFx5_ASAP7_75t_SL U48896 ( .A(n75958), .Y(n53310) );
  NOR2x1_ASAP7_75t_SL U48897 ( .A(n69119), .B(n68695), .Y(n68701) );
  INVx2_ASAP7_75t_SL U48898 ( .A(n68701), .Y(n58194) );
  BUFx5_ASAP7_75t_SL U48899 ( .A(n59464), .Y(n53311) );
  XNOR2xp5_ASAP7_75t_SL U48900 ( .A(n67590), .B(n57672), .Y(n58787) );
  AOI21x1_ASAP7_75t_SL U48901 ( .A1(n64974), .A2(n53312), .B(n64973), .Y(
        n65001) );
  XNOR2xp5_ASAP7_75t_SL U48902 ( .A(n64972), .B(n64971), .Y(n53312) );
  NAND2xp5_ASAP7_75t_SL U48903 ( .A(n64504), .B(n53313), .Y(n57531) );
  NAND3xp33_ASAP7_75t_SL U48904 ( .A(n57960), .B(n60918), .C(n60917), .Y(
        n53313) );
  INVx3_ASAP7_75t_SL U48905 ( .A(n67585), .Y(n68087) );
  BUFx5_ASAP7_75t_SL U48906 ( .A(n58686), .Y(n53314) );
  INVx4_ASAP7_75t_SL U48907 ( .A(n62614), .Y(n58056) );
  BUFx5_ASAP7_75t_SL U48908 ( .A(n59057), .Y(n53315) );
  NOR2x1p5_ASAP7_75t_SL U48909 ( .A(n61809), .B(n61808), .Y(n61914) );
  NAND3x1_ASAP7_75t_SL U48910 ( .A(n57592), .B(n57593), .C(n59256), .Y(n61808)
         );
  BUFx6f_ASAP7_75t_SL U48911 ( .A(n67906), .Y(n57362) );
  OR2x6_ASAP7_75t_SL U48912 ( .A(n57362), .B(n64040), .Y(n58491) );
  XNOR2x1_ASAP7_75t_SL U48913 ( .A(n58160), .B(n68452), .Y(n58159) );
  BUFx5_ASAP7_75t_SL U48914 ( .A(n76690), .Y(n53316) );
  XNOR2x2_ASAP7_75t_SL U48915 ( .A(n63640), .B(n63212), .Y(n63624) );
  INVx2_ASAP7_75t_SL U48916 ( .A(n63624), .Y(n57479) );
  BUFx5_ASAP7_75t_SL U48917 ( .A(n59507), .Y(n53317) );
  NAND2xp5_ASAP7_75t_SL U48918 ( .A(n57176), .B(n53318), .Y(n67312) );
  INVx1_ASAP7_75t_SL U48919 ( .A(n53319), .Y(n53318) );
  OAI21xp5_ASAP7_75t_SL U48920 ( .A1(n67311), .A2(n67310), .B(n67309), .Y(
        n53319) );
  BUFx5_ASAP7_75t_SL U48921 ( .A(n59611), .Y(n53320) );
  XOR2xp5_ASAP7_75t_SL U48922 ( .A(n58963), .B(n68065), .Y(n57487) );
  O2A1O1Ixp5_ASAP7_75t_SL U48923 ( .A1(n53321), .A2(n57830), .B(n68066), .C(
        n53338), .Y(n59061) );
  INVx1_ASAP7_75t_SL U48924 ( .A(n58963), .Y(n53321) );
  NAND2x2_ASAP7_75t_SL U48925 ( .A(n53323), .B(n53322), .Y(n67489) );
  NAND2x2_ASAP7_75t_SL U48926 ( .A(n67411), .B(n58025), .Y(n53322) );
  NAND2x2_ASAP7_75t_SL U48927 ( .A(n59171), .B(n67477), .Y(n53323) );
  XNOR2x1_ASAP7_75t_SL U48928 ( .A(n67488), .B(n67489), .Y(n57767) );
  INVx1_ASAP7_75t_SL U48929 ( .A(n53324), .Y(n68151) );
  O2A1O1Ixp5_ASAP7_75t_SL U48930 ( .A1(n75962), .A2(n59618), .B(n68092), .C(
        n68091), .Y(n53324) );
  INVx1_ASAP7_75t_SL U48931 ( .A(n68151), .Y(n68149) );
  INVx1_ASAP7_75t_SL U48932 ( .A(n67452), .Y(n62877) );
  AOI211x1_ASAP7_75t_SL U48933 ( .A1(n68098), .A2(n59651), .B(n68095), .C(
        n67452), .Y(n53325) );
  AOI21xp5_ASAP7_75t_SL U48934 ( .A1(n68101), .A2(n58015), .B(n68099), .Y(
        n53326) );
  INVx2_ASAP7_75t_SL U48935 ( .A(n66280), .Y(n75893) );
  INVx8_ASAP7_75t_SL U48936 ( .A(n59518), .Y(n75644) );
  NAND2xp5_ASAP7_75t_SL U48937 ( .A(n59657), .B(n67643), .Y(n67644) );
  NAND2xp5_ASAP7_75t_SL U48938 ( .A(n75894), .B(n75468), .Y(n67643) );
  AND2x2_ASAP7_75t_SL U48939 ( .A(n59518), .B(n66280), .Y(n75468) );
  INVx2_ASAP7_75t_SL U48940 ( .A(n53327), .Y(n67451) );
  NOR2x1p5_ASAP7_75t_SL U48941 ( .A(n59435), .B(n58211), .Y(n53327) );
  NAND2xp5_ASAP7_75t_SL U48942 ( .A(n57104), .B(n53327), .Y(n59409) );
  NOR2xp33_ASAP7_75t_SL U48943 ( .A(n76172), .B(n53328), .Y(n67867) );
  NOR2x1p5_ASAP7_75t_SL U48944 ( .A(n53329), .B(n67451), .Y(n53328) );
  INVx3_ASAP7_75t_SL U48945 ( .A(n68098), .Y(n53329) );
  AOI21xp5_ASAP7_75t_SL U48946 ( .A1(n62679), .A2(n53331), .B(n53330), .Y(
        n62774) );
  O2A1O1Ixp5_ASAP7_75t_SL U48947 ( .A1(n62678), .A2(n59620), .B(n62677), .C(
        n53331), .Y(n53330) );
  INVx1_ASAP7_75t_SL U48948 ( .A(n67451), .Y(n53331) );
  INVx2_ASAP7_75t_SL U48949 ( .A(n53332), .Y(n64366) );
  NOR2x1p5_ASAP7_75t_SL U48950 ( .A(n75438), .B(n67147), .Y(n53332) );
  NAND2x2_ASAP7_75t_SL U48951 ( .A(n56844), .B(n57176), .Y(n67147) );
  NAND2x2_ASAP7_75t_SL U48952 ( .A(n59488), .B(n64367), .Y(n75438) );
  NAND2x2_ASAP7_75t_SL U48953 ( .A(n53333), .B(n64366), .Y(n67464) );
  NAND2x1_ASAP7_75t_SL U48954 ( .A(n67634), .B(n53334), .Y(n53333) );
  INVx2_ASAP7_75t_SL U48955 ( .A(n67634), .Y(n66333) );
  INVx1_ASAP7_75t_SL U48956 ( .A(n57942), .Y(n58743) );
  INVx1_ASAP7_75t_SL U48957 ( .A(n67151), .Y(n53334) );
  NOR2x1_ASAP7_75t_SL U48958 ( .A(n58659), .B(n58660), .Y(n57942) );
  XOR2xp5_ASAP7_75t_SL U48959 ( .A(n53335), .B(n66966), .Y(n66967) );
  OA21x2_ASAP7_75t_SL U48960 ( .A1(n67871), .A2(n59302), .B(n53336), .Y(n66966) );
  INVx1_ASAP7_75t_SL U48961 ( .A(n66965), .Y(n53335) );
  NAND3xp33_ASAP7_75t_SL U48962 ( .A(n53616), .B(n53337), .C(n59299), .Y(
        n53336) );
  INVx1_ASAP7_75t_SL U48963 ( .A(n66729), .Y(n53337) );
  NAND2x1_ASAP7_75t_SL U48964 ( .A(n68150), .B(n57334), .Y(n59285) );
  AOI22x1_ASAP7_75t_SL U48965 ( .A1(n57478), .A2(n64384), .B1(n68086), .B2(
        n64383), .Y(n64439) );
  NOR2x2_ASAP7_75t_SL U48966 ( .A(n58819), .B(n58845), .Y(n57768) );
  NAND2x2_ASAP7_75t_SL U48967 ( .A(n67968), .B(n67967), .Y(n67969) );
  NOR2x1_ASAP7_75t_SL U48968 ( .A(n76077), .B(n57405), .Y(n66620) );
  NOR2x1_ASAP7_75t_SL U48969 ( .A(n59380), .B(n59376), .Y(n59375) );
  INVx1_ASAP7_75t_SL U48970 ( .A(n69007), .Y(n57784) );
  NAND2x1_ASAP7_75t_SL U48971 ( .A(n68730), .B(n57784), .Y(n69030) );
  NAND2xp5_ASAP7_75t_SL U48972 ( .A(n57179), .B(n75906), .Y(n67403) );
  OAI21x1_ASAP7_75t_SL U48973 ( .A1(n68087), .A2(n57179), .B(n67403), .Y(
        n67568) );
  XNOR2x2_ASAP7_75t_SL U48974 ( .A(n57154), .B(n64411), .Y(n64528) );
  NAND2xp5_ASAP7_75t_SL U48975 ( .A(n66758), .B(n57065), .Y(n66724) );
  OAI21x1_ASAP7_75t_SL U48976 ( .A1(n66758), .A2(n66993), .B(n66724), .Y(
        n58124) );
  NOR2x1_ASAP7_75t_SL U48977 ( .A(n57408), .B(n58845), .Y(n67414) );
  XNOR2x1_ASAP7_75t_SL U48978 ( .A(n53263), .B(n57612), .Y(n68160) );
  AOI21xp5_ASAP7_75t_SL U48979 ( .A1(n67902), .A2(n59662), .B(n67370), .Y(
        n67371) );
  OAI22x1_ASAP7_75t_SL U48980 ( .A1(n59067), .A2(n67369), .B1(n67368), .B2(
        n57253), .Y(n67373) );
  NAND2x1_ASAP7_75t_SL U48981 ( .A(n57402), .B(n59517), .Y(n67863) );
  INVx2_ASAP7_75t_SL U48982 ( .A(n67863), .Y(n57904) );
  XNOR2x2_ASAP7_75t_SL U48983 ( .A(n68179), .B(n58741), .Y(n68205) );
  INVx2_ASAP7_75t_SL U48984 ( .A(n68205), .Y(n68206) );
  BUFx6f_ASAP7_75t_SL U48985 ( .A(n59517), .Y(n57292) );
  AO21x2_ASAP7_75t_SL U48986 ( .A1(n57292), .A2(n75900), .B(n57510), .Y(n66933) );
  NAND2x2_ASAP7_75t_SL U48987 ( .A(n58505), .B(n67829), .Y(n58645) );
  INVx2_ASAP7_75t_SL U48988 ( .A(n58645), .Y(n58644) );
  NAND2xp5_ASAP7_75t_SL U48989 ( .A(n67845), .B(n57417), .Y(n63121) );
  NAND2x1p5_ASAP7_75t_SL U48990 ( .A(n68538), .B(n68537), .Y(n68955) );
  BUFx6f_ASAP7_75t_SL U48991 ( .A(n59454), .Y(n57165) );
  NAND2x2_ASAP7_75t_SL U48992 ( .A(n67947), .B(n66805), .Y(n67901) );
  XNOR2x1_ASAP7_75t_SL U48993 ( .A(n66606), .B(n66605), .Y(n68621) );
  NOR2x1p5_ASAP7_75t_SL U48994 ( .A(n68622), .B(n68621), .Y(n66607) );
  OAI21xp5_ASAP7_75t_SL U48995 ( .A1(n53207), .A2(n67704), .B(n67703), .Y(
        n67707) );
  AOI21x1_ASAP7_75t_SL U48996 ( .A1(n68722), .A2(n68723), .B(n68724), .Y(
        n58730) );
  BUFx6f_ASAP7_75t_SL U48997 ( .A(or1200_cpu_alu_op_2_), .Y(n59566) );
  NOR2x1p5_ASAP7_75t_SL U48998 ( .A(n59566), .B(n62561), .Y(n62554) );
  INVx2_ASAP7_75t_SL U48999 ( .A(n65002), .Y(n64975) );
  AOI21x1_ASAP7_75t_SL U49000 ( .A1(n68131), .A2(n57224), .B(n68130), .Y(
        n57289) );
  NOR2x1_ASAP7_75t_SL U49001 ( .A(n67884), .B(n56953), .Y(n57785) );
  XNOR2x2_ASAP7_75t_SL U49002 ( .A(n58722), .B(n58721), .Y(n58723) );
  OAI21x1_ASAP7_75t_SL U49003 ( .A1(n58483), .A2(n63082), .B(n68079), .Y(
        n58989) );
  NOR2xp67_ASAP7_75t_SL U49004 ( .A(n53338), .B(n67887), .Y(n67943) );
  NOR2x1_ASAP7_75t_SL U49005 ( .A(n68065), .B(n58963), .Y(n53338) );
  XOR2xp5_ASAP7_75t_SL U49006 ( .A(n68171), .B(n68170), .Y(n53339) );
  OAI22xp5_ASAP7_75t_SL U49007 ( .A1(n65041), .A2(n67627), .B1(n59612), .B2(
        n67946), .Y(n68172) );
  XNOR2xp5_ASAP7_75t_SL U49008 ( .A(n65038), .B(n65039), .Y(n68259) );
  XNOR2xp5_ASAP7_75t_SL U49009 ( .A(n65037), .B(n53340), .Y(n65039) );
  NAND2xp67_ASAP7_75t_SL U49010 ( .A(n53343), .B(n59357), .Y(n58719) );
  INVx1_ASAP7_75t_SL U49011 ( .A(n59483), .Y(n53343) );
  NAND2x2_ASAP7_75t_SL U49012 ( .A(n57636), .B(n53341), .Y(n57638) );
  INVx3_ASAP7_75t_SL U49013 ( .A(n59483), .Y(n53341) );
  NAND2xp5_ASAP7_75t_SL U49014 ( .A(n59483), .B(n57181), .Y(n56999) );
  OAI21xp5_ASAP7_75t_SL U49015 ( .A1(n59508), .A2(n53343), .B(n57638), .Y(
        n58197) );
  INVx2_ASAP7_75t_SL U49016 ( .A(n59067), .Y(n68414) );
  INVx1_ASAP7_75t_SL U49017 ( .A(n57253), .Y(n56967) );
  INVx1_ASAP7_75t_SL U49018 ( .A(n64582), .Y(n64457) );
  OAI21xp5_ASAP7_75t_SL U49019 ( .A1(n64455), .A2(n64456), .B(n64454), .Y(
        n64582) );
  NOR2x1_ASAP7_75t_SL U49020 ( .A(n53346), .B(n53344), .Y(n64454) );
  NOR2x1_ASAP7_75t_SL U49021 ( .A(n53345), .B(n57253), .Y(n53344) );
  INVx1_ASAP7_75t_SL U49022 ( .A(n64616), .Y(n53345) );
  NOR2xp33_ASAP7_75t_SL U49023 ( .A(n53347), .B(n59067), .Y(n53346) );
  INVx1_ASAP7_75t_SL U49024 ( .A(n64498), .Y(n53347) );
  NOR2x1_ASAP7_75t_SL U49025 ( .A(n64451), .B(n64450), .Y(n64455) );
  NOR2x1_ASAP7_75t_SL U49026 ( .A(n64445), .B(n67434), .Y(n64451) );
  NOR2x1_ASAP7_75t_SL U49027 ( .A(n53348), .B(n64447), .Y(n64456) );
  INVx1_ASAP7_75t_SL U49028 ( .A(n67885), .Y(n53349) );
  XNOR2x1_ASAP7_75t_SL U49029 ( .A(n53349), .B(n57862), .Y(n57627) );
  XNOR2xp5_ASAP7_75t_SL U49030 ( .A(n68191), .B(n57627), .Y(n68192) );
  NOR2x1_ASAP7_75t_SL U49031 ( .A(n57521), .B(n57520), .Y(n68264) );
  INVx1_ASAP7_75t_SL U49032 ( .A(n68201), .Y(n68212) );
  OAI211xp5_ASAP7_75t_SL U49033 ( .A1(n57520), .A2(n53351), .B(n53353), .C(
        n53350), .Y(n68201) );
  AO21x1_ASAP7_75t_SL U49034 ( .A1(n58891), .A2(n57438), .B(n68266), .Y(n53350) );
  NAND2xp5_ASAP7_75t_SL U49035 ( .A(n53352), .B(n58890), .Y(n53351) );
  INVx1_ASAP7_75t_SL U49036 ( .A(n57521), .Y(n53352) );
  NAND3xp33_ASAP7_75t_SL U49037 ( .A(n68128), .B(n68127), .C(n68126), .Y(
        n53353) );
  NAND3xp33_ASAP7_75t_SL U49038 ( .A(n53356), .B(n59249), .C(n53354), .Y(
        n52001) );
  NAND2xp5_ASAP7_75t_SL U49039 ( .A(n53355), .B(n58839), .Y(n53354) );
  INVx1_ASAP7_75t_SL U49040 ( .A(n58533), .Y(n53355) );
  NAND2xp5_ASAP7_75t_SL U49041 ( .A(n58450), .B(n53357), .Y(n53356) );
  INVx1_ASAP7_75t_SL U49042 ( .A(n58839), .Y(n53357) );
  NAND2x1_ASAP7_75t_SL U49043 ( .A(n67209), .B(n53386), .Y(n68673) );
  NOR2x1p5_ASAP7_75t_SL U49044 ( .A(n68648), .B(n58448), .Y(n53386) );
  NAND2x1_ASAP7_75t_SL U49045 ( .A(n59309), .B(n58894), .Y(n67209) );
  NOR2x1_ASAP7_75t_SL U49046 ( .A(n69295), .B(n69296), .Y(n68657) );
  A2O1A1Ixp33_ASAP7_75t_SL U49047 ( .A1(n68673), .A2(n68674), .B(n68653), .C(
        n53358), .Y(n69296) );
  NAND4xp25_ASAP7_75t_SL U49048 ( .A(n53361), .B(n58958), .C(n53359), .D(
        n68699), .Y(n53358) );
  NOR2x1_ASAP7_75t_SL U49049 ( .A(n69119), .B(n69038), .Y(n68699) );
  NOR2x1_ASAP7_75t_SL U49050 ( .A(n68648), .B(n53360), .Y(n53359) );
  INVx1_ASAP7_75t_SL U49051 ( .A(n68700), .Y(n53360) );
  INVx1_ASAP7_75t_SL U49052 ( .A(n58957), .Y(n53361) );
  OAI21x1_ASAP7_75t_SL U49053 ( .A1(n59596), .A2(n57169), .B(n53362), .Y(
        n59469) );
  INVx2_ASAP7_75t_SL U49054 ( .A(n57240), .Y(n53362) );
  NAND2x1_ASAP7_75t_SL U49055 ( .A(n64429), .B(n56836), .Y(n64462) );
  INVx1_ASAP7_75t_SL U49056 ( .A(n53363), .Y(n58341) );
  INVx1_ASAP7_75t_SL U49057 ( .A(n64590), .Y(n57143) );
  NAND2xp5_ASAP7_75t_SL U49058 ( .A(n53364), .B(n64460), .Y(n64590) );
  INVx1_ASAP7_75t_SL U49059 ( .A(n53368), .Y(n53364) );
  XNOR2x1_ASAP7_75t_SL U49060 ( .A(n53365), .B(n58341), .Y(n64689) );
  NOR2x1_ASAP7_75t_SL U49061 ( .A(n64458), .B(n64457), .Y(n53363) );
  XNOR2xp5_ASAP7_75t_SL U49062 ( .A(n57143), .B(n64587), .Y(n53365) );
  MAJIxp5_ASAP7_75t_SL U49063 ( .A(n64462), .B(n64464), .C(n64463), .Y(n64587)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U49064 ( .A1(n55485), .A2(n64427), .B(n64426), .C(
        n55486), .Y(n64463) );
  OAI21xp5_ASAP7_75t_SL U49065 ( .A1(n53366), .A2(n64423), .B(n64422), .Y(
        n64464) );
  INVx1_ASAP7_75t_SL U49066 ( .A(n53367), .Y(n53366) );
  NAND2xp5_ASAP7_75t_SL U49067 ( .A(n67911), .B(n64424), .Y(n53367) );
  NOR2x1_ASAP7_75t_SL U49068 ( .A(n64461), .B(n67974), .Y(n53368) );
  AOI21x1_ASAP7_75t_SL U49069 ( .A1(n53197), .A2(n53369), .B(n67482), .Y(
        n67684) );
  AOI21xp5_ASAP7_75t_SL U49070 ( .A1(n58755), .A2(n53369), .B(n67737), .Y(
        n68374) );
  NAND2x2_ASAP7_75t_SL U49071 ( .A(n53370), .B(n67479), .Y(n53369) );
  INVx2_ASAP7_75t_SL U49072 ( .A(n53371), .Y(n53370) );
  NOR2x1_ASAP7_75t_SL U49073 ( .A(n53303), .B(n59651), .Y(n53371) );
  NOR2x1_ASAP7_75t_SL U49074 ( .A(n62617), .B(n53372), .Y(n62619) );
  NOR2x1_ASAP7_75t_SL U49075 ( .A(n77278), .B(n53372), .Y(n62618) );
  NOR2x1_ASAP7_75t_SL U49076 ( .A(n59471), .B(n62616), .Y(n53372) );
  INVx1_ASAP7_75t_SL U49077 ( .A(n53373), .Y(n57571) );
  XNOR2xp5_ASAP7_75t_SL U49078 ( .A(n67770), .B(n67769), .Y(n53373) );
  MAJIxp5_ASAP7_75t_SL U49079 ( .A(n53373), .B(n53509), .C(n68038), .Y(n68041)
         );
  OAI22xp5_ASAP7_75t_SL U49080 ( .A1(n56958), .A2(n56957), .B1(n57099), .B2(
        n67390), .Y(n67504) );
  INVx1_ASAP7_75t_SL U49081 ( .A(n67399), .Y(n57094) );
  XNOR2xp5_ASAP7_75t_SL U49082 ( .A(n53556), .B(n53374), .Y(n67399) );
  XOR2xp5_ASAP7_75t_SL U49083 ( .A(n67505), .B(n67504), .Y(n53374) );
  NOR2x2_ASAP7_75t_SL U49084 ( .A(n57174), .B(n53375), .Y(n67845) );
  INVx3_ASAP7_75t_SL U49085 ( .A(n59200), .Y(n53375) );
  OAI21xp5_ASAP7_75t_SL U49086 ( .A1(n53375), .A2(n59616), .B(n67227), .Y(
        n63098) );
  AOI21xp5_ASAP7_75t_SL U49087 ( .A1(n53382), .A2(n57983), .B(n53376), .Y(
        n52006) );
  INVx1_ASAP7_75t_SL U49088 ( .A(n53377), .Y(n53376) );
  OAI21xp5_ASAP7_75t_SL U49089 ( .A1(n68716), .A2(n53381), .B(n68715), .Y(
        n53377) );
  NAND2xp5_ASAP7_75t_SL U49090 ( .A(n53379), .B(n53378), .Y(n57983) );
  INVx1_ASAP7_75t_SL U49091 ( .A(n53474), .Y(n53378) );
  NOR2x1_ASAP7_75t_SL U49092 ( .A(n53380), .B(n75109), .Y(n53379) );
  INVx1_ASAP7_75t_SL U49093 ( .A(n68714), .Y(n53380) );
  NOR2x1p5_ASAP7_75t_SL U49094 ( .A(n75109), .B(n53474), .Y(n53381) );
  NAND2xp5_ASAP7_75t_SL U49095 ( .A(n57982), .B(n53381), .Y(n57981) );
  NAND2xp5_ASAP7_75t_SL U49096 ( .A(n58769), .B(n53381), .Y(n58768) );
  AOI21xp5_ASAP7_75t_SL U49097 ( .A1(n53381), .A2(n75470), .B(n75090), .Y(
        n75094) );
  AOI21xp5_ASAP7_75t_SL U49098 ( .A1(n75282), .A2(n53381), .B(n75281), .Y(
        n75289) );
  INVx1_ASAP7_75t_SL U49099 ( .A(n68713), .Y(n53382) );
  NAND2xp5_ASAP7_75t_SL U49100 ( .A(n53383), .B(n69147), .Y(n59089) );
  NAND2xp5_ASAP7_75t_SL U49101 ( .A(n69141), .B(n67106), .Y(n53383) );
  INVxp33_ASAP7_75t_SL U49102 ( .A(n53383), .Y(n68697) );
  OR2x2_ASAP7_75t_SL U49103 ( .A(n53384), .B(n68697), .Y(n69149) );
  INVx1_ASAP7_75t_SL U49104 ( .A(n69143), .Y(n53384) );
  AND2x2_ASAP7_75t_SL U49105 ( .A(n53383), .B(n68695), .Y(n58448) );
  XNOR2xp5_ASAP7_75t_SL U49106 ( .A(n66946), .B(n66945), .Y(n66948) );
  XNOR2xp5_ASAP7_75t_SL U49107 ( .A(n66737), .B(n53385), .Y(n66946) );
  XNOR2xp5_ASAP7_75t_SL U49108 ( .A(n66738), .B(n66739), .Y(n53385) );
  AOI21xp5_ASAP7_75t_SL U49109 ( .A1(n57360), .A2(n59515), .B(n59238), .Y(
        n66737) );
  OAI21xp5_ASAP7_75t_SL U49110 ( .A1(n59391), .A2(n67209), .B(n53386), .Y(
        n59390) );
  NOR2x1p5_ASAP7_75t_SL U49111 ( .A(n58731), .B(n53387), .Y(n68724) );
  NOR2x1p5_ASAP7_75t_SL U49112 ( .A(n57870), .B(n57869), .Y(n53387) );
  INVx1_ASAP7_75t_SL U49113 ( .A(n53387), .Y(n68734) );
  NOR2x1_ASAP7_75t_SL U49114 ( .A(n53388), .B(n68734), .Y(n68559) );
  INVx1_ASAP7_75t_SL U49115 ( .A(n68735), .Y(n53388) );
  AOI21xp5_ASAP7_75t_SL U49116 ( .A1(n68750), .A2(n53387), .B(n68749), .Y(
        n68751) );
  OAI21xp33_ASAP7_75t_SL U49117 ( .A1(n68245), .A2(n68244), .B(n53389), .Y(
        n68141) );
  INVx1_ASAP7_75t_SL U49118 ( .A(n68246), .Y(n53389) );
  AND2x2_ASAP7_75t_SL U49119 ( .A(n58943), .B(n57894), .Y(n68246) );
  NOR2x1_ASAP7_75t_SL U49120 ( .A(n67084), .B(n53390), .Y(n63154) );
  NOR2xp33_ASAP7_75t_SL U49121 ( .A(n53390), .B(n63090), .Y(n63092) );
  XNOR2xp5_ASAP7_75t_SL U49122 ( .A(n53390), .B(n62764), .Y(n62765) );
  NOR2x1p5_ASAP7_75t_SL U49123 ( .A(n53392), .B(n53391), .Y(n53390) );
  INVx2_ASAP7_75t_SL U49124 ( .A(n57380), .Y(n53391) );
  INVx3_ASAP7_75t_SL U49125 ( .A(n59656), .Y(n53392) );
  NOR2xp67_ASAP7_75t_SL U49126 ( .A(n53397), .B(n53393), .Y(n66845) );
  NAND2x1_ASAP7_75t_SL U49127 ( .A(n66661), .B(n66662), .Y(n53393) );
  AOI21x1_ASAP7_75t_SL U49128 ( .A1(n56967), .A2(n66827), .B(n53394), .Y(
        n66662) );
  AOI21xp33_ASAP7_75t_SL U49129 ( .A1(n66657), .A2(n57104), .B(n53395), .Y(
        n53394) );
  NAND2x1_ASAP7_75t_SL U49130 ( .A(n53396), .B(n66658), .Y(n53395) );
  INVx2_ASAP7_75t_SL U49131 ( .A(n66656), .Y(n53396) );
  NAND2x1_ASAP7_75t_SL U49132 ( .A(n66655), .B(n53398), .Y(n66661) );
  NOR2x1p5_ASAP7_75t_SL U49133 ( .A(n66659), .B(n66660), .Y(n53397) );
  INVx2_ASAP7_75t_SL U49134 ( .A(n66654), .Y(n66660) );
  OAI22x1_ASAP7_75t_SL U49135 ( .A1(n66651), .A2(n58903), .B1(n67442), .B2(
        n66682), .Y(n66654) );
  NOR2x1p5_ASAP7_75t_SL U49136 ( .A(n66655), .B(n53398), .Y(n66659) );
  OAI22x1_ASAP7_75t_SL U49137 ( .A1(n64920), .A2(n59238), .B1(n66711), .B2(
        n59460), .Y(n53398) );
  OAI21x1_ASAP7_75t_SL U49138 ( .A1(n66767), .A2(n57410), .B(n57594), .Y(
        n66655) );
  NAND2xp33_ASAP7_75t_SL U49139 ( .A(n53399), .B(n53402), .Y(n53401) );
  NAND2x1_ASAP7_75t_SL U49140 ( .A(n68572), .B(n68573), .Y(n53399) );
  INVxp33_ASAP7_75t_SL U49141 ( .A(n53399), .Y(n68719) );
  NOR2x1_ASAP7_75t_SL U49142 ( .A(n53401), .B(n53400), .Y(n68913) );
  INVx1_ASAP7_75t_SL U49143 ( .A(n68909), .Y(n53400) );
  INVx1_ASAP7_75t_SL U49144 ( .A(n68961), .Y(n53402) );
  INVx1_ASAP7_75t_SL U49145 ( .A(n67739), .Y(n53403) );
  NAND2xp5_ASAP7_75t_SL U49146 ( .A(n75942), .B(n53403), .Y(n58041) );
  NOR2x1p5_ASAP7_75t_SL U49147 ( .A(n59455), .B(n63826), .Y(n67739) );
  OR2x2_ASAP7_75t_SL U49148 ( .A(n67604), .B(n67605), .Y(n75942) );
  XNOR2xp5_ASAP7_75t_SL U49149 ( .A(n68273), .B(n68272), .Y(n68274) );
  XNOR2xp5_ASAP7_75t_SL U49150 ( .A(n68215), .B(n53404), .Y(n68272) );
  XNOR2xp5_ASAP7_75t_SL U49151 ( .A(n57145), .B(n57329), .Y(n53404) );
  NOR2x1_ASAP7_75t_SL U49152 ( .A(n53406), .B(n68977), .Y(n68979) );
  O2A1O1Ixp5_ASAP7_75t_SL U49153 ( .A1(n68976), .A2(n53406), .B(n53405), .C(
        n53527), .Y(n53526) );
  NAND2xp5_ASAP7_75t_SL U49154 ( .A(n68967), .B(n53406), .Y(n53405) );
  OAI21xp5_ASAP7_75t_SL U49155 ( .A1(n68965), .A2(n68964), .B(n68963), .Y(
        n53406) );
  OAI21xp33_ASAP7_75t_SL U49156 ( .A1(n53621), .A2(n68733), .B(n53407), .Y(
        n51998) );
  AOI21xp33_ASAP7_75t_SL U49157 ( .A1(n53621), .A2(n56858), .B(n53408), .Y(
        n53407) );
  INVxp67_ASAP7_75t_SL U49158 ( .A(n53409), .Y(n53408) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U49159 ( .A1(n69030), .A2(n53411), .B(n68732), 
        .C(n53410), .Y(n53409) );
  NAND3x1_ASAP7_75t_SL U49160 ( .A(n69030), .B(n68732), .C(n69029), .Y(n53410)
         );
  INVxp67_ASAP7_75t_SL U49161 ( .A(n53412), .Y(n53411) );
  NAND2xp67_ASAP7_75t_SL U49162 ( .A(n69029), .B(n69032), .Y(n53412) );
  NOR2x1p5_ASAP7_75t_SL U49163 ( .A(n69003), .B(n53413), .Y(n53621) );
  NAND2x1_ASAP7_75t_SL U49164 ( .A(n53414), .B(n59425), .Y(n53413) );
  NAND2x1_ASAP7_75t_SL U49165 ( .A(n68725), .B(n59426), .Y(n59425) );
  O2A1O1Ixp33_ASAP7_75t_SL U49166 ( .A1(n68719), .A2(n68869), .B(n58371), .C(
        n57475), .Y(n53414) );
  NOR2x1p5_ASAP7_75t_SL U49167 ( .A(n68834), .B(n53415), .Y(n69003) );
  NAND2x1_ASAP7_75t_SL U49168 ( .A(n68974), .B(n68725), .Y(n53415) );
  NOR2x1p5_ASAP7_75t_SL U49169 ( .A(n68728), .B(n53547), .Y(n68834) );
  XOR2xp5_ASAP7_75t_SL U49170 ( .A(n66823), .B(n66824), .Y(n66769) );
  NOR2x1_ASAP7_75t_SL U49171 ( .A(n53417), .B(n53416), .Y(n66824) );
  NOR2x1_ASAP7_75t_SL U49172 ( .A(n66767), .B(n67434), .Y(n53416) );
  NOR2x1_ASAP7_75t_SL U49173 ( .A(n66768), .B(n57410), .Y(n53417) );
  OAI21xp33_ASAP7_75t_SL U49174 ( .A1(n53420), .A2(n53418), .B(n64712), .Y(
        n57497) );
  NOR3x1_ASAP7_75t_SL U49175 ( .A(n64709), .B(n53419), .C(n64710), .Y(n53418)
         );
  INVx2_ASAP7_75t_SL U49176 ( .A(n64718), .Y(n53419) );
  NAND2x2_ASAP7_75t_SL U49177 ( .A(n64047), .B(n58470), .Y(n64709) );
  A2O1A1Ixp33_ASAP7_75t_SL U49178 ( .A1(n59364), .A2(n64047), .B(n64718), .C(
        n64721), .Y(n53420) );
  XOR2x1_ASAP7_75t_SL U49179 ( .A(n64682), .B(n53421), .Y(n64718) );
  INVx2_ASAP7_75t_SL U49180 ( .A(n64683), .Y(n53421) );
  INVx2_ASAP7_75t_SL U49181 ( .A(n64717), .Y(n64047) );
  INVx1_ASAP7_75t_SL U49182 ( .A(n66980), .Y(n67039) );
  INVxp67_ASAP7_75t_SL U49183 ( .A(n69097), .Y(n67044) );
  NAND2xp5_ASAP7_75t_SL U49184 ( .A(n69096), .B(n69097), .Y(n69095) );
  XNOR2x1_ASAP7_75t_SL U49185 ( .A(n53423), .B(n53422), .Y(n69097) );
  XNOR2x1_ASAP7_75t_SL U49186 ( .A(n66983), .B(n66904), .Y(n53422) );
  XNOR2x1_ASAP7_75t_SL U49187 ( .A(n66982), .B(n66903), .Y(n53423) );
  AND2x2_ASAP7_75t_SL U49188 ( .A(n53424), .B(n67043), .Y(n69096) );
  OAI21xp5_ASAP7_75t_SL U49189 ( .A1(n66980), .A2(n66981), .B(n57052), .Y(
        n67043) );
  NAND2xp5_ASAP7_75t_SL U49190 ( .A(n53425), .B(n66980), .Y(n53424) );
  AOI21xp5_ASAP7_75t_SL U49191 ( .A1(n67041), .A2(n67042), .B(n67040), .Y(
        n53425) );
  OR2x2_ASAP7_75t_SL U49192 ( .A(n53427), .B(n68623), .Y(n68684) );
  NOR2x1_ASAP7_75t_SL U49193 ( .A(n66533), .B(n53426), .Y(n68623) );
  NOR2x1_ASAP7_75t_SL U49194 ( .A(n66532), .B(n66531), .Y(n53426) );
  NOR2x1_ASAP7_75t_SL U49195 ( .A(n66529), .B(n66530), .Y(n66533) );
  INVx1_ASAP7_75t_SL U49196 ( .A(n66534), .Y(n53427) );
  BUFx2_ASAP7_75t_SL U49197 ( .A(n58415), .Y(n53428) );
  INVx5_ASAP7_75t_SL U49198 ( .A(n58415), .Y(n57137) );
  NOR2x1_ASAP7_75t_SL U49199 ( .A(n63753), .B(n76577), .Y(n76589) );
  INVx8_ASAP7_75t_SL U49200 ( .A(n72516), .Y(n57125) );
  AND2x4_ASAP7_75t_SL U49201 ( .A(n59527), .B(n72367), .Y(n72516) );
  NAND2x1p5_ASAP7_75t_SL U49202 ( .A(n74162), .B(n76971), .Y(n77171) );
  INVx3_ASAP7_75t_SL U49203 ( .A(n77171), .Y(n77194) );
  INVx4_ASAP7_75t_SL U49204 ( .A(n77139), .Y(n74899) );
  NAND2x1p5_ASAP7_75t_SL U49205 ( .A(n58821), .B(n58820), .Y(n77139) );
  NOR2x1_ASAP7_75t_SL U49206 ( .A(n70761), .B(n70760), .Y(n70764) );
  INVx1_ASAP7_75t_SL U49207 ( .A(n70764), .Y(n70762) );
  O2A1O1Ixp5_ASAP7_75t_SL U49208 ( .A1(n70796), .A2(n70785), .B(n70795), .C(
        n70797), .Y(n55563) );
  NOR2x1_ASAP7_75t_SL U49209 ( .A(n70763), .B(n70762), .Y(n70796) );
  BUFx2_ASAP7_75t_SL U49210 ( .A(n60630), .Y(n53429) );
  NOR2x1_ASAP7_75t_SL U49211 ( .A(n53429), .B(n78182), .Y(n53430) );
  NOR2x1p5_ASAP7_75t_SL U49212 ( .A(n74025), .B(n76427), .Y(n78182) );
  HB1xp67_ASAP7_75t_SL U49213 ( .A(n65179), .Y(n53431) );
  AOI31xp33_ASAP7_75t_SL U49214 ( .A1(n68937), .A2(n68936), .A3(n68935), .B(
        n68934), .Y(n53432) );
  NOR2x1_ASAP7_75t_SL U49215 ( .A(n76663), .B(n62154), .Y(n77163) );
  NAND2x1p5_ASAP7_75t_SL U49216 ( .A(n22057), .B(n60330), .Y(n77954) );
  OAI22xp33_ASAP7_75t_SRAM U49217 ( .A1(or1200_cpu_or1200_except_n176), .A2(
        n57070), .B1(n77597), .B2(n77294), .Y(n76207) );
  OAI22xp33_ASAP7_75t_SRAM U49218 ( .A1(or1200_cpu_or1200_except_n168), .A2(
        n57070), .B1(n76508), .B2(n77294), .Y(n76246) );
  OAI22xp33_ASAP7_75t_SRAM U49219 ( .A1(or1200_cpu_or1200_except_n144), .A2(
        n57070), .B1(n75431), .B2(n77294), .Y(n75432) );
  OAI22xp33_ASAP7_75t_SRAM U49220 ( .A1(or1200_cpu_or1200_except_n152), .A2(
        n57070), .B1(n75302), .B2(n77294), .Y(n75303) );
  OAI22xp33_ASAP7_75t_SRAM U49221 ( .A1(or1200_cpu_or1200_except_n150), .A2(
        n57070), .B1(n74984), .B2(n77294), .Y(n74985) );
  OAI22xp33_ASAP7_75t_SRAM U49222 ( .A1(or1200_cpu_or1200_except_n140), .A2(
        n57070), .B1(n75620), .B2(n77294), .Y(n75621) );
  OAI22xp33_ASAP7_75t_SRAM U49223 ( .A1(or1200_cpu_or1200_except_n148), .A2(
        n57070), .B1(n74639), .B2(n77294), .Y(n74577) );
  NAND2x1p5_ASAP7_75t_SL U49224 ( .A(n59020), .B(n58407), .Y(n59361) );
  NAND2xp5_ASAP7_75t_SL U49225 ( .A(n62596), .B(n59020), .Y(n62805) );
  XNOR2x1_ASAP7_75t_SL U49226 ( .A(n70742), .B(n70743), .Y(n70753) );
  OAI21xp5_ASAP7_75t_SL U49227 ( .A1(n70800), .A2(n70799), .B(n70798), .Y(
        n70801) );
  OAI22xp5_ASAP7_75t_SL U49228 ( .A1(n53991), .A2(n53433), .B1(
        or1200_cpu_or1200_mult_mac_n40), .B2(n56274), .Y(
        or1200_cpu_or1200_mult_mac_n1515) );
  XNOR2xp5_ASAP7_75t_SL U49229 ( .A(or1200_cpu_or1200_mult_mac_n42), .B(n76056), .Y(n53433) );
  INVx1_ASAP7_75t_SL U49230 ( .A(n58600), .Y(n56274) );
  NOR2x1_ASAP7_75t_SL U49231 ( .A(n70090), .B(n70089), .Y(n70094) );
  OAI21x1_ASAP7_75t_SL U49232 ( .A1(n69791), .A2(n69790), .B(n69789), .Y(
        n69801) );
  NOR2x1_ASAP7_75t_SL U49233 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[25]), .B(n73519), .Y(
        n73874) );
  NOR2x1_ASAP7_75t_SL U49234 ( .A(n73575), .B(n73574), .Y(n73658) );
  NOR2x1p5_ASAP7_75t_SL U49235 ( .A(n76941), .B(n74887), .Y(n76963) );
  NOR2x1_ASAP7_75t_SL U49236 ( .A(n76945), .B(n74871), .Y(n76933) );
  INVx1_ASAP7_75t_SL U49237 ( .A(n74871), .Y(n76970) );
  NAND2x1p5_ASAP7_75t_SL U49238 ( .A(n76965), .B(n76934), .Y(n74871) );
  NOR2x1_ASAP7_75t_SL U49239 ( .A(n70700), .B(n70712), .Y(n70713) );
  HB1xp67_ASAP7_75t_SL U49240 ( .A(n70195), .Y(n53435) );
  NOR2x1_ASAP7_75t_SL U49241 ( .A(n73590), .B(n73660), .Y(n73610) );
  NOR2x2_ASAP7_75t_SL U49242 ( .A(n77451), .B(n62152), .Y(n77209) );
  INVx2_ASAP7_75t_SL U49243 ( .A(n62154), .Y(n62152) );
  NOR2x1_ASAP7_75t_SL U49244 ( .A(n70825), .B(n70824), .Y(n71162) );
  NOR2x1_ASAP7_75t_SL U49245 ( .A(n70823), .B(n59524), .Y(n70824) );
  NOR2x1p5_ASAP7_75t_SL U49246 ( .A(n70784), .B(n70783), .Y(n70795) );
  NOR2x1_ASAP7_75t_SL U49247 ( .A(n70774), .B(n70773), .Y(n70783) );
  AOI21x1_ASAP7_75t_SL U49248 ( .A1(n70836), .A2(n70819), .B(n70818), .Y(
        n70834) );
  OAI21x1_ASAP7_75t_SL U49249 ( .A1(n70797), .A2(n70795), .B(n70794), .Y(
        n70819) );
  NOR2x1_ASAP7_75t_SL U49250 ( .A(n70817), .B(n70816), .Y(n70836) );
  NOR2x1_ASAP7_75t_SL U49251 ( .A(n57111), .B(n57362), .Y(n62898) );
  INVx8_ASAP7_75t_SL U49252 ( .A(n58447), .Y(n57203) );
  OAI22xp5_ASAP7_75t_SL U49253 ( .A1(n57077), .A2(n76094), .B1(
        or1200_cpu_or1200_mult_mac_n30), .B2(n57105), .Y(
        or1200_cpu_or1200_mult_mac_n1510) );
  OAI22xp5_ASAP7_75t_SL U49254 ( .A1(n57077), .A2(n75987), .B1(
        or1200_cpu_or1200_mult_mac_n60), .B2(n57105), .Y(
        or1200_cpu_or1200_mult_mac_n1525) );
  OAI22xp5_ASAP7_75t_SL U49255 ( .A1(n57077), .A2(n76170), .B1(
        or1200_cpu_or1200_mult_mac_n12), .B2(n57105), .Y(
        or1200_cpu_or1200_mult_mac_n1501) );
  OAI22xp5_ASAP7_75t_SL U49256 ( .A1(n57077), .A2(n76121), .B1(
        or1200_cpu_or1200_mult_mac_n24), .B2(n57105), .Y(
        or1200_cpu_or1200_mult_mac_n1507) );
  OAI22xp5_ASAP7_75t_SL U49257 ( .A1(n57077), .A2(n76184), .B1(
        or1200_cpu_or1200_mult_mac_n6), .B2(n57105), .Y(
        or1200_cpu_or1200_mult_mac_n1498) );
  OAI22xp5_ASAP7_75t_SL U49258 ( .A1(n57077), .A2(n76180), .B1(
        or1200_cpu_or1200_mult_mac_n8), .B2(n57105), .Y(
        or1200_cpu_or1200_mult_mac_n1499) );
  BUFx3_ASAP7_75t_SL U49259 ( .A(n60523), .Y(n53436) );
  INVx3_ASAP7_75t_SL U49260 ( .A(n53436), .Y(n77379) );
  NOR2x1_ASAP7_75t_SL U49261 ( .A(n71152), .B(n71151), .Y(n71169) );
  INVx1_ASAP7_75t_SL U49262 ( .A(n71074), .Y(n70788) );
  OAI22xp5_ASAP7_75t_SL U49263 ( .A1(n57077), .A2(n76175), .B1(
        or1200_cpu_or1200_mult_mac_n10), .B2(n57105), .Y(
        or1200_cpu_or1200_mult_mac_n1500) );
  HB1xp67_ASAP7_75t_SL U49264 ( .A(n68795), .Y(n53437) );
  INVxp33_ASAP7_75t_SRAM U49265 ( .A(n69271), .Y(n69263) );
  OAI21x1_ASAP7_75t_SL U49266 ( .A1(n69255), .A2(n69254), .B(n69253), .Y(
        n69271) );
  OAI22xp5_ASAP7_75t_SL U49267 ( .A1(n57115), .A2(n70893), .B1(n70881), .B2(
        n70993), .Y(n71219) );
  NOR2x1_ASAP7_75t_SL U49268 ( .A(n70687), .B(n70993), .Y(n70688) );
  OAI22xp5_ASAP7_75t_SL U49269 ( .A1(n57115), .A2(n70911), .B1(n70910), .B2(
        n70993), .Y(n71244) );
  INVx1_ASAP7_75t_SL U49270 ( .A(n70993), .Y(n71013) );
  NOR2x1p5_ASAP7_75t_SL U49271 ( .A(n78197), .B(n74218), .Y(n74839) );
  NOR2x1p5_ASAP7_75t_SL U49272 ( .A(n76956), .B(n74839), .Y(n74901) );
  INVx8_ASAP7_75t_SL U49273 ( .A(n58291), .Y(n57115) );
  AND2x4_ASAP7_75t_SL U49274 ( .A(n70686), .B(n70721), .Y(n58291) );
  NOR2x1_ASAP7_75t_SL U49275 ( .A(n76588), .B(n76589), .Y(n76587) );
  BUFx4_ASAP7_75t_SL U49276 ( .A(n1667), .Y(n59535) );
  NAND2x1_ASAP7_75t_SL U49277 ( .A(n1667), .B(n1651), .Y(n59053) );
  NAND2xp5_ASAP7_75t_SL U49278 ( .A(n71315), .B(n71073), .Y(n70915) );
  INVx2_ASAP7_75t_SL U49279 ( .A(n76590), .Y(n53438) );
  INVx1_ASAP7_75t_SL U49280 ( .A(n53438), .Y(n53439) );
  INVx3_ASAP7_75t_SL U49281 ( .A(n53438), .Y(n53440) );
  AND2x2_ASAP7_75t_SL U49282 ( .A(n57100), .B(n53439), .Y(n53441) );
  NOR2x1_ASAP7_75t_SL U49283 ( .A(n77349), .B(n77341), .Y(n77352) );
  NAND2xp5_ASAP7_75t_SL U49284 ( .A(n77997), .B(n77998), .Y(n53442) );
  NAND2x1_ASAP7_75t_SL U49285 ( .A(n59945), .B(n77012), .Y(n77292) );
  NAND2x1_ASAP7_75t_SL U49286 ( .A(n77997), .B(n77998), .Y(n59875) );
  INVx13_ASAP7_75t_SL U49287 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_21_), .Y(
        n53443) );
  AND2x4_ASAP7_75t_SL U49288 ( .A(n74430), .B(n53444), .Y(n74441) );
  NOR2x1p5_ASAP7_75t_SL U49289 ( .A(n53443), .B(n74442), .Y(n53444) );
  NOR2x1p5_ASAP7_75t_SL U49290 ( .A(n74422), .B(n74423), .Y(n74430) );
  INVxp33_ASAP7_75t_SRAM U49291 ( .A(n75442), .Y(n53445) );
  INVx1_ASAP7_75t_SL U49292 ( .A(n53445), .Y(n53446) );
  NOR2x1_ASAP7_75t_SL U49293 ( .A(n59837), .B(n59838), .Y(n77998) );
  INVxp33_ASAP7_75t_SRAM U49294 ( .A(n63445), .Y(n55006) );
  INVx5_ASAP7_75t_SL U49295 ( .A(n59582), .Y(n78327) );
  NOR2x1_ASAP7_75t_SL U49296 ( .A(n75750), .B(n75751), .Y(n75749) );
  AND2x4_ASAP7_75t_SL U49297 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .B(
        n59527), .Y(n58447) );
  INVx4_ASAP7_75t_SL U49298 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .Y(
        n72367) );
  OAI21xp5_ASAP7_75t_SL U49299 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .A2(
        n72533), .B(n72525), .Y(n72529) );
  NOR2x1_ASAP7_75t_SL U49300 ( .A(n78200), .B(n78201), .Y(n74215) );
  OAI22xp5_ASAP7_75t_SL U49301 ( .A1(n57077), .A2(n76189), .B1(
        or1200_cpu_or1200_mult_mac_n4), .B2(n57105), .Y(
        or1200_cpu_or1200_mult_mac_n1497) );
  HB1xp67_ASAP7_75t_SL U49302 ( .A(n77347), .Y(n53447) );
  BUFx6f_ASAP7_75t_SL U49303 ( .A(n77336), .Y(n53448) );
  BUFx6f_ASAP7_75t_SL U49304 ( .A(n77336), .Y(n57136) );
  HB1xp67_ASAP7_75t_SL U49305 ( .A(n75673), .Y(n53449) );
  NOR2x1p5_ASAP7_75t_SL U49306 ( .A(n75672), .B(n75671), .Y(n75673) );
  AND2x2_ASAP7_75t_SL U49307 ( .A(n53450), .B(n77307), .Y(n77347) );
  OR2x2_ASAP7_75t_SL U49308 ( .A(n1853), .B(n77338), .Y(n53450) );
  INVx1_ASAP7_75t_SL U49309 ( .A(n77307), .Y(n77313) );
  NAND2x1p5_ASAP7_75t_SL U49310 ( .A(n70554), .B(n74288), .Y(n74369) );
  OAI21x1_ASAP7_75t_SL U49311 ( .A1(n70567), .A2(n70566), .B(n74284), .Y(
        n74288) );
  INVx3_ASAP7_75t_SL U49312 ( .A(n76004), .Y(n76158) );
  NAND2x1p5_ASAP7_75t_SL U49313 ( .A(n58302), .B(n58373), .Y(n70993) );
  NOR2x1_ASAP7_75t_SL U49314 ( .A(n53442), .B(n59874), .Y(n60210) );
  NAND2x1_ASAP7_75t_SL U49315 ( .A(n60282), .B(n77500), .Y(n77341) );
  NOR2x1_ASAP7_75t_SL U49316 ( .A(n69272), .B(n69271), .Y(n69326) );
  OAI21xp5_ASAP7_75t_SL U49317 ( .A1(n75778), .A2(n59847), .B(n59846), .Y(
        n59849) );
  NOR2x1p5_ASAP7_75t_SL U49318 ( .A(n63719), .B(n60221), .Y(n63706) );
  NOR2x2_ASAP7_75t_SL U49319 ( .A(n74925), .B(n63701), .Y(n62150) );
  NOR2x1_ASAP7_75t_SL U49320 ( .A(n62083), .B(n62082), .Y(n75306) );
  INVx1_ASAP7_75t_SL U49321 ( .A(n62501), .Y(n62082) );
  NAND2x1_ASAP7_75t_SL U49322 ( .A(n77353), .B(n77398), .Y(n59157) );
  INVx3_ASAP7_75t_SL U49323 ( .A(n59498), .Y(n61826) );
  NAND2x1_ASAP7_75t_SL U49324 ( .A(n73236), .B(n73480), .Y(n73478) );
  NAND2x1_ASAP7_75t_SL U49325 ( .A(n73482), .B(n73481), .Y(n73480) );
  AOI31xp67_ASAP7_75t_SL U49326 ( .A1(n73447), .A2(n73366), .A3(n73448), .B(
        n73321), .Y(n73360) );
  AO21x2_ASAP7_75t_SL U49327 ( .A1(n73301), .A2(n73436), .B(n73300), .Y(n73447) );
  OAI21xp33_ASAP7_75t_SRAM U49328 ( .A1(n74120), .A2(n75427), .B(n74119), .Y(
        n76228) );
  NAND2x1p5_ASAP7_75t_SL U49329 ( .A(n74926), .B(n63706), .Y(n63701) );
  NOR2x1_ASAP7_75t_SL U49330 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_10_), .B(n65385), .Y(
        n65244) );
  NOR2x1p5_ASAP7_75t_SL U49331 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_r_a), .B(n65363), .Y(
        n65318) );
  NAND2x1p5_ASAP7_75t_SL U49332 ( .A(n65361), .B(n65353), .Y(n65363) );
  NOR2x1_ASAP7_75t_SL U49333 ( .A(n63754), .B(n76587), .Y(n77268) );
  NOR2x2_ASAP7_75t_SL U49334 ( .A(n69747), .B(n69445), .Y(n70149) );
  AOI22xp5_ASAP7_75t_SL U49335 ( .A1(n70151), .A2(n70150), .B1(n70149), .B2(
        n70148), .Y(n70175) );
  INVx2_ASAP7_75t_SL U49336 ( .A(n70149), .Y(n70077) );
  NOR2x1_ASAP7_75t_SL U49337 ( .A(n62087), .B(n62086), .Y(n64147) );
  INVx1_ASAP7_75t_SL U49338 ( .A(n74627), .Y(n62086) );
  NOR2x2_ASAP7_75t_SL U49339 ( .A(n77308), .B(n77347), .Y(n77314) );
  OR3x2_ASAP7_75t_SL U49340 ( .A(n77314), .B(n59156), .C(n59158), .Y(n77336)
         );
  BUFx3_ASAP7_75t_SL U49341 ( .A(n58434), .Y(n58316) );
  NOR2x1p5_ASAP7_75t_SL U49342 ( .A(n77314), .B(n59157), .Y(n58434) );
  AOI31xp33_ASAP7_75t_SL U49343 ( .A1(n62150), .A2(n60300), .A3(n62148), .B(
        n60265), .Y(n77449) );
  NOR2x2_ASAP7_75t_SL U49344 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[0]), .B(
        n70104), .Y(n70110) );
  INVxp33_ASAP7_75t_SRAM U49345 ( .A(n70104), .Y(n70106) );
  OAI21x1_ASAP7_75t_SL U49346 ( .A1(n70131), .A2(n70130), .B(n70129), .Y(
        n70142) );
  NAND2x1p5_ASAP7_75t_SL U49347 ( .A(n69766), .B(n70104), .Y(n70054) );
  NOR2x2_ASAP7_75t_SL U49348 ( .A(n70124), .B(n70104), .Y(n70038) );
  NAND2xp5_ASAP7_75t_SL U49349 ( .A(n69948), .B(n70104), .Y(n69925) );
  NOR2xp33_ASAP7_75t_SL U49350 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[14]), .B(n70104), .Y(n69894) );
  NAND3x2_ASAP7_75t_SL U49351 ( .A(n75548), .B(n75449), .C(n75622), .Y(n75549)
         );
  NOR2x1p5_ASAP7_75t_SL U49352 ( .A(or1200_cpu_or1200_except_n530), .B(n64107), 
        .Y(n75548) );
  NOR2x1p5_ASAP7_75t_SL U49353 ( .A(n61839), .B(n75549), .Y(n64814) );
  NAND2x1_ASAP7_75t_SL U49354 ( .A(n73263), .B(n73469), .Y(n73453) );
  OAI21xp5_ASAP7_75t_SL U49355 ( .A1(n73291), .A2(n73410), .B(n73290), .Y(
        n73436) );
  NAND2x1_ASAP7_75t_SL U49356 ( .A(n59560), .B(n59570), .Y(n57578) );
  NOR2x1p5_ASAP7_75t_SL U49357 ( .A(n74311), .B(n74312), .Y(n74416) );
  NAND2x1p5_ASAP7_75t_SL U49358 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_18_), 
        .B(n74403), .Y(n74312) );
  NAND2x1p5_ASAP7_75t_SL U49359 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_22_), 
        .B(n74435), .Y(n74434) );
  NOR2x1p5_ASAP7_75t_SL U49360 ( .A(n74425), .B(n74426), .Y(n74435) );
  XOR2xp5_ASAP7_75t_SL U49361 ( .A(n53451), .B(n75300), .Y(n59733) );
  INVx13_ASAP7_75t_SL U49362 ( .A(or1200_dc_top_tag_5_), .Y(n53451) );
  NAND2x1p5_ASAP7_75t_SL U49363 ( .A(n69574), .B(n69431), .Y(n70118) );
  INVx3_ASAP7_75t_SL U49364 ( .A(n70118), .Y(n70078) );
  NOR2xp33_ASAP7_75t_SL U49365 ( .A(n70118), .B(n69808), .Y(n69434) );
  NAND2x1_ASAP7_75t_SL U49366 ( .A(n71267), .B(n71276), .Y(n71205) );
  NOR2x1p5_ASAP7_75t_SL U49367 ( .A(n74226), .B(n74434), .Y(n74227) );
  NAND2x1_ASAP7_75t_SL U49368 ( .A(n74270), .B(n74250), .Y(n74254) );
  OA21x2_ASAP7_75t_SL U49369 ( .A1(n63361), .A2(n58817), .B(n57889), .Y(n53452) );
  NAND2x1_ASAP7_75t_SL U49370 ( .A(n58816), .B(n58815), .Y(n63361) );
  HB1xp67_ASAP7_75t_SL U49371 ( .A(n74998), .Y(n53453) );
  NAND2xp5_ASAP7_75t_SL U49372 ( .A(n63399), .B(n63398), .Y(n63401) );
  INVx2_ASAP7_75t_SL U49373 ( .A(n59875), .Y(n59883) );
  NOR2x1p5_ASAP7_75t_SL U49374 ( .A(n60283), .B(n77352), .Y(n77796) );
  INVxp33_ASAP7_75t_SRAM U49375 ( .A(n53449), .Y(n54249) );
  NAND2x1_ASAP7_75t_SL U49376 ( .A(n69734), .B(n69735), .Y(n69762) );
  NOR2x1_ASAP7_75t_SL U49377 ( .A(n70098), .B(n70097), .Y(n70099) );
  NOR2x1_ASAP7_75t_SL U49378 ( .A(n70093), .B(n70094), .Y(n70097) );
  NAND2xp67_ASAP7_75t_SRAM U49379 ( .A(iwb_dat_i[21]), .B(n77373), .Y(n60429)
         );
  AOI21xp5_ASAP7_75t_SL U49380 ( .A1(n77765), .A2(n60295), .B(n60204), .Y(
        n60205) );
  INVx11_ASAP7_75t_SL U49381 ( .A(n57144), .Y(n59690) );
  NOR2x1_ASAP7_75t_SL U49382 ( .A(n70902), .B(n70903), .Y(n70938) );
  INVx2_ASAP7_75t_SL U49383 ( .A(n77943), .Y(n77966) );
  NOR2x1_ASAP7_75t_SL U49384 ( .A(n77943), .B(n61342), .Y(n61693) );
  NOR2xp33_ASAP7_75t_SL U49385 ( .A(n77943), .B(n64283), .Y(n75555) );
  NOR2x1p5_ASAP7_75t_SL U49386 ( .A(n59931), .B(n59930), .Y(n77943) );
  NAND2xp5_ASAP7_75t_SL U49387 ( .A(n76720), .B(n77852), .Y(n61755) );
  AOI22xp5_ASAP7_75t_SL U49388 ( .A1(n62318), .A2(n62409), .B1(n62317), .B2(
        n76720), .Y(n62381) );
  AOI21xp5_ASAP7_75t_SL U49389 ( .A1(n76720), .A2(n62237), .B(n62236), .Y(
        n77601) );
  NOR2x2_ASAP7_75t_SL U49390 ( .A(n77966), .B(n64283), .Y(n76720) );
  NAND2x1p5_ASAP7_75t_SL U49391 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_23_), .B(
        n74441), .Y(n74449) );
  NAND3x2_ASAP7_75t_SL U49392 ( .A(n59949), .B(n60273), .C(n59948), .Y(n22057)
         );
  AOI21x1_ASAP7_75t_SL U49393 ( .A1(n60274), .A2(n2759), .B(n57084), .Y(n59949) );
  INVx8_ASAP7_75t_SL U49394 ( .A(n58451), .Y(n57168) );
  AND2x4_ASAP7_75t_SL U49395 ( .A(n59968), .B(n77367), .Y(n58451) );
  O2A1O1Ixp5_ASAP7_75t_SL U49396 ( .A1(n58315), .A2(n70652), .B(n70651), .C(
        n58307), .Y(n70656) );
  OAI21x1_ASAP7_75t_SL U49397 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[11]), .A2(
        n73171), .B(n73063), .Y(n73075) );
  NAND2x1_ASAP7_75t_SL U49398 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[12]), .B(
        n73180), .Y(n73063) );
  INVx1_ASAP7_75t_SL U49399 ( .A(n76204), .Y(n76206) );
  INVxp33_ASAP7_75t_SRAM U49400 ( .A(n71024), .Y(n70979) );
  AO21x2_ASAP7_75t_SL U49401 ( .A1(n75953), .A2(n75959), .B(n75952), .Y(n76181) );
  NOR2x1_ASAP7_75t_SL U49402 ( .A(n75896), .B(n76136), .Y(n76143) );
  NOR2x1_ASAP7_75t_SL U49403 ( .A(n76133), .B(n76132), .Y(n76136) );
  NAND2x1_ASAP7_75t_SL U49404 ( .A(n75452), .B(n60575), .Y(n60833) );
  NAND2xp5_ASAP7_75t_SL U49405 ( .A(n61481), .B(n60575), .Y(n77165) );
  NAND2xp5_ASAP7_75t_SL U49406 ( .A(n77853), .B(n60575), .Y(n60576) );
  NOR2x1p5_ASAP7_75t_SL U49407 ( .A(n60550), .B(n59973), .Y(n60575) );
  NAND2x1_ASAP7_75t_SL U49408 ( .A(n77312), .B(n77313), .Y(n77398) );
  OA21x2_ASAP7_75t_SL U49409 ( .A1(n60731), .A2(n75478), .B(n76327), .Y(n53454) );
  OA21x2_ASAP7_75t_SL U49410 ( .A1(n60731), .A2(n75478), .B(n76327), .Y(n53455) );
  HB1xp67_ASAP7_75t_SL U49411 ( .A(n62501), .Y(n53456) );
  INVx8_ASAP7_75t_SL U49412 ( .A(n53454), .Y(n57120) );
  NOR2x1_ASAP7_75t_SL U49413 ( .A(n76946), .B(n74840), .Y(n74902) );
  NOR2x1_ASAP7_75t_SL U49414 ( .A(n78246), .B(n78203), .Y(n58663) );
  OAI21xp5_ASAP7_75t_SL U49415 ( .A1(n74166), .A2(n74190), .B(n74179), .Y(
        n74198) );
  OAI21xp5_ASAP7_75t_SL U49416 ( .A1(n70879), .A2(n70878), .B(n70877), .Y(
        n71055) );
  NOR2x1_ASAP7_75t_SL U49417 ( .A(n76117), .B(n75913), .Y(n75937) );
  NAND2xp5_ASAP7_75t_SL U49418 ( .A(n76109), .B(n75938), .Y(n75913) );
  OAI21xp5_ASAP7_75t_SL U49419 ( .A1(n76097), .A2(n76090), .B(n75936), .Y(
        n76095) );
  NAND2x1p5_ASAP7_75t_SL U49420 ( .A(n58304), .B(n73660), .Y(n73652) );
  INVx4_ASAP7_75t_SL U49421 ( .A(n73616), .Y(n73660) );
  NAND4xp75_ASAP7_75t_SL U49422 ( .A(n60186), .B(n60185), .C(n60184), .D(
        n60183), .Y(n60187) );
  INVx1_ASAP7_75t_SL U49423 ( .A(n64809), .Y(n53457) );
  NOR2x1p5_ASAP7_75t_SL U49424 ( .A(n63514), .B(n63513), .Y(n63539) );
  NOR2x1_ASAP7_75t_SL U49425 ( .A(n63518), .B(n63523), .Y(n63513) );
  OAI21x1_ASAP7_75t_SL U49426 ( .A1(n74937), .A2(n63710), .B(n75768), .Y(
        n62148) );
  AOI21xp5_ASAP7_75t_SL U49427 ( .A1(n53436), .A2(or1200_ic_top_from_icram[21]), .B(n60428), .Y(n60430) );
  NOR2x1p5_ASAP7_75t_SL U49428 ( .A(n76503), .B(n60231), .Y(n77212) );
  AOI21x1_ASAP7_75t_SL U49429 ( .A1(n77459), .A2(n61162), .B(n77429), .Y(
        n76835) );
  NAND2xp5_ASAP7_75t_SL U49430 ( .A(n73257), .B(n73053), .Y(n73058) );
  NAND2x1_ASAP7_75t_SL U49431 ( .A(n70835), .B(n70834), .Y(n70840) );
  XNOR2xp5_ASAP7_75t_SL U49432 ( .A(n62953), .B(n62952), .Y(n57044) );
  NOR2x2_ASAP7_75t_SL U49433 ( .A(n60337), .B(n77834), .Y(n78173) );
  INVx3_ASAP7_75t_SL U49434 ( .A(n78440), .Y(n77834) );
  NOR2x1_ASAP7_75t_SL U49435 ( .A(n57090), .B(n78006), .Y(n77373) );
  NOR2x1_ASAP7_75t_SL U49436 ( .A(n77406), .B(n78006), .Y(n77836) );
  NOR2x1p5_ASAP7_75t_SL U49437 ( .A(n53473), .B(n71229), .Y(n71245) );
  AOI22xp5_ASAP7_75t_SL U49438 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[18]), .A2(n70675), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[17]), .B2(
        n70674), .Y(n70679) );
  NAND2x2_ASAP7_75t_SL U49439 ( .A(n59702), .B(n76847), .Y(n77276) );
  NAND2x1p5_ASAP7_75t_SL U49440 ( .A(n77833), .B(n60330), .Y(n78006) );
  HB1xp67_ASAP7_75t_SL U49441 ( .A(n74418), .Y(n53460) );
  INVx2_ASAP7_75t_SL U49442 ( .A(n74313), .Y(n74444) );
  NAND2x1_ASAP7_75t_SL U49443 ( .A(n74270), .B(n74362), .Y(n74313) );
  OAI21xp33_ASAP7_75t_SRAM U49444 ( .A1(n73482), .A2(n73481), .B(n73480), .Y(
        n12864) );
  AOI21x1_ASAP7_75t_SL U49445 ( .A1(n69161), .A2(n69275), .B(n69277), .Y(
        n69213) );
  INVx6_ASAP7_75t_SL U49446 ( .A(n59712), .Y(n59711) );
  INVx4_ASAP7_75t_SL U49447 ( .A(n1725), .Y(n59712) );
  INVx4_ASAP7_75t_SL U49448 ( .A(n59712), .Y(n59710) );
  INVx2_ASAP7_75t_SL U49449 ( .A(n74254), .Y(n74437) );
  NOR2x2_ASAP7_75t_SL U49450 ( .A(n69348), .B(n69370), .Y(n77235) );
  BUFx5_ASAP7_75t_SL U49451 ( .A(n77289), .Y(n57135) );
  AOI22xp5_ASAP7_75t_SL U49452 ( .A1(n76114), .A2(n75938), .B1(n76095), .B2(
        n75937), .Y(n76123) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U49453 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[5]), .A2(
        n74502), .B(n73260), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[5]), .Y(
        n73261) );
  NAND2xp33_ASAP7_75t_SRAM U49454 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[5]), .B(
        n58284), .Y(n73223) );
  OAI22xp33_ASAP7_75t_SRAM U49455 ( .A1(n76818), .A2(n76817), .B1(n59703), 
        .B2(n76816), .Y(n76819) );
  AOI22xp33_ASAP7_75t_SRAM U49456 ( .A1(n59701), .A2(n63984), .B1(n63983), 
        .B2(n53440), .Y(n63985) );
  AOI22xp33_ASAP7_75t_SRAM U49457 ( .A1(n59701), .A2(n63987), .B1(n63986), 
        .B2(n53440), .Y(n63988) );
  AOI22xp33_ASAP7_75t_SRAM U49458 ( .A1(n59701), .A2(n75171), .B1(n75170), 
        .B2(n53440), .Y(n75172) );
  AOI22xp33_ASAP7_75t_SRAM U49459 ( .A1(n59701), .A2(n75174), .B1(n75173), 
        .B2(n53440), .Y(n75175) );
  AOI22xp33_ASAP7_75t_SRAM U49460 ( .A1(n59701), .A2(n75161), .B1(n75160), 
        .B2(n53440), .Y(n75162) );
  NAND2xp33_ASAP7_75t_SRAM U49461 ( .A(n76604), .B(n53440), .Y(n61176) );
  INVxp33_ASAP7_75t_SRAM U49462 ( .A(n53440), .Y(n76593) );
  BUFx2_ASAP7_75t_SL U49463 ( .A(n70667), .Y(n58300) );
  AOI31xp67_ASAP7_75t_SL U49464 ( .A1(n71303), .A2(n71302), .A3(n71301), .B(
        n71300), .Y(n71304) );
  NAND2x1p5_ASAP7_75t_SL U49465 ( .A(n59982), .B(n60116), .Y(n60114) );
  NAND2x1_ASAP7_75t_SL U49466 ( .A(n78183), .B(n4095), .Y(icqmem_adr_qmem[31])
         );
  NOR2x1_ASAP7_75t_SL U49467 ( .A(n59981), .B(n60041), .Y(n60116) );
  INVxp33_ASAP7_75t_SRAM U49468 ( .A(n58372), .Y(n53461) );
  INVx1_ASAP7_75t_SL U49469 ( .A(n53461), .Y(n53462) );
  NOR2x1p5_ASAP7_75t_SL U49470 ( .A(n74838), .B(n74875), .Y(n74204) );
  INVx2_ASAP7_75t_SL U49471 ( .A(n78243), .Y(n71512) );
  NAND2x1_ASAP7_75t_SL U49472 ( .A(n78366), .B(n69556), .Y(n69557) );
  NOR2x1_ASAP7_75t_SL U49473 ( .A(n70114), .B(n70113), .Y(n70123) );
  OAI22xp5_ASAP7_75t_SL U49474 ( .A1(n59698), .A2(n71261), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_39_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n220) );
  NOR2x1_ASAP7_75t_SL U49475 ( .A(n70765), .B(n70764), .Y(n70784) );
  HB1xp67_ASAP7_75t_SL U49476 ( .A(n73469), .Y(n53463) );
  NOR2x1_ASAP7_75t_SL U49477 ( .A(n61953), .B(n62497), .Y(n76257) );
  A2O1A1Ixp33_ASAP7_75t_SL U49478 ( .A1(n75996), .A2(n75995), .B(n75994), .C(
        n75998), .Y(n53464) );
  NAND3x1_ASAP7_75t_SL U49479 ( .A(n74215), .B(n58664), .C(n58663), .Y(n74218)
         );
  NOR2x1_ASAP7_75t_SL U49480 ( .A(n78202), .B(n74214), .Y(n58664) );
  NOR2x1p5_ASAP7_75t_SL U49481 ( .A(n77171), .B(n74901), .Y(n74872) );
  NOR2x1p5_ASAP7_75t_SL U49482 ( .A(n60421), .B(n57090), .Y(n76847) );
  NOR2x1_ASAP7_75t_SL U49483 ( .A(n63755), .B(n77266), .Y(n76602) );
  NOR2x1_ASAP7_75t_SL U49484 ( .A(n77267), .B(n77268), .Y(n77266) );
  NOR2x2_ASAP7_75t_SL U49485 ( .A(n58604), .B(n74966), .Y(n64162) );
  NOR2x1p5_ASAP7_75t_SL U49486 ( .A(n74967), .B(n74968), .Y(n74966) );
  NOR4xp75_ASAP7_75t_SL U49487 ( .A(n60187), .B(n60189), .C(n60188), .D(n60190), .Y(n60267) );
  AOI22xp5_ASAP7_75t_SL U49488 ( .A1(n77506), .A2(n77505), .B1(n58434), .B2(
        n77796), .Y(n77795) );
  INVx1_ASAP7_75t_SL U49489 ( .A(n62077), .Y(n62078) );
  AOI21xp5_ASAP7_75t_SL U49490 ( .A1(n76324), .A2(n2826), .B(n76321), .Y(
        n76332) );
  NOR2x1_ASAP7_75t_SL U49491 ( .A(n61986), .B(n75683), .Y(n75519) );
  XNOR2x1_ASAP7_75t_SL U49492 ( .A(n61987), .B(n75519), .Y(n76256) );
  NOR2x1_ASAP7_75t_SL U49493 ( .A(n61236), .B(n61237), .Y(n61397) );
  NOR2x1_ASAP7_75t_SL U49494 ( .A(n64188), .B(n76277), .Y(n75554) );
  NOR2x1_ASAP7_75t_SL U49495 ( .A(n64187), .B(n64197), .Y(n76277) );
  NOR2x1_ASAP7_75t_SL U49496 ( .A(n70938), .B(n70937), .Y(n70975) );
  AOI31xp33_ASAP7_75t_SL U49497 ( .A1(n71053), .A2(n71052), .A3(n71051), .B(
        n71050), .Y(n71054) );
  NAND2xp33_ASAP7_75t_SRAM U49498 ( .A(n71245), .B(n71331), .Y(n71246) );
  AOI22xp33_ASAP7_75t_SRAM U49499 ( .A1(n71245), .A2(n71074), .B1(n71087), 
        .B2(n71244), .Y(n70999) );
  AOI22xp33_ASAP7_75t_SRAM U49500 ( .A1(n71209), .A2(n71138), .B1(n71245), 
        .B2(n71192), .Y(n71285) );
  AOI22xp33_ASAP7_75t_SRAM U49501 ( .A1(n71245), .A2(n71115), .B1(n71087), 
        .B2(n71311), .Y(n71065) );
  AOI22xp33_ASAP7_75t_SRAM U49502 ( .A1(n71209), .A2(n71016), .B1(n71245), 
        .B2(n71085), .Y(n71017) );
  INVxp33_ASAP7_75t_SRAM U49503 ( .A(n71245), .Y(n70895) );
  NOR2x1_ASAP7_75t_SL U49504 ( .A(n75939), .B(n76145), .Y(n76162) );
  NOR2x1_ASAP7_75t_SL U49505 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_12_), .B(n65246), .Y(
        n65248) );
  AOI21x1_ASAP7_75t_SL U49506 ( .A1(n65275), .A2(n2865), .B(n78435), .Y(n65277) );
  NOR2x1p5_ASAP7_75t_SL U49507 ( .A(n65264), .B(n65263), .Y(n65275) );
  O2A1O1Ixp5_ASAP7_75t_SL U49508 ( .A1(n57185), .A2(n73239), .B(n54559), .C(
        n54560), .Y(n73248) );
  NOR2x1_ASAP7_75t_SL U49509 ( .A(n76258), .B(n76257), .Y(n76262) );
  INVx1_ASAP7_75t_SL U49510 ( .A(n63480), .Y(n53465) );
  INVx2_ASAP7_75t_SL U49511 ( .A(n53465), .Y(n53466) );
  AOI21x1_ASAP7_75t_SL U49512 ( .A1(n75988), .A2(
        or1200_cpu_or1200_mult_mac_n60), .B(n75989), .Y(n75996) );
  NOR2x1_ASAP7_75t_SL U49513 ( .A(n62079), .B(n62078), .Y(n64273) );
  OAI21x1_ASAP7_75t_SL U49514 ( .A1(n59863), .A2(n75427), .B(n59862), .Y(
        n75442) );
  NOR2x1_ASAP7_75t_SL U49515 ( .A(n61681), .B(n76541), .Y(n60221) );
  NAND2x2_ASAP7_75t_SL U49516 ( .A(n65400), .B(n74726), .Y(n65308) );
  NAND2x1p5_ASAP7_75t_SL U49517 ( .A(n65320), .B(n65318), .Y(n74726) );
  NAND4xp75_ASAP7_75t_SL U49518 ( .A(n60269), .B(n60268), .C(n60267), .D(
        n60266), .Y(n77307) );
  XNOR2xp5_ASAP7_75t_SL U49519 ( .A(n73247), .B(n73248), .Y(n73473) );
  NOR2x1_ASAP7_75t_SL U49520 ( .A(n73402), .B(n73403), .Y(n73401) );
  INVx1_ASAP7_75t_SL U49521 ( .A(n75299), .Y(n74981) );
  AOI22x1_ASAP7_75t_SL U49522 ( .A1(n71087), .A2(n70997), .B1(n70996), .B2(
        n71074), .Y(n70880) );
  OAI22x1_ASAP7_75t_SL U49523 ( .A1(n57115), .A2(n70709), .B1(n70705), .B2(
        n59524), .Y(n70997) );
  NOR2x1p5_ASAP7_75t_SL U49524 ( .A(n70772), .B(n70771), .Y(n70797) );
  INVx1_ASAP7_75t_SL U49525 ( .A(n70773), .Y(n70771) );
  NOR2x1_ASAP7_75t_SL U49526 ( .A(n70689), .B(n70688), .Y(n70882) );
  NOR2x1_ASAP7_75t_SL U49527 ( .A(n70691), .B(n57115), .Y(n70689) );
  AND2x2_ASAP7_75t_SL U49528 ( .A(n70996), .B(n70951), .Y(n53467) );
  AOI31xp67_ASAP7_75t_SL U49529 ( .A1(n69195), .A2(n69194), .A3(n69193), .B(
        n69192), .Y(n75295) );
  NOR2x1p5_ASAP7_75t_SL U49530 ( .A(n69086), .B(n69085), .Y(n69195) );
  OAI21x1_ASAP7_75t_SL U49531 ( .A1(n69206), .A2(n75295), .B(n69205), .Y(
        n69252) );
  INVx3_ASAP7_75t_SL U49532 ( .A(n59437), .Y(n59145) );
  NAND2x1_ASAP7_75t_SL U49533 ( .A(n70996), .B(n70951), .Y(n70768) );
  XNOR2xp5_ASAP7_75t_SL U49534 ( .A(n64674), .B(n64673), .Y(n64706) );
  NAND2x1p5_ASAP7_75t_SL U49535 ( .A(n70229), .B(n70371), .Y(n70528) );
  NOR2x2_ASAP7_75t_SL U49536 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_2_), .B(n70260), .Y(
        n70371) );
  NAND2xp5_ASAP7_75t_SL U49537 ( .A(n69594), .B(n69730), .Y(n69726) );
  NOR2x1_ASAP7_75t_SL U49538 ( .A(n59843), .B(n59726), .Y(n77012) );
  INVx5_ASAP7_75t_SL U49539 ( .A(n58315), .Y(n71314) );
  BUFx6f_ASAP7_75t_SL U49540 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_3_), .Y(n58315) );
  NAND2x1_ASAP7_75t_SL U49541 ( .A(n71255), .B(n71254), .Y(n71301) );
  INVxp33_ASAP7_75t_SRAM U49542 ( .A(n71053), .Y(n71034) );
  NOR2x1_ASAP7_75t_SL U49543 ( .A(n61398), .B(n61397), .Y(n61559) );
  AOI22xp5_ASAP7_75t_SL U49544 ( .A1(n70695), .A2(n70997), .B1(n71315), .B2(
        n53467), .Y(n70698) );
  INVxp33_ASAP7_75t_SRAM U49545 ( .A(n70880), .Y(n70852) );
  OAI22xp33_ASAP7_75t_SRAM U49546 ( .A1(n70880), .A2(n71335), .B1(n71284), 
        .B2(n71044), .Y(n70887) );
  AOI21xp5_ASAP7_75t_SL U49547 ( .A1(n68200), .A2(n68212), .B(n68199), .Y(
        n68140) );
  A2O1A1Ixp33_ASAP7_75t_SL U49548 ( .A1(n57133), .A2(n76080), .B(n54451), .C(
        n54453), .Y(n53469) );
  BUFx6f_ASAP7_75t_SL U49549 ( .A(n76187), .Y(n57133) );
  NAND2x2_ASAP7_75t_SL U49550 ( .A(n64163), .B(n64162), .Y(n65207) );
  NOR2x1_ASAP7_75t_SL U49551 ( .A(n58558), .B(n76600), .Y(n76815) );
  NOR2x1_ASAP7_75t_SL U49552 ( .A(n76601), .B(n76602), .Y(n76600) );
  OAI21x1_ASAP7_75t_SL U49553 ( .A1(n65208), .A2(n65207), .B(n65206), .Y(
        n65230) );
  AOI31xp67_ASAP7_75t_SL U49554 ( .A1(n59883), .A2(n60198), .A3(n60194), .B(
        n59880), .Y(n60213) );
  NOR2x1_ASAP7_75t_SL U49555 ( .A(n73271), .B(n73420), .Y(n73410) );
  A2O1A1Ixp33_ASAP7_75t_SL U49556 ( .A1(n62308), .A2(n62296), .B(n62309), .C(
        n60773), .Y(n53470) );
  INVx2_ASAP7_75t_SL U49557 ( .A(n67326), .Y(n67607) );
  XNOR2xp5_ASAP7_75t_SL U49558 ( .A(n63117), .B(n63116), .Y(n63118) );
  NAND2x1p5_ASAP7_75t_SL U49559 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_12_), 
        .B(n74328), .Y(n74340) );
  AOI21xp5_ASAP7_75t_SL U49560 ( .A1(n74321), .A2(n58283), .B(n74328), .Y(
        n74330) );
  NOR2x1p5_ASAP7_75t_SL U49561 ( .A(n74321), .B(n74322), .Y(n74328) );
  NAND2x1_ASAP7_75t_SL U49562 ( .A(n73870), .B(n74418), .Y(n73898) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U49563 ( .A1(n53460), .A2(n73875), .B(n73898), 
        .C(n74361), .Y(n73900) );
  NOR2xp33_ASAP7_75t_SL U49564 ( .A(n68981), .B(n68905), .Y(n58886) );
  NAND2x1p5_ASAP7_75t_SL U49565 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_22_), .B(n76933), 
        .Y(n74875) );
  NAND2xp5_ASAP7_75t_SL U49566 ( .A(n68973), .B(n58260), .Y(n68905) );
  OR2x6_ASAP7_75t_SL U49567 ( .A(n73379), .B(n73853), .Y(n58284) );
  XNOR2xp5_ASAP7_75t_SL U49568 ( .A(n67272), .B(n67508), .Y(n57523) );
  XOR2xp5_ASAP7_75t_SL U49569 ( .A(n68829), .B(n59208), .Y(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N34) );
  OAI21xp33_ASAP7_75t_SRAM U49570 ( .A1(n70819), .A2(n70841), .B(n70805), .Y(
        n70806) );
  NOR2x1p5_ASAP7_75t_SL U49571 ( .A(n70841), .B(n70840), .Y(n70876) );
  NOR2x1_ASAP7_75t_SL U49572 ( .A(n70811), .B(n70810), .Y(n71148) );
  NOR2x1_ASAP7_75t_SL U49573 ( .A(n71024), .B(n71025), .Y(n71033) );
  NAND2xp5_ASAP7_75t_SL U49574 ( .A(n57525), .B(n58892), .Y(n58657) );
  OAI21xp5_ASAP7_75t_SL U49575 ( .A1(n57525), .A2(n53251), .B(n58657), .Y(
        n67390) );
  INVx3_ASAP7_75t_SL U49576 ( .A(n59356), .Y(n58397) );
  NOR2x1_ASAP7_75t_SL U49577 ( .A(n68129), .B(n68131), .Y(n53522) );
  INVx1_ASAP7_75t_SL U49578 ( .A(n68239), .Y(n68230) );
  A2O1A1Ixp33_ASAP7_75t_SL U49579 ( .A1(n76165), .A2(n76166), .B(n75946), .C(
        n76163), .Y(n53471) );
  OR2x2_ASAP7_75t_SL U49580 ( .A(n53475), .B(n53618), .Y(n53472) );
  NAND2x1_ASAP7_75t_SL U49581 ( .A(n59595), .B(n59648), .Y(n68103) );
  NOR2x1_ASAP7_75t_SL U49582 ( .A(n59098), .B(n59434), .Y(n68807) );
  INVx2_ASAP7_75t_SL U49583 ( .A(n53501), .Y(n59434) );
  BUFx6f_ASAP7_75t_SL U49584 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_2_), .Y(n53473) );
  NAND2xp5_ASAP7_75t_SL U49585 ( .A(n59597), .B(n57912), .Y(n64684) );
  BUFx3_ASAP7_75t_SL U49586 ( .A(n53523), .Y(n53474) );
  NOR2x1_ASAP7_75t_SL U49587 ( .A(n69117), .B(n58677), .Y(n53523) );
  INVx1_ASAP7_75t_SL U49588 ( .A(n53523), .Y(n59427) );
  OA21x2_ASAP7_75t_SL U49589 ( .A1(n58910), .A2(n67400), .B(n58911), .Y(n53475) );
  INVxp33_ASAP7_75t_SRAM U49590 ( .A(n63993), .Y(n53476) );
  INVx1_ASAP7_75t_SL U49591 ( .A(n53476), .Y(n53477) );
  INVxp33_ASAP7_75t_SRAM U49592 ( .A(n75159), .Y(n53478) );
  INVx1_ASAP7_75t_SL U49593 ( .A(n53478), .Y(n53479) );
  AOI31xp67_ASAP7_75t_SL U49594 ( .A1(n63981), .A2(n63980), .A3(n63979), .B(
        n63978), .Y(n63993) );
  INVx3_ASAP7_75t_SL U49595 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .Y(n71229) );
  INVx1_ASAP7_75t_SL U49596 ( .A(n68328), .Y(n53480) );
  INVx2_ASAP7_75t_SL U49597 ( .A(n53480), .Y(n53481) );
  HB1xp67_ASAP7_75t_SL U49598 ( .A(n68740), .Y(n53482) );
  OAI21x1_ASAP7_75t_SL U49599 ( .A1(n67042), .A2(n67040), .B(n67041), .Y(
        n66981) );
  NOR2xp33_ASAP7_75t_SL U49600 ( .A(n68975), .B(n58887), .Y(n53529) );
  AOI21xp5_ASAP7_75t_SL U49601 ( .A1(n58885), .A2(n57086), .B(n58259), .Y(
        n58258) );
  XNOR2xp5_ASAP7_75t_SL U49602 ( .A(n66649), .B(n66648), .Y(n66775) );
  NOR2x1_ASAP7_75t_SL U49603 ( .A(n59518), .B(n66280), .Y(n67645) );
  XNOR2xp5_ASAP7_75t_SL U49604 ( .A(n68162), .B(n57891), .Y(n53483) );
  XNOR2xp5_ASAP7_75t_SL U49605 ( .A(n68162), .B(n57891), .Y(n68316) );
  NAND2x1_ASAP7_75t_SL U49606 ( .A(n58954), .B(n68159), .Y(n68162) );
  INVx1_ASAP7_75t_SL U49607 ( .A(n57026), .Y(n53484) );
  INVx2_ASAP7_75t_SL U49608 ( .A(n53484), .Y(n53485) );
  INVx2_ASAP7_75t_SL U49609 ( .A(n67842), .Y(n67315) );
  AOI22xp5_ASAP7_75t_SL U49610 ( .A1(n57380), .A2(n64467), .B1(n64466), .B2(
        n67842), .Y(n64471) );
  NOR2x1p5_ASAP7_75t_SL U49611 ( .A(n59487), .B(n59484), .Y(n67639) );
  NOR2x1p5_ASAP7_75t_SL U49612 ( .A(n58211), .B(n68098), .Y(n59408) );
  INVx1_ASAP7_75t_SL U49613 ( .A(n67602), .Y(n57849) );
  XOR2x1_ASAP7_75t_SL U49614 ( .A(n59247), .B(n64591), .Y(n58337) );
  AOI22x1_ASAP7_75t_SL U49615 ( .A1(n67476), .A2(n57273), .B1(n67475), .B2(
        n67700), .Y(n67686) );
  XNOR2xp5_ASAP7_75t_SL U49616 ( .A(n57943), .B(n57853), .Y(n53486) );
  XOR2x2_ASAP7_75t_SL U49617 ( .A(n67273), .B(n57854), .Y(n57853) );
  INVx1_ASAP7_75t_SL U49618 ( .A(n66497), .Y(n66505) );
  XNOR2x2_ASAP7_75t_SL U49619 ( .A(n66508), .B(n66513), .Y(n67111) );
  NAND2x1_ASAP7_75t_SL U49620 ( .A(n67448), .B(n67449), .Y(n67624) );
  HB1xp67_ASAP7_75t_SL U49621 ( .A(n68402), .Y(n53487) );
  INVx1_ASAP7_75t_SL U49622 ( .A(n53517), .Y(n53488) );
  INVx2_ASAP7_75t_SL U49623 ( .A(n57644), .Y(n53517) );
  AOI21x1_ASAP7_75t_SL U49624 ( .A1(n67446), .A2(n66852), .B(n57546), .Y(
        n67006) );
  OAI22x1_ASAP7_75t_SL U49625 ( .A1(n67284), .A2(n67283), .B1(n67282), .B2(
        n75032), .Y(n67472) );
  BUFx3_ASAP7_75t_SL U49626 ( .A(n64907), .Y(n58394) );
  NAND2x1_ASAP7_75t_SL U49627 ( .A(n58998), .B(n58997), .Y(n68916) );
  NAND2x1_ASAP7_75t_SL U49628 ( .A(n62688), .B(n58353), .Y(n75917) );
  NAND2x1_ASAP7_75t_SL U49629 ( .A(n59585), .B(n64779), .Y(n62688) );
  INVx2_ASAP7_75t_SL U49630 ( .A(n59514), .Y(n67850) );
  OAI22x1_ASAP7_75t_SL U49631 ( .A1(n66859), .A2(n57076), .B1(n67871), .B2(
        n67003), .Y(n67034) );
  INVx3_ASAP7_75t_SL U49632 ( .A(n67593), .Y(n67871) );
  XOR2x1_ASAP7_75t_SL U49633 ( .A(n68546), .B(n59016), .Y(n69036) );
  XNOR2x2_ASAP7_75t_SL U49634 ( .A(n66780), .B(n59086), .Y(n68546) );
  HB1xp67_ASAP7_75t_SL U49635 ( .A(n68251), .Y(n53489) );
  HB1xp67_ASAP7_75t_SL U49636 ( .A(n58324), .Y(n53490) );
  NOR2x1_ASAP7_75t_SL U49637 ( .A(n59101), .B(n66679), .Y(n66871) );
  NAND2x1p5_ASAP7_75t_SL U49638 ( .A(n57556), .B(n56980), .Y(n66263) );
  NOR2x1_ASAP7_75t_SL U49639 ( .A(n53314), .B(n57085), .Y(n68725) );
  XNOR2xp5_ASAP7_75t_SL U49640 ( .A(n57930), .B(n53491), .Y(n58255) );
  AOI21xp5_ASAP7_75t_SL U49641 ( .A1(n67833), .A2(n57069), .B(n67832), .Y(
        n53491) );
  NOR2x1_ASAP7_75t_SL U49642 ( .A(n75642), .B(n58775), .Y(n67340) );
  BUFx2_ASAP7_75t_SL U49643 ( .A(n59104), .Y(n53492) );
  NAND2x1_ASAP7_75t_SL U49644 ( .A(n67856), .B(n67857), .Y(n67873) );
  NAND2x1p5_ASAP7_75t_SL U49645 ( .A(n56972), .B(n58915), .Y(n67872) );
  INVx1_ASAP7_75t_SL U49646 ( .A(n64890), .Y(n54535) );
  AOI22xp33_ASAP7_75t_SRAM U49647 ( .A1(n59100), .A2(n67419), .B1(n67298), 
        .B2(n67229), .Y(n53493) );
  INVx8_ASAP7_75t_SL U49648 ( .A(n59506), .Y(n68079) );
  XNOR2x1_ASAP7_75t_SL U49649 ( .A(n58472), .B(n57512), .Y(n59294) );
  INVx2_ASAP7_75t_SL U49650 ( .A(n57468), .Y(n53494) );
  NAND2xp5_ASAP7_75t_SL U49651 ( .A(n67833), .B(n66994), .Y(n66995) );
  AOI21xp5_ASAP7_75t_SL U49652 ( .A1(n57069), .A2(n67833), .B(n67832), .Y(
        n67313) );
  NOR2x1_ASAP7_75t_SL U49653 ( .A(n57946), .B(n67350), .Y(n57945) );
  XNOR2x1_ASAP7_75t_SL U49654 ( .A(n57856), .B(n67291), .Y(n67486) );
  HB1xp67_ASAP7_75t_SL U49655 ( .A(n57522), .Y(n53495) );
  INVx2_ASAP7_75t_SL U49656 ( .A(n68034), .Y(n58739) );
  HB1xp67_ASAP7_75t_SL U49657 ( .A(n66972), .Y(n53496) );
  NAND2x1_ASAP7_75t_SL U49658 ( .A(n59506), .B(n57108), .Y(n67883) );
  XNOR2x1_ASAP7_75t_SL U49659 ( .A(n68072), .B(n68071), .Y(n58943) );
  BUFx2_ASAP7_75t_SL U49660 ( .A(n68037), .Y(n53497) );
  XNOR2xp5_ASAP7_75t_SL U49661 ( .A(n67782), .B(n59082), .Y(n68037) );
  XOR2x2_ASAP7_75t_SL U49662 ( .A(n59362), .B(n59363), .Y(n68294) );
  OAI21x1_ASAP7_75t_SL U49663 ( .A1(n59466), .A2(n59510), .B(n57717), .Y(
        n65061) );
  INVx4_ASAP7_75t_SL U49664 ( .A(n57709), .Y(n58884) );
  OAI22xp5_ASAP7_75t_SL U49665 ( .A1(n59238), .A2(n64920), .B1(n66711), .B2(
        n59460), .Y(n53498) );
  INVx1_ASAP7_75t_SL U49666 ( .A(n69139), .Y(n53499) );
  INVx1_ASAP7_75t_SL U49667 ( .A(n53499), .Y(n53500) );
  HB1xp67_ASAP7_75t_SL U49668 ( .A(n59433), .Y(n53501) );
  MAJx2_ASAP7_75t_SL U49669 ( .A(n68198), .B(n68194), .C(n68195), .Y(n53502)
         );
  XOR2x1_ASAP7_75t_SL U49670 ( .A(n57028), .B(n68114), .Y(n68195) );
  XOR2x2_ASAP7_75t_SL U49671 ( .A(n68549), .B(n68536), .Y(n58500) );
  HB1xp67_ASAP7_75t_SL U49672 ( .A(n68144), .Y(n53503) );
  INVx5_ASAP7_75t_SL U49673 ( .A(n59229), .Y(n59460) );
  XNOR2xp5_ASAP7_75t_SRAM U49674 ( .A(n68341), .B(n68344), .Y(n68293) );
  INVx1_ASAP7_75t_SL U49675 ( .A(n59243), .Y(n53504) );
  INVx1_ASAP7_75t_SL U49676 ( .A(n53504), .Y(n53505) );
  INVx1_ASAP7_75t_SL U49677 ( .A(n67739), .Y(n53506) );
  INVxp33_ASAP7_75t_SL U49678 ( .A(n64897), .Y(n53507) );
  NAND2xp5_ASAP7_75t_SL U49679 ( .A(n58851), .B(n53507), .Y(n59148) );
  NOR2x1_ASAP7_75t_SL U49680 ( .A(n53507), .B(n57311), .Y(n68377) );
  INVx1_ASAP7_75t_SL U49681 ( .A(n2508), .Y(n53508) );
  NOR2x1_ASAP7_75t_SL U49682 ( .A(n53508), .B(n59464), .Y(n59080) );
  INVxp33_ASAP7_75t_SL U49683 ( .A(n68720), .Y(n58371) );
  NAND2xp33_ASAP7_75t_SL U49684 ( .A(n68916), .B(n68717), .Y(n68720) );
  XNOR2x1_ASAP7_75t_SL U49685 ( .A(n67783), .B(n59083), .Y(n53509) );
  NAND2xp5_ASAP7_75t_SL U49686 ( .A(n68168), .B(n53510), .Y(n65029) );
  NAND2xp5_ASAP7_75t_SL U49687 ( .A(n53513), .B(n64898), .Y(n53510) );
  NOR2x1_ASAP7_75t_SL U49688 ( .A(n53512), .B(n53511), .Y(n64898) );
  INVx1_ASAP7_75t_SL U49689 ( .A(n58103), .Y(n53511) );
  INVx1_ASAP7_75t_SL U49690 ( .A(n65024), .Y(n53513) );
  NOR2xp33_ASAP7_75t_SL U49691 ( .A(n59505), .B(n59620), .Y(n63205) );
  NOR2x1_ASAP7_75t_SL U49692 ( .A(n59620), .B(n57179), .Y(n67412) );
  NOR2x1_ASAP7_75t_SL U49693 ( .A(n59620), .B(n59519), .Y(n68411) );
  INVx13_ASAP7_75t_SL U49694 ( .A(n75904), .Y(n59620) );
  AND2x6_ASAP7_75t_SL U49695 ( .A(n57811), .B(n59396), .Y(n75904) );
  XOR2x2_ASAP7_75t_SL U49696 ( .A(n57727), .B(n53514), .Y(n68202) );
  NAND2x2_ASAP7_75t_SL U49697 ( .A(n53587), .B(n53586), .Y(n53514) );
  NOR2x1_ASAP7_75t_SL U49698 ( .A(n67919), .B(n53514), .Y(n67929) );
  AOI21xp5_ASAP7_75t_SL U49699 ( .A1(n53514), .A2(n67919), .B(n53592), .Y(
        n67928) );
  XOR2x2_ASAP7_75t_SL U49700 ( .A(n53515), .B(n68292), .Y(n68342) );
  XNOR2xp5_ASAP7_75t_SL U49701 ( .A(n68302), .B(n68303), .Y(n53515) );
  MAJIxp5_ASAP7_75t_SL U49702 ( .A(n53516), .B(n68283), .C(n68282), .Y(n68303)
         );
  NOR2x1_ASAP7_75t_SL U49703 ( .A(n68287), .B(n58031), .Y(n68302) );
  XNOR2xp5_ASAP7_75t_SL U49704 ( .A(n68281), .B(n68280), .Y(n53516) );
  INVx1_ASAP7_75t_SL U49705 ( .A(n62748), .Y(n53519) );
  NAND2x2_ASAP7_75t_SL U49706 ( .A(n53518), .B(n62749), .Y(n57175) );
  OR2x2_ASAP7_75t_SL U49707 ( .A(n57644), .B(n53521), .Y(n62749) );
  OAI21x1_ASAP7_75t_SL U49708 ( .A1(n59553), .A2(n59591), .B(n53519), .Y(
        n53518) );
  BUFx6f_ASAP7_75t_SL U49709 ( .A(n57175), .Y(n53520) );
  INVx3_ASAP7_75t_SL U49710 ( .A(n57175), .Y(n67569) );
  INVx1_ASAP7_75t_SL U49711 ( .A(n57644), .Y(n62668) );
  INVxp67_ASAP7_75t_SL U49712 ( .A(n64389), .Y(n53521) );
  INVx1_ASAP7_75t_SL U49713 ( .A(n53522), .Y(n58692) );
  NOR2x1_ASAP7_75t_SL U49714 ( .A(n57289), .B(n53522), .Y(n68137) );
  OR2x2_ASAP7_75t_SL U49715 ( .A(n75107), .B(n53523), .Y(n58325) );
  OR2x2_ASAP7_75t_SL U49716 ( .A(n57130), .B(n53523), .Y(n58870) );
  NAND2xp5_ASAP7_75t_SL U49717 ( .A(n53524), .B(n58191), .Y(n58189) );
  NAND2xp5_ASAP7_75t_SL U49718 ( .A(n53525), .B(n59427), .Y(n53524) );
  NAND2xp5_ASAP7_75t_SL U49719 ( .A(n58190), .B(n58830), .Y(n53525) );
  OAI21xp5_ASAP7_75t_SL U49720 ( .A1(n53530), .A2(n68968), .B(n53526), .Y(
        n51993) );
  NOR3xp33_ASAP7_75t_SL U49721 ( .A(n58886), .B(n68978), .C(n53528), .Y(n53527) );
  INVx1_ASAP7_75t_SL U49722 ( .A(n53529), .Y(n53528) );
  INVx1_ASAP7_75t_SL U49723 ( .A(n53531), .Y(n53530) );
  NOR2x1_ASAP7_75t_SL U49724 ( .A(n68967), .B(n68966), .Y(n53531) );
  NAND2xp5_ASAP7_75t_SL U49725 ( .A(n53532), .B(n68140), .Y(n58218) );
  OAI21xp33_ASAP7_75t_SL U49726 ( .A1(n57774), .A2(n68140), .B(n53532), .Y(
        n68193) );
  NAND2x1_ASAP7_75t_SL U49727 ( .A(n58948), .B(n53623), .Y(n53532) );
  AND2x2_ASAP7_75t_SL U49728 ( .A(n1753), .B(n58717), .Y(n62571) );
  NAND2xp5_ASAP7_75t_SL U49729 ( .A(n62010), .B(n76678), .Y(n53533) );
  INVx1_ASAP7_75t_SL U49730 ( .A(n53536), .Y(n68473) );
  XOR2xp5_ASAP7_75t_SL U49731 ( .A(n53534), .B(n68478), .Y(n53536) );
  XNOR2xp5_ASAP7_75t_SL U49732 ( .A(n68477), .B(n68476), .Y(n53534) );
  MAJIxp5_ASAP7_75t_SL U49733 ( .A(n53536), .B(n68496), .C(n68495), .Y(n68523)
         );
  XNOR2xp5_ASAP7_75t_SL U49734 ( .A(n68457), .B(n53535), .Y(n68495) );
  XOR2xp5_ASAP7_75t_SL U49735 ( .A(n68456), .B(n68498), .Y(n53535) );
  XNOR2xp5_ASAP7_75t_SL U49736 ( .A(n58161), .B(n58159), .Y(n68456) );
  NAND2x1_ASAP7_75t_SL U49737 ( .A(n53538), .B(n53537), .Y(n67120) );
  OAI21xp5_ASAP7_75t_SL U49738 ( .A1(n53541), .A2(n67165), .B(n67168), .Y(
        n53537) );
  NAND2xp5_ASAP7_75t_SL U49739 ( .A(n53541), .B(n67165), .Y(n53538) );
  NAND2x1_ASAP7_75t_SL U49740 ( .A(n57615), .B(n57614), .Y(n57412) );
  XNOR2x1_ASAP7_75t_SL U49741 ( .A(n53539), .B(n67120), .Y(n57614) );
  XNOR2x1_ASAP7_75t_SL U49742 ( .A(n67118), .B(n53540), .Y(n53539) );
  XNOR2x2_ASAP7_75t_SL U49743 ( .A(n66504), .B(n66497), .Y(n67118) );
  INVx2_ASAP7_75t_SL U49744 ( .A(n67119), .Y(n53540) );
  INVx1_ASAP7_75t_SL U49745 ( .A(n67166), .Y(n53541) );
  XNOR2xp5_ASAP7_75t_SL U49746 ( .A(n53542), .B(n66591), .Y(n66600) );
  XOR2xp5_ASAP7_75t_SL U49747 ( .A(n53546), .B(n66589), .Y(n53542) );
  MAJIxp5_ASAP7_75t_SL U49748 ( .A(n66559), .B(n66557), .C(n66558), .Y(n66589)
         );
  OAI21xp5_ASAP7_75t_SL U49749 ( .A1(n66289), .A2(n59116), .B(n53543), .Y(
        n66558) );
  NAND2xp5_ASAP7_75t_SL U49750 ( .A(n53545), .B(n53544), .Y(n53543) );
  INVx1_ASAP7_75t_SL U49751 ( .A(n66561), .Y(n53544) );
  INVx1_ASAP7_75t_SL U49752 ( .A(n68119), .Y(n53545) );
  INVx1_ASAP7_75t_SL U49753 ( .A(n66590), .Y(n53546) );
  NOR2x1_ASAP7_75t_SL U49754 ( .A(n68903), .B(n53547), .Y(n68981) );
  OR2x2_ASAP7_75t_SL U49755 ( .A(n68727), .B(n68726), .Y(n53547) );
  INVx2_ASAP7_75t_SL U49756 ( .A(n68081), .Y(n67468) );
  INVx1_ASAP7_75t_SL U49757 ( .A(n67681), .Y(n67680) );
  OAI21xp5_ASAP7_75t_SL U49758 ( .A1(n53549), .A2(n67468), .B(n53548), .Y(
        n67681) );
  OAI21xp5_ASAP7_75t_SL U49759 ( .A1(n58672), .A2(n57241), .B(n67469), .Y(
        n53548) );
  NOR2x1_ASAP7_75t_SL U49760 ( .A(n53551), .B(n53550), .Y(n53549) );
  INVx1_ASAP7_75t_SL U49761 ( .A(n58412), .Y(n53550) );
  NOR2x1_ASAP7_75t_SL U49762 ( .A(n57108), .B(n53275), .Y(n53551) );
  A2O1A1Ixp33_ASAP7_75t_SL U49763 ( .A1(n58863), .A2(n57230), .B(n59038), .C(
        n53552), .Y(n59039) );
  OAI22xp33_ASAP7_75t_SL U49764 ( .A1(n67743), .A2(n67958), .B1(n53552), .B2(
        n57099), .Y(n65038) );
  INVx1_ASAP7_75t_SL U49765 ( .A(n64937), .Y(n53552) );
  XNOR2xp5_ASAP7_75t_SL U49766 ( .A(n59511), .B(n57525), .Y(n64937) );
  INVx2_ASAP7_75t_SL U49767 ( .A(n53553), .Y(n63177) );
  NAND3xp33_ASAP7_75t_SL U49768 ( .A(n58428), .B(n53553), .C(n57206), .Y(
        n57574) );
  NOR2x1p5_ASAP7_75t_SL U49769 ( .A(n57576), .B(n57575), .Y(n53553) );
  NOR2x1_ASAP7_75t_SL U49770 ( .A(n63177), .B(n53554), .Y(n61207) );
  INVx1_ASAP7_75t_SL U49771 ( .A(n58428), .Y(n53554) );
  NOR2x1_ASAP7_75t_SL U49772 ( .A(n59306), .B(n59305), .Y(n67501) );
  XNOR2x1_ASAP7_75t_SL U49773 ( .A(n53557), .B(n53555), .Y(n67391) );
  OAI21x1_ASAP7_75t_SL U49774 ( .A1(n67388), .A2(n59064), .B(n56959), .Y(
        n67505) );
  XOR2xp5_ASAP7_75t_SL U49775 ( .A(n67391), .B(n67399), .Y(n67392) );
  INVx1_ASAP7_75t_SL U49776 ( .A(n67503), .Y(n53556) );
  INVx1_ASAP7_75t_SL U49777 ( .A(n57001), .Y(n53557) );
  INVx1_ASAP7_75t_SL U49778 ( .A(n53558), .Y(n59217) );
  XNOR2xp5_ASAP7_75t_SL U49779 ( .A(n56998), .B(n57381), .Y(n53558) );
  XNOR2xp5_ASAP7_75t_SL U49780 ( .A(n59217), .B(n67990), .Y(n67991) );
  INVx2_ASAP7_75t_SL U49781 ( .A(or1200_cpu_or1200_except_ex_freeze_prev), .Y(
        n76673) );
  AO21x1_ASAP7_75t_SL U49782 ( .A1(n53563), .A2(n67882), .B(n53559), .Y(n68111) );
  OAI22xp5_ASAP7_75t_SL U49783 ( .A1(n53562), .A2(n67883), .B1(n68079), .B2(
        n53560), .Y(n53559) );
  INVx1_ASAP7_75t_SL U49784 ( .A(n53561), .Y(n53560) );
  NOR2x1_ASAP7_75t_SL U49785 ( .A(n59648), .B(n57108), .Y(n53561) );
  INVx1_ASAP7_75t_SL U49786 ( .A(n59648), .Y(n53562) );
  NOR2x1_ASAP7_75t_SL U49787 ( .A(n59506), .B(n57563), .Y(n67882) );
  INVx1_ASAP7_75t_SL U49788 ( .A(n67882), .Y(n57075) );
  NOR2x1_ASAP7_75t_SL U49789 ( .A(n68109), .B(n68111), .Y(n59037) );
  INVx1_ASAP7_75t_SL U49790 ( .A(n58093), .Y(n53563) );
  XNOR2x1_ASAP7_75t_SL U49791 ( .A(n53564), .B(n58153), .Y(n57541) );
  MAJx2_ASAP7_75t_SL U49792 ( .A(n68400), .B(n68401), .C(n68399), .Y(n58153)
         );
  INVx1_ASAP7_75t_SL U49793 ( .A(n68398), .Y(n53564) );
  OR2x2_ASAP7_75t_SL U49794 ( .A(n59314), .B(n53565), .Y(n58965) );
  NAND2xp5_ASAP7_75t_SL U49795 ( .A(n57651), .B(n57652), .Y(n53565) );
  OAI21xp5_ASAP7_75t_SL U49796 ( .A1(n59479), .A2(n53568), .B(n53566), .Y(
        n57924) );
  NAND2xp5_ASAP7_75t_SL U49797 ( .A(n53567), .B(n59479), .Y(n53566) );
  INVx1_ASAP7_75t_SL U49798 ( .A(n57128), .Y(n53567) );
  NAND2xp5_ASAP7_75t_SL U49799 ( .A(n57128), .B(n59588), .Y(n53568) );
  AOI22x1_ASAP7_75t_SL U49800 ( .A1(n53571), .A2(n53570), .B1(n53572), .B2(
        n53569), .Y(n68155) );
  INVx1_ASAP7_75t_SL U49801 ( .A(n65063), .Y(n53569) );
  NAND2xp5_ASAP7_75t_SL U49802 ( .A(n58851), .B(n57366), .Y(n53570) );
  NAND2xp5_ASAP7_75t_SL U49803 ( .A(n59659), .B(n67632), .Y(n53571) );
  XNOR2x1_ASAP7_75t_SL U49804 ( .A(n68153), .B(n68154), .Y(n53573) );
  AOI22x1_ASAP7_75t_SL U49805 ( .A1(n67842), .A2(n65061), .B1(n57380), .B2(
        n65062), .Y(n68154) );
  INVx1_ASAP7_75t_SL U49806 ( .A(n58991), .Y(n53572) );
  XNOR2xp5_ASAP7_75t_SL U49807 ( .A(n53574), .B(n68270), .Y(n65064) );
  XNOR2xp5_ASAP7_75t_SL U49808 ( .A(n53573), .B(n68155), .Y(n68270) );
  INVx1_ASAP7_75t_SL U49809 ( .A(n68269), .Y(n53574) );
  MAJIxp5_ASAP7_75t_SL U49810 ( .A(n65058), .B(n65057), .C(n65056), .Y(n68269)
         );
  OAI21xp5_ASAP7_75t_SL U49811 ( .A1(n53575), .A2(n64916), .B(n64915), .Y(
        n65058) );
  INVx1_ASAP7_75t_SL U49812 ( .A(n53576), .Y(n53575) );
  NAND2xp5_ASAP7_75t_SL U49813 ( .A(n57484), .B(n57065), .Y(n53576) );
  BUFx6f_ASAP7_75t_SL U49814 ( .A(n53582), .Y(n53577) );
  INVx2_ASAP7_75t_SL U49815 ( .A(n53582), .Y(n67948) );
  NAND3x2_ASAP7_75t_SL U49816 ( .A(n64032), .B(n63827), .C(n67586), .Y(n53582)
         );
  NOR2x1_ASAP7_75t_SL U49817 ( .A(n59511), .B(n53577), .Y(n59033) );
  NOR2x1_ASAP7_75t_SL U49818 ( .A(n75901), .B(n53577), .Y(n65015) );
  NAND2xp5_ASAP7_75t_SL U49819 ( .A(n67955), .B(n53577), .Y(n67954) );
  INVx1_ASAP7_75t_SL U49820 ( .A(n53578), .Y(n67848) );
  NOR2x1_ASAP7_75t_SL U49821 ( .A(n67948), .B(n53579), .Y(n53578) );
  INVx1_ASAP7_75t_SL U49822 ( .A(n57167), .Y(n53579) );
  NAND2xp5_ASAP7_75t_SL U49823 ( .A(n75903), .B(n53577), .Y(n58105) );
  NAND2xp5_ASAP7_75t_SL U49824 ( .A(n59651), .B(n53577), .Y(n58257) );
  OR2x2_ASAP7_75t_SL U49825 ( .A(n53580), .B(n67948), .Y(n68379) );
  INVx1_ASAP7_75t_SL U49826 ( .A(n58753), .Y(n53580) );
  NOR2x1_ASAP7_75t_SL U49827 ( .A(n53581), .B(n67948), .Y(n58525) );
  INVx1_ASAP7_75t_SL U49828 ( .A(n59668), .Y(n53581) );
  NAND2xp5_ASAP7_75t_SL U49829 ( .A(n59190), .B(n53577), .Y(n66880) );
  OAI21xp5_ASAP7_75t_SL U49830 ( .A1(n67288), .A2(n53613), .B(n53583), .Y(
        n64450) );
  NAND2xp5_ASAP7_75t_SL U49831 ( .A(n53584), .B(n67948), .Y(n53583) );
  INVx1_ASAP7_75t_SL U49832 ( .A(n58431), .Y(n53584) );
  NAND2xp5_ASAP7_75t_SL U49833 ( .A(n53585), .B(n58541), .Y(n68929) );
  NOR2x1_ASAP7_75t_SL U49834 ( .A(n68927), .B(n53585), .Y(n68910) );
  O2A1O1Ixp5_ASAP7_75t_SL U49835 ( .A1(n68981), .A2(n68905), .B(n58885), .C(
        n56205), .Y(n53585) );
  NAND2x1_ASAP7_75t_SL U49836 ( .A(n58025), .B(n57730), .Y(n53586) );
  NAND2xp5_ASAP7_75t_SL U49837 ( .A(n59171), .B(n67907), .Y(n53587) );
  NOR2x1_ASAP7_75t_SL U49838 ( .A(n67929), .B(n67928), .Y(n67983) );
  XNOR2x1_ASAP7_75t_SL U49839 ( .A(n57109), .B(n59647), .Y(n53588) );
  OAI22x1_ASAP7_75t_SL U49840 ( .A1(n59074), .A2(n59073), .B1(n67974), .B2(
        n53588), .Y(n67616) );
  A2O1A1Ixp33_ASAP7_75t_SL U49841 ( .A1(n75996), .A2(n75995), .B(n75994), .C(
        n75998), .Y(n76012) );
  NOR2x1_ASAP7_75t_SL U49842 ( .A(n59513), .B(n75921), .Y(n75989) );
  NOR2x1_ASAP7_75t_SL U49843 ( .A(n75920), .B(n75919), .Y(n75921) );
  AOI21xp5_ASAP7_75t_SL U49844 ( .A1(n67304), .A2(n58900), .B(n53589), .Y(
        n57800) );
  OAI21xp33_ASAP7_75t_SL U49845 ( .A1(n57104), .A2(n67302), .B(n67301), .Y(
        n53590) );
  O2A1O1Ixp5_ASAP7_75t_SL U49846 ( .A1(n57110), .A2(n67736), .B(n67299), .C(
        n68079), .Y(n53591) );
  INVx1_ASAP7_75t_SL U49847 ( .A(n67303), .Y(n58900) );
  AOI21xp5_ASAP7_75t_SL U49848 ( .A1(n67298), .A2(n59656), .B(n59638), .Y(
        n67304) );
  XNOR2xp5_ASAP7_75t_SL U49849 ( .A(n53592), .B(n57728), .Y(n57727) );
  NAND2xp5_ASAP7_75t_SL U49850 ( .A(n57729), .B(n59134), .Y(n53592) );
  AND2x2_ASAP7_75t_SL U49851 ( .A(n53475), .B(n53618), .Y(n67756) );
  AOI21x1_ASAP7_75t_SL U49852 ( .A1(n59245), .A2(n58648), .B(n66864), .Y(
        n53595) );
  NAND2xp5_ASAP7_75t_SL U49853 ( .A(n53594), .B(n53593), .Y(n66336) );
  NAND2xp5_ASAP7_75t_SL U49854 ( .A(n67743), .B(n53595), .Y(n53593) );
  INVx1_ASAP7_75t_SL U49855 ( .A(n66334), .Y(n53594) );
  OAI21xp5_ASAP7_75t_SL U49856 ( .A1(n53595), .A2(n67266), .B(n67265), .Y(
        n67352) );
  OAI21x1_ASAP7_75t_SL U49857 ( .A1(n58966), .A2(n67624), .B(n58967), .Y(
        n67652) );
  XNOR2xp5_ASAP7_75t_SL U49858 ( .A(n67654), .B(n53596), .Y(n67770) );
  XNOR2xp5_ASAP7_75t_SL U49859 ( .A(n53597), .B(n67652), .Y(n53596) );
  NAND2xp5_ASAP7_75t_SL U49860 ( .A(n58969), .B(n53598), .Y(n53597) );
  NAND2xp5_ASAP7_75t_SL U49861 ( .A(n67620), .B(n57033), .Y(n53598) );
  OR2x2_ASAP7_75t_SL U49862 ( .A(n67619), .B(n67618), .Y(n57033) );
  MAJIxp5_ASAP7_75t_SL U49863 ( .A(n67774), .B(n67773), .C(n53599), .Y(n67654)
         );
  INVx1_ASAP7_75t_SL U49864 ( .A(n67776), .Y(n53599) );
  NAND2xp5_ASAP7_75t_SL U49865 ( .A(n67436), .B(n67437), .Y(n67773) );
  NAND2xp5_ASAP7_75t_SL U49866 ( .A(n67433), .B(n57319), .Y(n67774) );
  OAI21xp5_ASAP7_75t_SL U49867 ( .A1(n59516), .A2(n59594), .B(n53600), .Y(
        n65054) );
  NAND2xp5_ASAP7_75t_SL U49868 ( .A(n59594), .B(n67741), .Y(n53600) );
  OAI22xp5_ASAP7_75t_SL U49869 ( .A1(n59594), .A2(n53602), .B1(n67741), .B2(
        n53601), .Y(n53605) );
  INVx1_ASAP7_75t_SL U49870 ( .A(n59594), .Y(n53601) );
  INVx1_ASAP7_75t_SL U49871 ( .A(n59516), .Y(n53602) );
  INVx2_ASAP7_75t_SL U49872 ( .A(n64607), .Y(n57097) );
  NAND2x2_ASAP7_75t_SL U49873 ( .A(n68011), .B(n58141), .Y(n64607) );
  NOR2xp67_ASAP7_75t_SL U49874 ( .A(n68102), .B(n68093), .Y(n53603) );
  OAI21x1_ASAP7_75t_SL U49875 ( .A1(n59594), .A2(n66800), .B(n53604), .Y(
        n68093) );
  NAND2x2_ASAP7_75t_SL U49876 ( .A(n59594), .B(n58753), .Y(n53604) );
  AND2x2_ASAP7_75t_SL U49877 ( .A(n59043), .B(n58718), .Y(n66800) );
  A2O1A1Ixp33_ASAP7_75t_SL U49878 ( .A1(n57277), .A2(n58275), .B(n67533), .C(
        n53606), .Y(n67692) );
  A2O1A1Ixp33_ASAP7_75t_SL U49879 ( .A1(n57484), .A2(n67532), .B(n53607), .C(
        n67531), .Y(n53606) );
  INVx1_ASAP7_75t_SL U49880 ( .A(n67530), .Y(n53607) );
  NAND2xp5_ASAP7_75t_SL U49881 ( .A(n59644), .B(n75930), .Y(n67530) );
  XNOR2x2_ASAP7_75t_SL U49882 ( .A(n66894), .B(n66990), .Y(n66895) );
  XNOR2x1_ASAP7_75t_SL U49883 ( .A(n66896), .B(n66895), .Y(n66985) );
  NOR2x1p5_ASAP7_75t_SL U49884 ( .A(n62723), .B(n62722), .Y(n67965) );
  NAND2x1_ASAP7_75t_SL U49885 ( .A(n68015), .B(n59619), .Y(n68023) );
  AND3x4_ASAP7_75t_SL U49886 ( .A(n57960), .B(n59555), .C(n59571), .Y(n62589)
         );
  AND2x2_ASAP7_75t_SL U49887 ( .A(n67227), .B(n59518), .Y(n59399) );
  NOR2x2_ASAP7_75t_SL U49888 ( .A(n59348), .B(n59349), .Y(n75642) );
  INVx1_ASAP7_75t_SL U49889 ( .A(n75642), .Y(n59643) );
  OAI21x1_ASAP7_75t_SL U49890 ( .A1(n66966), .A2(n66747), .B(n66746), .Y(
        n66779) );
  INVx1_ASAP7_75t_SL U49891 ( .A(n66968), .Y(n66747) );
  NOR2x1_ASAP7_75t_SL U49892 ( .A(n57347), .B(n58944), .Y(n67605) );
  NAND2x1_ASAP7_75t_SL U49893 ( .A(n68737), .B(n59433), .Y(n58728) );
  XOR2x1_ASAP7_75t_SL U49894 ( .A(n57525), .B(n67228), .Y(n67970) );
  INVx2_ASAP7_75t_SL U49895 ( .A(n57569), .Y(n58137) );
  AND2x2_ASAP7_75t_SL U49896 ( .A(n58190), .B(n58830), .Y(n53608) );
  NAND2x1_ASAP7_75t_SL U49897 ( .A(n53609), .B(n53610), .Y(n53611) );
  NAND2xp5_ASAP7_75t_SL U49898 ( .A(n53611), .B(n66312), .Y(n66309) );
  INVx1_ASAP7_75t_SL U49899 ( .A(n66306), .Y(n53609) );
  INVx1_ASAP7_75t_SL U49900 ( .A(n66305), .Y(n53610) );
  INVx1_ASAP7_75t_SL U49901 ( .A(n66304), .Y(n66306) );
  NAND2xp5_ASAP7_75t_SL U49902 ( .A(n59165), .B(n64609), .Y(n53612) );
  NAND2xp5_ASAP7_75t_SL U49903 ( .A(n59165), .B(n64609), .Y(n53613) );
  XNOR2x1_ASAP7_75t_SL U49904 ( .A(n53497), .B(n57582), .Y(n68062) );
  XNOR2x1_ASAP7_75t_SL U49905 ( .A(n57461), .B(n68036), .Y(n57582) );
  NAND2xp5_ASAP7_75t_SL U49906 ( .A(n59165), .B(n64609), .Y(n67562) );
  NAND2xp5_ASAP7_75t_SL U49907 ( .A(n66241), .B(n66242), .Y(n53614) );
  NAND2x1p5_ASAP7_75t_SL U49908 ( .A(n66241), .B(n66242), .Y(n78167) );
  NAND2x1_ASAP7_75t_SL U49909 ( .A(n62615), .B(n58277), .Y(n59235) );
  AOI21x1_ASAP7_75t_SL U49910 ( .A1(n68735), .A2(n68338), .B(n68337), .Y(
        n68723) );
  OAI21x1_ASAP7_75t_SL U49911 ( .A1(n64947), .A2(n64946), .B(n64945), .Y(
        n64979) );
  BUFx2_ASAP7_75t_SL U49912 ( .A(n65000), .Y(n57489) );
  XNOR2x2_ASAP7_75t_SL U49913 ( .A(n63198), .B(n58876), .Y(n63162) );
  AOI21x1_ASAP7_75t_SL U49914 ( .A1(n67375), .A2(n67376), .B(n67374), .Y(
        n67614) );
  INVx1_ASAP7_75t_SL U49915 ( .A(n67237), .Y(n67536) );
  NOR2x2_ASAP7_75t_SL U49916 ( .A(n67237), .B(n57941), .Y(n67463) );
  NOR2x1_ASAP7_75t_SL U49917 ( .A(n64568), .B(n64567), .Y(n64518) );
  INVx2_ASAP7_75t_SL U49918 ( .A(n64569), .Y(n64567) );
  NAND2xp5_ASAP7_75t_SL U49919 ( .A(n59657), .B(n64567), .Y(n64478) );
  NOR2x1_ASAP7_75t_SL U49920 ( .A(n59462), .B(n60623), .Y(n75477) );
  NOR2x1p5_ASAP7_75t_SL U49921 ( .A(n67395), .B(n67394), .Y(n57832) );
  BUFx2_ASAP7_75t_SL U49922 ( .A(n68054), .Y(n59176) );
  NOR2x1p5_ASAP7_75t_SL U49923 ( .A(n58644), .B(n58643), .Y(n67817) );
  INVx6_ASAP7_75t_SL U49924 ( .A(n59606), .Y(n59466) );
  NAND2x1p5_ASAP7_75t_SL U49925 ( .A(n68756), .B(n68754), .Y(n57869) );
  NAND2x1_ASAP7_75t_SL U49926 ( .A(n65038), .B(n65039), .Y(n68128) );
  NOR2x1p5_ASAP7_75t_SL U49927 ( .A(n58756), .B(n64633), .Y(n64884) );
  NOR2x1_ASAP7_75t_SL U49928 ( .A(n64589), .B(n64588), .Y(n58995) );
  XNOR2x2_ASAP7_75t_SL U49929 ( .A(n64638), .B(n57378), .Y(n64589) );
  INVx8_ASAP7_75t_SL U49930 ( .A(n67365), .Y(n75962) );
  AOI22xp5_ASAP7_75t_SL U49931 ( .A1(n68409), .A2(n67365), .B1(n57260), .B2(
        n66568), .Y(n66552) );
  OR2x6_ASAP7_75t_SL U49932 ( .A(n66287), .B(n66286), .Y(n67365) );
  INVx2_ASAP7_75t_SL U49933 ( .A(n66244), .Y(n53615) );
  INVx1_ASAP7_75t_SL U49934 ( .A(n66244), .Y(n63814) );
  INVx1_ASAP7_75t_SL U49935 ( .A(n56141), .Y(n53616) );
  INVx1_ASAP7_75t_SL U49936 ( .A(n59300), .Y(n56141) );
  HB1xp67_ASAP7_75t_SL U49937 ( .A(n59256), .Y(n53617) );
  NOR2x1p5_ASAP7_75t_SL U49938 ( .A(n56955), .B(n56954), .Y(n59256) );
  INVx1_ASAP7_75t_SL U49939 ( .A(n59589), .Y(n57629) );
  INVx1_ASAP7_75t_SL U49940 ( .A(n59318), .Y(n53618) );
  OAI22xp5_ASAP7_75t_SL U49941 ( .A1(n67415), .A2(n67414), .B1(n67413), .B2(
        n59042), .Y(n53619) );
  AOI21xp5_ASAP7_75t_SL U49942 ( .A1(n59620), .A2(n59517), .B(n67412), .Y(
        n67415) );
  NAND2xp5_ASAP7_75t_SL U49943 ( .A(n58383), .B(n76049), .Y(n57702) );
  INVx4_ASAP7_75t_SL U49944 ( .A(n67845), .Y(n68383) );
  INVx4_ASAP7_75t_SL U49945 ( .A(n67228), .Y(n75922) );
  NOR2x1_ASAP7_75t_SL U49946 ( .A(n59576), .B(n66257), .Y(n66259) );
  NOR2x1p5_ASAP7_75t_SL U49947 ( .A(n57912), .B(n67151), .Y(n67242) );
  INVx5_ASAP7_75t_SL U49948 ( .A(n59314), .Y(n59613) );
  NAND2x2_ASAP7_75t_SL U49949 ( .A(n67636), .B(n59599), .Y(n67151) );
  NAND2x1_ASAP7_75t_SL U49950 ( .A(n68853), .B(n68718), .Y(n68578) );
  OAI21xp33_ASAP7_75t_SRAM U49951 ( .A1(n58433), .A2(n66298), .B(n66297), .Y(
        n67604) );
  INVx5_ASAP7_75t_SL U49952 ( .A(n58433), .Y(n57186) );
  NAND2x1_ASAP7_75t_SL U49953 ( .A(n77735), .B(n58433), .Y(n66375) );
  AND2x4_ASAP7_75t_SL U49954 ( .A(n59470), .B(n59507), .Y(n62648) );
  OAI22x1_ASAP7_75t_SL U49955 ( .A1(n59037), .A2(n58713), .B1(n59035), .B2(
        n68113), .Y(n59036) );
  NAND2x1_ASAP7_75t_SL U49956 ( .A(n59448), .B(n64651), .Y(n59144) );
  INVx5_ASAP7_75t_SL U49957 ( .A(n58786), .Y(n59448) );
  OR2x2_ASAP7_75t_SL U49958 ( .A(n59042), .B(n59002), .Y(n53620) );
  NAND2x1p5_ASAP7_75t_SL U49959 ( .A(n53620), .B(n59430), .Y(n65024) );
  XOR2x2_ASAP7_75t_SL U49960 ( .A(n67227), .B(n59607), .Y(n59002) );
  NAND2x1_ASAP7_75t_SL U49961 ( .A(n59003), .B(n65024), .Y(n68168) );
  NAND2xp67_ASAP7_75t_SRAM U49962 ( .A(n53280), .B(n67364), .Y(n63115) );
  XNOR2x1_ASAP7_75t_SL U49963 ( .A(n63609), .B(n63605), .Y(n63241) );
  XOR2x2_ASAP7_75t_SL U49964 ( .A(n63643), .B(n63642), .Y(n63605) );
  INVx1_ASAP7_75t_SL U49965 ( .A(n65072), .Y(n59291) );
  NOR2x1_ASAP7_75t_SL U49966 ( .A(n65072), .B(n57184), .Y(n58789) );
  XNOR2x1_ASAP7_75t_SL U49967 ( .A(n64519), .B(n64584), .Y(n64588) );
  XNOR2xp5_ASAP7_75t_SL U49968 ( .A(n58953), .B(n67033), .Y(n58459) );
  XNOR2x1_ASAP7_75t_SL U49969 ( .A(n58951), .B(n67034), .Y(n58953) );
  NAND2x1p5_ASAP7_75t_SL U49970 ( .A(n58021), .B(n67634), .Y(n66373) );
  INVx2_ASAP7_75t_SL U49971 ( .A(n59448), .Y(n58021) );
  MAJIxp5_ASAP7_75t_SL U49972 ( .A(n68330), .B(n57420), .C(n58918), .Y(n53622)
         );
  XNOR2xp5_ASAP7_75t_SL U49973 ( .A(n57741), .B(n57740), .Y(n53623) );
  XOR2x2_ASAP7_75t_SL U49974 ( .A(n68137), .B(n68138), .Y(n57740) );
  NAND2xp5_ASAP7_75t_SL U49975 ( .A(n63181), .B(n59400), .Y(n53624) );
  INVx1_ASAP7_75t_SL U49976 ( .A(n58219), .Y(n53625) );
  NAND2x1_ASAP7_75t_SL U49977 ( .A(n63181), .B(n59400), .Y(n59339) );
  INVx1_ASAP7_75t_SL U49978 ( .A(n68974), .Y(n58219) );
  NOR2x1_ASAP7_75t_SL U49979 ( .A(n58543), .B(n69160), .Y(n58868) );
  XNOR2x2_ASAP7_75t_SL U49980 ( .A(n67835), .B(n58255), .Y(n67934) );
  NOR2x1_ASAP7_75t_SL U49981 ( .A(n60445), .B(n60444), .Y(n77364) );
  INVx1_ASAP7_75t_SL U49982 ( .A(n60468), .Y(n60444) );
  NAND2xp5_ASAP7_75t_SL U49983 ( .A(n61044), .B(n61040), .Y(n60445) );
  NOR2x1_ASAP7_75t_SL U49984 ( .A(n61293), .B(n60210), .Y(n60214) );
  NOR2x1_ASAP7_75t_SL U49985 ( .A(n59849), .B(n59848), .Y(n75427) );
  NOR2x1_ASAP7_75t_SL U49986 ( .A(n59847), .B(n75777), .Y(n59848) );
  AOI31xp67_ASAP7_75t_SL U49987 ( .A1(n69363), .A2(n69364), .A3(n59873), .B(
        n59872), .Y(n75671) );
  XNOR2xp5_ASAP7_75t_SRAM U49988 ( .A(n59461), .B(n68335), .Y(n68228) );
  NAND2x1p5_ASAP7_75t_SL U49989 ( .A(n66253), .B(n66258), .Y(n57556) );
  XNOR2xp5_ASAP7_75t_SL U49990 ( .A(n53626), .B(n68145), .Y(n68827) );
  XNOR2xp5_ASAP7_75t_SL U49991 ( .A(n68143), .B(n68144), .Y(n53626) );
  NAND2x1p5_ASAP7_75t_SL U49992 ( .A(n68902), .B(n68736), .Y(n68560) );
  INVx4_ASAP7_75t_SL U49993 ( .A(n67421), .Y(n67424) );
  NAND2x2_ASAP7_75t_SL U49994 ( .A(n58458), .B(n59361), .Y(n67421) );
  NAND3x1_ASAP7_75t_SL U49995 ( .A(n57790), .B(n57789), .C(n61965), .Y(n66297)
         );
  OAI21x1_ASAP7_75t_SL U49996 ( .A1(n58519), .A2(n67261), .B(n67260), .Y(
        n67351) );
  NAND2x1_ASAP7_75t_SL U49997 ( .A(n62601), .B(n62600), .Y(n67610) );
  INVx5_ASAP7_75t_SL U49998 ( .A(n59649), .Y(n59647) );
  XNOR2x2_ASAP7_75t_SL U49999 ( .A(n53498), .B(n66652), .Y(n66774) );
  INVx1_ASAP7_75t_SL U50000 ( .A(n57567), .Y(n53627) );
  NOR2x1_ASAP7_75t_SL U50001 ( .A(n66248), .B(n76430), .Y(n67422) );
  NAND2x1p5_ASAP7_75t_SL U50002 ( .A(n65113), .B(n65115), .Y(n68736) );
  NOR2x1_ASAP7_75t_SL U50003 ( .A(n63102), .B(n63101), .Y(n63498) );
  NOR2x1_ASAP7_75t_SL U50004 ( .A(n63243), .B(n63498), .Y(n63883) );
  NOR2x1_ASAP7_75t_SL U50005 ( .A(n70707), .B(n70706), .Y(n70896) );
  NOR2x1_ASAP7_75t_SL U50006 ( .A(n70691), .B(n59524), .Y(n70706) );
  NOR2x1_ASAP7_75t_SL U50007 ( .A(n70871), .B(n70870), .Y(n70906) );
  NAND2x1p5_ASAP7_75t_SL U50008 ( .A(n58302), .B(n58372), .Y(n59524) );
  NAND2x1p5_ASAP7_75t_SL U50009 ( .A(n58221), .B(n57118), .Y(n58220) );
  INVx2_ASAP7_75t_SL U50010 ( .A(n62589), .Y(n62646) );
  INVx2_ASAP7_75t_SL U50011 ( .A(n67274), .Y(n57854) );
  NOR2x1p5_ASAP7_75t_SL U50012 ( .A(n61157), .B(n58146), .Y(n76677) );
  INVx2_ASAP7_75t_SL U50013 ( .A(or1200_cpu_or1200_except_n690), .Y(n61157) );
  AOI31xp67_ASAP7_75t_SL U50014 ( .A1(n63403), .A2(n63402), .A3(n63401), .B(
        n63400), .Y(n63428) );
  NOR2x1_ASAP7_75t_SL U50015 ( .A(or1200_cpu_or1200_mult_mac_n287), .B(n63270), 
        .Y(n63274) );
  INVx2_ASAP7_75t_SL U50016 ( .A(or1200_cpu_or1200_mult_mac_n141), .Y(n63270)
         );
  NOR2x1p5_ASAP7_75t_SL U50017 ( .A(n63429), .B(n63428), .Y(n63782) );
  NOR2x1_ASAP7_75t_SL U50018 ( .A(n70606), .B(n70605), .Y(n70607) );
  NOR2x1_ASAP7_75t_SL U50019 ( .A(n70592), .B(n70586), .Y(n70603) );
  NOR2x1p5_ASAP7_75t_SL U50020 ( .A(DP_OP_742J1_130_9702_n59), .B(n74457), .Y(
        n70600) );
  NAND2x1p5_ASAP7_75t_SL U50021 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_25_), .B(
        n74458), .Y(n74457) );
  NAND2x1p5_ASAP7_75t_SL U50022 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_11_), .B(
        n74324), .Y(n74337) );
  NOR2x1p5_ASAP7_75t_SL U50023 ( .A(n74318), .B(n74319), .Y(n74324) );
  NOR2x1p5_ASAP7_75t_SL U50024 ( .A(n74448), .B(n74449), .Y(n74458) );
  NAND2x1p5_ASAP7_75t_SL U50025 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_9_), .B(
        n74353), .Y(n74319) );
  NOR2x2_ASAP7_75t_SL U50026 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39), .B(n74466), .Y(n74465) );
  NAND2x1p5_ASAP7_75t_SL U50027 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_45_), .B(
        n74450), .Y(n74466) );
  NAND2x1p5_ASAP7_75t_SL U50028 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_41_), .B(
        n74424), .Y(n74433) );
  NOR2x1p5_ASAP7_75t_SL U50029 ( .A(n74414), .B(n74415), .Y(n74424) );
  AOI22xp5_ASAP7_75t_SL U50030 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_4_), .A2(
        n72549), .B1(n72565), .B2(n72548), .Y(n74292) );
  NAND2x1p5_ASAP7_75t_SL U50031 ( .A(n72534), .B(n72533), .Y(n72547) );
  NOR2x2_ASAP7_75t_SL U50032 ( .A(n74265), .B(n57203), .Y(n72533) );
  NOR2x1_ASAP7_75t_SL U50033 ( .A(n74314), .B(n74315), .Y(n74320) );
  NAND2x1p5_ASAP7_75t_SL U50034 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_29_), .B(
        n74355), .Y(n74315) );
  NOR2x1p5_ASAP7_75t_SL U50035 ( .A(n74356), .B(n74370), .Y(n74355) );
  NAND2x1p5_ASAP7_75t_SL U50036 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_27_), .B(
        n74371), .Y(n74370) );
  NOR2xp33_ASAP7_75t_SL U50037 ( .A(n57111), .B(n59065), .Y(n58131) );
  XNOR2xp5_ASAP7_75t_SL U50038 ( .A(n59504), .B(n58865), .Y(n67869) );
  OAI21xp5_ASAP7_75t_SL U50039 ( .A1(n67872), .A2(n68119), .B(n67873), .Y(
        n57936) );
  NOR2xp33_ASAP7_75t_SL U50040 ( .A(n67861), .B(n57904), .Y(n58914) );
  INVx1_ASAP7_75t_SL U50041 ( .A(n67528), .Y(n57929) );
  INVx1_ASAP7_75t_SL U50042 ( .A(n67275), .Y(n57943) );
  NOR2xp33_ASAP7_75t_SL U50043 ( .A(n66481), .B(n57165), .Y(n57885) );
  AO21x1_ASAP7_75t_SL U50044 ( .A1(n59012), .A2(n57735), .B(n57734), .Y(n63090) );
  BUFx3_ASAP7_75t_SL U50045 ( .A(n64625), .Y(n57900) );
  NAND2xp5_ASAP7_75t_SL U50046 ( .A(n63122), .B(n57706), .Y(n57705) );
  XNOR2xp5_ASAP7_75t_SL U50047 ( .A(n63820), .B(n64678), .Y(n63821) );
  INVx1_ASAP7_75t_SL U50048 ( .A(n64619), .Y(n58240) );
  BUFx2_ASAP7_75t_SL U50049 ( .A(n64617), .Y(n57424) );
  INVx1_ASAP7_75t_SL U50050 ( .A(n67628), .Y(n57669) );
  XNOR2xp5_ASAP7_75t_SL U50051 ( .A(n57109), .B(n75895), .Y(n67907) );
  OAI22xp5_ASAP7_75t_SL U50052 ( .A1(n67383), .A2(n57485), .B1(n53342), .B2(
        n67467), .Y(n67628) );
  HB1xp67_ASAP7_75t_SL U50053 ( .A(n67986), .Y(n57235) );
  INVx1_ASAP7_75t_SL U50054 ( .A(n67593), .Y(n59277) );
  NOR2xp33_ASAP7_75t_SL U50055 ( .A(n59603), .B(n67408), .Y(n58261) );
  NOR2xp33_ASAP7_75t_SL U50056 ( .A(n59659), .B(n57505), .Y(n57690) );
  BUFx2_ASAP7_75t_SL U50057 ( .A(n67130), .Y(n58333) );
  BUFx2_ASAP7_75t_SL U50058 ( .A(n68017), .Y(n57375) );
  NOR2xp33_ASAP7_75t_SL U50059 ( .A(n64035), .B(n58903), .Y(n57759) );
  NAND2x1p5_ASAP7_75t_SL U50060 ( .A(n59657), .B(n57414), .Y(n63818) );
  INVx1_ASAP7_75t_SL U50061 ( .A(n57225), .Y(n57224) );
  NOR2xp33_ASAP7_75t_SL U50062 ( .A(n53275), .B(n67234), .Y(n67236) );
  INVx1_ASAP7_75t_SL U50063 ( .A(n66667), .Y(n59238) );
  NOR2xp33_ASAP7_75t_SL U50064 ( .A(n66456), .B(n59636), .Y(n66457) );
  OAI22xp5_ASAP7_75t_SL U50065 ( .A1(n53271), .A2(n58016), .B1(n76176), .B2(
        n59600), .Y(n66481) );
  NAND2xp5_ASAP7_75t_SL U50066 ( .A(n67481), .B(n67963), .Y(n66782) );
  OAI21xp5_ASAP7_75t_SL U50067 ( .A1(n63840), .A2(n58961), .B(n59619), .Y(
        n58179) );
  XNOR2xp5_ASAP7_75t_SL U50068 ( .A(n59381), .B(n68098), .Y(n64408) );
  INVx1_ASAP7_75t_SL U50069 ( .A(n67242), .Y(n57667) );
  BUFx2_ASAP7_75t_SL U50070 ( .A(n67864), .Y(n57422) );
  INVx1_ASAP7_75t_SL U50071 ( .A(n63055), .Y(n57708) );
  NOR2x1_ASAP7_75t_SL U50072 ( .A(n58995), .B(n58993), .Y(n64909) );
  OAI21xp5_ASAP7_75t_SL U50073 ( .A1(n68031), .A2(n68030), .B(n68029), .Y(
        n68064) );
  NOR2x1_ASAP7_75t_SL U50074 ( .A(n58206), .B(n63177), .Y(n60914) );
  OAI21xp5_ASAP7_75t_SL U50075 ( .A1(n57362), .A2(n64628), .B(n64627), .Y(
        n64962) );
  BUFx3_ASAP7_75t_SL U50076 ( .A(n67845), .Y(n57380) );
  BUFx6f_ASAP7_75t_SL U50077 ( .A(n58397), .Y(n57414) );
  OAI21xp5_ASAP7_75t_SL U50078 ( .A1(n68079), .A2(n68021), .B(n68020), .Y(
        n68076) );
  NAND2x1_ASAP7_75t_SL U50079 ( .A(n67402), .B(n67401), .Y(n58747) );
  NAND2xp5_ASAP7_75t_SL U50080 ( .A(n58397), .B(n64611), .Y(n57910) );
  NOR2x1_ASAP7_75t_SL U50081 ( .A(n63661), .B(n63669), .Y(n63175) );
  XNOR2xp5_ASAP7_75t_SL U50082 ( .A(n63869), .B(n64062), .Y(n63870) );
  XNOR2xp5_ASAP7_75t_SL U50083 ( .A(n63848), .B(n63847), .Y(n64021) );
  HB1xp67_ASAP7_75t_SL U50084 ( .A(n65067), .Y(n57290) );
  NOR2x1_ASAP7_75t_SL U50085 ( .A(n65005), .B(n65004), .Y(n68221) );
  NAND2xp5_ASAP7_75t_SL U50086 ( .A(n67920), .B(n59607), .Y(n57605) );
  NOR2x1_ASAP7_75t_SL U50087 ( .A(n59607), .B(n75927), .Y(n58776) );
  NAND2xp5_ASAP7_75t_SL U50088 ( .A(n59284), .B(n68156), .Y(n58652) );
  NAND2xp5_ASAP7_75t_SL U50089 ( .A(n67906), .B(n67249), .Y(n59376) );
  INVx1_ASAP7_75t_SL U50090 ( .A(n59353), .Y(n64513) );
  AO21x1_ASAP7_75t_SL U50091 ( .A1(n58185), .A2(n63049), .B(n58184), .Y(n63104) );
  HB1xp67_ASAP7_75t_SL U50092 ( .A(n69004), .Y(n57475) );
  NAND2x1_ASAP7_75t_SL U50093 ( .A(n67110), .B(n67109), .Y(n69148) );
  NAND2xp5_ASAP7_75t_SL U50094 ( .A(n57248), .B(n57247), .Y(n67603) );
  OAI21xp5_ASAP7_75t_SL U50095 ( .A1(n59664), .A2(n67601), .B(n67600), .Y(
        n57248) );
  NAND2x1p5_ASAP7_75t_SL U50096 ( .A(n59711), .B(n59707), .Y(n60747) );
  BUFx3_ASAP7_75t_SL U50097 ( .A(n61909), .Y(n57466) );
  NOR2x1_ASAP7_75t_SL U50098 ( .A(n53481), .B(n68327), .Y(n68740) );
  OAI21xp5_ASAP7_75t_SL U50099 ( .A1(n58383), .A2(n59510), .B(n57702), .Y(
        n67438) );
  INVx1_ASAP7_75t_SL U50100 ( .A(n63675), .Y(n56863) );
  XNOR2xp5_ASAP7_75t_SL U50101 ( .A(n58402), .B(n59504), .Y(n64445) );
  INVx2_ASAP7_75t_SL U50102 ( .A(n58884), .Y(n58755) );
  NAND2x1_ASAP7_75t_SL U50103 ( .A(n68086), .B(n57669), .Y(n57670) );
  NAND2xp5_ASAP7_75t_SL U50104 ( .A(n59452), .B(n67907), .Y(n57998) );
  NAND2xp5_ASAP7_75t_SL U50105 ( .A(n58891), .B(n57438), .Y(n58890) );
  AOI22xp5_ASAP7_75t_SL U50106 ( .A1(n59670), .A2(n67428), .B1(n59476), .B2(
        n67621), .Y(n67642) );
  INVx1_ASAP7_75t_SL U50107 ( .A(n67682), .Y(n58271) );
  XNOR2xp5_ASAP7_75t_SL U50108 ( .A(n59030), .B(n59029), .Y(n59031) );
  NOR2xp33_ASAP7_75t_SL U50109 ( .A(n58851), .B(n58148), .Y(n59146) );
  AOI22xp5_ASAP7_75t_SL U50110 ( .A1(n67078), .A2(n67446), .B1(n59447), .B2(
        n66474), .Y(n67122) );
  HB1xp67_ASAP7_75t_SL U50111 ( .A(n67962), .Y(n57244) );
  XNOR2xp5_ASAP7_75t_SL U50112 ( .A(n64579), .B(n64580), .Y(n64584) );
  NOR2xp33_ASAP7_75t_SL U50113 ( .A(n58919), .B(n57366), .Y(n58163) );
  HB1xp67_ASAP7_75t_SL U50114 ( .A(n56830), .Y(n57329) );
  NAND2xp5_ASAP7_75t_SL U50115 ( .A(n68002), .B(n59613), .Y(n57872) );
  INVx1_ASAP7_75t_SL U50116 ( .A(n67401), .Y(n57873) );
  NOR2xp33_ASAP7_75t_SL U50117 ( .A(n67998), .B(n68000), .Y(n57954) );
  INVx1_ASAP7_75t_SL U50118 ( .A(n67999), .Y(n57953) );
  INVx1_ASAP7_75t_SL U50119 ( .A(n68368), .Y(n57618) );
  NOR2xp33_ASAP7_75t_SL U50120 ( .A(n57912), .B(n67467), .Y(n57911) );
  AOI22xp5_ASAP7_75t_SL U50121 ( .A1(n67306), .A2(n67031), .B1(n57161), .B2(
        n67032), .Y(n67068) );
  NOR2xp33_ASAP7_75t_SL U50122 ( .A(n59614), .B(n67432), .Y(n64397) );
  NOR2x1_ASAP7_75t_SL U50123 ( .A(n58514), .B(n59596), .Y(n58660) );
  NAND2xp5_ASAP7_75t_SL U50124 ( .A(n57662), .B(n59468), .Y(n59359) );
  NOR2x1_ASAP7_75t_SL U50125 ( .A(n64369), .B(n58658), .Y(n57499) );
  BUFx2_ASAP7_75t_SL U50126 ( .A(n67151), .Y(n57242) );
  OAI21xp5_ASAP7_75t_SL U50127 ( .A1(n64883), .A2(n64882), .B(n64881), .Y(
        n65049) );
  NAND2xp5_ASAP7_75t_SL U50128 ( .A(n57265), .B(n57861), .Y(n67885) );
  XOR2xp5_ASAP7_75t_SL U50129 ( .A(n67788), .B(n57725), .Y(n68040) );
  NOR2xp33_ASAP7_75t_SL U50130 ( .A(n58711), .B(n67706), .Y(n66629) );
  HB1xp67_ASAP7_75t_SL U50131 ( .A(n68442), .Y(n57220) );
  NOR2x1_ASAP7_75t_SL U50132 ( .A(n57493), .B(n58452), .Y(n68239) );
  AOI22xp5_ASAP7_75t_SL U50133 ( .A1(n59670), .A2(n66863), .B1(n64567), .B2(
        n58634), .Y(n58633) );
  HB1xp67_ASAP7_75t_SL U50134 ( .A(n58406), .Y(n57441) );
  OAI21xp5_ASAP7_75t_SL U50135 ( .A1(n64393), .A2(n58356), .B(n64392), .Y(
        n64540) );
  NOR2x1_ASAP7_75t_SL U50136 ( .A(n62806), .B(n57538), .Y(n64966) );
  BUFx2_ASAP7_75t_SL U50137 ( .A(n67951), .Y(n57359) );
  NOR2x1p5_ASAP7_75t_SL U50138 ( .A(n67971), .B(n58931), .Y(n58026) );
  INVx2_ASAP7_75t_SL U50139 ( .A(n59616), .Y(n57516) );
  XNOR2xp5_ASAP7_75t_SL U50140 ( .A(n67115), .B(n67114), .Y(n67116) );
  NAND2xp5_ASAP7_75t_SL U50141 ( .A(n66758), .B(n67428), .Y(n64572) );
  NOR2xp33_ASAP7_75t_SL U50142 ( .A(n62699), .B(n59515), .Y(n62691) );
  NAND2xp5_ASAP7_75t_SL U50143 ( .A(n62750), .B(n57358), .Y(n57707) );
  HB1xp67_ASAP7_75t_SL U50144 ( .A(n68052), .Y(n57305) );
  XNOR2xp5_ASAP7_75t_SL U50145 ( .A(n66909), .B(n66908), .Y(n58721) );
  XNOR2xp5_ASAP7_75t_SL U50146 ( .A(n66777), .B(n66776), .Y(n68548) );
  INVx1_ASAP7_75t_SL U50147 ( .A(n59594), .Y(n57630) );
  AOI21xp5_ASAP7_75t_SL U50148 ( .A1(n64408), .A2(n58802), .B(n64407), .Y(
        n64598) );
  XNOR2xp5_ASAP7_75t_SL U50149 ( .A(n57109), .B(n57107), .Y(n68084) );
  HB1xp67_ASAP7_75t_SL U50150 ( .A(n68171), .Y(n57231) );
  NAND2xp5_ASAP7_75t_SL U50151 ( .A(n59190), .B(n67883), .Y(n59189) );
  NAND2xp5_ASAP7_75t_SL U50152 ( .A(n76049), .B(n59607), .Y(n66917) );
  NOR2xp33_ASAP7_75t_SL U50153 ( .A(n57219), .B(n59387), .Y(n57593) );
  BUFx2_ASAP7_75t_SL U50154 ( .A(n57799), .Y(n57798) );
  NAND2xp5_ASAP7_75t_SL U50155 ( .A(n57384), .B(n57383), .Y(n58461) );
  XOR2xp5_ASAP7_75t_SL U50156 ( .A(n63629), .B(n63195), .Y(n63643) );
  HB1xp67_ASAP7_75t_SL U50157 ( .A(n68901), .Y(n57481) );
  INVx2_ASAP7_75t_SL U50158 ( .A(n56947), .Y(n75275) );
  NOR2xp33_ASAP7_75t_SL U50159 ( .A(n59561), .B(n58496), .Y(n58241) );
  INVx1_ASAP7_75t_SL U50160 ( .A(n60914), .Y(n60596) );
  NAND2xp5_ASAP7_75t_SL U50161 ( .A(n2939), .B(n2006), .Y(n60919) );
  HB1xp67_ASAP7_75t_SL U50162 ( .A(n66283), .Y(n57506) );
  NAND2xp5_ASAP7_75t_SL U50163 ( .A(n59578), .B(n58853), .Y(n66452) );
  AND2x2_ASAP7_75t_SL U50164 ( .A(n57630), .B(n67230), .Y(n67535) );
  BUFx3_ASAP7_75t_SL U50165 ( .A(n59483), .Y(n57352) );
  NOR2xp33_ASAP7_75t_SL U50166 ( .A(n59515), .B(n67581), .Y(n67582) );
  NAND2xp5_ASAP7_75t_SL U50167 ( .A(n58861), .B(n67580), .Y(n58862) );
  NOR2xp33_ASAP7_75t_SL U50168 ( .A(n1868), .B(n59591), .Y(n57261) );
  BUFx6f_ASAP7_75t_SL U50169 ( .A(n59516), .Y(n57394) );
  INVx3_ASAP7_75t_SL U50170 ( .A(n75967), .Y(n59669) );
  AOI21xp5_ASAP7_75t_SL U50171 ( .A1(n57186), .A2(n67423), .B(n59582), .Y(
        n75967) );
  NOR2xp33_ASAP7_75t_SL U50172 ( .A(n62561), .B(n59322), .Y(n59321) );
  NAND2xp5_ASAP7_75t_SL U50173 ( .A(n62581), .B(n59655), .Y(n62675) );
  NOR2x1_ASAP7_75t_SL U50174 ( .A(n59614), .B(n67629), .Y(n67268) );
  NOR2x1_ASAP7_75t_SL U50175 ( .A(n59591), .B(n66634), .Y(n66636) );
  INVxp33_ASAP7_75t_SRAM U50176 ( .A(n70695), .Y(n70737) );
  NAND2xp5_ASAP7_75t_SL U50177 ( .A(n63242), .B(n63257), .Y(n63243) );
  XOR2xp5_ASAP7_75t_SL U50178 ( .A(n64021), .B(n63874), .Y(n63875) );
  NAND2xp5_ASAP7_75t_SL U50179 ( .A(n57909), .B(n57908), .Y(n68828) );
  HB1xp67_ASAP7_75t_SL U50180 ( .A(n53399), .Y(n57421) );
  NAND2xp5_ASAP7_75t_SL U50181 ( .A(n74562), .B(n74563), .Y(n75287) );
  BUFx6f_ASAP7_75t_SL U50182 ( .A(n59669), .Y(n57456) );
  NAND2xp5_ASAP7_75t_SL U50183 ( .A(n2544), .B(n59540), .Y(n76547) );
  NOR2x1_ASAP7_75t_SL U50184 ( .A(n64229), .B(n61854), .Y(n75245) );
  NAND2xp5_ASAP7_75t_SL U50185 ( .A(n59538), .B(n59540), .Y(n60607) );
  NAND2xp5_ASAP7_75t_SL U50186 ( .A(n59560), .B(n59570), .Y(n57591) );
  BUFx2_ASAP7_75t_SL U50187 ( .A(n59462), .Y(n57407) );
  INVx1_ASAP7_75t_SL U50188 ( .A(n62476), .Y(n62477) );
  INVx1_ASAP7_75t_SL U50189 ( .A(dc_en), .Y(n61289) );
  NAND2xp5_ASAP7_75t_SL U50190 ( .A(n57126), .B(n76763), .Y(n77101) );
  INVx1_ASAP7_75t_SL U50191 ( .A(n77686), .Y(n77748) );
  NAND2x1p5_ASAP7_75t_SL U50192 ( .A(n67837), .B(n59436), .Y(n59356) );
  INVx2_ASAP7_75t_SL U50193 ( .A(n59435), .Y(n57106) );
  NAND2x1p5_ASAP7_75t_SL U50194 ( .A(n57212), .B(n57119), .Y(n57802) );
  NAND2x1p5_ASAP7_75t_SL U50195 ( .A(n59455), .B(n63182), .Y(n66805) );
  BUFx2_ASAP7_75t_SL U50196 ( .A(n67912), .Y(n57358) );
  INVx2_ASAP7_75t_SL U50197 ( .A(n58172), .Y(n57880) );
  NAND2x1p5_ASAP7_75t_SL U50198 ( .A(n67424), .B(n59231), .Y(n67598) );
  NOR2xp33_ASAP7_75t_SL U50199 ( .A(n1626), .B(n58176), .Y(n58494) );
  INVx1_ASAP7_75t_SL U50200 ( .A(n64515), .Y(n59351) );
  NAND2xp5_ASAP7_75t_SL U50201 ( .A(n57117), .B(n63673), .Y(n58045) );
  AO21x1_ASAP7_75t_SL U50202 ( .A1(n78004), .A2(n58433), .B(n62621), .Y(n62601) );
  HB1xp67_ASAP7_75t_SL U50203 ( .A(n1686), .Y(n57331) );
  BUFx2_ASAP7_75t_SL U50204 ( .A(n58856), .Y(n57246) );
  BUFx2_ASAP7_75t_SL U50205 ( .A(n65102), .Y(n57332) );
  INVx1_ASAP7_75t_SL U50206 ( .A(n64984), .Y(n64869) );
  BUFx2_ASAP7_75t_SL U50207 ( .A(n68805), .Y(n57269) );
  NOR2xp33_ASAP7_75t_SL U50208 ( .A(n58840), .B(n58842), .Y(n57606) );
  NAND2xp33_ASAP7_75t_SRAM U50209 ( .A(n77850), .B(n59686), .Y(n77929) );
  BUFx2_ASAP7_75t_SL U50210 ( .A(n75477), .Y(n57318) );
  NOR2xp33_ASAP7_75t_SL U50211 ( .A(dbg_we_i), .B(n78439), .Y(n77847) );
  NOR2xp33_ASAP7_75t_SL U50212 ( .A(dbg_we_i), .B(n77581), .Y(n77675) );
  BUFx2_ASAP7_75t_SL U50213 ( .A(n1770), .Y(n57404) );
  BUFx2_ASAP7_75t_SL U50214 ( .A(n59566), .Y(n57483) );
  NAND2xp5_ASAP7_75t_SL U50215 ( .A(n59661), .B(n68098), .Y(n67459) );
  INVx3_ASAP7_75t_SL U50216 ( .A(n68119), .Y(n57163) );
  NAND2x1p5_ASAP7_75t_SL U50217 ( .A(n63654), .B(n64930), .Y(n63809) );
  INVx5_ASAP7_75t_SL U50218 ( .A(n59570), .Y(n57128) );
  NAND2x1_ASAP7_75t_SL U50219 ( .A(n56861), .B(n59559), .Y(n57648) );
  XOR2xp5_ASAP7_75t_SL U50220 ( .A(n58955), .B(n57792), .Y(n68320) );
  NAND2x1p5_ASAP7_75t_SL U50221 ( .A(n59532), .B(n59536), .Y(n61807) );
  NOR2xp33_ASAP7_75t_SL U50222 ( .A(n57219), .B(n57214), .Y(n58212) );
  BUFx2_ASAP7_75t_SL U50223 ( .A(n59437), .Y(n57272) );
  BUFx2_ASAP7_75t_SL U50224 ( .A(n75895), .Y(n57311) );
  BUFx2_ASAP7_75t_SL U50225 ( .A(n62591), .Y(n57448) );
  NAND3xp33_ASAP7_75t_SL U50226 ( .A(n56944), .B(n56942), .C(n56941), .Y(
        n51997) );
  NAND2xp5_ASAP7_75t_SL U50227 ( .A(n56859), .B(n58262), .Y(n56941) );
  INVx1_ASAP7_75t_SL U50228 ( .A(dbg_stb_i), .Y(n78439) );
  AOI211xp5_ASAP7_75t_SL U50229 ( .A1(n57101), .A2(n58871), .B(n67541), .C(
        n58196), .Y(n67545) );
  NAND2xp5_ASAP7_75t_SL U50230 ( .A(n59599), .B(n57662), .Y(n67289) );
  NOR2xp33_ASAP7_75t_SL U50231 ( .A(n68383), .B(n67382), .Y(n59305) );
  NOR2xp33_ASAP7_75t_SL U50232 ( .A(n59418), .B(n67740), .Y(n57232) );
  NAND2xp5_ASAP7_75t_SL U50233 ( .A(n59649), .B(n67428), .Y(n57542) );
  NAND2xp5_ASAP7_75t_SL U50234 ( .A(n59666), .B(n67364), .Y(n67375) );
  NOR2xp33_ASAP7_75t_SL U50235 ( .A(n67962), .B(n59605), .Y(n67960) );
  NOR2xp33_ASAP7_75t_SL U50236 ( .A(n64934), .B(n58658), .Y(n64935) );
  INVx1_ASAP7_75t_SL U50237 ( .A(n59557), .Y(n57576) );
  NAND2x1p5_ASAP7_75t_SL U50238 ( .A(n1796), .B(n59555), .Y(n58808) );
  NOR2xp33_ASAP7_75t_SL U50239 ( .A(n67343), .B(n75894), .Y(n67286) );
  NOR2xp33_ASAP7_75t_SL U50240 ( .A(n57312), .B(n59591), .Y(n57661) );
  NOR2xp33_ASAP7_75t_SL U50241 ( .A(n59617), .B(n75912), .Y(n57816) );
  NOR2xp33_ASAP7_75t_SL U50242 ( .A(n59662), .B(n57821), .Y(n67370) );
  NOR2xp33_ASAP7_75t_SL U50243 ( .A(n58851), .B(n67511), .Y(n58196) );
  NAND2x1p5_ASAP7_75t_SL U50244 ( .A(n59555), .B(n57960), .Y(n62615) );
  XOR2xp5_ASAP7_75t_SL U50245 ( .A(n57691), .B(n67616), .Y(n57268) );
  HB1xp67_ASAP7_75t_SL U50246 ( .A(n62805), .Y(n57462) );
  HB1xp67_ASAP7_75t_SL U50247 ( .A(n62804), .Y(n57443) );
  BUFx2_ASAP7_75t_SL U50248 ( .A(n67356), .Y(n57428) );
  O2A1O1Ixp33_ASAP7_75t_SL U50249 ( .A1(n66374), .A2(n66378), .B(n67306), .C(
        n53630), .Y(n66350) );
  INVx1_ASAP7_75t_SL U50250 ( .A(n66545), .Y(n53631) );
  HAxp5_ASAP7_75t_SL U50251 ( .A(n61946), .B(n59531), .CON(), .SN(n62074) );
  A2O1A1Ixp33_ASAP7_75t_SL U50252 ( .A1(n67227), .A2(n67580), .B(n53633), .C(
        n62717), .Y(n53634) );
  A2O1A1Ixp33_ASAP7_75t_SL U50253 ( .A1(n62719), .A2(n62720), .B(n62718), .C(
        n53634), .Y(n62734) );
  INVxp33_ASAP7_75t_SRAM U50254 ( .A(n75073), .Y(n53635) );
  O2A1O1Ixp33_ASAP7_75t_SL U50255 ( .A1(n59636), .A2(n53635), .B(n53636), .C(
        n53637), .Y(n75081) );
  INVx1_ASAP7_75t_SL U50256 ( .A(n60962), .Y(n53638) );
  INVxp33_ASAP7_75t_SRAM U50257 ( .A(n65082), .Y(n53652) );
  INVxp33_ASAP7_75t_SRAM U50258 ( .A(n65089), .Y(n53653) );
  INVxp33_ASAP7_75t_SRAM U50259 ( .A(n1891), .Y(n53655) );
  INVxp33_ASAP7_75t_SRAM U50260 ( .A(n76860), .Y(n53657) );
  INVx1_ASAP7_75t_SL U50261 ( .A(n53667), .Y(n61425) );
  INVxp33_ASAP7_75t_SRAM U50262 ( .A(n73889), .Y(n53668) );
  INVx1_ASAP7_75t_SL U50263 ( .A(n74269), .Y(n53669) );
  OAI21xp33_ASAP7_75t_SL U50264 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[1]), 
        .A2(n53669), .B(n53668), .Y(n53670) );
  A2O1A1Ixp33_ASAP7_75t_SL U50265 ( .A1(n74269), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[1]), .B(
        n53668), .C(n53670), .Y(n53671) );
  INVxp33_ASAP7_75t_SRAM U50266 ( .A(n72641), .Y(n53673) );
  INVxp33_ASAP7_75t_SRAM U50267 ( .A(n75661), .Y(n53687) );
  INVxp33_ASAP7_75t_SRAM U50268 ( .A(n75659), .Y(n53689) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50269 ( .A1(n75664), .A2(n53687), .B(n53691), 
        .C(n75663), .Y(n76895) );
  INVxp33_ASAP7_75t_SRAM U50270 ( .A(n69284), .Y(n53692) );
  INVx1_ASAP7_75t_SL U50271 ( .A(n69176), .Y(n53693) );
  INVxp33_ASAP7_75t_SRAM U50272 ( .A(n63245), .Y(n53694) );
  INVx1_ASAP7_75t_SL U50273 ( .A(n53696), .Y(n53697) );
  INVx1_ASAP7_75t_SL U50274 ( .A(n74071), .Y(n53699) );
  INVxp33_ASAP7_75t_SRAM U50275 ( .A(n74884), .Y(n53700) );
  INVx1_ASAP7_75t_SL U50276 ( .A(n64329), .Y(n53701) );
  INVxp33_ASAP7_75t_SRAM U50277 ( .A(n65203), .Y(n53708) );
  INVxp33_ASAP7_75t_SRAM U50278 ( .A(n3100), .Y(n53711) );
  INVxp33_ASAP7_75t_SRAM U50279 ( .A(n70240), .Y(n53715) );
  INVxp33_ASAP7_75t_SRAM U50280 ( .A(n66085), .Y(n53718) );
  NAND3xp33_ASAP7_75t_SL U50281 ( .A(n53720), .B(n71179), .C(n71271), .Y(
        n53721) );
  A2O1A1Ixp33_ASAP7_75t_SL U50282 ( .A1(n71179), .A2(n71271), .B(n53720), .C(
        n53721), .Y(n53722) );
  INVxp33_ASAP7_75t_SRAM U50283 ( .A(n59698), .Y(n53723) );
  INVxp33_ASAP7_75t_SRAM U50284 ( .A(n74276), .Y(n53739) );
  OAI21xp33_ASAP7_75t_SRAM U50285 ( .A1(n74265), .A2(n74264), .B(n53739), .Y(
        n53740) );
  A2O1A1Ixp33_ASAP7_75t_SL U50286 ( .A1(n74264), .A2(n74265), .B(n53740), .C(
        n74275), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n55) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50287 ( .A1(n78166), .A2(n78165), .B(n3090), .C(
        n78164), .Y(or1200_dc_top_dcfsm_tag_we) );
  INVxp33_ASAP7_75t_SRAM U50288 ( .A(n69050), .Y(n53762) );
  INVxp33_ASAP7_75t_SRAM U50289 ( .A(n63319), .Y(n53773) );
  AOI21xp33_ASAP7_75t_SRAM U50290 ( .A1(n63316), .A2(n53773), .B(n76897), .Y(
        n53774) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50291 ( .A1(n63316), .A2(n53773), .B(n53774), 
        .C(n53772), .Y(n53775) );
  OAI21xp33_ASAP7_75t_SRAM U50292 ( .A1(n63399), .A2(n63320), .B(n59674), .Y(
        n53776) );
  A2O1A1Ixp33_ASAP7_75t_SL U50293 ( .A1(n63320), .A2(n63399), .B(n53776), .C(
        n53775), .Y(n53777) );
  INVx1_ASAP7_75t_SL U50294 ( .A(n53777), .Y(n53778) );
  INVxp33_ASAP7_75t_SRAM U50295 ( .A(n53440), .Y(n53779) );
  INVxp33_ASAP7_75t_SRAM U50296 ( .A(n74973), .Y(n53783) );
  A2O1A1Ixp33_ASAP7_75t_SL U50297 ( .A1(n74984), .A2(n77287), .B(n53782), .C(
        n53783), .Y(or1200_pic_N65) );
  INVxp33_ASAP7_75t_SRAM U50298 ( .A(n57144), .Y(n53786) );
  INVx1_ASAP7_75t_SL U50299 ( .A(n65400), .Y(n53794) );
  INVxp33_ASAP7_75t_SRAM U50300 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_4_), .Y(n53798) );
  INVx1_ASAP7_75t_SL U50301 ( .A(n57202), .Y(n53801) );
  INVxp33_ASAP7_75t_SRAM U50302 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[26]), .Y(n53805) );
  A2O1A1Ixp33_ASAP7_75t_SL U50303 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[26]), .A2(n53804), 
        .B(n59621), .C(n53806), .Y(n2439) );
  INVxp33_ASAP7_75t_SRAM U50304 ( .A(n57144), .Y(n53808) );
  INVx1_ASAP7_75t_SL U50305 ( .A(n60726), .Y(n53811) );
  INVxp33_ASAP7_75t_SRAM U50306 ( .A(n2649), .Y(n53814) );
  NAND2xp33_ASAP7_75t_SRAM U50307 ( .A(iwb_dat_i[9]), .B(n59496), .Y(n60396)
         );
  INVx1_ASAP7_75t_SL U50308 ( .A(n67992), .Y(n53826) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50309 ( .A1(n64951), .A2(n53455), .B(n53828), 
        .C(n64950), .Y(n61966) );
  O2A1O1Ixp33_ASAP7_75t_SL U50310 ( .A1(n67232), .A2(n67264), .B(n53829), .C(
        n53830), .Y(n63062) );
  INVxp33_ASAP7_75t_SRAM U50311 ( .A(n66430), .Y(n53831) );
  INVxp33_ASAP7_75t_SRAM U50312 ( .A(n66535), .Y(n53832) );
  INVxp33_ASAP7_75t_SRAM U50313 ( .A(n66378), .Y(n53833) );
  INVxp33_ASAP7_75t_SRAM U50314 ( .A(n59554), .Y(n53838) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50315 ( .A1(n59511), .A2(n59503), .B(n67424), 
        .C(n57246), .Y(n53844) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50316 ( .A1(n67424), .A2(n53843), .B(n57246), 
        .C(n53844), .Y(n53845) );
  O2A1O1Ixp33_ASAP7_75t_SL U50317 ( .A1(n67343), .A2(n67601), .B(n53842), .C(
        n53845), .Y(n62866) );
  INVxp33_ASAP7_75t_SRAM U50318 ( .A(n75082), .Y(n53846) );
  INVxp33_ASAP7_75t_SRAM U50319 ( .A(n62295), .Y(n53847) );
  INVxp33_ASAP7_75t_SRAM U50320 ( .A(n76087), .Y(n53854) );
  INVx1_ASAP7_75t_SL U50321 ( .A(n72945), .Y(n53855) );
  INVxp33_ASAP7_75t_SRAM U50322 ( .A(n60656), .Y(n53860) );
  AOI22xp33_ASAP7_75t_SRAM U50323 ( .A1(n75570), .A2(
        or1200_dc_top_from_dcram_19_), .B1(dwb_dat_i[19]), .B2(n75569), .Y(
        n61553) );
  INVxp33_ASAP7_75t_SRAM U50324 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .Y(
        n53863) );
  A2O1A1Ixp33_ASAP7_75t_SL U50325 ( .A1(n70189), .A2(n53863), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[6]), .C(
        n53864), .Y(n70201) );
  INVx1_ASAP7_75t_SL U50326 ( .A(n72621), .Y(n53865) );
  INVx1_ASAP7_75t_SL U50327 ( .A(n71213), .Y(n53879) );
  INVx1_ASAP7_75t_SL U50328 ( .A(n74082), .Y(n53886) );
  A2O1A1Ixp33_ASAP7_75t_SL U50329 ( .A1(n69111), .A2(n69112), .B(n53888), .C(
        n53889), .Y(n69125) );
  INVxp33_ASAP7_75t_SRAM U50330 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_12_), .Y(n53900)
         );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50331 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_14_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_13_), .B(n53899), 
        .C(n53901), .Y(n53902) );
  A2O1A1Ixp33_ASAP7_75t_SL U50332 ( .A1(n76943), .A2(n76944), .B(n76942), .C(
        n53902), .Y(n53903) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50333 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_0_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_1_), .B(n53898), 
        .C(n53903), .Y(n53904) );
  INVxp33_ASAP7_75t_SRAM U50334 ( .A(n73888), .Y(n53908) );
  INVx1_ASAP7_75t_SL U50335 ( .A(n74101), .Y(n53909) );
  OAI21xp5_ASAP7_75t_SL U50336 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[3]), 
        .A2(n53909), .B(n53908), .Y(n53910) );
  A2O1A1Ixp33_ASAP7_75t_SL U50337 ( .A1(n74101), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[3]), .B(
        n53908), .C(n53910), .Y(n74257) );
  INVx1_ASAP7_75t_SL U50338 ( .A(n73571), .Y(n53912) );
  A2O1A1Ixp33_ASAP7_75t_SL U50339 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_5_), .A2(n66166), 
        .B(n66165), .C(n66164), .Y(n53929) );
  A2O1A1Ixp33_ASAP7_75t_SL U50340 ( .A1(n71122), .A2(n53931), .B(n59699), .C(
        n53932), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n190) );
  A2O1A1Ixp33_ASAP7_75t_SL U50341 ( .A1(n71030), .A2(n71023), .B(n59698), .C(
        n70992), .Y(n53936) );
  A2O1A1Ixp33_ASAP7_75t_SL U50342 ( .A1(n71023), .A2(n53935), .B(n70992), .C(
        n53936), .Y(n53937) );
  INVxp33_ASAP7_75t_SRAM U50343 ( .A(n72534), .Y(n53939) );
  INVxp33_ASAP7_75t_SRAM U50344 ( .A(n72544), .Y(n53946) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50345 ( .A1(n72329), .A2(n72499), .B(n72474), 
        .C(n53948), .Y(n53949) );
  A2O1A1Ixp33_ASAP7_75t_SL U50346 ( .A1(n72331), .A2(n53944), .B(n53949), .C(
        n72330), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n67) );
  A2O1A1Ixp33_ASAP7_75t_SL U50347 ( .A1(n74099), .A2(n74100), .B(n74233), .C(
        n74239), .Y(n53950) );
  INVxp33_ASAP7_75t_SRAM U50348 ( .A(n890), .Y(n78030) );
  A2O1A1Ixp33_ASAP7_75t_SL U50349 ( .A1(n57080), .A2(n53958), .B(n53961), .C(
        n53963), .Y(n53964) );
  INVxp33_ASAP7_75t_SRAM U50350 ( .A(n63509), .Y(n53965) );
  INVxp33_ASAP7_75t_SRAM U50351 ( .A(n63534), .Y(n53973) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50352 ( .A1(n63511), .A2(n53974), .B(n63513), 
        .C(n63516), .Y(n53975) );
  INVxp33_ASAP7_75t_SRAM U50353 ( .A(n63269), .Y(n53980) );
  INVx1_ASAP7_75t_SL U50354 ( .A(n62032), .Y(n53985) );
  INVxp33_ASAP7_75t_SRAM U50355 ( .A(n76631), .Y(n53991) );
  A2O1A1Ixp33_ASAP7_75t_SL U50356 ( .A1(or1200_cpu_or1200_mult_mac_n60), .A2(
        n53990), .B(n53993), .C(n53994), .Y(or1200_cpu_or1200_mult_mac_n1524)
         );
  INVxp33_ASAP7_75t_SRAM U50357 ( .A(n53440), .Y(n53995) );
  INVx1_ASAP7_75t_SL U50358 ( .A(n77287), .Y(n53999) );
  INVxp33_ASAP7_75t_SRAM U50359 ( .A(n77207), .Y(n54003) );
  OAI22xp33_ASAP7_75t_SRAM U50360 ( .A1(n2549), .A2(n59679), .B1(n59548), .B2(
        n57074), .Y(n75803) );
  INVxp33_ASAP7_75t_SRAM U50361 ( .A(n65391), .Y(n54009) );
  A2O1A1Ixp33_ASAP7_75t_SL U50362 ( .A1(n65393), .A2(n65394), .B(n65392), .C(
        n54010), .Y(n54011) );
  INVxp33_ASAP7_75t_SRAM U50363 ( .A(ex_insn[16]), .Y(n54017) );
  NAND2xp33_ASAP7_75t_SRAM U50364 ( .A(iwb_dat_i[8]), .B(n59495), .Y(n60390)
         );
  INVx1_ASAP7_75t_SL U50365 ( .A(n64084), .Y(n54022) );
  O2A1O1Ixp33_ASAP7_75t_SL U50366 ( .A1(n54023), .A2(n64336), .B(n64340), .C(
        n54024), .Y(n54025) );
  XNOR2xp5_ASAP7_75t_SL U50367 ( .A(n64337), .B(n54025), .Y(n64665) );
  INVx1_ASAP7_75t_SL U50368 ( .A(n67752), .Y(n54026) );
  INVxp33_ASAP7_75t_SRAM U50369 ( .A(n53229), .Y(n54029) );
  O2A1O1Ixp33_ASAP7_75t_SL U50370 ( .A1(n59578), .A2(n57120), .B(n54028), .C(
        n54029), .Y(n61962) );
  INVx1_ASAP7_75t_SL U50371 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[4]), .Y(
        n54032) );
  INVxp33_ASAP7_75t_SRAM U50372 ( .A(n70864), .Y(n54033) );
  INVxp33_ASAP7_75t_SRAM U50373 ( .A(n75034), .Y(n54034) );
  AOI21xp33_ASAP7_75t_SRAM U50374 ( .A1(n77011), .A2(n59811), .B(n77014), .Y(
        n59792) );
  INVxp33_ASAP7_75t_SRAM U50375 ( .A(n76124), .Y(n54040) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50376 ( .A1(n59614), .A2(n67227), .B(n62835), 
        .C(n68079), .Y(n54041) );
  INVx1_ASAP7_75t_SL U50377 ( .A(n64755), .Y(n54044) );
  INVxp33_ASAP7_75t_SRAM U50378 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[1]), .Y(
        n54051) );
  INVxp33_ASAP7_75t_SRAM U50379 ( .A(n65408), .Y(n54053) );
  INVx1_ASAP7_75t_SL U50380 ( .A(n66092), .Y(n54062) );
  INVx1_ASAP7_75t_SL U50381 ( .A(n54063), .Y(n54064) );
  INVx1_ASAP7_75t_SL U50382 ( .A(n54066), .Y(n70818) );
  INVx1_ASAP7_75t_SL U50383 ( .A(n74236), .Y(n54071) );
  INVxp33_ASAP7_75t_SRAM U50384 ( .A(n69209), .Y(n54075) );
  INVx1_ASAP7_75t_SL U50385 ( .A(dbg_dat_i[26]), .Y(n54080) );
  O2A1O1Ixp33_ASAP7_75t_SL U50386 ( .A1(n76548), .A2(n54081), .B(n54084), .C(
        n54085), .Y(n77970) );
  A2O1A1Ixp33_ASAP7_75t_SL U50387 ( .A1(n2569), .A2(n77752), .B(n3423), .C(
        n54093), .Y(n54094) );
  INVxp33_ASAP7_75t_SRAM U50388 ( .A(n61292), .Y(n54096) );
  INVxp33_ASAP7_75t_SRAM U50389 ( .A(n71156), .Y(n54098) );
  INVxp33_ASAP7_75t_SRAM U50390 ( .A(n71157), .Y(n54099) );
  INVxp33_ASAP7_75t_SRAM U50391 ( .A(n71601), .Y(n54107) );
  INVxp33_ASAP7_75t_SRAM U50392 ( .A(n72472), .Y(n54118) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50393 ( .A1(n72474), .A2(n72473), .B(n54122), 
        .C(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .Y(
        n54123) );
  INVxp33_ASAP7_75t_SRAM U50394 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .Y(
        n54124) );
  INVxp33_ASAP7_75t_SRAM U50395 ( .A(n1345), .Y(n77497) );
  INVxp33_ASAP7_75t_SRAM U50396 ( .A(n77495), .Y(n77496) );
  INVxp33_ASAP7_75t_SRAM U50397 ( .A(n63385), .Y(n54132) );
  INVxp33_ASAP7_75t_SRAM U50398 ( .A(n63394), .Y(n54133) );
  INVxp33_ASAP7_75t_SRAM U50399 ( .A(n53440), .Y(n54143) );
  INVxp33_ASAP7_75t_SRAM U50400 ( .A(n1220), .Y(n78097) );
  INVxp33_ASAP7_75t_SRAM U50401 ( .A(n78089), .Y(n78091) );
  INVxp33_ASAP7_75t_SRAM U50402 ( .A(n76856), .Y(n54147) );
  A2O1A1Ixp33_ASAP7_75t_SL U50403 ( .A1(n77591), .A2(n77287), .B(n54146), .C(
        n54147), .Y(or1200_pic_N50) );
  INVx1_ASAP7_75t_SL U50404 ( .A(n78435), .Y(n54160) );
  NAND3xp33_ASAP7_75t_SL U50405 ( .A(n54160), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_0_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_1_), .Y(n54161) );
  A2O1A1Ixp33_ASAP7_75t_SL U50406 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_0_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_1_), .B(n54160), .C(
        n54161), .Y(n1729) );
  INVxp33_ASAP7_75t_SRAM U50407 ( .A(n59680), .Y(n54163) );
  INVxp33_ASAP7_75t_SRAM U50408 ( .A(n2009), .Y(n54166) );
  INVxp33_ASAP7_75t_SRAM U50409 ( .A(n69788), .Y(n54167) );
  INVxp33_ASAP7_75t_SRAM U50410 ( .A(n70515), .Y(n54168) );
  AOI22xp33_ASAP7_75t_SRAM U50411 ( .A1(n70515), .A2(n69788), .B1(n54167), 
        .B2(n54168), .Y(n54169) );
  A2O1A1Ixp33_ASAP7_75t_SL U50412 ( .A1(n70372), .A2(n54168), .B(n70502), .C(
        n54171), .Y(n54172) );
  A2O1A1Ixp33_ASAP7_75t_SL U50413 ( .A1(n69801), .A2(n54169), .B(n54170), .C(
        n54172), .Y(n2297) );
  INVx1_ASAP7_75t_SL U50414 ( .A(n57202), .Y(n54174) );
  INVxp33_ASAP7_75t_SRAM U50415 ( .A(n70469), .Y(n54179) );
  A2O1A1Ixp33_ASAP7_75t_SL U50416 ( .A1(n60344), .A2(n60343), .B(n62003), .C(
        n61155), .Y(n54191) );
  INVxp33_ASAP7_75t_SRAM U50417 ( .A(n2662), .Y(n54192) );
  NAND2xp33_ASAP7_75t_SRAM U50418 ( .A(iwb_dat_i[7]), .B(n78021), .Y(n60384)
         );
  OAI22xp33_ASAP7_75t_SRAM U50419 ( .A1(n2555), .A2(n77463), .B1(n59575), .B2(
        n57073), .Y(n76853) );
  AOI21xp33_ASAP7_75t_SRAM U50420 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[29]), .B(n76853), .Y(n76854) );
  A2O1A1Ixp33_ASAP7_75t_SL U50421 ( .A1(n75158), .A2(n53479), .B(n75180), .C(
        n59694), .Y(n54197) );
  INVxp33_ASAP7_75t_SRAM U50422 ( .A(n70576), .Y(n54198) );
  INVxp33_ASAP7_75t_SRAM U50423 ( .A(n67821), .Y(n54206) );
  INVx1_ASAP7_75t_SL U50424 ( .A(n62094), .Y(n54207) );
  INVxp33_ASAP7_75t_SRAM U50425 ( .A(n63210), .Y(n54209) );
  A2O1A1Ixp33_ASAP7_75t_SL U50426 ( .A1(n59594), .A2(n67920), .B(n54212), .C(
        n67609), .Y(n54213) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50427 ( .A1(n57365), .A2(n59668), .B(n54214), 
        .C(n54215), .Y(n75037) );
  A2O1A1Ixp33_ASAP7_75t_SL U50428 ( .A1(n54216), .A2(n54218), .B(n60979), .C(
        n54219), .Y(n76291) );
  INVxp33_ASAP7_75t_SRAM U50429 ( .A(n75426), .Y(n54221) );
  AOI22xp33_ASAP7_75t_SRAM U50430 ( .A1(dwb_dat_i[22]), .A2(n61548), .B1(
        n75569), .B2(dwb_dat_i[30]), .Y(n60838) );
  INVx1_ASAP7_75t_SL U50431 ( .A(n54236), .Y(n54237) );
  A2O1A1Ixp33_ASAP7_75t_SL U50432 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_), 
        .A2(n72309), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_), 
        .C(n72308), .Y(n54241) );
  INVxp33_ASAP7_75t_SRAM U50433 ( .A(n63759), .Y(n54259) );
  INVxp33_ASAP7_75t_SRAM U50434 ( .A(n57211), .Y(n54262) );
  A2O1A1Ixp33_ASAP7_75t_SL U50435 ( .A1(n71130), .A2(n59523), .B(n71099), .C(
        n54264), .Y(n54265) );
  INVxp33_ASAP7_75t_SRAM U50436 ( .A(n72482), .Y(n54267) );
  INVxp33_ASAP7_75t_SRAM U50437 ( .A(n899), .Y(n78031) );
  INVxp33_ASAP7_75t_SRAM U50438 ( .A(n69255), .Y(n54282) );
  A2O1A1Ixp33_ASAP7_75t_SL U50439 ( .A1(n59672), .A2(n54281), .B(n54284), .C(
        n54286), .Y(n54287) );
  A2O1A1Ixp33_ASAP7_75t_SL U50440 ( .A1(n69000), .A2(n54289), .B(n68995), .C(
        n57079), .Y(n54303) );
  INVxp33_ASAP7_75t_SRAM U50441 ( .A(n53440), .Y(n54309) );
  INVx1_ASAP7_75t_SL U50442 ( .A(n77287), .Y(n54315) );
  INVxp33_ASAP7_75t_SRAM U50443 ( .A(n76993), .Y(n54319) );
  NAND2xp33_ASAP7_75t_SRAM U50444 ( .A(n59678), .B(n77872), .Y(n64807) );
  INVx1_ASAP7_75t_SL U50445 ( .A(n77675), .Y(n54326) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50446 ( .A1(n54329), .A2(n65391), .B(n65400), 
        .C(n65401), .Y(n54330) );
  A2O1A1Ixp33_ASAP7_75t_SL U50447 ( .A1(n65400), .A2(n54331), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_5_), .C(n54332), .Y(
        n1839) );
  INVxp33_ASAP7_75t_SRAM U50448 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_5_), .Y(n54329) );
  INVxp33_ASAP7_75t_SRAM U50449 ( .A(n65391), .Y(n54331) );
  INVx1_ASAP7_75t_SL U50450 ( .A(n54330), .Y(n54332) );
  INVx1_ASAP7_75t_SL U50451 ( .A(n54333), .Y(n54334) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50452 ( .A1(n62047), .A2(n62048), .B(n62046), 
        .C(n54337), .Y(n54338) );
  INVxp33_ASAP7_75t_SRAM U50453 ( .A(n62000), .Y(n54339) );
  INVxp33_ASAP7_75t_SRAM U50454 ( .A(n2676), .Y(n54343) );
  NAND2xp33_ASAP7_75t_SRAM U50455 ( .A(iwb_dat_i[6]), .B(n59496), .Y(n61023)
         );
  INVx1_ASAP7_75t_SL U50456 ( .A(n72762), .Y(n54345) );
  INVxp33_ASAP7_75t_SRAM U50457 ( .A(n74460), .Y(n54351) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50458 ( .A1(n74463), .A2(n54351), .B(n74716), 
        .C(n74462), .Y(n54352) );
  OAI22xp33_ASAP7_75t_SRAM U50459 ( .A1(n2958), .A2(n77463), .B1(n59579), .B2(
        n57074), .Y(n76987) );
  AOI21xp33_ASAP7_75t_SRAM U50460 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[31]), .B(n76987), .Y(n76988) );
  INVxp33_ASAP7_75t_SRAM U50461 ( .A(n57144), .Y(n54354) );
  A2O1A1Ixp33_ASAP7_75t_SL U50462 ( .A1(n75157), .A2(n54354), .B(n75156), .C(
        n54355), .Y(n54356) );
  INVxp33_ASAP7_75t_SRAM U50463 ( .A(n70597), .Y(n54357) );
  INVx1_ASAP7_75t_SL U50464 ( .A(n59478), .Y(n54359) );
  O2A1O1Ixp33_ASAP7_75t_SL U50465 ( .A1(n68024), .A2(n68117), .B(n68023), .C(
        n54359), .Y(n54360) );
  O2A1O1Ixp5_ASAP7_75t_SL U50466 ( .A1(n58811), .A2(n59478), .B(n68076), .C(
        n54360), .Y(n68203) );
  A2O1A1Ixp33_ASAP7_75t_SL U50467 ( .A1(n75046), .A2(n59190), .B(n54366), .C(
        n54367), .Y(n75063) );
  INVx1_ASAP7_75t_SL U50468 ( .A(n2583), .Y(n54374) );
  INVxp33_ASAP7_75t_SRAM U50469 ( .A(n74118), .Y(n54375) );
  AOI22xp33_ASAP7_75t_SRAM U50470 ( .A1(n75570), .A2(
        or1200_dc_top_from_dcram_16_), .B1(dwb_dat_i[16]), .B2(n75569), .Y(
        n60593) );
  NAND2xp33_ASAP7_75t_SRAM U50471 ( .A(n77752), .B(n60592), .Y(n60594) );
  INVxp33_ASAP7_75t_SRAM U50472 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[4]), .Y(
        n54391) );
  INVxp33_ASAP7_75t_SRAM U50473 ( .A(n74138), .Y(n54392) );
  INVxp33_ASAP7_75t_SRAM U50474 ( .A(n76519), .Y(n54398) );
  A2O1A1Ixp33_ASAP7_75t_SL U50475 ( .A1(n70941), .A2(n70978), .B(n59699), .C(
        n54405), .Y(n54406) );
  A2O1A1Ixp33_ASAP7_75t_SL U50476 ( .A1(n70978), .A2(n54402), .B(n54405), .C(
        n54406), .Y(n54407) );
  A2O1A1Ixp33_ASAP7_75t_SL U50477 ( .A1(n70729), .A2(n70720), .B(n59698), .C(
        n70732), .Y(n54411) );
  A2O1A1Ixp33_ASAP7_75t_SL U50478 ( .A1(n70720), .A2(n54410), .B(n70732), .C(
        n54411), .Y(n54412) );
  INVxp33_ASAP7_75t_SRAM U50479 ( .A(or1200_cpu_or1200_mult_mac_n161), .Y(
        n54441) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50480 ( .A1(n63439), .A2(n63531), .B(n54440), 
        .C(n54449), .Y(n54450) );
  INVxp33_ASAP7_75t_SRAM U50481 ( .A(n76077), .Y(n54451) );
  INVx1_ASAP7_75t_SL U50482 ( .A(n57133), .Y(n54452) );
  OAI21xp5_ASAP7_75t_SL U50483 ( .A1(n76080), .A2(n54452), .B(n54451), .Y(
        n54453) );
  OAI21xp5_ASAP7_75t_SL U50484 ( .A1(or1200_cpu_or1200_mult_mac_n36), .A2(
        n53469), .B(n76631), .Y(n54455) );
  A2O1A1Ixp33_ASAP7_75t_SL U50485 ( .A1(or1200_cpu_or1200_mult_mac_n36), .A2(
        n53469), .B(n54455), .C(n54454), .Y(or1200_cpu_or1200_mult_mac_n1512)
         );
  INVxp33_ASAP7_75t_SRAM U50486 ( .A(n53440), .Y(n54456) );
  INVxp33_ASAP7_75t_SRAM U50487 ( .A(n59680), .Y(n54472) );
  INVxp33_ASAP7_75t_SRAM U50488 ( .A(n77199), .Y(n54473) );
  A2O1A1Ixp33_ASAP7_75t_SL U50489 ( .A1(n77162), .A2(n54474), .B(n77161), .C(
        n1985), .Y(n54475) );
  INVxp33_ASAP7_75t_SRAM U50490 ( .A(n65400), .Y(n54478) );
  INVxp33_ASAP7_75t_SRAM U50491 ( .A(n69780), .Y(n54480) );
  INVx1_ASAP7_75t_SL U50492 ( .A(n57202), .Y(n54490) );
  INVxp33_ASAP7_75t_SRAM U50493 ( .A(n70483), .Y(n54505) );
  INVxp33_ASAP7_75t_SRAM U50494 ( .A(n77408), .Y(n54510) );
  NAND2xp33_ASAP7_75t_SRAM U50495 ( .A(iwb_dat_i[5]), .B(n78021), .Y(n61590)
         );
  AOI22xp33_ASAP7_75t_SRAM U50496 ( .A1(n76653), .A2(n57144), .B1(n76652), 
        .B2(n77279), .Y(n76656) );
  INVxp33_ASAP7_75t_SRAM U50497 ( .A(n74875), .Y(n54515) );
  A2O1A1Ixp33_ASAP7_75t_SL U50498 ( .A1(n74876), .A2(n54514), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_22_), .C(n54516), 
        .Y(n52504) );
  INVx1_ASAP7_75t_SL U50499 ( .A(n70602), .Y(n54525) );
  A2O1A1Ixp33_ASAP7_75t_SL U50500 ( .A1(n54524), .A2(n54525), .B(n70594), .C(
        n54526), .Y(n51980) );
  O2A1O1Ixp33_ASAP7_75t_SL U50501 ( .A1(n73424), .A2(n73425), .B(n73416), .C(
        n54534), .Y(n78215) );
  O2A1O1Ixp33_ASAP7_75t_SL U50502 ( .A1(n64893), .A2(n54535), .B(n65026), .C(
        n65025), .Y(n64901) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50503 ( .A1(n58711), .A2(n59659), .B(n54537), 
        .C(n57260), .Y(n54538) );
  NOR3xp33_ASAP7_75t_SL U50504 ( .A(n54540), .B(n64974), .C(n64973), .Y(n54541) );
  O2A1O1Ixp33_ASAP7_75t_SL U50505 ( .A1(n54540), .A2(n64973), .B(n64974), .C(
        n54541), .Y(n64904) );
  INVx1_ASAP7_75t_SL U50506 ( .A(n61966), .Y(n54542) );
  INVx1_ASAP7_75t_SL U50507 ( .A(n54543), .Y(n59259) );
  NAND2xp33_ASAP7_75t_SRAM U50508 ( .A(n59809), .B(n59945), .Y(n59812) );
  INVx1_ASAP7_75t_SL U50509 ( .A(n62599), .Y(n54545) );
  INVx1_ASAP7_75t_SL U50510 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[4]), .Y(
        n54547) );
  INVxp33_ASAP7_75t_SRAM U50511 ( .A(n65170), .Y(n54550) );
  AOI22xp33_ASAP7_75t_SRAM U50512 ( .A1(dwb_dat_i[20]), .A2(n61548), .B1(
        n75569), .B2(dwb_dat_i[28]), .Y(n61402) );
  INVx1_ASAP7_75t_SL U50513 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .Y(
        n55293) );
  INVxp33_ASAP7_75t_SRAM U50514 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .Y(n54565) );
  INVxp33_ASAP7_75t_SRAM U50515 ( .A(n69321), .Y(n54584) );
  INVx1_ASAP7_75t_SL U50516 ( .A(or1200_cpu_or1200_mult_mac_n379), .Y(n54585)
         );
  INVxp33_ASAP7_75t_SRAM U50517 ( .A(n76031), .Y(n54589) );
  INVx1_ASAP7_75t_SL U50518 ( .A(dbg_dat_i[30]), .Y(n54592) );
  INVx1_ASAP7_75t_SL U50519 ( .A(dbg_dat_i[24]), .Y(n54593) );
  INVx1_ASAP7_75t_SL U50520 ( .A(n4067), .Y(n54594) );
  INVxp33_ASAP7_75t_SRAM U50521 ( .A(n75423), .Y(n54595) );
  INVxp33_ASAP7_75t_SRAM U50522 ( .A(n59694), .Y(n54601) );
  INVx1_ASAP7_75t_SL U50523 ( .A(n73887), .Y(n54602) );
  INVxp33_ASAP7_75t_SRAM U50524 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_1_), 
        .Y(n54604) );
  A2O1A1Ixp33_ASAP7_75t_SL U50525 ( .A1(n74305), .A2(n54605), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_3_), 
        .C(n74304), .Y(n74737) );
  INVxp33_ASAP7_75t_SRAM U50526 ( .A(n71513), .Y(n54606) );
  INVxp33_ASAP7_75t_SRAM U50527 ( .A(n59698), .Y(n54607) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50528 ( .A1(n72497), .A2(n72496), .B(n72495), 
        .C(n54618), .Y(n54619) );
  A2O1A1Ixp33_ASAP7_75t_SL U50529 ( .A1(n74253), .A2(n54622), .B(n74276), .C(
        n74275), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n52) );
  INVxp33_ASAP7_75t_SRAM U50530 ( .A(n944), .Y(n78036) );
  INVxp33_ASAP7_75t_SRAM U50531 ( .A(n69130), .Y(n54627) );
  INVxp33_ASAP7_75t_SRAM U50532 ( .A(n69164), .Y(n54628) );
  A2O1A1Ixp33_ASAP7_75t_SL U50533 ( .A1(n57080), .A2(n54627), .B(n54630), .C(
        n54633), .Y(n54634) );
  INVxp33_ASAP7_75t_SRAM U50534 ( .A(n68845), .Y(n54636) );
  INVxp33_ASAP7_75t_SRAM U50535 ( .A(n63303), .Y(n54645) );
  INVxp33_ASAP7_75t_SRAM U50536 ( .A(or1200_cpu_or1200_mult_mac_div_free), .Y(
        n54652) );
  INVxp33_ASAP7_75t_SRAM U50537 ( .A(n53440), .Y(n54655) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50538 ( .A1(n1345), .A2(n1343), .B(n77488), .C(
        n77487), .Y(n54658) );
  INVxp33_ASAP7_75t_SRAM U50539 ( .A(n1343), .Y(n54660) );
  A2O1A1Ixp33_ASAP7_75t_SL U50540 ( .A1(n1790), .A2(n54667), .B(n59680), .C(
        n54668), .Y(or1200_du_N106) );
  INVxp33_ASAP7_75t_SRAM U50541 ( .A(n77133), .Y(n54669) );
  INVxp33_ASAP7_75t_SRAM U50542 ( .A(n70484), .Y(n54671) );
  A2O1A1Ixp33_ASAP7_75t_SL U50543 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[10]), .A2(n54676), 
        .B(n54677), .C(n2456), .Y(n2443) );
  INVxp33_ASAP7_75t_SRAM U50544 ( .A(n61140), .Y(n54678) );
  INVxp33_ASAP7_75t_SRAM U50545 ( .A(n60351), .Y(n54680) );
  OAI21xp33_ASAP7_75t_SRAM U50546 ( .A1(n54681), .A2(n61028), .B(n54678), .Y(
        n54683) );
  A2O1A1Ixp33_ASAP7_75t_SL U50547 ( .A1(n61028), .A2(n54682), .B(n54678), .C(
        n54683), .Y(n54684) );
  INVx1_ASAP7_75t_SL U50548 ( .A(n57072), .Y(n54686) );
  INVxp33_ASAP7_75t_SRAM U50549 ( .A(n65400), .Y(n54688) );
  INVxp33_ASAP7_75t_SRAM U50550 ( .A(n2683), .Y(n54692) );
  NAND2xp33_ASAP7_75t_SRAM U50551 ( .A(iwb_dat_i[4]), .B(n59495), .Y(n60892)
         );
  INVx1_ASAP7_75t_SL U50552 ( .A(n72720), .Y(n54698) );
  OAI22xp33_ASAP7_75t_SRAM U50553 ( .A1(n2558), .A2(n77463), .B1(n59576), .B2(
        n57074), .Y(n77464) );
  AOI21xp33_ASAP7_75t_SRAM U50554 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[30]), .B(n77464), .Y(n77466) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50555 ( .A1(n74871), .A2(n76956), .B(n76935), 
        .C(n77171), .Y(n54700) );
  INVxp33_ASAP7_75t_SRAM U50556 ( .A(n65224), .Y(n54703) );
  NOR3xp33_ASAP7_75t_SL U50557 ( .A(n54703), .B(n65226), .C(n54704), .Y(n54705) );
  O2A1O1Ixp33_ASAP7_75t_SL U50558 ( .A1(n54703), .A2(n54704), .B(n65226), .C(
        n54705), .Y(n54706) );
  A2O1A1Ixp33_ASAP7_75t_SL U50559 ( .A1(n59689), .A2(n76528), .B(n76529), .C(
        n54710), .Y(n54711) );
  INVxp33_ASAP7_75t_SRAM U50560 ( .A(n77705), .Y(n54715) );
  NAND3xp33_ASAP7_75t_SL U50561 ( .A(n54715), .B(n57120), .C(n64026), .Y(
        n54716) );
  A2O1A1Ixp33_ASAP7_75t_SL U50562 ( .A1(n57120), .A2(n64026), .B(n54715), .C(
        n54716), .Y(n61938) );
  INVxp33_ASAP7_75t_SRAM U50563 ( .A(n66483), .Y(n54717) );
  INVxp33_ASAP7_75t_SRAM U50564 ( .A(n57292), .Y(n54718) );
  A2O1A1Ixp33_ASAP7_75t_SL U50565 ( .A1(n75641), .A2(n54719), .B(n54720), .C(
        n66349), .Y(n54721) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50566 ( .A1(n66373), .A2(n54717), .B(n66350), 
        .C(n54721), .Y(n54722) );
  INVxp33_ASAP7_75t_SRAM U50567 ( .A(n77011), .Y(n54730) );
  INVxp33_ASAP7_75t_SRAM U50568 ( .A(n62002), .Y(n54745) );
  INVxp33_ASAP7_75t_SRAM U50569 ( .A(n75120), .Y(n54746) );
  INVxp33_ASAP7_75t_SRAM U50570 ( .A(n76095), .Y(n54747) );
  INVxp33_ASAP7_75t_SRAM U50571 ( .A(n62898), .Y(n54748) );
  INVxp33_ASAP7_75t_SRAM U50572 ( .A(n63242), .Y(n54750) );
  INVxp33_ASAP7_75t_SRAM U50573 ( .A(n76637), .Y(n54752) );
  INVxp33_ASAP7_75t_SRAM U50574 ( .A(n76615), .Y(n54753) );
  INVx1_ASAP7_75t_SL U50575 ( .A(n54758), .Y(n54759) );
  A2O1A1Ixp33_ASAP7_75t_SL U50576 ( .A1(n66096), .A2(n66093), .B(n66158), .C(
        n54776), .Y(n54777) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50577 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_3_), .A2(n66136), 
        .B(n66135), .C(n66138), .Y(n54784) );
  O2A1O1Ixp33_ASAP7_75t_SL U50578 ( .A1(n54785), .A2(n71404), .B(n71389), .C(
        n59698), .Y(n54786) );
  OAI31xp33_ASAP7_75t_SL U50579 ( .A1(n71389), .A2(n54785), .A3(n71404), .B(
        n54786), .Y(n54787) );
  INVxp33_ASAP7_75t_SRAM U50580 ( .A(n71790), .Y(n54788) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50581 ( .A1(n71793), .A2(n54788), .B(n71792), 
        .C(n71791), .Y(n54789) );
  INVxp33_ASAP7_75t_SRAM U50582 ( .A(n926), .Y(n78034) );
  A2O1A1Ixp33_ASAP7_75t_SL U50583 ( .A1(n74117), .A2(n57079), .B(n54798), .C(
        n54800), .Y(n54801) );
  INVxp33_ASAP7_75t_SRAM U50584 ( .A(n53440), .Y(n54806) );
  O2A1O1Ixp5_ASAP7_75t_SL U50585 ( .A1(n1119), .A2(n1121), .B(n54809), .C(
        n54810), .Y(n54811) );
  INVxp33_ASAP7_75t_SRAM U50586 ( .A(n1119), .Y(n54812) );
  A2O1A1Ixp33_ASAP7_75t_SL U50587 ( .A1(n1345), .A2(n77489), .B(n54814), .C(
        n54815), .Y(n9346) );
  INVx1_ASAP7_75t_SL U50588 ( .A(n77287), .Y(n54817) );
  INVxp33_ASAP7_75t_SRAM U50589 ( .A(n76610), .Y(n54821) );
  INVx1_ASAP7_75t_SL U50590 ( .A(n77287), .Y(n54822) );
  INVx1_ASAP7_75t_SL U50591 ( .A(pic_ints_i[0]), .Y(n54826) );
  INVxp33_ASAP7_75t_SRAM U50592 ( .A(n62071), .Y(n54829) );
  INVx1_ASAP7_75t_SL U50593 ( .A(n77761), .Y(n54831) );
  INVx1_ASAP7_75t_SL U50594 ( .A(n57202), .Y(n54844) );
  INVx1_ASAP7_75t_SL U50595 ( .A(n57202), .Y(n54848) );
  INVxp33_ASAP7_75t_SRAM U50596 ( .A(n70384), .Y(n54851) );
  A2O1A1Ixp33_ASAP7_75t_SL U50597 ( .A1(n59621), .A2(n54852), .B(n54853), .C(
        n2456), .Y(n2445) );
  INVxp33_ASAP7_75t_SRAM U50598 ( .A(n2657), .Y(n54854) );
  NAND2xp33_ASAP7_75t_SRAM U50599 ( .A(iwb_dat_i[3]), .B(n59496), .Y(n60353)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U50600 ( .A1(n77680), .A2(n77683), .B(n77285), .C(
        n77233), .Y(n54857) );
  INVx1_ASAP7_75t_SL U50601 ( .A(n77138), .Y(n54861) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50602 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_15_), .A2(n77171), 
        .B(n77139), .C(n54861), .Y(n52503) );
  NAND2xp33_ASAP7_75t_SRAM U50603 ( .A(n59678), .B(n77876), .Y(n64331) );
  OAI22xp33_ASAP7_75t_SRAM U50604 ( .A1(n2564), .A2(n59679), .B1(n59578), .B2(
        n57074), .Y(n64328) );
  A2O1A1Ixp33_ASAP7_75t_SL U50605 ( .A1(n75417), .A2(n75416), .B(n75415), .C(
        n75414), .Y(n54862) );
  A2O1A1Ixp33_ASAP7_75t_SL U50606 ( .A1(n75419), .A2(n54862), .B(n59695), .C(
        n54863), .Y(n3007) );
  INVxp33_ASAP7_75t_SRAM U50607 ( .A(n73654), .Y(n54871) );
  O2A1O1Ixp5_ASAP7_75t_SL U50608 ( .A1(n73434), .A2(n54874), .B(n73433), .C(
        n73432), .Y(n78213) );
  O2A1O1Ixp33_ASAP7_75t_SL U50609 ( .A1(n64350), .A2(n64351), .B(n57819), .C(
        n54875), .Y(n54876) );
  INVx1_ASAP7_75t_SL U50610 ( .A(n61962), .Y(n54877) );
  A2O1A1Ixp33_ASAP7_75t_SL U50611 ( .A1(n67264), .A2(n53612), .B(n54879), .C(
        n54880), .Y(n68165) );
  INVxp33_ASAP7_75t_SRAM U50612 ( .A(n76258), .Y(n54884) );
  A2O1A1Ixp33_ASAP7_75t_SL U50613 ( .A1(n62498), .A2(n54885), .B(n62499), .C(
        n62500), .Y(n54886) );
  INVxp33_ASAP7_75t_SRAM U50614 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .Y(
        n54893) );
  AOI22xp33_ASAP7_75t_SRAM U50615 ( .A1(dwb_dat_i[19]), .A2(n61548), .B1(
        n75569), .B2(dwb_dat_i[27]), .Y(n61549) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50616 ( .A1(n59526), .A2(n71223), .B(n54904), 
        .C(n71413), .Y(n71270) );
  A2O1A1Ixp33_ASAP7_75t_SL U50617 ( .A1(n71675), .A2(n71677), .B(n54918), .C(
        n71679), .Y(n54919) );
  INVxp33_ASAP7_75t_SRAM U50618 ( .A(n78149), .Y(n54921) );
  INVxp33_ASAP7_75t_SRAM U50619 ( .A(n77435), .Y(n54922) );
  INVx1_ASAP7_75t_SL U50620 ( .A(n63893), .Y(n54923) );
  INVxp33_ASAP7_75t_SRAM U50621 ( .A(n76059), .Y(n54927) );
  INVx1_ASAP7_75t_SL U50622 ( .A(dbg_dat_i[31]), .Y(n54930) );
  INVxp33_ASAP7_75t_SRAM U50623 ( .A(n74124), .Y(n54932) );
  A2O1A1Ixp33_ASAP7_75t_SL U50624 ( .A1(n54932), .A2(n54933), .B(n74125), .C(
        n54934), .Y(n78121) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50625 ( .A1(n76548), .A2(n76550), .B(n76549), 
        .C(n54935), .Y(n77964) );
  INVxp33_ASAP7_75t_SRAM U50626 ( .A(n76636), .Y(n54936) );
  FAx1_ASAP7_75t_SL U50627 ( .A(n59569), .B(n2119), .CI(n54937), .CON(), .SN(
        n77985) );
  A2O1A1Ixp33_ASAP7_75t_SL U50628 ( .A1(n69913), .A2(n69914), .B(n54940), .C(
        n69912), .Y(n69915) );
  XOR2xp5_ASAP7_75t_SL U50629 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_9_), 
        .B(n74358), .Y(n74365) );
  A2O1A1Ixp33_ASAP7_75t_SL U50630 ( .A1(n65658), .A2(n54958), .B(n65660), .C(
        n65659), .Y(n54959) );
  INVxp33_ASAP7_75t_SRAM U50631 ( .A(n70872), .Y(n54960) );
  A2O1A1Ixp33_ASAP7_75t_SL U50632 ( .A1(n70872), .A2(n54962), .B(n59698), .C(
        n54963), .Y(n54964) );
  A2O1A1Ixp33_ASAP7_75t_SL U50633 ( .A1(n54961), .A2(n54962), .B(n54963), .C(
        n54964), .Y(n54965) );
  INVx1_ASAP7_75t_SL U50634 ( .A(n70720), .Y(n54971) );
  A2O1A1Ixp33_ASAP7_75t_SL U50635 ( .A1(n70733), .A2(n70729), .B(n70715), .C(
        n57211), .Y(n54974) );
  INVxp33_ASAP7_75t_SRAM U50636 ( .A(n74727), .Y(n54987) );
  A2O1A1Ixp33_ASAP7_75t_SL U50637 ( .A1(n74730), .A2(n54987), .B(n74729), .C(
        n74728), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n56) );
  INVx1_ASAP7_75t_SL U50638 ( .A(n57137), .Y(n54988) );
  INVxp33_ASAP7_75t_SRAM U50639 ( .A(n76906), .Y(n54995) );
  INVxp33_ASAP7_75t_SRAM U50640 ( .A(n69019), .Y(n55000) );
  OAI21xp33_ASAP7_75t_SL U50641 ( .A1(n54996), .A2(n69017), .B(n54995), .Y(
        n55005) );
  A2O1A1Ixp33_ASAP7_75t_SL U50642 ( .A1(n69017), .A2(n54996), .B(n55005), .C(
        n55004), .Y(or1200_cpu_or1200_mult_mac_n1616) );
  INVxp33_ASAP7_75t_SRAM U50643 ( .A(n53440), .Y(n55009) );
  OAI22xp33_ASAP7_75t_SRAM U50644 ( .A1(n59706), .A2(n77779), .B1(n57083), 
        .B2(n1327), .Y(n1328) );
  INVx1_ASAP7_75t_SL U50645 ( .A(n77287), .Y(n55013) );
  INVxp33_ASAP7_75t_SRAM U50646 ( .A(n77286), .Y(n55017) );
  INVxp33_ASAP7_75t_SRAM U50647 ( .A(n77587), .Y(n55022) );
  O2A1O1Ixp33_ASAP7_75t_SL U50648 ( .A1(n1737), .A2(n55022), .B(n77588), .C(
        n77645), .Y(n55023) );
  INVxp33_ASAP7_75t_SRAM U50649 ( .A(n57144), .Y(n55025) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50650 ( .A1(n55039), .A2(n70477), .B(n70530), 
        .C(n27447), .Y(n55040) );
  INVxp33_ASAP7_75t_SRAM U50651 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_8_), .Y(n55042) );
  A2O1A1Ixp33_ASAP7_75t_SL U50652 ( .A1(n65400), .A2(n55041), .B(n65401), .C(
        n55044), .Y(n2478) );
  OAI22xp33_ASAP7_75t_SRAM U50653 ( .A1(n57090), .A2(n60478), .B1(n2623), .B2(
        n77454), .Y(n9594) );
  NAND2xp33_ASAP7_75t_SRAM U50654 ( .A(iwb_dat_i[2]), .B(n59496), .Y(n60346)
         );
  INVxp33_ASAP7_75t_SRAM U50655 ( .A(n74887), .Y(n55052) );
  A2O1A1Ixp33_ASAP7_75t_SL U50656 ( .A1(n77197), .A2(n55051), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_14_), .C(n55053), 
        .Y(n52490) );
  OAI22xp33_ASAP7_75t_SRAM U50657 ( .A1(n2941), .A2(n77463), .B1(n59577), .B2(
        n57073), .Y(n75436) );
  AOI21xp33_ASAP7_75t_SRAM U50658 ( .A1(or1200_cpu_spr_dat_rf[21]), .A2(n77465), .B(n75436), .Y(n75437) );
  O2A1O1Ixp33_ASAP7_75t_SL U50659 ( .A1(n75541), .A2(n55056), .B(n75543), .C(
        n55057), .Y(n55058) );
  A2O1A1Ixp33_ASAP7_75t_SL U50660 ( .A1(n63952), .A2(n55060), .B(n59695), .C(
        n55061), .Y(n3040) );
  A2O1A1Ixp33_ASAP7_75t_SL U50661 ( .A1(n3088), .A2(n77469), .B(n61318), .C(
        n61317), .Y(n55062) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50662 ( .A1(n73658), .A2(n73659), .B(n73657), 
        .C(n55066), .Y(n55067) );
  INVxp33_ASAP7_75t_SRAM U50663 ( .A(n73826), .Y(n55070) );
  INVxp33_ASAP7_75t_SRAM U50664 ( .A(n72667), .Y(n55072) );
  INVx1_ASAP7_75t_SL U50665 ( .A(n55075), .Y(n55076) );
  O2A1O1Ixp33_ASAP7_75t_SL U50666 ( .A1(n67432), .A2(n59618), .B(n55077), .C(
        n55078), .Y(n63646) );
  INVxp33_ASAP7_75t_SRAM U50667 ( .A(n64756), .Y(n55081) );
  INVxp33_ASAP7_75t_SRAM U50668 ( .A(n75039), .Y(n55085) );
  XOR2xp5_ASAP7_75t_SL U50669 ( .A(n61620), .B(n61619), .Y(n76293) );
  INVx1_ASAP7_75t_SL U50670 ( .A(n55088), .Y(n55089) );
  INVxp33_ASAP7_75t_SRAM U50671 ( .A(n71685), .Y(n55094) );
  INVx1_ASAP7_75t_SL U50672 ( .A(n55095), .Y(n71030) );
  INVxp33_ASAP7_75t_SRAM U50673 ( .A(or1200_cpu_or1200_except_n290), .Y(n55109) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50674 ( .A1(n77438), .A2(n55109), .B(n77440), 
        .C(n77430), .Y(n55110) );
  INVxp33_ASAP7_75t_SRAM U50675 ( .A(n65172), .Y(n55112) );
  INVxp33_ASAP7_75t_SRAM U50676 ( .A(n76074), .Y(n55116) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50677 ( .A1(n76076), .A2(n76088), .B(n76075), 
        .C(n55116), .Y(n76080) );
  INVxp33_ASAP7_75t_SRAM U50678 ( .A(n76122), .Y(n55117) );
  INVxp33_ASAP7_75t_SRAM U50679 ( .A(n63311), .Y(n55118) );
  INVxp33_ASAP7_75t_SRAM U50680 ( .A(n63497), .Y(n55119) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50681 ( .A1(n75298), .A2(n74981), .B(n74982), 
        .C(n55125), .Y(n78129) );
  INVxp33_ASAP7_75t_SRAM U50682 ( .A(n2966), .Y(n55126) );
  INVxp33_ASAP7_75t_SRAM U50683 ( .A(n74754), .Y(n55127) );
  INVxp33_ASAP7_75t_SRAM U50684 ( .A(n71529), .Y(n55132) );
  INVxp33_ASAP7_75t_SRAM U50685 ( .A(n66097), .Y(n55144) );
  INVxp33_ASAP7_75t_SRAM U50686 ( .A(n66147), .Y(n55145) );
  INVxp33_ASAP7_75t_SRAM U50687 ( .A(n66113), .Y(n55147) );
  INVxp33_ASAP7_75t_SRAM U50688 ( .A(n66122), .Y(n55148) );
  INVxp33_ASAP7_75t_SRAM U50689 ( .A(n66137), .Y(n55156) );
  INVxp33_ASAP7_75t_SRAM U50690 ( .A(n74253), .Y(n55157) );
  INVxp33_ASAP7_75t_SRAM U50691 ( .A(n962), .Y(n78038) );
  HAxp5_ASAP7_75t_SL U50692 ( .A(or1200_cpu_or1200_mult_mac_n259), .B(
        or1200_cpu_or1200_mult_mac_n405), .CON(), .SN(n55172) );
  INVxp33_ASAP7_75t_SRAM U50693 ( .A(n69060), .Y(n55181) );
  O2A1O1Ixp33_ASAP7_75t_SL U50694 ( .A1(n76906), .A2(n69020), .B(n55188), .C(
        n55189), .Y(n55190) );
  A2O1A1Ixp33_ASAP7_75t_SL U50695 ( .A1(n57080), .A2(n68861), .B(n55197), .C(
        n55199), .Y(n55200) );
  A2O1A1Ixp33_ASAP7_75t_SL U50696 ( .A1(or1200_cpu_or1200_mult_mac_div_cntr_2_), .A2(n76631), .B(n61811), .C(n55203), .Y(or1200_cpu_or1200_mult_mac_n1104) );
  INVxp33_ASAP7_75t_SRAM U50697 ( .A(n53440), .Y(n55204) );
  INVx1_ASAP7_75t_SL U50698 ( .A(n57142), .Y(n55208) );
  INVx1_ASAP7_75t_SL U50699 ( .A(n57142), .Y(n55211) );
  INVx1_ASAP7_75t_SL U50700 ( .A(n77675), .Y(n55217) );
  OAI22xp33_ASAP7_75t_SRAM U50701 ( .A1(n1776), .A2(n77463), .B1(n59538), .B2(
        n57074), .Y(n77230) );
  INVxp33_ASAP7_75t_SRAM U50702 ( .A(n77026), .Y(n55220) );
  INVx1_ASAP7_75t_SL U50703 ( .A(n57202), .Y(n55226) );
  INVx1_ASAP7_75t_SL U50704 ( .A(n59621), .Y(n55230) );
  INVxp33_ASAP7_75t_SRAM U50705 ( .A(n57144), .Y(n55232) );
  OAI22xp33_ASAP7_75t_SRAM U50706 ( .A1(n57090), .A2(n60487), .B1(n2630), .B2(
        n77454), .Y(n9593) );
  INVxp33_ASAP7_75t_SRAM U50707 ( .A(n2669), .Y(n55235) );
  INVx1_ASAP7_75t_SL U50708 ( .A(n60272), .Y(n55237) );
  O2A1O1Ixp33_ASAP7_75t_SL U50709 ( .A1(n2775), .A2(n77402), .B(n57084), .C(
        n55239), .Y(n78181) );
  A2O1A1Ixp33_ASAP7_75t_SL U50710 ( .A1(n77196), .A2(n77197), .B(n55240), .C(
        n77195), .Y(n52508) );
  INVxp33_ASAP7_75t_SRAM U50711 ( .A(n77457), .Y(n55241) );
  A2O1A1Ixp33_ASAP7_75t_SL U50712 ( .A1(n77462), .A2(n55242), .B(n77461), .C(
        n55243), .Y(n9458) );
  FAx1_ASAP7_75t_SL U50713 ( .A(n70104), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[0]), .CI(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[0]), .CON(), 
        .SN(n55250) );
  XOR2xp5_ASAP7_75t_SL U50714 ( .A(n70109), .B(n55250), .Y(n12874) );
  INVxp33_ASAP7_75t_SRAM U50715 ( .A(n73827), .Y(n55253) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50716 ( .A1(n73474), .A2(n73475), .B(n73476), 
        .C(n55254), .Y(n12861) );
  A2O1A1Ixp33_ASAP7_75t_SL U50717 ( .A1(n63861), .A2(n63860), .B(n57108), .C(
        n57566), .Y(n55255) );
  INVx1_ASAP7_75t_SL U50718 ( .A(n55255), .Y(n64030) );
  INVxp33_ASAP7_75t_SRAM U50719 ( .A(n58746), .Y(n55256) );
  INVxp33_ASAP7_75t_SRAM U50720 ( .A(n75076), .Y(n55259) );
  INVx1_ASAP7_75t_SL U50721 ( .A(n57110), .Y(n55262) );
  OAI21xp33_ASAP7_75t_SRAM U50722 ( .A1(n59620), .A2(n55262), .B(n59506), .Y(
        n55264) );
  A2O1A1Ixp33_ASAP7_75t_SL U50723 ( .A1(n59620), .A2(n55262), .B(n55264), .C(
        n55263), .Y(n55265) );
  INVx1_ASAP7_75t_SL U50724 ( .A(n55265), .Y(n63200) );
  INVx1_ASAP7_75t_SL U50725 ( .A(n67194), .Y(n55266) );
  INVx1_ASAP7_75t_SL U50726 ( .A(n67196), .Y(n55267) );
  NAND3xp33_ASAP7_75t_SL U50727 ( .A(n55267), .B(n67195), .C(n55266), .Y(
        n55268) );
  A2O1A1Ixp33_ASAP7_75t_SL U50728 ( .A1(n67195), .A2(n55266), .B(n55267), .C(
        n55268), .Y(n67203) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50729 ( .A1(n57120), .A2(n59549), .B(n55270), 
        .C(n66249), .Y(n61985) );
  XNOR2x2_ASAP7_75t_SL U50730 ( .A(n68621), .B(n68622), .Y(n69228) );
  O2A1O1Ixp5_ASAP7_75t_SL U50731 ( .A1(n57141), .A2(n57057), .B(n55272), .C(
        n64669), .Y(n64091) );
  INVx1_ASAP7_75t_SL U50732 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[21]), .Y(
        n55274) );
  INVx1_ASAP7_75t_SL U50733 ( .A(n74598), .Y(n55275) );
  A2O1A1Ixp33_ASAP7_75t_SL U50734 ( .A1(n57194), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[15]), .B(n55276), 
        .C(n65782), .Y(n55277) );
  INVxp33_ASAP7_75t_SRAM U50735 ( .A(n59526), .Y(n55278) );
  O2A1O1Ixp5_ASAP7_75t_SL U50736 ( .A1(n58672), .A2(n75467), .B(n55282), .C(
        n55283), .Y(n75469) );
  INVx1_ASAP7_75t_SL U50737 ( .A(n59870), .Y(n55285) );
  HAxp5_ASAP7_75t_SL U50738 ( .A(n61237), .B(n61236), .CON(), .SN(n76290) );
  INVxp33_ASAP7_75t_SRAM U50739 ( .A(n61353), .Y(n55286) );
  INVxp33_ASAP7_75t_SRAM U50740 ( .A(n75322), .Y(n55287) );
  INVx1_ASAP7_75t_SL U50741 ( .A(n61799), .Y(n55290) );
  NAND3xp33_ASAP7_75t_SL U50742 ( .A(n61676), .B(n55291), .C(n61671), .Y(
        n55292) );
  A2O1A1Ixp33_ASAP7_75t_SL U50743 ( .A1(n55291), .A2(n61676), .B(n61671), .C(
        n55292), .Y(n76307) );
  FAx1_ASAP7_75t_SL U50744 ( .A(n70189), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[6]), .CI(
        n55293), .CON(), .SN(n70197) );
  INVx1_ASAP7_75t_SL U50745 ( .A(n55294), .Y(n71081) );
  INVxp33_ASAP7_75t_SRAM U50746 ( .A(n71583), .Y(n55295) );
  INVx1_ASAP7_75t_SL U50747 ( .A(or1200_cpu_or1200_mult_mac_n357), .Y(n55309)
         );
  INVx1_ASAP7_75t_SL U50748 ( .A(dbg_dat_i[16]), .Y(n55314) );
  INVxp33_ASAP7_75t_SRAM U50749 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_3_), .Y(
        n55318) );
  INVxp33_ASAP7_75t_SRAM U50750 ( .A(n69817), .Y(n55321) );
  INVxp33_ASAP7_75t_SRAM U50751 ( .A(n66165), .Y(n55335) );
  O2A1O1Ixp33_ASAP7_75t_SL U50752 ( .A1(n72544), .A2(n72387), .B(n55349), .C(
        n55350), .Y(n55351) );
  INVxp33_ASAP7_75t_SRAM U50753 ( .A(or1200_cpu_or1200_except_n555), .Y(n55354) );
  INVxp33_ASAP7_75t_SRAM U50754 ( .A(n2691), .Y(n55357) );
  INVxp33_ASAP7_75t_SRAM U50755 ( .A(n2970), .Y(n55358) );
  A2O1A1Ixp33_ASAP7_75t_SL U50756 ( .A1(n2970), .A2(n55356), .B(n77685), .C(
        n2691), .Y(n55359) );
  A2O1A1Ixp33_ASAP7_75t_SL U50757 ( .A1(n55358), .A2(n55356), .B(n77685), .C(
        n55357), .Y(n55360) );
  NAND2xp33_ASAP7_75t_SL U50758 ( .A(n55359), .B(n55360), .Y(n55361) );
  A2O1A1Ixp33_ASAP7_75t_SL U50759 ( .A1(n55355), .A2(n55363), .B(n57343), .C(
        n55366), .Y(n55367) );
  INVxp33_ASAP7_75t_SRAM U50760 ( .A(n980), .Y(n78040) );
  INVxp33_ASAP7_75t_SRAM U50761 ( .A(or1200_cpu_or1200_mult_mac_n253), .Y(
        n55374) );
  INVxp33_ASAP7_75t_SRAM U50762 ( .A(or1200_cpu_or1200_mult_mac_n399), .Y(
        n55377) );
  AOI22xp33_ASAP7_75t_SRAM U50763 ( .A1(or1200_cpu_or1200_mult_mac_n253), .A2(
        or1200_cpu_or1200_mult_mac_n399), .B1(n55377), .B2(n55374), .Y(n55378)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U50764 ( .A1(n57080), .A2(n69310), .B(n55379), .C(
        n55381), .Y(n55382) );
  INVxp33_ASAP7_75t_SRAM U50765 ( .A(n76883), .Y(n55385) );
  INVxp33_ASAP7_75t_SRAM U50766 ( .A(n76885), .Y(n55387) );
  A2O1A1Ixp33_ASAP7_75t_SL U50767 ( .A1(n57080), .A2(n55386), .B(n55389), .C(
        n55391), .Y(n55392) );
  INVxp33_ASAP7_75t_SRAM U50768 ( .A(n63273), .Y(n55393) );
  INVxp33_ASAP7_75t_SRAM U50769 ( .A(n53440), .Y(n55413) );
  INVx1_ASAP7_75t_SL U50770 ( .A(icqmem_adr_qmem[19]), .Y(n55416) );
  A2O1A1Ixp33_ASAP7_75t_SL U50771 ( .A1(n1121), .A2(n76891), .B(n55417), .C(
        n55418), .Y(n9246) );
  INVxp33_ASAP7_75t_SRAM U50772 ( .A(n77141), .Y(n55420) );
  A2O1A1Ixp33_ASAP7_75t_SL U50773 ( .A1(n77287), .A2(n77646), .B(n55419), .C(
        n55420), .Y(or1200_pic_N62) );
  INVx1_ASAP7_75t_SL U50774 ( .A(n77287), .Y(n55421) );
  INVxp33_ASAP7_75t_SRAM U50775 ( .A(n76694), .Y(n55425) );
  INVx1_ASAP7_75t_SL U50776 ( .A(n77287), .Y(n55427) );
  INVxp33_ASAP7_75t_SRAM U50777 ( .A(n76687), .Y(n55431) );
  INVxp33_ASAP7_75t_SRAM U50778 ( .A(n2564), .Y(n75457) );
  INVxp33_ASAP7_75t_SRAM U50779 ( .A(n69344), .Y(n55440) );
  INVxp33_ASAP7_75t_SRAM U50780 ( .A(n57144), .Y(n55443) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50781 ( .A1(n55463), .A2(n65396), .B(n65400), 
        .C(n65401), .Y(n55464) );
  A2O1A1Ixp33_ASAP7_75t_SL U50782 ( .A1(n65400), .A2(n55465), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_2_), .C(n55466), .Y(
        n2480) );
  INVxp33_ASAP7_75t_SRAM U50783 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_2_), .Y(n55463) );
  INVxp33_ASAP7_75t_SRAM U50784 ( .A(n65396), .Y(n55465) );
  INVx1_ASAP7_75t_SL U50785 ( .A(n55464), .Y(n55466) );
  OAI22xp33_ASAP7_75t_SRAM U50786 ( .A1(n57090), .A2(n60488), .B1(n2637), .B2(
        n77454), .Y(n9592) );
  NAND2xp33_ASAP7_75t_SRAM U50787 ( .A(iwb_dat_i[1]), .B(n59496), .Y(n60374)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U50788 ( .A1(n53628), .A2(n77142), .B(n77401), .C(
        n55470), .Y(or1200_cpu_to_sr[4]) );
  INVxp33_ASAP7_75t_SRAM U50789 ( .A(n57144), .Y(n55471) );
  NAND3xp33_ASAP7_75t_SL U50790 ( .A(n77479), .B(n77484), .C(n77485), .Y(n9383) );
  INVx1_ASAP7_75t_SL U50791 ( .A(n73401), .Y(n55478) );
  NAND3xp33_ASAP7_75t_SL U50792 ( .A(n73378), .B(n55478), .C(n74502), .Y(
        n55479) );
  A2O1A1Ixp33_ASAP7_75t_SL U50793 ( .A1(n55478), .A2(n73378), .B(n74502), .C(
        n55479), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_27_)
         );
  INVxp33_ASAP7_75t_SRAM U50794 ( .A(n72673), .Y(n55480) );
  INVx1_ASAP7_75t_SL U50795 ( .A(n67446), .Y(n55483) );
  A2O1A1Ixp33_ASAP7_75t_SL U50796 ( .A1(n59041), .A2(n59614), .B(n64425), .C(
        n59506), .Y(n55486) );
  INVx1_ASAP7_75t_SL U50797 ( .A(n59230), .Y(n55487) );
  OAI21xp33_ASAP7_75t_SRAM U50798 ( .A1(n59662), .A2(n55487), .B(n67912), .Y(
        n55489) );
  A2O1A1Ixp33_ASAP7_75t_SL U50799 ( .A1(n59662), .A2(n55487), .B(n55489), .C(
        n55488), .Y(n68452) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50800 ( .A1(n64482), .A2(n53232), .B(n57120), 
        .C(n55490), .Y(n61947) );
  INVx1_ASAP7_75t_SL U50801 ( .A(n57682), .Y(n55491) );
  INVx1_ASAP7_75t_SL U50802 ( .A(n55492), .Y(n55493) );
  INVx1_ASAP7_75t_SL U50803 ( .A(n55495), .Y(n76437) );
  INVxp33_ASAP7_75t_SRAM U50804 ( .A(n78384), .Y(n55496) );
  INVxp33_ASAP7_75t_SRAM U50805 ( .A(n71204), .Y(n55497) );
  INVx1_ASAP7_75t_SL U50806 ( .A(or1200_cpu_or1200_mult_mac_n405), .Y(n55498)
         );
  INVxp33_ASAP7_75t_SRAM U50807 ( .A(n847), .Y(n55501) );
  INVxp33_ASAP7_75t_SRAM U50808 ( .A(n61323), .Y(n55502) );
  INVx1_ASAP7_75t_SL U50809 ( .A(n61674), .Y(n55503) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50810 ( .A1(n59559), .A2(n75227), .B(n76775), 
        .C(n59567), .Y(n55504) );
  INVx1_ASAP7_75t_SL U50811 ( .A(n63176), .Y(n55508) );
  O2A1O1Ixp33_ASAP7_75t_SL U50812 ( .A1(n71894), .A2(n72197), .B(n55519), .C(
        n55520), .Y(n72072) );
  INVxp33_ASAP7_75t_SRAM U50813 ( .A(n78000), .Y(n55525) );
  INVxp33_ASAP7_75t_SRAM U50814 ( .A(n68778), .Y(n55526) );
  INVx1_ASAP7_75t_SL U50815 ( .A(n63898), .Y(n55527) );
  INVxp33_ASAP7_75t_SRAM U50816 ( .A(n63526), .Y(n55528) );
  INVxp33_ASAP7_75t_SRAM U50817 ( .A(n75072), .Y(n55530) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50818 ( .A1(n59670), .A2(n75070), .B(n75069), 
        .C(n59116), .Y(n55532) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50819 ( .A1(n55531), .A2(n55532), .B(n75071), 
        .C(n75065), .Y(n55533) );
  INVx1_ASAP7_75t_SL U50820 ( .A(dbg_dat_i[17]), .Y(n55536) );
  INVxp33_ASAP7_75t_SRAM U50821 ( .A(n845), .Y(n55537) );
  INVxp33_ASAP7_75t_SRAM U50822 ( .A(n74652), .Y(n55539) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50823 ( .A1(n74741), .A2(n55545), .B(n55546), 
        .C(n55547), .Y(n55548) );
  INVxp33_ASAP7_75t_SRAM U50824 ( .A(n70638), .Y(n55551) );
  INVxp33_ASAP7_75t_SRAM U50825 ( .A(n71080), .Y(n55553) );
  A2O1A1Ixp33_ASAP7_75t_SL U50826 ( .A1(n71063), .A2(n71080), .B(n59698), .C(
        n55555), .Y(n55556) );
  A2O1A1Ixp33_ASAP7_75t_SL U50827 ( .A1(n71063), .A2(n55554), .B(n55555), .C(
        n55556), .Y(n55557) );
  A2O1A1Ixp33_ASAP7_75t_SL U50828 ( .A1(n70849), .A2(n55558), .B(n55559), .C(
        n55560), .Y(n55561) );
  INVxp33_ASAP7_75t_SRAM U50829 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .Y(n55573) );
  INVxp33_ASAP7_75t_SRAM U50830 ( .A(n71633), .Y(n55574) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50831 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_36_), 
        .A2(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_), .B(n71542), .C(n55575), .Y(n55576) );
  INVxp33_ASAP7_75t_SRAM U50832 ( .A(n57192), .Y(n55588) );
  O2A1O1Ixp33_ASAP7_75t_SL U50833 ( .A1(n72510), .A2(n72391), .B(n55587), .C(
        n55590), .Y(n55591) );
  A2O1A1Ixp33_ASAP7_75t_SL U50834 ( .A1(n74493), .A2(n55592), .B(n74238), .C(
        n74274), .Y(n55593) );
  INVxp33_ASAP7_75t_SRAM U50835 ( .A(n76671), .Y(n55595) );
  INVxp33_ASAP7_75t_SRAM U50836 ( .A(or1200_cpu_or1200_except_n290), .Y(n55605) );
  INVx1_ASAP7_75t_SL U50837 ( .A(n74572), .Y(n55607) );
  NAND2xp33_ASAP7_75t_SL U50838 ( .A(n57080), .B(n55609), .Y(n55610) );
  A2O1A1Ixp33_ASAP7_75t_SL U50839 ( .A1(n57080), .A2(n55609), .B(
        or1200_cpu_or1200_mult_mac_n243), .C(or1200_cpu_or1200_mult_mac_n389), 
        .Y(n55611) );
  A2O1A1Ixp33_ASAP7_75t_SL U50840 ( .A1(or1200_cpu_or1200_mult_mac_n243), .A2(
        n55610), .B(or1200_cpu_or1200_mult_mac_n389), .C(n55611), .Y(n55612)
         );
  XOR2xp5_ASAP7_75t_SL U50841 ( .A(or1200_cpu_or1200_mult_mac_n243), .B(
        or1200_cpu_or1200_mult_mac_n389), .Y(n55614) );
  INVx1_ASAP7_75t_SL U50842 ( .A(n55608), .Y(n55616) );
  A2O1A1Ixp33_ASAP7_75t_SL U50843 ( .A1(n59672), .A2(n55608), .B(n55612), .C(
        n55618), .Y(n55619) );
  INVxp33_ASAP7_75t_SRAM U50844 ( .A(n69106), .Y(n55622) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50845 ( .A1(n59671), .A2(n55624), .B(n69093), 
        .C(n55626), .Y(n55627) );
  INVxp33_ASAP7_75t_SRAM U50846 ( .A(n68940), .Y(n55633) );
  INVxp33_ASAP7_75t_SRAM U50847 ( .A(n68939), .Y(n55636) );
  A2O1A1Ixp33_ASAP7_75t_SL U50848 ( .A1(n68935), .A2(n55635), .B(n59671), .C(
        n55637), .Y(n55638) );
  A2O1A1Ixp33_ASAP7_75t_SL U50849 ( .A1(n57080), .A2(n55634), .B(n55638), .C(
        n55640), .Y(n55641) );
  INVx1_ASAP7_75t_SL U50850 ( .A(n76226), .Y(n55642) );
  INVxp33_ASAP7_75t_SRAM U50851 ( .A(n53440), .Y(n55646) );
  INVxp33_ASAP7_75t_SRAM U50852 ( .A(n1190), .Y(n78065) );
  OAI22xp33_ASAP7_75t_SRAM U50853 ( .A1(n59706), .A2(n77785), .B1(n57083), 
        .B2(n1297), .Y(n1298) );
  INVx1_ASAP7_75t_SL U50854 ( .A(n57142), .Y(n55650) );
  INVxp33_ASAP7_75t_SRAM U50855 ( .A(n76635), .Y(n55654) );
  A2O1A1Ixp33_ASAP7_75t_SL U50856 ( .A1(n76828), .A2(n77287), .B(n55653), .C(
        n55654), .Y(or1200_pic_N55) );
  INVxp33_ASAP7_75t_SRAM U50857 ( .A(n74830), .Y(n55656) );
  INVxp33_ASAP7_75t_SRAM U50858 ( .A(n1642), .Y(n76875) );
  INVx1_ASAP7_75t_SL U50859 ( .A(n74934), .Y(n55659) );
  A2O1A1Ixp33_ASAP7_75t_SL U50860 ( .A1(n77233), .A2(n1963), .B(n55663), .C(
        n55664), .Y(n18256) );
  INVx1_ASAP7_75t_SL U50861 ( .A(n57202), .Y(n55668) );
  INVxp33_ASAP7_75t_SRAM U50862 ( .A(n70289), .Y(n55671) );
  INVx1_ASAP7_75t_SL U50863 ( .A(n65257), .Y(n55672) );
  INVxp33_ASAP7_75t_SRAM U50864 ( .A(n2579), .Y(n55676) );
  OAI22xp33_ASAP7_75t_SRAM U50865 ( .A1(n57090), .A2(n60477), .B1(n3392), .B2(
        n77454), .Y(n9590) );
  NAND2xp33_ASAP7_75t_SRAM U50866 ( .A(iwb_dat_i[0]), .B(n59495), .Y(n60364)
         );
  INVxp33_ASAP7_75t_SRAM U50867 ( .A(ex_insn[28]), .Y(n55677) );
  INVxp33_ASAP7_75t_SRAM U50868 ( .A(n77388), .Y(n55683) );
  INVxp33_ASAP7_75t_SRAM U50869 ( .A(n75181), .Y(n55684) );
  A2O1A1Ixp33_ASAP7_75t_SL U50870 ( .A1(n75181), .A2(n59694), .B(n55682), .C(
        n77388), .Y(n55685) );
  A2O1A1Ixp33_ASAP7_75t_SL U50871 ( .A1(n55684), .A2(n59694), .B(n55682), .C(
        n55683), .Y(n55686) );
  NAND2xp33_ASAP7_75t_SL U50872 ( .A(n55685), .B(n55686), .Y(n2986) );
  A2O1A1Ixp33_ASAP7_75t_SL U50873 ( .A1(n75417), .A2(n59694), .B(n75416), .C(
        n55689), .Y(n55690) );
  INVx1_ASAP7_75t_SL U50874 ( .A(n77414), .Y(n55691) );
  OAI22xp33_ASAP7_75t_SRAM U50875 ( .A1(n77408), .A2(n77025), .B1(n59580), 
        .B2(n57074), .Y(n76559) );
  INVx1_ASAP7_75t_SL U50876 ( .A(n55692), .Y(n55693) );
  INVxp33_ASAP7_75t_SRAM U50877 ( .A(n72614), .Y(n55695) );
  INVx1_ASAP7_75t_SL U50878 ( .A(n73474), .Y(n55701) );
  INVx1_ASAP7_75t_SL U50879 ( .A(n55703), .Y(n55704) );
  INVx1_ASAP7_75t_SL U50880 ( .A(n59446), .Y(n55705) );
  INVx1_ASAP7_75t_SL U50881 ( .A(n59440), .Y(n55706) );
  OAI21xp33_ASAP7_75t_SRAM U50882 ( .A1(n58865), .A2(n75899), .B(n55705), .Y(
        n55708) );
  A2O1A1Ixp33_ASAP7_75t_SL U50883 ( .A1(n75899), .A2(n58865), .B(n55708), .C(
        n55707), .Y(n67159) );
  A2O1A1Ixp33_ASAP7_75t_SL U50884 ( .A1(n58851), .A2(n67457), .B(n55709), .C(
        n55710), .Y(n64889) );
  A2O1A1Ixp33_ASAP7_75t_SL U50885 ( .A1(n75045), .A2(n55711), .B(n75077), .C(
        n75075), .Y(n75053) );
  INVx1_ASAP7_75t_SL U50886 ( .A(n61947), .Y(n55712) );
  INVxp33_ASAP7_75t_SRAM U50887 ( .A(n60742), .Y(n55713) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50888 ( .A1(n60744), .A2(n55713), .B(n57082), 
        .C(n60745), .Y(n61671) );
  INVxp33_ASAP7_75t_SRAM U50889 ( .A(n61724), .Y(n55715) );
  INVx1_ASAP7_75t_SL U50890 ( .A(n55728), .Y(n63345) );
  INVxp33_ASAP7_75t_SRAM U50891 ( .A(n59922), .Y(n55729) );
  INVxp33_ASAP7_75t_SRAM U50892 ( .A(n74689), .Y(n55730) );
  INVxp33_ASAP7_75t_SRAM U50893 ( .A(n73999), .Y(n55731) );
  INVxp33_ASAP7_75t_SRAM U50894 ( .A(n61201), .Y(n55732) );
  INVx1_ASAP7_75t_SL U50895 ( .A(n70138), .Y(n55734) );
  INVxp33_ASAP7_75t_SRAM U50896 ( .A(n66024), .Y(n55736) );
  INVxp33_ASAP7_75t_SRAM U50897 ( .A(n71234), .Y(n55742) );
  INVxp33_ASAP7_75t_SRAM U50898 ( .A(n71541), .Y(n55744) );
  A2O1A1Ixp33_ASAP7_75t_SL U50899 ( .A1(n71628), .A2(n55743), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_22_), 
        .C(n55744), .Y(n71633) );
  A2O1A1Ixp33_ASAP7_75t_SL U50900 ( .A1(n74235), .A2(n74237), .B(n74234), .C(
        n74233), .Y(n55748) );
  INVx1_ASAP7_75t_SL U50901 ( .A(n3136), .Y(n55752) );
  INVx1_ASAP7_75t_SL U50902 ( .A(or1200_cpu_or1200_mult_mac_n355), .Y(n55753)
         );
  INVxp33_ASAP7_75t_SRAM U50903 ( .A(n74997), .Y(n55754) );
  INVxp33_ASAP7_75t_SRAM U50904 ( .A(n65094), .Y(n55755) );
  INVxp33_ASAP7_75t_SRAM U50905 ( .A(n63455), .Y(n55756) );
  A2O1A1Ixp33_ASAP7_75t_SL U50906 ( .A1(n63460), .A2(n63461), .B(n63458), .C(
        n55756), .Y(n63435) );
  INVxp33_ASAP7_75t_SRAM U50907 ( .A(n63384), .Y(n55757) );
  INVx1_ASAP7_75t_SL U50908 ( .A(n76060), .Y(n55758) );
  INVxp33_ASAP7_75t_SRAM U50909 ( .A(n76147), .Y(n55760) );
  INVxp33_ASAP7_75t_SRAM U50910 ( .A(n74994), .Y(n55761) );
  INVx1_ASAP7_75t_SL U50911 ( .A(dbg_dat_i[28]), .Y(n55762) );
  INVxp33_ASAP7_75t_SRAM U50912 ( .A(n75192), .Y(n55764) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50913 ( .A1(n75195), .A2(n75194), .B(n75193), 
        .C(n75192), .Y(n55766) );
  O2A1O1Ixp33_ASAP7_75t_SL U50914 ( .A1(n75196), .A2(n77175), .B(n55765), .C(
        n55766), .Y(n78076) );
  INVx1_ASAP7_75t_SL U50915 ( .A(n55768), .Y(n77494) );
  INVx1_ASAP7_75t_SL U50916 ( .A(n70200), .Y(n55769) );
  INVx1_ASAP7_75t_SL U50917 ( .A(n72605), .Y(n55770) );
  INVx1_ASAP7_75t_SL U50918 ( .A(n55780), .Y(n67544) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50919 ( .A1(n72322), .A2(n72482), .B(n57192), 
        .C(n72500), .Y(n55786) );
  A2O1A1Ixp33_ASAP7_75t_SL U50920 ( .A1(n72323), .A2(n72324), .B(n72546), .C(
        n55787), .Y(n55788) );
  INVxp33_ASAP7_75t_SRAM U50921 ( .A(n74491), .Y(n55789) );
  INVxp33_ASAP7_75t_SRAM U50922 ( .A(n74490), .Y(n55791) );
  INVxp33_ASAP7_75t_SRAM U50923 ( .A(n71799), .Y(n55797) );
  A2O1A1Ixp33_ASAP7_75t_SL U50924 ( .A1(n77248), .A2(n77445), .B(n77451), .C(
        n55804), .Y(or1200_cpu_or1200_except_n1733) );
  INVxp33_ASAP7_75t_SRAM U50925 ( .A(n881), .Y(n78029) );
  INVxp33_ASAP7_75t_SRAM U50926 ( .A(n989), .Y(n78041) );
  INVxp33_ASAP7_75t_SRAM U50927 ( .A(n1025), .Y(n78045) );
  INVxp33_ASAP7_75t_SRAM U50928 ( .A(n75652), .Y(n55805) );
  O2A1O1Ixp33_ASAP7_75t_SL U50929 ( .A1(n75141), .A2(n55805), .B(n55806), .C(
        n55810), .Y(n55811) );
  A2O1A1Ixp33_ASAP7_75t_SL U50930 ( .A1(n69213), .A2(n57079), .B(
        or1200_cpu_or1200_mult_mac_n381), .C(or1200_cpu_or1200_mult_mac_n235), 
        .Y(n55817) );
  A2O1A1Ixp33_ASAP7_75t_SL U50931 ( .A1(or1200_cpu_or1200_mult_mac_n381), .A2(
        n55816), .B(or1200_cpu_or1200_mult_mac_n235), .C(n55817), .Y(n55818)
         );
  INVxp33_ASAP7_75t_SRAM U50932 ( .A(or1200_cpu_or1200_mult_mac_n235), .Y(
        n55819) );
  INVxp33_ASAP7_75t_SRAM U50933 ( .A(n76190), .Y(n55841) );
  A2O1A1Ixp33_ASAP7_75t_SL U50934 ( .A1(or1200_cpu_or1200_mult_mac_n6), .A2(
        n76192), .B(n76191), .C(n57321), .Y(n55842) );
  A2O1A1Ixp33_ASAP7_75t_SL U50935 ( .A1(n76194), .A2(n55843), .B(n55844), .C(
        n76631), .Y(n55845) );
  OAI22xp33_ASAP7_75t_SRAM U50936 ( .A1(n59700), .A2(n77827), .B1(n57084), 
        .B2(n959), .Y(n960) );
  INVx1_ASAP7_75t_SL U50937 ( .A(n77287), .Y(n55847) );
  A2O1A1Ixp33_ASAP7_75t_SL U50938 ( .A1(n75646), .A2(n75030), .B(n75647), .C(
        n76891), .Y(n55852) );
  INVx1_ASAP7_75t_SL U50939 ( .A(n57142), .Y(n55854) );
  OAI22xp33_ASAP7_75t_SRAM U50940 ( .A1(n59706), .A2(n77782), .B1(n57083), 
        .B2(n1312), .Y(n1313) );
  A2O1A1Ixp33_ASAP7_75t_SL U50941 ( .A1(n77763), .A2(n3418), .B(n77762), .C(
        n57083), .Y(n55856) );
  INVx1_ASAP7_75t_SL U50942 ( .A(n77287), .Y(n55857) );
  INVxp33_ASAP7_75t_SRAM U50943 ( .A(n75773), .Y(n55861) );
  INVx1_ASAP7_75t_SL U50944 ( .A(n77287), .Y(n55862) );
  INVxp33_ASAP7_75t_SRAM U50945 ( .A(n76243), .Y(n55866) );
  INVxp33_ASAP7_75t_SRAM U50946 ( .A(n77671), .Y(n55870) );
  INVx1_ASAP7_75t_SL U50947 ( .A(n77761), .Y(n55872) );
  INVx1_ASAP7_75t_SL U50948 ( .A(n61126), .Y(n55876) );
  INVxp33_ASAP7_75t_SRAM U50949 ( .A(n69727), .Y(n55879) );
  INVx1_ASAP7_75t_SL U50950 ( .A(n57202), .Y(n55890) );
  INVxp33_ASAP7_75t_SRAM U50951 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_12_), .Y(n55893) );
  INVxp33_ASAP7_75t_SRAM U50952 ( .A(n2819), .Y(n55896) );
  INVxp33_ASAP7_75t_SRAM U50953 ( .A(n76950), .Y(n55902) );
  A2O1A1Ixp33_ASAP7_75t_SL U50954 ( .A1(n63980), .A2(n63967), .B(n63966), .C(
        n63965), .Y(n55904) );
  A2O1A1Ixp33_ASAP7_75t_SL U50955 ( .A1(n63982), .A2(n55904), .B(n59695), .C(
        n55905), .Y(n3031) );
  A2O1A1Ixp33_ASAP7_75t_SL U50956 ( .A1(n76840), .A2(n59690), .B(n76841), .C(
        n55908), .Y(n55909) );
  INVxp33_ASAP7_75t_SRAM U50957 ( .A(n3107), .Y(n55911) );
  NAND3x1_ASAP7_75t_SL U50958 ( .A(n60431), .B(n60430), .C(n60429), .Y(n9584)
         );
  INVxp33_ASAP7_75t_SRAM U50959 ( .A(n70575), .Y(n55918) );
  INVxp33_ASAP7_75t_SRAM U50960 ( .A(n70580), .Y(n55920) );
  A2O1A1Ixp33_ASAP7_75t_SL U50961 ( .A1(n70579), .A2(n70582), .B(n55921), .C(
        n55922), .Y(n55923) );
  A2O1A1Ixp33_ASAP7_75t_SL U50962 ( .A1(n73830), .A2(n59704), .B(n55929), .C(
        n73834), .Y(n3284) );
  INVx1_ASAP7_75t_SL U50963 ( .A(n67020), .Y(n55930) );
  INVx1_ASAP7_75t_SL U50964 ( .A(n67190), .Y(n55933) );
  NOR2x1_ASAP7_75t_SL U50965 ( .A(or1200_dc_top_tag_13_), .B(n59760), .Y(
        n59762) );
  XOR2xp5_ASAP7_75t_SL U50966 ( .A(n61978), .B(n57212), .Y(n64812) );
  INVx1_ASAP7_75t_SL U50967 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[25]), .Y(
        n55936) );
  INVx1_ASAP7_75t_SL U50968 ( .A(n73991), .Y(n55939) );
  INVxp33_ASAP7_75t_SRAM U50969 ( .A(n74007), .Y(n55940) );
  INVx1_ASAP7_75t_SL U50970 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[2]), .Y(
        n55941) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50971 ( .A1(n57185), .A2(n73265), .B(n55942), 
        .C(n55943), .Y(n73267) );
  INVxp33_ASAP7_75t_SRAM U50972 ( .A(or1200_cpu_or1200_mult_mac_n385), .Y(
        n55949) );
  INVxp33_ASAP7_75t_SRAM U50973 ( .A(n74041), .Y(n55951) );
  INVxp33_ASAP7_75t_SRAM U50974 ( .A(n62760), .Y(n55954) );
  INVxp33_ASAP7_75t_SRAM U50975 ( .A(n75548), .Y(n55955) );
  INVxp33_ASAP7_75t_SRAM U50976 ( .A(n77082), .Y(n55956) );
  OAI21xp33_ASAP7_75t_SL U50977 ( .A1(or1200_cpu_or1200_except_n532), .A2(
        n55956), .B(n55955), .Y(n55957) );
  A2O1A1Ixp33_ASAP7_75t_SL U50978 ( .A1(n77082), .A2(
        or1200_cpu_or1200_except_n532), .B(n55955), .C(n55957), .Y(n64330) );
  INVx1_ASAP7_75t_SL U50979 ( .A(n67534), .Y(n55959) );
  INVx1_ASAP7_75t_SL U50980 ( .A(n71145), .Y(n55965) );
  INVxp33_ASAP7_75t_SRAM U50981 ( .A(n72595), .Y(n55972) );
  INVx1_ASAP7_75t_SL U50982 ( .A(or1200_cpu_or1200_mult_mac_n371), .Y(n55975)
         );
  INVxp33_ASAP7_75t_SRAM U50983 ( .A(n68992), .Y(n55976) );
  INVxp33_ASAP7_75t_SRAM U50984 ( .A(n68816), .Y(n55979) );
  INVxp33_ASAP7_75t_SRAM U50985 ( .A(n63530), .Y(n55980) );
  INVxp33_ASAP7_75t_SRAM U50986 ( .A(n63345), .Y(n55981) );
  HAxp5_ASAP7_75t_SL U50987 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_4_), .B(n74143), 
        .CON(), .SN(n55991) );
  INVx1_ASAP7_75t_SL U50988 ( .A(n58919), .Y(n55996) );
  INVx1_ASAP7_75t_SL U50989 ( .A(n76009), .Y(n55997) );
  INVx1_ASAP7_75t_SL U50990 ( .A(n62609), .Y(n55998) );
  INVxp33_ASAP7_75t_SRAM U50991 ( .A(n66075), .Y(n55999) );
  INVxp33_ASAP7_75t_SRAM U50992 ( .A(n59699), .Y(n56000) );
  OAI21xp33_ASAP7_75t_SRAM U50993 ( .A1(n59699), .A2(n71110), .B(n71109), .Y(
        n56001) );
  A2O1A1Ixp33_ASAP7_75t_SL U50994 ( .A1(n71110), .A2(n56000), .B(n71109), .C(
        n56001), .Y(n56002) );
  INVxp33_ASAP7_75t_SRAM U50995 ( .A(n70967), .Y(n56003) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U50996 ( .A1(n56003), .A2(n70906), .B(n70982), 
        .C(n59699), .Y(n56004) );
  OAI31xp33_ASAP7_75t_SL U50997 ( .A1(n70982), .A2(n56003), .A3(n70906), .B(
        n56004), .Y(n56005) );
  INVxp33_ASAP7_75t_SRAM U50998 ( .A(n71467), .Y(n56006) );
  A2O1A1Ixp33_ASAP7_75t_SL U50999 ( .A1(n71787), .A2(n71786), .B(n71793), .C(
        n71785), .Y(n56007) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51000 ( .A1(n72279), .A2(n72280), .B(n72495), 
        .C(n56022), .Y(n56023) );
  NAND2xp5_ASAP7_75t_SL U51001 ( .A(n59687), .B(n78068), .Y(n565) );
  INVxp33_ASAP7_75t_SRAM U51002 ( .A(n863), .Y(n78027) );
  INVxp33_ASAP7_75t_SRAM U51003 ( .A(n872), .Y(n78028) );
  A2O1A1Ixp33_ASAP7_75t_SL U51004 ( .A1(n75141), .A2(n75661), .B(n75660), .C(
        n57079), .Y(n56039) );
  INVxp33_ASAP7_75t_SRAM U51005 ( .A(n65073), .Y(n56050) );
  INVxp33_ASAP7_75t_SRAM U51006 ( .A(n65131), .Y(n56052) );
  A2O1A1Ixp33_ASAP7_75t_SL U51007 ( .A1(n57080), .A2(n56051), .B(n56054), .C(
        n56056), .Y(n56057) );
  A2O1A1Ixp33_ASAP7_75t_SL U51008 ( .A1(n63297), .A2(n63298), .B(n63296), .C(
        n63299), .Y(n56064) );
  FAx1_ASAP7_75t_SL U51009 ( .A(n53466), .B(n63476), .CI(n63477), .CON(), .SN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N13) );
  XOR2xp5_ASAP7_75t_SL U51010 ( .A(n63686), .B(n63685), .Y(n56065) );
  INVx1_ASAP7_75t_SL U51011 ( .A(n56065), .Y(n56067) );
  A2O1A1Ixp33_ASAP7_75t_SL U51012 ( .A1(n58281), .A2(n63257), .B(n56066), .C(
        n56068), .Y(n52050) );
  INVxp33_ASAP7_75t_SRAM U51013 ( .A(n53440), .Y(n56069) );
  INVx1_ASAP7_75t_SL U51014 ( .A(icqmem_adr_qmem[18]), .Y(n56072) );
  INVx1_ASAP7_75t_SL U51015 ( .A(icqmem_adr_qmem[24]), .Y(n56073) );
  INVxp33_ASAP7_75t_SRAM U51016 ( .A(n1125), .Y(n56074) );
  A2O1A1Ixp33_ASAP7_75t_SL U51017 ( .A1(n75029), .A2(n56075), .B(n75647), .C(
        n56076), .Y(n9248) );
  OAI22xp33_ASAP7_75t_SRAM U51018 ( .A1(n59706), .A2(n77783), .B1(n57083), 
        .B2(n1307), .Y(n1308) );
  INVx1_ASAP7_75t_SL U51019 ( .A(n57142), .Y(n56078) );
  INVxp33_ASAP7_75t_SRAM U51020 ( .A(n77761), .Y(n56084) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51021 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n70389), .B(n56105), .C(n70483), .Y(n56106) );
  INVxp33_ASAP7_75t_SRAM U51022 ( .A(n61155), .Y(n56115) );
  A2O1A1Ixp33_ASAP7_75t_SL U51023 ( .A1(n74845), .A2(n56119), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_5_), .C(n56120), 
        .Y(n52493) );
  A2O1A1Ixp33_ASAP7_75t_SL U51024 ( .A1(n63995), .A2(n63996), .B(n64001), .C(
        n59694), .Y(n56121) );
  OAI22xp33_ASAP7_75t_SRAM U51025 ( .A1(n3068), .A2(n59679), .B1(n59581), .B2(
        n57074), .Y(n76808) );
  INVxp33_ASAP7_75t_SRAM U51026 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[1]), .Y(
        n56127) );
  A2O1A1Ixp33_ASAP7_75t_SL U51027 ( .A1(n71539), .A2(n78383), .B(n56131), .C(
        n71538), .Y(n3265) );
  INVx1_ASAP7_75t_SL U51028 ( .A(n71519), .Y(n56132) );
  A2O1A1Ixp33_ASAP7_75t_SL U51029 ( .A1(n71518), .A2(n56132), .B(n71520), .C(
        n56133), .Y(n12875) );
  INVxp33_ASAP7_75t_SRAM U51030 ( .A(n73651), .Y(n56134) );
  A2O1A1Ixp33_ASAP7_75t_SL U51031 ( .A1(n73835), .A2(n59704), .B(n56135), .C(
        n73834), .Y(n3283) );
  A2O1A1Ixp33_ASAP7_75t_SL U51032 ( .A1(n73472), .A2(n73477), .B(n73473), .C(
        n56136), .Y(n21879) );
  INVxp33_ASAP7_75t_SRAM U51033 ( .A(n72676), .Y(n56137) );
  INVx1_ASAP7_75t_SL U51034 ( .A(n66720), .Y(n56140) );
  INVx1_ASAP7_75t_SL U51035 ( .A(n66481), .Y(n56143) );
  INVxp33_ASAP7_75t_SRAM U51036 ( .A(n66288), .Y(n56145) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51037 ( .A1(n59548), .A2(n57120), .B(n56144), 
        .C(n56145), .Y(n61982) );
  XNOR2x1_ASAP7_75t_SL U51038 ( .A(n64554), .B(n64552), .Y(n57555) );
  O2A1O1Ixp33_ASAP7_75t_SL U51039 ( .A1(n59614), .A2(n57394), .B(n56146), .C(
        n68079), .Y(n68080) );
  INVxp33_ASAP7_75t_SRAM U51040 ( .A(n75103), .Y(n56147) );
  O2A1O1Ixp33_ASAP7_75t_SL U51041 ( .A1(n75106), .A2(n75105), .B(n75104), .C(
        n56147), .Y(n75114) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51042 ( .A1(n59807), .A2(n69356), .B(
        or1200_dc_top_tag_12_), .C(n59806), .Y(n59808) );
  INVxp33_ASAP7_75t_SRAM U51043 ( .A(n72928), .Y(n56148) );
  INVxp33_ASAP7_75t_SRAM U51044 ( .A(n73986), .Y(n56149) );
  INVx1_ASAP7_75t_SL U51045 ( .A(or1200_cpu_or1200_mult_mac_n407), .Y(n56151)
         );
  INVxp33_ASAP7_75t_SRAM U51046 ( .A(n69140), .Y(n56155) );
  O2A1O1Ixp33_ASAP7_75t_SL U51047 ( .A1(n76765), .A2(n61353), .B(n56158), .C(
        n75872), .Y(n61089) );
  XNOR2xp5_ASAP7_75t_SL U51048 ( .A(n61400), .B(n56159), .Y(n76295) );
  AOI22xp33_ASAP7_75t_SRAM U51049 ( .A1(n75570), .A2(
        or1200_dc_top_from_dcram_21_), .B1(dwb_dat_i[21]), .B2(n75569), .Y(
        n61625) );
  INVxp33_ASAP7_75t_SRAM U51050 ( .A(n3095), .Y(n56160) );
  A2O1A1Ixp33_ASAP7_75t_SL U51051 ( .A1(n59442), .A2(n61492), .B(n61876), .C(
        n56161), .Y(n77102) );
  INVxp33_ASAP7_75t_SRAM U51052 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[2]), .Y(
        n56162) );
  INVxp33_ASAP7_75t_SRAM U51053 ( .A(n71682), .Y(n56164) );
  INVx1_ASAP7_75t_SL U51054 ( .A(n56171), .Y(n71297) );
  INVx1_ASAP7_75t_SL U51055 ( .A(n71020), .Y(n56172) );
  INVxp33_ASAP7_75t_SRAM U51056 ( .A(or1200_cpu_or1200_mult_mac_n395), .Y(
        n56197) );
  INVxp33_ASAP7_75t_SRAM U51057 ( .A(n69173), .Y(n56200) );
  INVxp33_ASAP7_75t_SRAM U51058 ( .A(n68942), .Y(n56201) );
  INVxp33_ASAP7_75t_SRAM U51059 ( .A(or1200_cpu_or1200_mult_mac_n185), .Y(
        n56202) );
  INVxp33_ASAP7_75t_SRAM U51060 ( .A(n63432), .Y(n56203) );
  INVxp33_ASAP7_75t_SRAM U51061 ( .A(n76098), .Y(n56204) );
  INVxp33_ASAP7_75t_SRAM U51062 ( .A(n68957), .Y(n56205) );
  INVxp33_ASAP7_75t_SRAM U51063 ( .A(n57398), .Y(n56206) );
  INVx1_ASAP7_75t_SL U51064 ( .A(dbg_dat_i[29]), .Y(n56212) );
  INVxp33_ASAP7_75t_SRAM U51065 ( .A(n69365), .Y(n56214) );
  INVxp33_ASAP7_75t_SRAM U51066 ( .A(n74702), .Y(n56218) );
  INVxp33_ASAP7_75t_SRAM U51067 ( .A(n70010), .Y(n56223) );
  INVxp33_ASAP7_75t_SRAM U51068 ( .A(n69785), .Y(n56224) );
  INVxp33_ASAP7_75t_SRAM U51069 ( .A(n66080), .Y(n56227) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51070 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_1_), .A2(n59697), 
        .B(n56228), .C(n70690), .Y(n56229) );
  INVxp33_ASAP7_75t_SRAM U51071 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_1_), .Y(n56231) );
  INVxp33_ASAP7_75t_SRAM U51072 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_0_), .Y(
        n56233) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51073 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39), .A2(n56233), .B(n74063), .C(n74097), .Y(n56234) );
  INVxp33_ASAP7_75t_SRAM U51074 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39), .Y(n56235) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51075 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_0_), .A2(
        n56235), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_1_), .C(
        n74098), .Y(n56236) );
  INVxp33_ASAP7_75t_SRAM U51076 ( .A(n908), .Y(n78032) );
  INVxp33_ASAP7_75t_SRAM U51077 ( .A(n935), .Y(n78035) );
  INVxp33_ASAP7_75t_SRAM U51078 ( .A(n953), .Y(n78037) );
  INVxp33_ASAP7_75t_SRAM U51079 ( .A(n998), .Y(n78042) );
  NAND2xp33_ASAP7_75t_SRAM U51080 ( .A(n57079), .B(n75118), .Y(n56246) );
  A2O1A1Ixp33_ASAP7_75t_SL U51081 ( .A1(n57079), .A2(n75118), .B(
        or1200_cpu_or1200_mult_mac_n257), .C(or1200_cpu_or1200_mult_mac_n403), 
        .Y(n56247) );
  A2O1A1Ixp33_ASAP7_75t_SL U51082 ( .A1(or1200_cpu_or1200_mult_mac_n257), .A2(
        n56246), .B(or1200_cpu_or1200_mult_mac_n403), .C(n56247), .Y(n56248)
         );
  XOR2xp5_ASAP7_75t_SL U51083 ( .A(or1200_cpu_or1200_mult_mac_n257), .B(
        or1200_cpu_or1200_mult_mac_n403), .Y(n56250) );
  INVxp33_ASAP7_75t_SRAM U51084 ( .A(n63535), .Y(n56255) );
  INVx1_ASAP7_75t_SL U51085 ( .A(n76633), .Y(n56268) );
  INVxp33_ASAP7_75t_SRAM U51086 ( .A(n76148), .Y(n56271) );
  AOI21xp33_ASAP7_75t_SRAM U51087 ( .A1(n76146), .A2(n58753), .B(n56271), .Y(
        n56272) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51088 ( .A1(n76146), .A2(n58753), .B(n56272), 
        .C(n76150), .Y(n56273) );
  INVxp33_ASAP7_75t_SRAM U51089 ( .A(n63368), .Y(n56278) );
  FAx1_ASAP7_75t_SL U51090 ( .A(n63367), .B(n56277), .CI(n56278), .CON(), .SN(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N9) );
  NOR3xp33_ASAP7_75t_SL U51091 ( .A(n65104), .B(n56279), .C(n64700), .Y(n56280) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51092 ( .A1(n65104), .A2(n64700), .B(n56279), 
        .C(n56280), .Y(n56281) );
  INVx1_ASAP7_75t_SL U51093 ( .A(n56281), .Y(n52052) );
  OAI22xp33_ASAP7_75t_SRAM U51094 ( .A1(n59700), .A2(n77816), .B1(n57084), 
        .B2(n860), .Y(n861) );
  OAI22xp33_ASAP7_75t_SRAM U51095 ( .A1(n59700), .A2(n77817), .B1(n57084), 
        .B2(n869), .Y(n870) );
  INVx1_ASAP7_75t_SL U51096 ( .A(icqmem_adr_qmem[16]), .Y(n56282) );
  INVx1_ASAP7_75t_SL U51097 ( .A(icqmem_adr_qmem[17]), .Y(n56283) );
  OAI22xp33_ASAP7_75t_SRAM U51098 ( .A1(n59700), .A2(n77823), .B1(n57084), 
        .B2(n923), .Y(n924) );
  OAI22xp33_ASAP7_75t_SRAM U51099 ( .A1(n59700), .A2(n77825), .B1(n57084), 
        .B2(n941), .Y(n942) );
  OAI22xp33_ASAP7_75t_SRAM U51100 ( .A1(n59700), .A2(n77829), .B1(n57084), 
        .B2(n1013), .Y(n1014) );
  OAI22xp33_ASAP7_75t_SRAM U51101 ( .A1(n59706), .A2(n77778), .B1(n57083), 
        .B2(n1332), .Y(n1333) );
  INVx1_ASAP7_75t_SL U51102 ( .A(n77287), .Y(n56284) );
  INVx1_ASAP7_75t_SL U51103 ( .A(pic_ints_i[1]), .Y(n56288) );
  INVxp33_ASAP7_75t_SRAM U51104 ( .A(n1520), .Y(n56290) );
  INVxp33_ASAP7_75t_SRAM U51105 ( .A(n72696), .Y(n56291) );
  INVxp33_ASAP7_75t_SRAM U51106 ( .A(n77761), .Y(n56296) );
  INVx1_ASAP7_75t_SL U51107 ( .A(n75148), .Y(n56301) );
  INVxp33_ASAP7_75t_SRAM U51108 ( .A(n2394), .Y(n56303) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51109 ( .A1(n74706), .A2(n70536), .B(n56307), 
        .C(n70535), .Y(n56308) );
  INVxp33_ASAP7_75t_SRAM U51110 ( .A(n61153), .Y(n56321) );
  OAI22xp33_ASAP7_75t_SRAM U51111 ( .A1(n57090), .A2(n60479), .B1(n2644), .B2(
        n77454), .Y(n9591) );
  INVxp33_ASAP7_75t_SRAM U51112 ( .A(n3068), .Y(n77280) );
  INVxp33_ASAP7_75t_SRAM U51113 ( .A(n2853), .Y(n56326) );
  A2O1A1Ixp33_ASAP7_75t_SL U51114 ( .A1(n74845), .A2(n74844), .B(n56330), .C(
        n77195), .Y(n52492) );
  FAx1_ASAP7_75t_SL U51115 ( .A(n65219), .B(id_insn_22_), .CI(
        or1200_cpu_or1200_except_n649), .CON(), .SN(n56331) );
  XOR2xp5_ASAP7_75t_SL U51116 ( .A(n2098), .B(n63967), .Y(n56338) );
  INVx1_ASAP7_75t_SL U51117 ( .A(n56338), .Y(n56339) );
  A2O1A1Ixp33_ASAP7_75t_SL U51118 ( .A1(n59693), .A2(n56338), .B(
        or1200_cpu_or1200_except_n613), .C(n56341), .Y(n56342) );
  A2O1A1Ixp33_ASAP7_75t_SL U51119 ( .A1(n76588), .A2(n76589), .B(n76587), .C(
        n59694), .Y(n56343) );
  INVxp33_ASAP7_75t_SRAM U51120 ( .A(n57090), .Y(n56344) );
  INVxp33_ASAP7_75t_SRAM U51121 ( .A(n77368), .Y(n56350) );
  INVxp33_ASAP7_75t_SRAM U51122 ( .A(n71530), .Y(n56356) );
  NOR3xp33_ASAP7_75t_SL U51123 ( .A(n73399), .B(n73400), .C(n73398), .Y(n56359) );
  O2A1O1Ixp33_ASAP7_75t_SL U51124 ( .A1(n73399), .A2(n73398), .B(n73400), .C(
        n56359), .Y(n78218) );
  INVxp33_ASAP7_75t_SRAM U51125 ( .A(n66373), .Y(n56360) );
  INVxp33_ASAP7_75t_SRAM U51126 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[3]), .Y(n56365)
         );
  NAND2xp33_ASAP7_75t_SRAM U51127 ( .A(n59815), .B(n75299), .Y(n59819) );
  INVxp33_ASAP7_75t_SRAM U51128 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[10]), .Y(n56368) );
  INVx1_ASAP7_75t_SL U51129 ( .A(n53430), .Y(n56369) );
  INVxp33_ASAP7_75t_SRAM U51130 ( .A(n71390), .Y(n56376) );
  INVxp33_ASAP7_75t_SRAM U51131 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_39_), .Y(n56377) );
  XOR2x2_ASAP7_75t_SL U51132 ( .A(n68494), .B(n58358), .Y(n68520) );
  INVxp33_ASAP7_75t_SRAM U51133 ( .A(n75278), .Y(n56379) );
  INVxp33_ASAP7_75t_SRAM U51134 ( .A(n1145), .Y(n56381) );
  INVx1_ASAP7_75t_SL U51135 ( .A(n72943), .Y(n56382) );
  INVx1_ASAP7_75t_SL U51136 ( .A(n56383), .Y(n76433) );
  INVxp33_ASAP7_75t_SRAM U51137 ( .A(n67213), .Y(n56388) );
  INVx1_ASAP7_75t_SL U51138 ( .A(n56389), .Y(n68263) );
  OAI21xp33_ASAP7_75t_SL U51139 ( .A1(n53221), .A2(n57110), .B(n56390), .Y(
        n56393) );
  A2O1A1Ixp33_ASAP7_75t_SL U51140 ( .A1(n57110), .A2(n53221), .B(n56393), .C(
        n56392), .Y(n67295) );
  INVx1_ASAP7_75t_SL U51141 ( .A(n56398), .Y(n71029) );
  INVxp33_ASAP7_75t_SRAM U51142 ( .A(n70803), .Y(n56399) );
  INVxp33_ASAP7_75t_SRAM U51143 ( .A(n69246), .Y(n56405) );
  INVx1_ASAP7_75t_SL U51144 ( .A(n74569), .Y(n56406) );
  INVxp33_ASAP7_75t_SRAM U51145 ( .A(n69112), .Y(n56407) );
  INVxp33_ASAP7_75t_SRAM U51146 ( .A(n68988), .Y(n56408) );
  INVxp33_ASAP7_75t_SRAM U51147 ( .A(n68876), .Y(n56409) );
  INVxp33_ASAP7_75t_SRAM U51148 ( .A(n63487), .Y(n56411) );
  INVxp33_ASAP7_75t_SRAM U51149 ( .A(n63337), .Y(n56412) );
  INVx1_ASAP7_75t_SL U51150 ( .A(n69098), .Y(n56413) );
  A2O1A1Ixp33_ASAP7_75t_SL U51151 ( .A1(n59637), .A2(n75466), .B(n56414), .C(
        n59635), .Y(n56415) );
  INVx1_ASAP7_75t_SL U51152 ( .A(dbg_dat_i[27]), .Y(n56416) );
  INVx1_ASAP7_75t_SL U51153 ( .A(dbg_dat_i[22]), .Y(n56417) );
  INVxp33_ASAP7_75t_SRAM U51154 ( .A(n74666), .Y(n56419) );
  INVxp33_ASAP7_75t_SRAM U51155 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[25]), .Y(n56422) );
  INVxp33_ASAP7_75t_SRAM U51156 ( .A(n69958), .Y(n56423) );
  INVx1_ASAP7_75t_SL U51157 ( .A(n77416), .Y(n56424) );
  INVxp33_ASAP7_75t_SRAM U51158 ( .A(n70123), .Y(n56426) );
  INVxp33_ASAP7_75t_SRAM U51159 ( .A(n71536), .Y(n56428) );
  A2O1A1Ixp33_ASAP7_75t_SL U51160 ( .A1(n57205), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[18]), .B(n56431), .C(
        n56432), .Y(n73763) );
  INVxp33_ASAP7_75t_SRAM U51161 ( .A(n66081), .Y(n56433) );
  A2O1A1Ixp33_ASAP7_75t_SL U51162 ( .A1(n58302), .A2(n56434), .B(n59699), .C(
        n70703), .Y(n56435) );
  A2O1A1Ixp33_ASAP7_75t_SL U51163 ( .A1(n70694), .A2(n56434), .B(n70703), .C(
        n56435), .Y(n56436) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51164 ( .A1(n72544), .A2(n72404), .B(n56452), 
        .C(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .Y(
        n56453) );
  A2O1A1Ixp33_ASAP7_75t_SL U51165 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .A2(
        n72369), .B(n56453), .C(n56454), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n58) );
  INVxp33_ASAP7_75t_SRAM U51166 ( .A(n835), .Y(n77510) );
  NAND2xp33_ASAP7_75t_SRAM U51167 ( .A(n77510), .B(n57189), .Y(n8750) );
  INVxp33_ASAP7_75t_SRAM U51168 ( .A(n1007), .Y(n78043) );
  INVxp33_ASAP7_75t_SRAM U51169 ( .A(n65132), .Y(n56490) );
  A2O1A1Ixp33_ASAP7_75t_SL U51170 ( .A1(n57080), .A2(n65126), .B(n56492), .C(
        n56494), .Y(n56495) );
  INVxp33_ASAP7_75t_SRAM U51171 ( .A(or1200_cpu_or1200_mult_mac_div_cntr_0_), 
        .Y(n56496) );
  INVxp33_ASAP7_75t_SRAM U51172 ( .A(n63365), .Y(n56503) );
  A2O1A1Ixp33_ASAP7_75t_SL U51173 ( .A1(n63364), .A2(n56506), .B(n57044), .C(
        n56507), .Y(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N10) );
  XOR2x2_ASAP7_75t_SL U51174 ( .A(n63481), .B(n63482), .Y(n56508) );
  A2O1A1Ixp33_ASAP7_75t_SL U51175 ( .A1(n57245), .A2(n56509), .B(n56508), .C(
        n56510), .Y(or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N15) );
  INVxp33_ASAP7_75t_SRAM U51176 ( .A(n64699), .Y(n56512) );
  A2O1A1Ixp33_ASAP7_75t_SL U51177 ( .A1(n63886), .A2(n63885), .B(n56511), .C(
        n56513), .Y(n52051) );
  NAND3xp33_ASAP7_75t_SL U51178 ( .A(n68345), .B(n68761), .C(n68337), .Y(
        n56514) );
  A2O1A1Ixp33_ASAP7_75t_SL U51179 ( .A1(n68761), .A2(n68345), .B(n68337), .C(
        n56514), .Y(n52056) );
  INVx1_ASAP7_75t_SL U51180 ( .A(icqmem_adr_qmem[14]), .Y(n56515) );
  OAI22xp33_ASAP7_75t_SRAM U51181 ( .A1(n59700), .A2(n77818), .B1(n57084), 
        .B2(n878), .Y(n879) );
  OAI22xp33_ASAP7_75t_SRAM U51182 ( .A1(n59700), .A2(n77819), .B1(n57084), 
        .B2(n887), .Y(n888) );
  OAI22xp33_ASAP7_75t_SRAM U51183 ( .A1(n59700), .A2(n77821), .B1(n57084), 
        .B2(n905), .Y(n906) );
  INVx1_ASAP7_75t_SL U51184 ( .A(icqmem_adr_qmem[20]), .Y(n56516) );
  OAI22xp33_ASAP7_75t_SRAM U51185 ( .A1(n59700), .A2(n77824), .B1(n57084), 
        .B2(n932), .Y(n933) );
  OAI22xp33_ASAP7_75t_SRAM U51186 ( .A1(n59700), .A2(n77826), .B1(n57084), 
        .B2(n950), .Y(n951) );
  OAI22xp33_ASAP7_75t_SRAM U51187 ( .A1(n59700), .A2(n77828), .B1(n57084), 
        .B2(n977), .Y(n978) );
  INVx1_ASAP7_75t_SL U51188 ( .A(icqmem_adr_qmem[28]), .Y(n56517) );
  INVx1_ASAP7_75t_SL U51189 ( .A(icqmem_adr_qmem[30]), .Y(n56518) );
  OAI22xp33_ASAP7_75t_SRAM U51190 ( .A1(n59700), .A2(n77830), .B1(n57084), 
        .B2(n1022), .Y(n1023) );
  INVxp33_ASAP7_75t_SRAM U51191 ( .A(n2843), .Y(n56519) );
  A2O1A1Ixp33_ASAP7_75t_SL U51192 ( .A1(n59687), .A2(n56519), .B(n56520), .C(
        n57083), .Y(n56521) );
  INVx1_ASAP7_75t_SL U51193 ( .A(n57142), .Y(n56523) );
  INVx1_ASAP7_75t_SL U51194 ( .A(n57142), .Y(n56526) );
  OAI22xp33_ASAP7_75t_SRAM U51195 ( .A1(n59706), .A2(n77780), .B1(n57083), 
        .B2(n1322), .Y(n1323) );
  INVx1_ASAP7_75t_SL U51196 ( .A(n57142), .Y(n56529) );
  INVx1_ASAP7_75t_SL U51197 ( .A(n77287), .Y(n56533) );
  INVx1_ASAP7_75t_SL U51198 ( .A(n77287), .Y(n56539) );
  INVx1_ASAP7_75t_SL U51199 ( .A(n77287), .Y(n56544) );
  INVxp33_ASAP7_75t_SRAM U51200 ( .A(n77010), .Y(n56548) );
  INVx1_ASAP7_75t_SL U51201 ( .A(n77287), .Y(n56549) );
  INVxp33_ASAP7_75t_SRAM U51202 ( .A(n76197), .Y(n56553) );
  INVxp33_ASAP7_75t_SRAM U51203 ( .A(n1631), .Y(n56557) );
  INVxp33_ASAP7_75t_SRAM U51204 ( .A(n1645), .Y(n56559) );
  INVxp33_ASAP7_75t_SRAM U51205 ( .A(n1661), .Y(n56560) );
  INVxp33_ASAP7_75t_SRAM U51206 ( .A(n1677), .Y(n56561) );
  INVxp33_ASAP7_75t_SRAM U51207 ( .A(n1695), .Y(n56562) );
  INVx1_ASAP7_75t_SL U51208 ( .A(n56568), .Y(n56569) );
  INVx1_ASAP7_75t_SL U51209 ( .A(n59621), .Y(n56576) );
  INVxp33_ASAP7_75t_SRAM U51210 ( .A(n69756), .Y(n56578) );
  A2O1A1Ixp33_ASAP7_75t_SL U51211 ( .A1(n69772), .A2(n56578), .B(n69790), .C(
        n59621), .Y(n56579) );
  INVxp33_ASAP7_75t_SRAM U51212 ( .A(n2322), .Y(n56583) );
  INVxp33_ASAP7_75t_SRAM U51213 ( .A(n2326), .Y(n56584) );
  INVxp33_ASAP7_75t_SRAM U51214 ( .A(n2338), .Y(n56585) );
  INVxp33_ASAP7_75t_SRAM U51215 ( .A(n2342), .Y(n56586) );
  INVxp33_ASAP7_75t_SRAM U51216 ( .A(n2348), .Y(n56587) );
  INVxp33_ASAP7_75t_SRAM U51217 ( .A(n2352), .Y(n56588) );
  INVxp33_ASAP7_75t_SRAM U51218 ( .A(n2362), .Y(n56589) );
  INVxp33_ASAP7_75t_SRAM U51219 ( .A(n2368), .Y(n56590) );
  INVxp33_ASAP7_75t_SRAM U51220 ( .A(n2378), .Y(n56591) );
  INVxp33_ASAP7_75t_SRAM U51221 ( .A(n2388), .Y(n56592) );
  INVxp33_ASAP7_75t_SRAM U51222 ( .A(n2404), .Y(n56593) );
  INVxp33_ASAP7_75t_SRAM U51223 ( .A(n2423), .Y(n56594) );
  INVxp33_ASAP7_75t_SRAM U51224 ( .A(n2427), .Y(n56595) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51225 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .A2(
        n70548), .B(n70547), .C(n56596), .Y(n56597) );
  INVxp33_ASAP7_75t_SRAM U51226 ( .A(n62022), .Y(n56607) );
  INVxp33_ASAP7_75t_SRAM U51227 ( .A(n57072), .Y(n56608) );
  INVxp33_ASAP7_75t_SRAM U51228 ( .A(n76991), .Y(n56611) );
  A2O1A1Ixp33_ASAP7_75t_SL U51229 ( .A1(n2794), .A2(n56612), .B(n59680), .C(
        n56613), .Y(n76992) );
  INVxp33_ASAP7_75t_SRAM U51230 ( .A(n2824), .Y(n56615) );
  INVx1_ASAP7_75t_SL U51231 ( .A(n57202), .Y(n56618) );
  INVxp33_ASAP7_75t_SRAM U51232 ( .A(n2549), .Y(n73954) );
  INVxp33_ASAP7_75t_SRAM U51233 ( .A(n77170), .Y(n56621) );
  INVxp33_ASAP7_75t_SRAM U51234 ( .A(n1615), .Y(n56622) );
  INVx1_ASAP7_75t_SL U51235 ( .A(n57202), .Y(n56624) );
  FAx1_ASAP7_75t_SL U51236 ( .A(n2685), .B(or1200_cpu_or1200_except_n643), 
        .CI(n75542), .CON(), .SN(n56627) );
  A2O1A1Ixp33_ASAP7_75t_SL U51237 ( .A1(n64009), .A2(n64010), .B(n64012), .C(
        n59694), .Y(n56629) );
  A2O1A1Ixp33_ASAP7_75t_SL U51238 ( .A1(n76601), .A2(n76602), .B(n76600), .C(
        n59694), .Y(n56630) );
  A2O1A1Ixp33_ASAP7_75t_SL U51239 ( .A1(n76578), .A2(n76579), .B(n76577), .C(
        n59694), .Y(n56631) );
  INVxp33_ASAP7_75t_SRAM U51240 ( .A(n57072), .Y(n56632) );
  O2A1O1Ixp33_ASAP7_75t_SL U51241 ( .A1(n77364), .A2(n56641), .B(n56642), .C(
        n56643), .Y(n9195) );
  XNOR2xp5_ASAP7_75t_SL U51242 ( .A(n78244), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .Y(n56826) );
  INVxp33_ASAP7_75t_SRAM U51243 ( .A(n73465), .Y(n56646) );
  XOR2xp5_ASAP7_75t_SL U51244 ( .A(n73458), .B(n73457), .Y(n56648) );
  A2O1A1Ixp33_ASAP7_75t_SL U51245 ( .A1(n73460), .A2(n56647), .B(n56648), .C(
        n56649), .Y(n53189) );
  INVxp33_ASAP7_75t_SRAM U51246 ( .A(n73483), .Y(n56650) );
  A2O1A1Ixp33_ASAP7_75t_SL U51247 ( .A1(n64401), .A2(n59283), .B(n56651), .C(
        n59012), .Y(n56652) );
  INVx1_ASAP7_75t_SL U51248 ( .A(n56654), .Y(n76455) );
  INVx1_ASAP7_75t_SL U51249 ( .A(n57069), .Y(n56655) );
  FAx1_ASAP7_75t_SL U51250 ( .A(n67113), .B(n67112), .CI(n67111), .CON(), .SN(
        n67213) );
  A2O1A1Ixp33_ASAP7_75t_SL U51251 ( .A1(n73965), .A2(n76336), .B(n77066), .C(
        n56660), .Y(n64234) );
  INVx1_ASAP7_75t_SL U51252 ( .A(iwb_err_i), .Y(n56661) );
  INVx1_ASAP7_75t_SL U51253 ( .A(n56668), .Y(n70873) );
  INVx1_ASAP7_75t_SL U51254 ( .A(or1200_cpu_or1200_mult_mac_n403), .Y(n56680)
         );
  INVx1_ASAP7_75t_SL U51255 ( .A(n69059), .Y(n56681) );
  INVx1_ASAP7_75t_SL U51256 ( .A(or1200_cpu_or1200_mult_mac_n193), .Y(n56682)
         );
  INVx1_ASAP7_75t_SL U51257 ( .A(n63774), .Y(n56683) );
  INVx1_ASAP7_75t_SL U51258 ( .A(or1200_cpu_or1200_mult_mac_n153), .Y(n56684)
         );
  INVx1_ASAP7_75t_SL U51259 ( .A(n63390), .Y(n56685) );
  INVx1_ASAP7_75t_SL U51260 ( .A(n75988), .Y(n56686) );
  INVx1_ASAP7_75t_SL U51261 ( .A(n76025), .Y(n56687) );
  INVx1_ASAP7_75t_SL U51262 ( .A(n68755), .Y(n56688) );
  INVx1_ASAP7_75t_SL U51263 ( .A(n74112), .Y(n56689) );
  XOR2xp5_ASAP7_75t_SL U51264 ( .A(n77174), .B(n77175), .Y(n78080) );
  XOR2xp5_ASAP7_75t_SL U51265 ( .A(n74574), .B(n74575), .Y(n78125) );
  INVx1_ASAP7_75t_SL U51266 ( .A(n77016), .Y(n56694) );
  INVx1_ASAP7_75t_SL U51267 ( .A(n69987), .Y(n56696) );
  INVx1_ASAP7_75t_SL U51268 ( .A(n65298), .Y(n56699) );
  O2A1O1Ixp33_ASAP7_75t_SL U51269 ( .A1(n65256), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .B(n56698), .C(
        n56699), .Y(n65302) );
  INVx1_ASAP7_75t_SL U51270 ( .A(n62024), .Y(n56700) );
  INVx1_ASAP7_75t_SL U51271 ( .A(n70186), .Y(n56708) );
  A2O1A1Ixp33_ASAP7_75t_SL U51272 ( .A1(n70766), .A2(n70785), .B(n70775), .C(
        n57211), .Y(n56715) );
  A2O1A1Ixp33_ASAP7_75t_SL U51273 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[0]), .A2(n53462), 
        .B(n71186), .C(n56716), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n103) );
  INVx1_ASAP7_75t_SL U51274 ( .A(n74274), .Y(n56717) );
  FAx1_ASAP7_75t_SL U51275 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_7_), .B(
        n74273), .CI(n56717), .CON(), .SN(n56718) );
  INVx1_ASAP7_75t_SL U51276 ( .A(n1600), .Y(n56723) );
  INVx1_ASAP7_75t_SL U51277 ( .A(n74568), .Y(n56725) );
  AOI21xp33_ASAP7_75t_SL U51278 ( .A1(n69198), .A2(n74572), .B(n76897), .Y(
        n56730) );
  O2A1O1Ixp33_ASAP7_75t_SL U51279 ( .A1(n69198), .A2(n74572), .B(n56730), .C(
        n56729), .Y(n56731) );
  INVx1_ASAP7_75t_SL U51280 ( .A(n65161), .Y(n56732) );
  INVx1_ASAP7_75t_SL U51281 ( .A(n65164), .Y(n56735) );
  AOI21xp33_ASAP7_75t_SL U51282 ( .A1(n65150), .A2(n56736), .B(n76897), .Y(
        n56737) );
  O2A1O1Ixp33_ASAP7_75t_SL U51283 ( .A1(n65150), .A2(n56736), .B(n56737), .C(
        n56734), .Y(n56738) );
  OAI21xp33_ASAP7_75t_SL U51284 ( .A1(n56733), .A2(n65149), .B(n59674), .Y(
        n56739) );
  A2O1A1Ixp33_ASAP7_75t_SL U51285 ( .A1(n65149), .A2(n56733), .B(n56739), .C(
        n56738), .Y(n56740) );
  INVx1_ASAP7_75t_SL U51286 ( .A(n56740), .Y(n56741) );
  INVx1_ASAP7_75t_SL U51287 ( .A(n76633), .Y(n56742) );
  INVx1_ASAP7_75t_SL U51288 ( .A(n57133), .Y(n56745) );
  NAND3xp33_ASAP7_75t_SL U51289 ( .A(n76160), .B(n76161), .C(n57104), .Y(
        n56746) );
  A2O1A1Ixp33_ASAP7_75t_SL U51290 ( .A1(n76161), .A2(n76160), .B(n57104), .C(
        n56746), .Y(n56747) );
  O2A1O1Ixp33_ASAP7_75t_SL U51291 ( .A1(n56745), .A2(n56747), .B(
        or1200_cpu_or1200_mult_mac_n16), .C(n57077), .Y(n56748) );
  OAI31xp33_ASAP7_75t_SL U51292 ( .A1(or1200_cpu_or1200_mult_mac_n16), .A2(
        n56745), .A3(n56747), .B(n56748), .Y(n56749) );
  INVx1_ASAP7_75t_SL U51293 ( .A(n58389), .Y(n56750) );
  INVx1_ASAP7_75t_SL U51294 ( .A(n68857), .Y(n56751) );
  INVx1_ASAP7_75t_SL U51295 ( .A(icqmem_adr_qmem[15]), .Y(n56754) );
  INVx1_ASAP7_75t_SL U51296 ( .A(icqmem_adr_qmem[21]), .Y(n56755) );
  INVx1_ASAP7_75t_SL U51297 ( .A(icqmem_adr_qmem[22]), .Y(n56756) );
  INVx1_ASAP7_75t_SL U51298 ( .A(icqmem_adr_qmem[23]), .Y(n56757) );
  INVx1_ASAP7_75t_SL U51299 ( .A(icqmem_adr_qmem[26]), .Y(n56758) );
  INVx1_ASAP7_75t_SL U51300 ( .A(icqmem_adr_qmem[27]), .Y(n56759) );
  INVx1_ASAP7_75t_SL U51301 ( .A(icqmem_adr_qmem[29]), .Y(n56760) );
  INVx1_ASAP7_75t_SL U51302 ( .A(icqmem_adr_qmem[31]), .Y(n56761) );
  INVx1_ASAP7_75t_SL U51303 ( .A(n53441), .Y(n56762) );
  A2O1A1Ixp33_ASAP7_75t_SL U51304 ( .A1(n77770), .A2(n59687), .B(n56765), .C(
        n57083), .Y(n56766) );
  INVx1_ASAP7_75t_SL U51305 ( .A(n76428), .Y(n56771) );
  INVx1_ASAP7_75t_SL U51306 ( .A(n77671), .Y(n56772) );
  INVx1_ASAP7_75t_SL U51307 ( .A(n1733), .Y(n56774) );
  INVx1_ASAP7_75t_SL U51308 ( .A(n69892), .Y(n56777) );
  INVx1_ASAP7_75t_SL U51309 ( .A(n70496), .Y(n56780) );
  OAI21xp33_ASAP7_75t_SL U51310 ( .A1(n56778), .A2(n69909), .B(n59621), .Y(
        n56782) );
  A2O1A1Ixp33_ASAP7_75t_SL U51311 ( .A1(n69909), .A2(n56778), .B(n56782), .C(
        n56781), .Y(n2283) );
  INVx1_ASAP7_75t_SL U51312 ( .A(n59621), .Y(n56787) );
  OAI21xp33_ASAP7_75t_SL U51313 ( .A1(n69718), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_0_), .B(n59621), .Y(
        n56789) );
  A2O1A1Ixp33_ASAP7_75t_SL U51314 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_0_), .A2(n69718), 
        .B(n56789), .C(n56788), .Y(n2313) );
  INVx1_ASAP7_75t_SL U51315 ( .A(n74341), .Y(n56790) );
  INVx1_ASAP7_75t_SL U51316 ( .A(n62146), .Y(n56792) );
  A2O1A1Ixp33_ASAP7_75t_SL U51317 ( .A1(n74967), .A2(n74968), .B(n74966), .C(
        n59694), .Y(n56800) );
  A2O1A1Ixp33_ASAP7_75t_SL U51318 ( .A1(n64003), .A2(n64004), .B(n64008), .C(
        n59694), .Y(n56801) );
  A2O1A1Ixp33_ASAP7_75t_SL U51319 ( .A1(n63982), .A2(n56802), .B(n53477), .C(
        n59694), .Y(n56803) );
  A2O1A1Ixp33_ASAP7_75t_SL U51320 ( .A1(n76814), .A2(n76815), .B(n76813), .C(
        n59694), .Y(n56804) );
  A2O1A1Ixp33_ASAP7_75t_SL U51321 ( .A1(n77267), .A2(n77268), .B(n77266), .C(
        n59694), .Y(n56805) );
  INVx1_ASAP7_75t_SL U51322 ( .A(n2491), .Y(n56809) );
  A2O1A1Ixp33_ASAP7_75t_SL U51323 ( .A1(n74752), .A2(n56817), .B(n56818), .C(
        n74751), .Y(n56819) );
  INVx1_ASAP7_75t_SL U51324 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[0]), .Y(
        n56822) );
  NAND3xp33_ASAP7_75t_SL U51325 ( .A(n56822), .B(n70570), .C(n74457), .Y(
        n56823) );
  A2O1A1Ixp33_ASAP7_75t_SL U51326 ( .A1(n70570), .A2(n74457), .B(n56822), .C(
        n56823), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_N586) );
  INVx1_ASAP7_75t_SL U51327 ( .A(n69824), .Y(n56825) );
  A2O1A1Ixp33_ASAP7_75t_SL U51328 ( .A1(n70077), .A2(n69825), .B(n56824), .C(
        n56825), .Y(n52524) );
  FAx1_ASAP7_75t_SL U51329 ( .A(n70142), .B(n70140), .CI(n53434), .CON(), .SN(
        n27047) );
  FAx1_ASAP7_75t_SL U51330 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_), 
        .B(n78243), .CI(n56826), .CON(), .SN(n12876) );
  FAx1_ASAP7_75t_SL U51331 ( .A(n72681), .B(n72679), .CI(n72680), .CON(), .SN(
        n27979) );
  AND2x4_ASAP7_75t_SL U51332 ( .A(n57663), .B(n58002), .Y(n57662) );
  OR2x6_ASAP7_75t_SL U51333 ( .A(n59592), .B(n63836), .Y(n56827) );
  BUFx6f_ASAP7_75t_SL U51334 ( .A(n76078), .Y(n57315) );
  AND2x6_ASAP7_75t_SL U51335 ( .A(n57665), .B(n56974), .Y(n58402) );
  AND2x4_ASAP7_75t_SL U51336 ( .A(n59537), .B(n59572), .Y(n56828) );
  INVx3_ASAP7_75t_SL U51337 ( .A(n59599), .Y(n57176) );
  INVx4_ASAP7_75t_SL U51338 ( .A(n57182), .Y(n59606) );
  BUFx6f_ASAP7_75t_SL U51339 ( .A(n68090), .Y(n59509) );
  NAND2x1p5_ASAP7_75t_SL U51340 ( .A(n76679), .B(n67424), .Y(n68090) );
  BUFx3_ASAP7_75t_SL U51341 ( .A(n1690), .Y(n57312) );
  INVx2_ASAP7_75t_SL U51342 ( .A(n64609), .Y(n67898) );
  NOR2x1p5_ASAP7_75t_SL U51343 ( .A(n63825), .B(n64034), .Y(n64609) );
  INVx6_ASAP7_75t_SL U51344 ( .A(n76172), .Y(n75947) );
  INVx6_ASAP7_75t_SL U51345 ( .A(n59644), .Y(n59641) );
  INVx8_ASAP7_75t_SL U51346 ( .A(n59615), .Y(n59614) );
  INVx5_ASAP7_75t_SL U51347 ( .A(n57537), .Y(n59615) );
  INVx2_ASAP7_75t_SL U51348 ( .A(n59535), .Y(n75378) );
  BUFx6f_ASAP7_75t_SL U51349 ( .A(n3130), .Y(n59582) );
  OAI21x1_ASAP7_75t_SL U51350 ( .A1(n77769), .A2(n77768), .B(n58399), .Y(
        n56829) );
  INVx3_ASAP7_75t_SL U51351 ( .A(n59050), .Y(n59649) );
  AO31x2_ASAP7_75t_SL U51352 ( .A1(n59613), .A2(n58761), .A3(n57025), .B(
        n58760), .Y(n56830) );
  AND4x1_ASAP7_75t_SL U51353 ( .A(n58215), .B(n59256), .C(n61908), .D(n58212), 
        .Y(n56831) );
  MAJx2_ASAP7_75t_SL U51354 ( .A(n67685), .B(n67686), .C(n67684), .Y(n56832)
         );
  XOR2xp5_ASAP7_75t_SL U51355 ( .A(n58332), .B(n57545), .Y(n56833) );
  OR2x2_ASAP7_75t_SL U51356 ( .A(n59599), .B(n76049), .Y(n56834) );
  INVx3_ASAP7_75t_SL U51357 ( .A(n64353), .Y(n59020) );
  AND2x2_ASAP7_75t_SL U51358 ( .A(n67463), .B(n58642), .Y(n56835) );
  OR2x2_ASAP7_75t_SL U51359 ( .A(n58499), .B(n58903), .Y(n56836) );
  OR2x2_ASAP7_75t_SL U51360 ( .A(n63177), .B(n57645), .Y(n56837) );
  BUFx3_ASAP7_75t_SL U51361 ( .A(n67897), .Y(n59455) );
  INVx3_ASAP7_75t_SL U51362 ( .A(n67897), .Y(n67738) );
  INVx2_ASAP7_75t_SL U51363 ( .A(n59242), .Y(n59165) );
  AO21x1_ASAP7_75t_SL U51364 ( .A1(n66258), .A2(n77242), .B(n59183), .Y(n56838) );
  NOR2x1_ASAP7_75t_SL U51365 ( .A(n75956), .B(n75955), .Y(n76191) );
  INVx6_ASAP7_75t_SL U51366 ( .A(n59099), .Y(n76049) );
  OR2x2_ASAP7_75t_SL U51367 ( .A(n59664), .B(n68413), .Y(n56839) );
  BUFx3_ASAP7_75t_SL U51368 ( .A(n59655), .Y(n57465) );
  AND2x2_ASAP7_75t_SL U51369 ( .A(n58204), .B(n62640), .Y(n56840) );
  AND2x2_ASAP7_75t_SL U51370 ( .A(n64651), .B(n57184), .Y(n56841) );
  HB1xp67_ASAP7_75t_SL U51371 ( .A(n59608), .Y(n57485) );
  BUFx6f_ASAP7_75t_SL U51372 ( .A(n57181), .Y(n57257) );
  MAJx2_ASAP7_75t_SL U51373 ( .A(n67470), .B(n67471), .C(n67472), .Y(n56842)
         );
  INVx2_ASAP7_75t_SL U51374 ( .A(n67639), .Y(n58711) );
  XOR2x2_ASAP7_75t_SL U51375 ( .A(n65008), .B(n57293), .Y(n56843) );
  AND2x2_ASAP7_75t_SL U51376 ( .A(n64038), .B(n64037), .Y(n56844) );
  INVx1_ASAP7_75t_SL U51377 ( .A(n56828), .Y(n57755) );
  OR2x2_ASAP7_75t_SL U51378 ( .A(n68102), .B(n63636), .Y(n56845) );
  OR2x2_ASAP7_75t_SL U51379 ( .A(n59446), .B(n57603), .Y(n56846) );
  OR2x2_ASAP7_75t_SL U51380 ( .A(n68720), .B(n68913), .Y(n56847) );
  INVx5_ASAP7_75t_SL U51381 ( .A(n58353), .Y(n57122) );
  INVx5_ASAP7_75t_SL U51382 ( .A(n58353), .Y(n59654) );
  INVx8_ASAP7_75t_SL U51383 ( .A(n58439), .Y(n59618) );
  OR2x6_ASAP7_75t_SL U51384 ( .A(n76679), .B(n62649), .Y(n58439) );
  OR2x2_ASAP7_75t_SL U51385 ( .A(n67517), .B(n57076), .Y(n56848) );
  BUFx3_ASAP7_75t_SL U51386 ( .A(n2547), .Y(n59438) );
  OR2x2_ASAP7_75t_SL U51387 ( .A(n67568), .B(n57165), .Y(n56849) );
  INVx6_ASAP7_75t_SL U51388 ( .A(n57628), .Y(n59456) );
  OR2x2_ASAP7_75t_SL U51389 ( .A(n75032), .B(n59139), .Y(n56850) );
  AND2x2_ASAP7_75t_SL U51390 ( .A(n53207), .B(n63068), .Y(n56851) );
  INVx2_ASAP7_75t_SL U51391 ( .A(n67965), .Y(n57113) );
  NOR2x1_ASAP7_75t_SL U51392 ( .A(n68102), .B(n67534), .Y(n67494) );
  INVx5_ASAP7_75t_SL U51393 ( .A(n59605), .Y(n59602) );
  INVx2_ASAP7_75t_SL U51394 ( .A(n67457), .Y(n67232) );
  INVx11_ASAP7_75t_SL U51395 ( .A(n59707), .Y(n59709) );
  INVx1_ASAP7_75t_SL U51396 ( .A(n59708), .Y(n59398) );
  INVx6_ASAP7_75t_SL U51397 ( .A(n57181), .Y(n59609) );
  AND2x2_ASAP7_75t_SL U51398 ( .A(n57913), .B(n59260), .Y(n56852) );
  INVx4_ASAP7_75t_SL U51399 ( .A(n59454), .Y(n67306) );
  INVx1_ASAP7_75t_SL U51400 ( .A(n64701), .Y(n64705) );
  XNOR2x1_ASAP7_75t_SL U51401 ( .A(n64435), .B(n64434), .Y(n64701) );
  INVx4_ASAP7_75t_SL U51402 ( .A(n57107), .Y(n59653) );
  AND3x1_ASAP7_75t_SL U51403 ( .A(n67701), .B(n62725), .C(n62767), .Y(n56853)
         );
  INVx1_ASAP7_75t_SL U51404 ( .A(n67898), .Y(n58155) );
  AO21x1_ASAP7_75t_SL U51405 ( .A1(n59655), .A2(n63063), .B(n57213), .Y(n56854) );
  INVx2_ASAP7_75t_SL U51406 ( .A(n61931), .Y(n61912) );
  AND2x2_ASAP7_75t_SL U51407 ( .A(n67410), .B(n59604), .Y(n56855) );
  NAND2xp5_ASAP7_75t_SL U51408 ( .A(n69015), .B(n69014), .Y(n56856) );
  AND2x2_ASAP7_75t_SL U51409 ( .A(n59662), .B(n57720), .Y(n56857) );
  BUFx6f_ASAP7_75t_SL U51410 ( .A(n1796), .Y(n59541) );
  INVx4_ASAP7_75t_SL U51411 ( .A(n59541), .Y(n58206) );
  INVx3_ASAP7_75t_SL U51412 ( .A(n70528), .Y(n70103) );
  INVx2_ASAP7_75t_SL U51413 ( .A(n67906), .Y(n67251) );
  HB1xp67_ASAP7_75t_SL U51414 ( .A(n75287), .Y(n57474) );
  AOI21x1_ASAP7_75t_SL U51415 ( .A1(n63711), .A2(n74931), .B(n63713), .Y(
        n76926) );
  BUFx3_ASAP7_75t_SL U51416 ( .A(n75035), .Y(n57436) );
  BUFx3_ASAP7_75t_SL U51417 ( .A(n58353), .Y(n57347) );
  AND2x4_ASAP7_75t_SL U51418 ( .A(n59197), .B(n64516), .Y(n67227) );
  INVx3_ASAP7_75t_SL U51419 ( .A(n67227), .Y(n67638) );
  AND2x6_ASAP7_75t_SL U51420 ( .A(n74502), .B(n73853), .Y(n73382) );
  INVx8_ASAP7_75t_SL U51421 ( .A(n73382), .Y(n59631) );
  INVx8_ASAP7_75t_SL U51422 ( .A(n73382), .Y(n59630) );
  OR2x4_ASAP7_75t_SL U51423 ( .A(n63714), .B(n63713), .Y(n63715) );
  INVx1_ASAP7_75t_SL U51424 ( .A(n63571), .Y(n59583) );
  OR2x4_ASAP7_75t_SL U51425 ( .A(n59711), .B(n59442), .Y(n63571) );
  BUFx3_ASAP7_75t_SL U51426 ( .A(n57184), .Y(n57491) );
  INVx1_ASAP7_75t_SL U51427 ( .A(n59536), .Y(n77711) );
  BUFx6f_ASAP7_75t_SL U51428 ( .A(n1672), .Y(n59536) );
  INVx6_ASAP7_75t_SL U51429 ( .A(n77298), .Y(n59681) );
  NAND2x1p5_ASAP7_75t_SL U51430 ( .A(n56838), .B(n59361), .Y(n62649) );
  INVx2_ASAP7_75t_SL U51431 ( .A(n58424), .Y(n57881) );
  AND2x2_ASAP7_75t_SL U51432 ( .A(n68732), .B(n68731), .Y(n56858) );
  BUFx3_ASAP7_75t_SL U51433 ( .A(n59502), .Y(n57284) );
  AND2x2_ASAP7_75t_SL U51434 ( .A(n69007), .B(n69011), .Y(n56859) );
  INVx4_ASAP7_75t_SL U51435 ( .A(n59563), .Y(n75628) );
  BUFx6f_ASAP7_75t_SL U51436 ( .A(n2011), .Y(n59563) );
  INVx4_ASAP7_75t_SL U51437 ( .A(n59572), .Y(n57210) );
  INVx3_ASAP7_75t_SL U51438 ( .A(n59554), .Y(n56954) );
  INVx3_ASAP7_75t_SL U51439 ( .A(n59559), .Y(n59182) );
  AND2x2_ASAP7_75t_SL U51440 ( .A(n74556), .B(n74555), .Y(n56860) );
  INVx2_ASAP7_75t_SL U51441 ( .A(n77362), .Y(n59685) );
  INVx2_ASAP7_75t_SL U51442 ( .A(n77362), .Y(n57071) );
  INVx1_ASAP7_75t_SL U51443 ( .A(n77362), .Y(n59684) );
  INVx2_ASAP7_75t_SL U51444 ( .A(n59576), .Y(n75740) );
  BUFx6f_ASAP7_75t_SL U51445 ( .A(n2902), .Y(n59576) );
  INVx8_ASAP7_75t_SL U51446 ( .A(n73047), .Y(n59629) );
  NAND2xp5_ASAP7_75t_SL U51447 ( .A(n59535), .B(n59533), .Y(n74005) );
  INVx1_ASAP7_75t_SL U51448 ( .A(n59053), .Y(n57753) );
  BUFx6f_ASAP7_75t_SL U51449 ( .A(n3351), .Y(n59702) );
  INVx11_ASAP7_75t_SL U51450 ( .A(n59702), .Y(n59703) );
  INVx8_ASAP7_75t_SL U51451 ( .A(n75872), .Y(n57126) );
  OR2x6_ASAP7_75t_SL U51452 ( .A(n60686), .B(n60685), .Y(n75872) );
  NOR2x1_ASAP7_75t_SL U51453 ( .A(n58595), .B(n74165), .Y(n76956) );
  INVx2_ASAP7_75t_SL U51454 ( .A(n3309), .Y(n59705) );
  INVx5_ASAP7_75t_SL U51455 ( .A(n70502), .Y(n57081) );
  OR2x6_ASAP7_75t_SL U51456 ( .A(n2455), .B(n70477), .Y(n70502) );
  INVx1_ASAP7_75t_SL U51457 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_state), .Y(n59699) );
  NAND2x1p5_ASAP7_75t_SL U51458 ( .A(n60658), .B(n59166), .Y(n66253) );
  XNOR2x1_ASAP7_75t_SL U51459 ( .A(n67198), .B(n67199), .Y(n67066) );
  AOI22x1_ASAP7_75t_SL U51460 ( .A1(n57478), .A2(n67721), .B1(n59171), .B2(
        n67720), .Y(n68384) );
  INVx5_ASAP7_75t_SL U51461 ( .A(n58384), .Y(n57912) );
  AOI21x1_ASAP7_75t_SL U51462 ( .A1(n68248), .A2(n68247), .B(n68246), .Y(
        n58638) );
  INVxp33_ASAP7_75t_SRAM U51463 ( .A(n57556), .Y(n58940) );
  BUFx3_ASAP7_75t_SL U51464 ( .A(n2016), .Y(n56861) );
  XNOR2x1_ASAP7_75t_SL U51465 ( .A(n68469), .B(n59151), .Y(n68435) );
  HB1xp67_ASAP7_75t_SL U51466 ( .A(n68956), .Y(n57477) );
  OAI21x1_ASAP7_75t_SL U51467 ( .A1(n57352), .A2(n62687), .B(n62686), .Y(
        n67701) );
  XNOR2x1_ASAP7_75t_SL U51468 ( .A(n64979), .B(n64978), .Y(n64980) );
  INVx1_ASAP7_75t_SL U51469 ( .A(n68160), .Y(n57892) );
  AOI22xp5_ASAP7_75t_SL U51470 ( .A1(n64937), .A2(n67306), .B1(n67970), .B2(
        n57161), .Y(n58690) );
  HB1xp67_ASAP7_75t_SL U51471 ( .A(n53290), .Y(n57333) );
  XOR2x2_ASAP7_75t_SL U51472 ( .A(n67667), .B(n67665), .Y(n67573) );
  HB1xp67_ASAP7_75t_SL U51473 ( .A(n68249), .Y(n57423) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51474 ( .A1(n67736), .A2(n59456), .B(n67735), 
        .C(n59012), .Y(n67737) );
  NOR2x1p5_ASAP7_75t_SL U51475 ( .A(n59456), .B(n57656), .Y(n67441) );
  XNOR2x2_ASAP7_75t_SL U51476 ( .A(n59076), .B(n67754), .Y(n68368) );
  HB1xp67_ASAP7_75t_SL U51477 ( .A(n66260), .Y(n57504) );
  BUFx3_ASAP7_75t_SL U51478 ( .A(n59613), .Y(n57463) );
  BUFx3_ASAP7_75t_SL U51479 ( .A(n66398), .Y(n57302) );
  INVx2_ASAP7_75t_SL U51480 ( .A(n64034), .Y(n63827) );
  BUFx2_ASAP7_75t_SL U51481 ( .A(n68131), .Y(n57438) );
  NAND2xp5_ASAP7_75t_SL U51482 ( .A(n68073), .B(n68074), .Y(n68048) );
  NAND2x1p5_ASAP7_75t_SL U51483 ( .A(n56834), .B(n59055), .Y(n67589) );
  HB1xp67_ASAP7_75t_SL U51484 ( .A(n68860), .Y(n58389) );
  INVxp33_ASAP7_75t_SRAM U51485 ( .A(n68860), .Y(n58087) );
  BUFx3_ASAP7_75t_SL U51486 ( .A(n67339), .Y(n56862) );
  NAND2xp5_ASAP7_75t_SL U51487 ( .A(n75643), .B(n59487), .Y(n67339) );
  NOR2x1_ASAP7_75t_SL U51488 ( .A(n62669), .B(n60777), .Y(n60744) );
  NOR2x1_ASAP7_75t_SL U51489 ( .A(n59580), .B(n62667), .Y(n62669) );
  INVxp33_ASAP7_75t_SRAM U51490 ( .A(n67980), .Y(n58072) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51491 ( .A1(n59182), .A2(n60655), .B(n59545), 
        .C(n76627), .Y(n60684) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U51492 ( .A1(n59545), .A2(n62590), .B(n60930), 
        .C(n77242), .Y(n60931) );
  BUFx2_ASAP7_75t_SL U51493 ( .A(n56861), .Y(n59564) );
  INVx4_ASAP7_75t_SL U51494 ( .A(n59564), .Y(n59183) );
  INVxp33_ASAP7_75t_SRAM U51495 ( .A(n68173), .Y(n68169) );
  HB1xp67_ASAP7_75t_SL U51496 ( .A(n59297), .Y(n57241) );
  XNOR2xp5_ASAP7_75t_SL U51497 ( .A(n58484), .B(n57745), .Y(n58726) );
  XNOR2x1_ASAP7_75t_SL U51498 ( .A(n58080), .B(n57315), .Y(n66696) );
  OAI22x1_ASAP7_75t_SL U51499 ( .A1(n67512), .A2(n58903), .B1(n68383), .B2(
        n67693), .Y(n67682) );
  NAND2x1p5_ASAP7_75t_SL U51500 ( .A(n59482), .B(n58071), .Y(n59474) );
  NAND2x1p5_ASAP7_75t_SL U51501 ( .A(n58234), .B(n58235), .Y(n62611) );
  INVx5_ASAP7_75t_SL U51502 ( .A(n59669), .Y(n59668) );
  AOI22xp33_ASAP7_75t_SRAM U51503 ( .A1(n59634), .A2(n66572), .B1(n68594), 
        .B2(n57067), .Y(n68595) );
  XNOR2x2_ASAP7_75t_SL U51504 ( .A(n68135), .B(n68134), .Y(n68210) );
  XOR2xp5_ASAP7_75t_SL U51505 ( .A(n68132), .B(n68133), .Y(n68134) );
  INVx1_ASAP7_75t_SL U51506 ( .A(n58143), .Y(n59517) );
  AND2x2_ASAP7_75t_SL U51507 ( .A(n58143), .B(n58789), .Y(n58845) );
  XNOR2x1_ASAP7_75t_SL U51508 ( .A(n64977), .B(n64976), .Y(n64999) );
  XNOR2x1_ASAP7_75t_SL U51509 ( .A(n64975), .B(n65001), .Y(n64976) );
  NOR2x1p5_ASAP7_75t_SL U51510 ( .A(n57589), .B(n57588), .Y(n63179) );
  NAND3x1_ASAP7_75t_SL U51511 ( .A(n59555), .B(n59569), .C(n1796), .Y(n57588)
         );
  INVxp33_ASAP7_75t_SRAM U51512 ( .A(n75107), .Y(n57982) );
  INVx1_ASAP7_75t_SL U51513 ( .A(n56863), .Y(n56864) );
  NAND2xp5_ASAP7_75t_SL U51514 ( .A(n77709), .B(n64081), .Y(n63675) );
  NOR2x1p5_ASAP7_75t_SL U51515 ( .A(n68573), .B(n68572), .Y(n58088) );
  NAND2xp5_ASAP7_75t_SL U51516 ( .A(n59595), .B(n67276), .Y(n64605) );
  XNOR2x2_ASAP7_75t_SL U51517 ( .A(n58495), .B(n68318), .Y(n59330) );
  BUFx2_ASAP7_75t_SL U51518 ( .A(n67421), .Y(n57486) );
  NAND2x1p5_ASAP7_75t_SL U51519 ( .A(n67421), .B(n57698), .Y(n68097) );
  INVxp33_ASAP7_75t_SRAM U51520 ( .A(n68906), .Y(n58259) );
  INVxp33_ASAP7_75t_SRAM U51521 ( .A(n68229), .Y(n68238) );
  XNOR2x1_ASAP7_75t_SL U51522 ( .A(n68404), .B(n57541), .Y(n68397) );
  HB1xp67_ASAP7_75t_SL U51523 ( .A(n68051), .Y(n57482) );
  HB1xp67_ASAP7_75t_SL U51524 ( .A(or1200_cpu_or1200_except_ex_freeze_prev), 
        .Y(n57343) );
  TIELOx1_ASAP7_75t_SL U51525 ( .L(pm_lvolt_o) );
  TIEHIx1_ASAP7_75t_SL U51526 ( .H(pm_wakeup_o) );
  TIELOx1_ASAP7_75t_SL U51527 ( .L(pm_cpu_gate_o) );
  TIELOx1_ASAP7_75t_SL U51528 ( .L(pm_tt_gate_o) );
  TIELOx1_ASAP7_75t_SL U51529 ( .L(pm_immu_gate_o) );
  TIELOx1_ASAP7_75t_SL U51530 ( .L(pm_dmmu_gate_o) );
  TIELOx1_ASAP7_75t_SL U51531 ( .L(pm_ic_gate_o) );
  TIELOx1_ASAP7_75t_SL U51532 ( .L(pm_dc_gate_o) );
  TIELOx1_ASAP7_75t_SL U51533 ( .L(pm_clksd_o[0]) );
  TIELOx1_ASAP7_75t_SL U51534 ( .L(pm_clksd_o[1]) );
  TIELOx1_ASAP7_75t_SL U51535 ( .L(pm_clksd_o[2]) );
  TIELOx1_ASAP7_75t_SL U51536 ( .L(pm_clksd_o[3]) );
  TIELOx1_ASAP7_75t_SL U51537 ( .L(dbg_wp_o[0]) );
  TIELOx1_ASAP7_75t_SL U51538 ( .L(dbg_wp_o[1]) );
  TIELOx1_ASAP7_75t_SL U51539 ( .L(dbg_wp_o[2]) );
  TIELOx1_ASAP7_75t_SL U51540 ( .L(dbg_wp_o[3]) );
  TIELOx1_ASAP7_75t_SL U51541 ( .L(dbg_wp_o[4]) );
  TIELOx1_ASAP7_75t_SL U51542 ( .L(dbg_wp_o[5]) );
  TIELOx1_ASAP7_75t_SL U51543 ( .L(dbg_wp_o[6]) );
  TIELOx1_ASAP7_75t_SL U51544 ( .L(dbg_wp_o[7]) );
  TIELOx1_ASAP7_75t_SL U51545 ( .L(dbg_wp_o[8]) );
  TIELOx1_ASAP7_75t_SL U51546 ( .L(dbg_wp_o[9]) );
  TIELOx1_ASAP7_75t_SL U51547 ( .L(dbg_wp_o[10]) );
  TIELOx1_ASAP7_75t_SL U51548 ( .L(dbg_lss_o[0]) );
  TIELOx1_ASAP7_75t_SL U51549 ( .L(dbg_lss_o[1]) );
  TIELOx1_ASAP7_75t_SL U51550 ( .L(dbg_lss_o[2]) );
  TIELOx1_ASAP7_75t_SL U51551 ( .L(dbg_lss_o[3]) );
  TIEHIx1_ASAP7_75t_SL U51552 ( .H(dwb_bte_o[0]) );
  TIELOx1_ASAP7_75t_SL U51553 ( .L(dwb_bte_o[1]) );
  TIEHIx1_ASAP7_75t_SL U51554 ( .H(dwb_cti_o[0]) );
  TIEHIx1_ASAP7_75t_SL U51555 ( .H(dwb_cti_o[1]) );
  TIEHIx1_ASAP7_75t_SL U51556 ( .H(dwb_cti_o[2]) );
  TIEHIx1_ASAP7_75t_SL U51557 ( .H(iwb_bte_o[0]) );
  TIELOx1_ASAP7_75t_SL U51558 ( .L(iwb_bte_o[1]) );
  TIEHIx1_ASAP7_75t_SL U51559 ( .H(iwb_cti_o[0]) );
  TIEHIx1_ASAP7_75t_SL U51560 ( .H(iwb_cti_o[1]) );
  TIEHIx1_ASAP7_75t_SL U51561 ( .H(iwb_cti_o[2]) );
  TIELOx1_ASAP7_75t_SL U51562 ( .L(iwb_dat_o[0]) );
  TIELOx1_ASAP7_75t_SL U51563 ( .L(iwb_dat_o[1]) );
  TIELOx1_ASAP7_75t_SL U51564 ( .L(iwb_dat_o[2]) );
  TIELOx1_ASAP7_75t_SL U51565 ( .L(iwb_dat_o[3]) );
  TIELOx1_ASAP7_75t_SL U51566 ( .L(iwb_dat_o[4]) );
  TIELOx1_ASAP7_75t_SL U51567 ( .L(iwb_dat_o[5]) );
  TIELOx1_ASAP7_75t_SL U51568 ( .L(iwb_dat_o[6]) );
  TIELOx1_ASAP7_75t_SL U51569 ( .L(iwb_dat_o[7]) );
  TIELOx1_ASAP7_75t_SL U51570 ( .L(iwb_dat_o[8]) );
  TIELOx1_ASAP7_75t_SL U51571 ( .L(iwb_dat_o[9]) );
  TIELOx1_ASAP7_75t_SL U51572 ( .L(iwb_dat_o[10]) );
  TIELOx1_ASAP7_75t_SL U51573 ( .L(iwb_dat_o[11]) );
  TIELOx1_ASAP7_75t_SL U51574 ( .L(iwb_dat_o[12]) );
  TIELOx1_ASAP7_75t_SL U51575 ( .L(iwb_dat_o[13]) );
  TIELOx1_ASAP7_75t_SL U51576 ( .L(iwb_dat_o[14]) );
  TIELOx1_ASAP7_75t_SL U51577 ( .L(iwb_dat_o[15]) );
  TIELOx1_ASAP7_75t_SL U51578 ( .L(iwb_dat_o[16]) );
  TIELOx1_ASAP7_75t_SL U51579 ( .L(iwb_dat_o[17]) );
  TIELOx1_ASAP7_75t_SL U51580 ( .L(iwb_dat_o[18]) );
  TIELOx1_ASAP7_75t_SL U51581 ( .L(iwb_dat_o[19]) );
  TIELOx1_ASAP7_75t_SL U51582 ( .L(iwb_dat_o[20]) );
  TIELOx1_ASAP7_75t_SL U51583 ( .L(iwb_dat_o[21]) );
  TIELOx1_ASAP7_75t_SL U51584 ( .L(iwb_dat_o[22]) );
  TIELOx1_ASAP7_75t_SL U51585 ( .L(iwb_dat_o[23]) );
  TIELOx1_ASAP7_75t_SL U51586 ( .L(iwb_dat_o[24]) );
  TIELOx1_ASAP7_75t_SL U51587 ( .L(iwb_dat_o[25]) );
  TIELOx1_ASAP7_75t_SL U51588 ( .L(iwb_dat_o[26]) );
  TIELOx1_ASAP7_75t_SL U51589 ( .L(iwb_dat_o[27]) );
  TIELOx1_ASAP7_75t_SL U51590 ( .L(iwb_dat_o[28]) );
  TIELOx1_ASAP7_75t_SL U51591 ( .L(iwb_dat_o[29]) );
  TIELOx1_ASAP7_75t_SL U51592 ( .L(iwb_dat_o[30]) );
  TIELOx1_ASAP7_75t_SL U51593 ( .L(iwb_dat_o[31]) );
  TIEHIx1_ASAP7_75t_SL U51594 ( .H(iwb_sel_o[0]) );
  TIEHIx1_ASAP7_75t_SL U51595 ( .H(iwb_sel_o[1]) );
  TIEHIx1_ASAP7_75t_SL U51596 ( .H(iwb_sel_o[2]) );
  TIEHIx1_ASAP7_75t_SL U51597 ( .H(iwb_sel_o[3]) );
  TIELOx1_ASAP7_75t_SL U51598 ( .L(iwb_we_o) );
  TIELOx1_ASAP7_75t_SL U51599 ( .L(iwb_adr_o[0]) );
  TIELOx1_ASAP7_75t_SL U51600 ( .L(iwb_adr_o[1]) );
  O2A1O1Ixp33_ASAP7_75t_SL U51601 ( .A1(n56943), .A2(n69003), .B(n56859), .C(
        n69013), .Y(n56942) );
  INVxp67_ASAP7_75t_SL U51602 ( .A(n69015), .Y(n56943) );
  INVxp67_ASAP7_75t_SL U51603 ( .A(n56945), .Y(n56944) );
  NOR3xp33_ASAP7_75t_SL U51604 ( .A(n58262), .B(n69003), .C(n56856), .Y(n56945) );
  INVx1_ASAP7_75t_SL U51605 ( .A(n56946), .Y(n57940) );
  NAND3xp33_ASAP7_75t_SL U51606 ( .A(n56946), .B(n76176), .C(n67326), .Y(
        n58641) );
  NOR2x1p5_ASAP7_75t_SL U51607 ( .A(n57941), .B(n57162), .Y(n56946) );
  NAND2xp5_ASAP7_75t_SL U51608 ( .A(n58482), .B(n56946), .Y(n59134) );
  XOR2xp5_ASAP7_75t_SL U51609 ( .A(n67190), .B(n67191), .Y(n56950) );
  OAI21xp5_ASAP7_75t_SL U51610 ( .A1(n56951), .A2(n56950), .B(n56948), .Y(
        n67204) );
  NAND2xp5_ASAP7_75t_SL U51611 ( .A(n56949), .B(n56950), .Y(n56948) );
  INVx1_ASAP7_75t_SL U51612 ( .A(n58635), .Y(n56949) );
  MAJx2_ASAP7_75t_SL U51613 ( .A(n67204), .B(n67203), .C(n67202), .Y(n56947)
         );
  NOR2x1_ASAP7_75t_SL U51614 ( .A(n67193), .B(n67192), .Y(n56951) );
  INVx1_ASAP7_75t_SL U51615 ( .A(n67197), .Y(n56952) );
  MAJIxp5_ASAP7_75t_SL U51616 ( .A(n67049), .B(n67047), .C(n67048), .Y(n67197)
         );
  AOI21xp5_ASAP7_75t_SL U51617 ( .A1(n66683), .A2(n58336), .B(n59174), .Y(
        n66771) );
  A2O1A1Ixp33_ASAP7_75t_SL U51618 ( .A1(n75466), .A2(n59641), .B(n75068), .C(
        n53205), .Y(n75066) );
  AOI22xp5_ASAP7_75t_SL U51619 ( .A1(n57163), .A2(n75077), .B1(n53205), .B2(
        n68604), .Y(n66566) );
  XOR2xp5_ASAP7_75t_SL U51620 ( .A(n56953), .B(n67884), .Y(n56966) );
  NOR2x1p5_ASAP7_75t_SL U51621 ( .A(n57849), .B(n57848), .Y(n56953) );
  NAND2xp5_ASAP7_75t_SL U51622 ( .A(n59580), .B(n59256), .Y(n58532) );
  NAND2xp5_ASAP7_75t_SL U51623 ( .A(n1802), .B(n59543), .Y(n56955) );
  NAND2xp5_ASAP7_75t_SL U51624 ( .A(n67387), .B(n58397), .Y(n56959) );
  NAND2xp5_ASAP7_75t_SL U51625 ( .A(n67389), .B(n56956), .Y(n67708) );
  INVx1_ASAP7_75t_SL U51626 ( .A(n56958), .Y(n56956) );
  NAND2xp5_ASAP7_75t_SL U51627 ( .A(n67306), .B(n67389), .Y(n56957) );
  NOR2x1_ASAP7_75t_SL U51628 ( .A(n67569), .B(n59600), .Y(n56958) );
  OAI211xp5_ASAP7_75t_SL U51629 ( .A1(n53621), .A2(n69047), .B(n56960), .C(
        n69046), .Y(n52009) );
  NAND2xp5_ASAP7_75t_SL U51630 ( .A(n58527), .B(n53621), .Y(n56960) );
  NAND2xp5_ASAP7_75t_SL U51631 ( .A(n68852), .B(n68859), .Y(n68839) );
  AO21x1_ASAP7_75t_SL U51632 ( .A1(n68721), .A2(n68834), .B(n56961), .Y(n68859) );
  OAI21xp5_ASAP7_75t_SL U51633 ( .A1(n68920), .A2(n68974), .B(n58637), .Y(
        n56961) );
  NOR2x1_ASAP7_75t_SL U51634 ( .A(n57481), .B(n68900), .Y(n68974) );
  NAND2xp5_ASAP7_75t_SL U51635 ( .A(n56963), .B(n56962), .Y(n67163) );
  NAND2xp5_ASAP7_75t_SL U51636 ( .A(n67157), .B(n58682), .Y(n56962) );
  OAI21xp5_ASAP7_75t_SL U51637 ( .A1(n67174), .A2(n67157), .B(n56964), .Y(
        n56963) );
  INVx1_ASAP7_75t_SL U51638 ( .A(n67175), .Y(n56964) );
  XNOR2xp5_ASAP7_75t_SL U51639 ( .A(n67142), .B(n56965), .Y(n67157) );
  XNOR2xp5_ASAP7_75t_SL U51640 ( .A(n67141), .B(n67140), .Y(n56965) );
  MAJIxp5_ASAP7_75t_SL U51641 ( .A(n57664), .B(n67144), .C(n67145), .Y(n67175)
         );
  INVx2_ASAP7_75t_SL U51642 ( .A(n59545), .Y(n57575) );
  XNOR2xp5_ASAP7_75t_SL U51643 ( .A(n57458), .B(n56966), .Y(n68116) );
  NOR2x2_ASAP7_75t_SL U51644 ( .A(n63169), .B(n58872), .Y(n59453) );
  NOR2x2_ASAP7_75t_SL U51645 ( .A(n67017), .B(n59057), .Y(n58872) );
  XOR2xp5_ASAP7_75t_SL U51646 ( .A(n58089), .B(n58355), .Y(n67205) );
  NOR2x1p5_ASAP7_75t_SL U51647 ( .A(n67861), .B(n66625), .Y(n67593) );
  XNOR2x1_ASAP7_75t_SL U51648 ( .A(n53485), .B(n58921), .Y(n67578) );
  XNOR2x1_ASAP7_75t_SL U51649 ( .A(n67351), .B(n58922), .Y(n67579) );
  BUFx6f_ASAP7_75t_SL U51650 ( .A(n2519), .Y(n59464) );
  NOR2x1_ASAP7_75t_SL U51651 ( .A(n59530), .B(n64894), .Y(n57808) );
  NOR2x1_ASAP7_75t_SL U51652 ( .A(n62761), .B(n64894), .Y(n59394) );
  XNOR2xp5_ASAP7_75t_SL U51653 ( .A(n57529), .B(n68533), .Y(n68521) );
  NAND2xp5_ASAP7_75t_SL U51654 ( .A(n66258), .B(n57439), .Y(n64364) );
  NOR2xp33_ASAP7_75t_SL U51655 ( .A(n57209), .B(n64357), .Y(n57439) );
  OAI21xp5_ASAP7_75t_SL U51656 ( .A1(n68242), .A2(n68241), .B(n68240), .Y(
        n68251) );
  HB1xp67_ASAP7_75t_SL U51657 ( .A(n62572), .Y(n56968) );
  INVx3_ASAP7_75t_SL U51658 ( .A(n59253), .Y(n58746) );
  NAND2xp5_ASAP7_75t_SL U51659 ( .A(n64752), .B(n68560), .Y(n64870) );
  XNOR2xp5_ASAP7_75t_SL U51660 ( .A(n64675), .B(n57877), .Y(n63629) );
  XOR2xp5_ASAP7_75t_SL U51661 ( .A(n56969), .B(n57602), .Y(n52005) );
  AND2x2_ASAP7_75t_SL U51662 ( .A(n69094), .B(n69102), .Y(n56969) );
  NOR2xp33_ASAP7_75t_SL U51663 ( .A(n57537), .B(n64966), .Y(n67300) );
  XNOR2x1_ASAP7_75t_SL U51664 ( .A(n68448), .B(n57338), .Y(n57620) );
  OAI21xp5_ASAP7_75t_SL U51665 ( .A1(n66800), .A2(n57112), .B(n64624), .Y(
        n64952) );
  XNOR2x2_ASAP7_75t_SL U51666 ( .A(n57112), .B(n68104), .Y(n64954) );
  AOI211xp5_ASAP7_75t_SL U51667 ( .A1(n59662), .A2(n57112), .B(n67451), .C(
        n67316), .Y(n67317) );
  NAND2xp5_ASAP7_75t_SL U51668 ( .A(n58753), .B(n57112), .Y(n64624) );
  NOR2x1_ASAP7_75t_SL U51669 ( .A(n57112), .B(n75962), .Y(n67595) );
  NAND2x1p5_ASAP7_75t_SL U51670 ( .A(n57112), .B(n59435), .Y(n67864) );
  INVx6_ASAP7_75t_SL U51671 ( .A(n57112), .Y(n68098) );
  INVx6_ASAP7_75t_SL U51672 ( .A(n58173), .Y(n57112) );
  NAND2x1_ASAP7_75t_SL U51673 ( .A(n64734), .B(n64733), .Y(n74993) );
  INVx4_ASAP7_75t_SL U51674 ( .A(n67972), .Y(n67911) );
  NAND2x1_ASAP7_75t_SL U51675 ( .A(n59532), .B(n63807), .Y(n63808) );
  XNOR2x1_ASAP7_75t_SL U51676 ( .A(n56970), .B(n57460), .Y(n68036) );
  XNOR2x1_ASAP7_75t_SL U51677 ( .A(n58455), .B(n67772), .Y(n56970) );
  XOR2xp5_ASAP7_75t_SL U51678 ( .A(n68062), .B(n68061), .Y(n68063) );
  OR2x2_ASAP7_75t_SL U51679 ( .A(n59549), .B(n57186), .Y(n56971) );
  INVx8_ASAP7_75t_SL U51680 ( .A(n59661), .Y(n59662) );
  OR2x2_ASAP7_75t_SL U51681 ( .A(n59644), .B(n59514), .Y(n56972) );
  NAND2x1_ASAP7_75t_SL U51682 ( .A(n62721), .B(n58905), .Y(n59467) );
  INVx3_ASAP7_75t_SL U51683 ( .A(n59511), .Y(n58701) );
  OR2x2_ASAP7_75t_SL U51684 ( .A(n59512), .B(n59641), .Y(n56973) );
  INVx8_ASAP7_75t_SL U51685 ( .A(n58639), .Y(n59597) );
  INVx2_ASAP7_75t_SL U51686 ( .A(n58402), .Y(n57696) );
  INVx2_ASAP7_75t_SL U51687 ( .A(n59617), .Y(n57827) );
  INVx6_ASAP7_75t_SL U51688 ( .A(n59617), .Y(n59616) );
  OR2x2_ASAP7_75t_SL U51689 ( .A(n59394), .B(n57666), .Y(n56974) );
  INVx5_ASAP7_75t_SL U51690 ( .A(n76028), .Y(n57169) );
  HB1xp67_ASAP7_75t_SL U51691 ( .A(n67636), .Y(n57221) );
  INVx3_ASAP7_75t_SL U51692 ( .A(n59639), .Y(n59638) );
  NOR2x1_ASAP7_75t_SL U51693 ( .A(n59710), .B(n59591), .Y(n75916) );
  BUFx6f_ASAP7_75t_SL U51694 ( .A(n75916), .Y(n59656) );
  INVx4_ASAP7_75t_SL U51695 ( .A(n59663), .Y(n59665) );
  OR2x2_ASAP7_75t_SL U51696 ( .A(n75930), .B(n67826), .Y(n56975) );
  OR2x2_ASAP7_75t_SL U51697 ( .A(n67481), .B(n57113), .Y(n56976) );
  AND2x2_ASAP7_75t_SL U51698 ( .A(n59641), .B(n67360), .Y(n56977) );
  OR2x2_ASAP7_75t_SL U51699 ( .A(n59239), .B(n66806), .Y(n56978) );
  AO21x1_ASAP7_75t_SL U51700 ( .A1(n62645), .A2(n62646), .B(n58220), .Y(n56979) );
  AND2x2_ASAP7_75t_SL U51701 ( .A(n57215), .B(n59590), .Y(n56980) );
  INVx8_ASAP7_75t_SL U51702 ( .A(n58404), .Y(n59670) );
  BUFx3_ASAP7_75t_SL U51703 ( .A(n58404), .Y(n57321) );
  OR2x2_ASAP7_75t_SL U51704 ( .A(n58015), .B(n53271), .Y(n56981) );
  INVx6_ASAP7_75t_SL U51705 ( .A(n67922), .Y(n59600) );
  AND2x2_ASAP7_75t_SL U51706 ( .A(n64516), .B(n59352), .Y(n56982) );
  AND2x2_ASAP7_75t_SL U51707 ( .A(n57179), .B(n75947), .Y(n56983) );
  OAI21x1_ASAP7_75t_SL U51708 ( .A1(n64514), .A2(n64513), .B(n59351), .Y(
        n59350) );
  AO21x1_ASAP7_75t_SL U51709 ( .A1(n75906), .A2(n58863), .B(n58864), .Y(n56984) );
  OR2x2_ASAP7_75t_SL U51710 ( .A(n66616), .B(n66615), .Y(n56985) );
  XOR2x2_ASAP7_75t_SL U51711 ( .A(n58919), .B(n57436), .Y(n56987) );
  OR2x2_ASAP7_75t_SL U51712 ( .A(n56984), .B(n59446), .Y(n56988) );
  OR2x2_ASAP7_75t_SL U51713 ( .A(n67822), .B(n59042), .Y(n56989) );
  AO21x1_ASAP7_75t_SL U51714 ( .A1(n59282), .A2(n57409), .B(n67245), .Y(n56990) );
  INVx4_ASAP7_75t_SL U51715 ( .A(n59659), .Y(n59658) );
  INVx2_ASAP7_75t_SL U51716 ( .A(n59590), .Y(n58176) );
  NAND2x2_ASAP7_75t_SL U51717 ( .A(n64395), .B(n64394), .Y(n76078) );
  OR2x2_ASAP7_75t_SL U51718 ( .A(n67740), .B(n67741), .Y(n56991) );
  OR2x2_ASAP7_75t_SL U51719 ( .A(n58672), .B(n67463), .Y(n56992) );
  INVx4_ASAP7_75t_SL U51720 ( .A(n67230), .Y(n57941) );
  OA21x2_ASAP7_75t_SL U51721 ( .A1(n67607), .A2(n58432), .B(n68011), .Y(n56993) );
  OR2x2_ASAP7_75t_SL U51722 ( .A(n75922), .B(n59519), .Y(n56994) );
  NOR2x1_ASAP7_75t_SL U51723 ( .A(n75032), .B(n67454), .Y(n58706) );
  AND2x2_ASAP7_75t_SL U51724 ( .A(n57260), .B(n66696), .Y(n56995) );
  AND2x2_ASAP7_75t_SL U51725 ( .A(n57284), .B(n67713), .Y(n56996) );
  NAND2x1_ASAP7_75t_SL U51726 ( .A(n75032), .B(n67641), .Y(n75076) );
  INVx2_ASAP7_75t_SL U51727 ( .A(n67641), .Y(n67284) );
  AOI21xp33_ASAP7_75t_SRAM U51728 ( .A1(n59510), .A2(n68409), .B(n66629), .Y(
        n56997) );
  OR2x2_ASAP7_75t_SL U51729 ( .A(n58706), .B(n67894), .Y(n56998) );
  INVx6_ASAP7_75t_SL U51730 ( .A(n67959), .Y(n59605) );
  OR2x2_ASAP7_75t_SL U51731 ( .A(n59012), .B(n66701), .Y(n57000) );
  OA21x2_ASAP7_75t_SL U51732 ( .A1(n58884), .A2(n67384), .B(n57002), .Y(n57001) );
  OR2x2_ASAP7_75t_SL U51733 ( .A(n67515), .B(n59012), .Y(n57002) );
  AO22x1_ASAP7_75t_SL U51734 ( .A1(n67829), .A2(n66931), .B1(n57706), .B2(
        n66930), .Y(n57003) );
  INVx1_ASAP7_75t_SL U51735 ( .A(n59012), .Y(n57706) );
  INVx1_ASAP7_75t_SL U51736 ( .A(n57698), .Y(n59231) );
  OR2x2_ASAP7_75t_SL U51737 ( .A(n62576), .B(n62579), .Y(n58856) );
  AND2x4_ASAP7_75t_SL U51738 ( .A(n64354), .B(n58238), .Y(n58786) );
  AND2x2_ASAP7_75t_SL U51739 ( .A(n59656), .B(n67071), .Y(n57004) );
  AO21x1_ASAP7_75t_SL U51740 ( .A1(n58439), .A2(n67736), .B(n64919), .Y(n57005) );
  AO21x1_ASAP7_75t_SL U51741 ( .A1(n57180), .A2(n59653), .B(n63658), .Y(n57006) );
  OR2x2_ASAP7_75t_SL U51742 ( .A(n59504), .B(n67866), .Y(n57007) );
  XOR2xp5_ASAP7_75t_SL U51743 ( .A(n67805), .B(n59450), .Y(n57008) );
  INVxp33_ASAP7_75t_SRAM U51744 ( .A(n67642), .Y(n67803) );
  AND2x2_ASAP7_75t_SL U51745 ( .A(n67551), .B(n67550), .Y(n57009) );
  INVx2_ASAP7_75t_SL U51746 ( .A(n68097), .Y(n58211) );
  AND2x2_ASAP7_75t_SL U51747 ( .A(n57336), .B(n68101), .Y(n57010) );
  OR2x2_ASAP7_75t_SL U51748 ( .A(n67819), .B(n68119), .Y(n57011) );
  OA21x2_ASAP7_75t_SL U51749 ( .A1(n67819), .A2(n57076), .B(n67602), .Y(n57012) );
  AND2x2_ASAP7_75t_SL U51750 ( .A(n66684), .B(n58336), .Y(n57013) );
  OA22x2_ASAP7_75t_SL U51751 ( .A1(n59116), .A2(n66730), .B1(n68119), .B2(
        n58507), .Y(n57014) );
  OA21x2_ASAP7_75t_SL U51752 ( .A1(n57720), .A2(n58861), .B(n58862), .Y(n57015) );
  OAI22x1_ASAP7_75t_SL U51753 ( .A1(n68014), .A2(n59460), .B1(n68013), .B2(
        n59515), .Y(n59478) );
  BUFx2_ASAP7_75t_SL U51754 ( .A(n59460), .Y(n57360) );
  INVx1_ASAP7_75t_SL U51755 ( .A(n75048), .Y(n75036) );
  OR2x2_ASAP7_75t_SL U51756 ( .A(n56987), .B(n57096), .Y(n57016) );
  AND2x2_ASAP7_75t_SL U51757 ( .A(n66471), .B(n57067), .Y(n57017) );
  OR2x2_ASAP7_75t_SL U51758 ( .A(n59652), .B(n67300), .Y(n57018) );
  AND2x2_ASAP7_75t_SL U51759 ( .A(n77278), .B(n66271), .Y(n57019) );
  NAND2x1p5_ASAP7_75t_SL U51760 ( .A(n59456), .B(n57656), .Y(n63120) );
  XOR2x2_ASAP7_75t_SL U51761 ( .A(n63134), .B(n63100), .Y(n57020) );
  OA21x2_ASAP7_75t_SL U51762 ( .A1(n67227), .A2(n63099), .B(n63098), .Y(n57021) );
  OR2x2_ASAP7_75t_SL U51763 ( .A(n64647), .B(n68383), .Y(n57022) );
  OR2x2_ASAP7_75t_SL U51764 ( .A(n63666), .B(n57759), .Y(n57024) );
  OR2x2_ASAP7_75t_SL U51765 ( .A(n58383), .B(n57484), .Y(n57025) );
  INVx8_ASAP7_75t_SL U51766 ( .A(n58383), .Y(n59601) );
  OA21x2_ASAP7_75t_SL U51767 ( .A1(n67242), .A2(n57111), .B(n64370), .Y(n57027) );
  XOR2x2_ASAP7_75t_SL U51768 ( .A(n68110), .B(n68109), .Y(n57028) );
  BUFx6f_ASAP7_75t_SL U51769 ( .A(n75438), .Y(n57505) );
  AND2x2_ASAP7_75t_SL U51770 ( .A(n58851), .B(n68418), .Y(n57029) );
  OR2x2_ASAP7_75t_SL U51771 ( .A(n57099), .B(n67708), .Y(n57030) );
  INVx4_ASAP7_75t_SL U51772 ( .A(n57099), .Y(n57161) );
  AO21x1_ASAP7_75t_SL U51773 ( .A1(n64567), .A2(n66483), .B(n66501), .Y(n57031) );
  XNOR2x2_ASAP7_75t_SL U51774 ( .A(n68184), .B(n68183), .Y(n58352) );
  AND2x2_ASAP7_75t_SL U51775 ( .A(n58486), .B(n66810), .Y(n57032) );
  XOR2xp5_ASAP7_75t_SL U51776 ( .A(n67794), .B(n67795), .Y(n57034) );
  BUFx3_ASAP7_75t_SL U51777 ( .A(n57567), .Y(n59171) );
  OR2x2_ASAP7_75t_SL U51778 ( .A(n58059), .B(n57156), .Y(n57035) );
  INVx2_ASAP7_75t_SL U51779 ( .A(n59171), .Y(n59073) );
  INVx3_ASAP7_75t_SL U51780 ( .A(n59507), .Y(n75761) );
  OR2x2_ASAP7_75t_SL U51781 ( .A(n59656), .B(n57108), .Y(n57036) );
  OR2x2_ASAP7_75t_SL U51782 ( .A(n64646), .B(n64645), .Y(n57037) );
  AND2x2_ASAP7_75t_SL U51783 ( .A(n59664), .B(n67883), .Y(n57038) );
  AND2x2_ASAP7_75t_SL U51784 ( .A(n59506), .B(n67750), .Y(n57039) );
  XOR2xp5_ASAP7_75t_SL U51785 ( .A(n53317), .B(n59650), .Y(n57040) );
  XOR2x2_ASAP7_75t_SL U51786 ( .A(n63109), .B(n58111), .Y(n57041) );
  OR2x2_ASAP7_75t_SL U51787 ( .A(n67271), .B(n67974), .Y(n57042) );
  OA21x2_ASAP7_75t_SL U51788 ( .A1(n57041), .A2(n58182), .B(n58181), .Y(n57043) );
  INVx2_ASAP7_75t_SL U51789 ( .A(n67974), .Y(n57157) );
  INVx2_ASAP7_75t_SL U51790 ( .A(n64743), .Y(n64744) );
  XNOR2x2_ASAP7_75t_SL U51791 ( .A(n68279), .B(n68280), .Y(n57045) );
  XNOR2x1_ASAP7_75t_SL U51792 ( .A(n62992), .B(n63004), .Y(n62995) );
  OR2x2_ASAP7_75t_SL U51793 ( .A(n67898), .B(n67097), .Y(n57046) );
  NAND2x1_ASAP7_75t_SL U51794 ( .A(n64043), .B(n64076), .Y(n64677) );
  AND2x2_ASAP7_75t_SL U51795 ( .A(n57111), .B(n66623), .Y(n57047) );
  AND2x2_ASAP7_75t_SL U51796 ( .A(n67483), .B(n67484), .Y(n57048) );
  XNOR2x2_ASAP7_75t_SL U51797 ( .A(n68374), .B(n67745), .Y(n68372) );
  XOR2x2_ASAP7_75t_SL U51798 ( .A(n67586), .B(n75908), .Y(n57049) );
  NOR2x1p5_ASAP7_75t_SL U51799 ( .A(n57152), .B(n58904), .Y(n57877) );
  XOR2xp5_ASAP7_75t_SL U51800 ( .A(n57472), .B(n57471), .Y(n57050) );
  AND2x2_ASAP7_75t_SL U51801 ( .A(n66902), .B(n66901), .Y(n57051) );
  XOR2xp5_ASAP7_75t_SL U51802 ( .A(n57051), .B(n66838), .Y(n57052) );
  OA21x2_ASAP7_75t_SL U51803 ( .A1(n53487), .A2(n58151), .B(n58150), .Y(n57053) );
  NAND2xp5_ASAP7_75t_SL U51804 ( .A(n57369), .B(n53206), .Y(n69115) );
  INVx2_ASAP7_75t_SL U51805 ( .A(n57902), .Y(n69233) );
  XOR2xp5_ASAP7_75t_SL U51806 ( .A(n67160), .B(n57658), .Y(n57054) );
  OA21x2_ASAP7_75t_SL U51807 ( .A1(n58740), .A2(n58739), .B(n58738), .Y(n57055) );
  AND2x2_ASAP7_75t_SL U51808 ( .A(n58689), .B(n59221), .Y(n57056) );
  AND2x2_ASAP7_75t_SL U51809 ( .A(n64667), .B(n64089), .Y(n57057) );
  XNOR2x2_ASAP7_75t_SL U51810 ( .A(n59372), .B(n68168), .Y(n68283) );
  AOI21x1_ASAP7_75t_SL U51811 ( .A1(n68300), .A2(n68298), .B(n68297), .Y(
        n68323) );
  AO21x1_ASAP7_75t_SL U51812 ( .A1(n57495), .A2(n66808), .B(n66807), .Y(n57058) );
  NOR2xp33_ASAP7_75t_SL U51813 ( .A(n68677), .B(n59449), .Y(n57059) );
  AND2x2_ASAP7_75t_SL U51814 ( .A(n69028), .B(n69029), .Y(n57060) );
  NOR2x1p5_ASAP7_75t_SL U51815 ( .A(n68835), .B(n68826), .Y(n68904) );
  INVx1_ASAP7_75t_SL U51816 ( .A(n58887), .Y(n58885) );
  AND2x2_ASAP7_75t_SL U51817 ( .A(n58258), .B(n68865), .Y(n57061) );
  MAJx2_ASAP7_75t_SL U51818 ( .A(n68228), .B(n68334), .C(n68227), .Y(n57062)
         );
  AND3x1_ASAP7_75t_SL U51819 ( .A(n58349), .B(n59063), .C(n68806), .Y(n57063)
         );
  INVx1_ASAP7_75t_SL U51820 ( .A(n63477), .Y(n63478) );
  XNOR2x2_ASAP7_75t_SL U51821 ( .A(n63042), .B(n63037), .Y(n63477) );
  HB1xp67_ASAP7_75t_SL U51822 ( .A(n57808), .Y(n57434) );
  NAND2xp5_ASAP7_75t_SL U51823 ( .A(n66939), .B(n66941), .Y(n66973) );
  BUFx2_ASAP7_75t_SL U51824 ( .A(n64892), .Y(n57064) );
  NOR2xp33_ASAP7_75t_SL U51825 ( .A(n68107), .B(n68000), .Y(n67933) );
  XNOR2x2_ASAP7_75t_SL U51826 ( .A(n67406), .B(n67405), .Y(n67259) );
  BUFx2_ASAP7_75t_SL U51827 ( .A(n67567), .Y(n57065) );
  NAND3xp33_ASAP7_75t_SL U51828 ( .A(n67837), .B(n59599), .C(n59436), .Y(
        n67567) );
  INVx1_ASAP7_75t_SL U51829 ( .A(n63475), .Y(n76224) );
  NOR2x1_ASAP7_75t_SL U51830 ( .A(n63047), .B(n63046), .Y(n63475) );
  HB1xp67_ASAP7_75t_SL U51831 ( .A(n68915), .Y(n57335) );
  XNOR2x1_ASAP7_75t_SL U51832 ( .A(n57516), .B(n59381), .Y(n67314) );
  XNOR2x1_ASAP7_75t_SL U51833 ( .A(n63831), .B(n63830), .Y(n64087) );
  NOR2x1p5_ASAP7_75t_SL U51834 ( .A(n59136), .B(n59137), .Y(n67772) );
  OAI22xp5_ASAP7_75t_SL U51835 ( .A1(n67220), .A2(n67219), .B1(n68586), .B2(
        n68585), .Y(n67221) );
  NAND2x1p5_ASAP7_75t_SL U51836 ( .A(n68586), .B(n74557), .Y(n68648) );
  NOR2x1_ASAP7_75t_SL U51837 ( .A(n74554), .B(n68692), .Y(n68586) );
  INVx8_ASAP7_75t_SL U51838 ( .A(n58788), .Y(n59440) );
  NOR2x1_ASAP7_75t_SL U51839 ( .A(n67819), .B(n57076), .Y(n57848) );
  OAI22xp5_ASAP7_75t_SL U51840 ( .A1(n67872), .A2(n57076), .B1(n67852), .B2(
        n68119), .Y(n57225) );
  NOR2x1p5_ASAP7_75t_SL U51841 ( .A(n66307), .B(n66302), .Y(n75643) );
  XNOR2xp5_ASAP7_75t_SL U51842 ( .A(n56842), .B(n67699), .Y(n57545) );
  AOI22x1_ASAP7_75t_SL U51843 ( .A1(n64953), .A2(n64952), .B1(n64954), .B2(
        n67251), .Y(n65011) );
  BUFx2_ASAP7_75t_SL U51844 ( .A(n59444), .Y(n57066) );
  BUFx6f_ASAP7_75t_SL U51845 ( .A(n59444), .Y(n57067) );
  NOR2x1p5_ASAP7_75t_SL U51846 ( .A(n58676), .B(n66301), .Y(n59348) );
  XNOR2x1_ASAP7_75t_SL U51847 ( .A(n67796), .B(n57034), .Y(n58963) );
  NAND2xp5_ASAP7_75t_SL U51848 ( .A(n59619), .B(n63149), .Y(n63093) );
  INVx6_ASAP7_75t_SL U51849 ( .A(n58070), .Y(n57099) );
  BUFx3_ASAP7_75t_SL U51850 ( .A(n64504), .Y(n59400) );
  BUFx3_ASAP7_75t_SL U51851 ( .A(n1606), .Y(n57068) );
  BUFx6f_ASAP7_75t_SL U51852 ( .A(n1949), .Y(n59554) );
  NAND2xp67_ASAP7_75t_SRAM U51853 ( .A(n59664), .B(n67864), .Y(n67318) );
  NOR2x1p5_ASAP7_75t_SL U51854 ( .A(n77715), .B(n64930), .Y(n64509) );
  NAND2x2_ASAP7_75t_SL U51855 ( .A(n59276), .B(n58056), .Y(n64930) );
  NOR2x1_ASAP7_75t_SL U51856 ( .A(n59374), .B(n65023), .Y(n68167) );
  NAND2x2_ASAP7_75t_SL U51857 ( .A(n67328), .B(n57098), .Y(n59229) );
  NAND2xp5_ASAP7_75t_SL U51858 ( .A(n57210), .B(n66244), .Y(n57666) );
  HB1xp67_ASAP7_75t_SL U51859 ( .A(n59188), .Y(n57493) );
  XOR2x2_ASAP7_75t_SL U51860 ( .A(n67979), .B(n58488), .Y(n57980) );
  BUFx2_ASAP7_75t_SL U51861 ( .A(n59356), .Y(n57508) );
  BUFx2_ASAP7_75t_SL U51862 ( .A(n67834), .Y(n57069) );
  NOR2x1p5_ASAP7_75t_SL U51863 ( .A(n58828), .B(n63175), .Y(n67897) );
  NAND2x1p5_ASAP7_75t_SL U51864 ( .A(n59462), .B(n62562), .Y(n57250) );
  OAI21x1_ASAP7_75t_SL U51865 ( .A1(n66768), .A2(n67434), .B(n57046), .Y(
        n66874) );
  NOR2x2_ASAP7_75t_SL U51866 ( .A(n57653), .B(n58176), .Y(n58173) );
  NAND2xp5_ASAP7_75t_SL U51867 ( .A(n58484), .B(n58652), .Y(n58651) );
  BUFx2_ASAP7_75t_SL U51868 ( .A(n59360), .Y(n58715) );
  XNOR2x1_ASAP7_75t_SL U51869 ( .A(n67684), .B(n67685), .Y(n59160) );
  HB1xp67_ASAP7_75t_SL U51870 ( .A(n68394), .Y(n58366) );
  NAND2x1_ASAP7_75t_SL U51871 ( .A(n67108), .B(n67107), .Y(n69143) );
  XNOR2x2_ASAP7_75t_SL U51872 ( .A(n59596), .B(n53241), .Y(n66412) );
  NOR2x1_ASAP7_75t_SL U51873 ( .A(n67242), .B(n67635), .Y(n67945) );
  INVx2_ASAP7_75t_SL U51874 ( .A(n68396), .Y(n59024) );
  XNOR2x2_ASAP7_75t_SL U51875 ( .A(n58880), .B(n58924), .Y(n68340) );
  XNOR2x1_ASAP7_75t_SL U51876 ( .A(n57374), .B(n67811), .Y(n57668) );
  NOR2x1_ASAP7_75t_SL U51877 ( .A(n62594), .B(n59482), .Y(n62636) );
  XNOR2xp5_ASAP7_75t_SL U51878 ( .A(n67680), .B(n59159), .Y(n67698) );
  NOR2x1_ASAP7_75t_SL U51879 ( .A(n68850), .B(n68860), .Y(n68906) );
  NOR2xp33_ASAP7_75t_SL U51880 ( .A(n68850), .B(n58088), .Y(n58086) );
  XOR2x1_ASAP7_75t_SL U51881 ( .A(n57597), .B(n63164), .Y(n63160) );
  NAND2x1p5_ASAP7_75t_SL U51882 ( .A(n69083), .B(n69082), .Y(n58881) );
  AOI21x1_ASAP7_75t_SL U51883 ( .A1(n58267), .A2(n57145), .B(n58266), .Y(
        n68148) );
  XNOR2x1_ASAP7_75t_SL U51884 ( .A(n67100), .B(n67010), .Y(n67105) );
  NAND2xp5_ASAP7_75t_SL U51885 ( .A(n69116), .B(n58881), .Y(n57602) );
  NOR2xp33_ASAP7_75t_SL U51886 ( .A(n74558), .B(n75287), .Y(n75285) );
  AOI21xp33_ASAP7_75t_SL U51887 ( .A1(n69152), .A2(n69151), .B(n69150), .Y(
        n69153) );
  INVxp67_ASAP7_75t_SL U51888 ( .A(n68923), .Y(n68926) );
  NOR2xp33_ASAP7_75t_SL U51889 ( .A(n58085), .B(n68908), .Y(n68957) );
  OAI21xp33_ASAP7_75t_SL U51890 ( .A1(or1200_cpu_or1200_mult_mac_n128), .A2(
        n57105), .B(n76196), .Y(or1200_cpu_or1200_mult_mac_n1527) );
  AOI21xp33_ASAP7_75t_SL U51891 ( .A1(n69227), .A2(n57087), .B(n69225), .Y(
        n69231) );
  NAND2x1_ASAP7_75t_SL U51892 ( .A(n57062), .B(n59480), .Y(n68973) );
  HB1xp67_ASAP7_75t_SL U51893 ( .A(n68667), .Y(n57376) );
  HB1xp67_ASAP7_75t_SL U51894 ( .A(n53296), .Y(n57341) );
  NAND2xp5_ASAP7_75t_SL U51895 ( .A(n68634), .B(n68633), .Y(n68667) );
  OAI21xp33_ASAP7_75t_SL U51896 ( .A1(n1025), .A2(n53448), .B(n77318), .Y(
        n9678) );
  OAI21xp33_ASAP7_75t_SL U51897 ( .A1(n962), .A2(n53448), .B(n77330), .Y(n9685) );
  AOI21xp5_ASAP7_75t_SL U51898 ( .A1(n57135), .A2(n75200), .B(n75199), .Y(
        n75201) );
  OAI21xp33_ASAP7_75t_SL U51899 ( .A1(n953), .A2(n53448), .B(n77329), .Y(n9686) );
  AOI21xp5_ASAP7_75t_SL U51900 ( .A1(n57135), .A2(n77227), .B(n77226), .Y(
        n77228) );
  AOI21xp5_ASAP7_75t_SL U51901 ( .A1(n57135), .A2(n77179), .B(n77178), .Y(
        n77180) );
  AOI21xp5_ASAP7_75t_SL U51902 ( .A1(n57135), .A2(n75686), .B(n75676), .Y(
        n75677) );
  OAI21xp33_ASAP7_75t_SL U51903 ( .A1(n1016), .A2(n53448), .B(n77326), .Y(
        n9679) );
  OAI21xp33_ASAP7_75t_SL U51904 ( .A1(n944), .A2(n53448), .B(n77333), .Y(n9687) );
  AOI21xp5_ASAP7_75t_SL U51905 ( .A1(n57135), .A2(n77021), .B(n77020), .Y(
        n77022) );
  OAI21xp33_ASAP7_75t_SL U51906 ( .A1(n935), .A2(n53448), .B(n77320), .Y(n9688) );
  AOI21xp5_ASAP7_75t_SL U51907 ( .A1(n57135), .A2(n77153), .B(n77152), .Y(
        n77154) );
  OAI21xp33_ASAP7_75t_SL U51908 ( .A1(n1007), .A2(n53448), .B(n77319), .Y(
        n9680) );
  AOI21xp5_ASAP7_75t_SL U51909 ( .A1(n57135), .A2(n76232), .B(n76231), .Y(
        n76233) );
  AOI21xp5_ASAP7_75t_SL U51910 ( .A1(n57135), .A2(n75798), .B(n75797), .Y(
        n75799) );
  OAI21xp33_ASAP7_75t_SL U51911 ( .A1(n998), .A2(n53448), .B(n77331), .Y(n9681) );
  OAI21xp33_ASAP7_75t_SL U51912 ( .A1(n971), .A2(n53448), .B(n77328), .Y(n9684) );
  AOI21xp5_ASAP7_75t_SL U51913 ( .A1(n57135), .A2(n69373), .B(n69372), .Y(
        n69374) );
  OAI21xp33_ASAP7_75t_SL U51914 ( .A1(n989), .A2(n53448), .B(n77325), .Y(n9682) );
  AOI21xp5_ASAP7_75t_SL U51915 ( .A1(n57135), .A2(n74081), .B(n74080), .Y(
        n74086) );
  AOI21xp5_ASAP7_75t_SL U51916 ( .A1(n57135), .A2(n74129), .B(n74128), .Y(
        n74130) );
  AOI21xp5_ASAP7_75t_SL U51917 ( .A1(n57135), .A2(n74047), .B(n74046), .Y(
        n74048) );
  AOI21xp5_ASAP7_75t_SL U51918 ( .A1(n57135), .A2(n75449), .B(n75448), .Y(
        n75450) );
  OAI21xp33_ASAP7_75t_SL U51919 ( .A1(n980), .A2(n53448), .B(n77324), .Y(n9683) );
  AOI21xp5_ASAP7_75t_SL U51920 ( .A1(n57135), .A2(n76999), .B(n76998), .Y(
        n77000) );
  AOI21xp5_ASAP7_75t_SL U51921 ( .A1(n57135), .A2(n77277), .B(n76207), .Y(
        n76208) );
  OAI21xp33_ASAP7_75t_SL U51922 ( .A1(n881), .A2(n53448), .B(n77317), .Y(n9694) );
  OAI21xp33_ASAP7_75t_SL U51923 ( .A1(n863), .A2(n53448), .B(n77334), .Y(n9696) );
  OAI21xp33_ASAP7_75t_SL U51924 ( .A1(n917), .A2(n53448), .B(n77321), .Y(n9690) );
  AOI21xp5_ASAP7_75t_SL U51925 ( .A1(n57135), .A2(n76619), .B(n76618), .Y(
        n76620) );
  OAI21xp33_ASAP7_75t_SL U51926 ( .A1(n890), .A2(n53448), .B(n77332), .Y(n9693) );
  OAI21xp33_ASAP7_75t_SL U51927 ( .A1(n852), .A2(n53448), .B(n77316), .Y(n9697) );
  AOI21xp5_ASAP7_75t_SL U51928 ( .A1(n57135), .A2(n76704), .B(n76697), .Y(
        n76698) );
  AOI21xp5_ASAP7_75t_SL U51929 ( .A1(n57135), .A2(n76851), .B(n76640), .Y(
        n76641) );
  OAI21xp33_ASAP7_75t_SL U51930 ( .A1(n899), .A2(n53448), .B(n77335), .Y(n9692) );
  OAI21xp33_ASAP7_75t_SL U51931 ( .A1(n872), .A2(n53448), .B(n77327), .Y(n9695) );
  AOI21xp5_ASAP7_75t_SL U51932 ( .A1(n57135), .A2(n76253), .B(n76246), .Y(
        n76247) );
  OAI21xp33_ASAP7_75t_SL U51933 ( .A1(n908), .A2(n53448), .B(n77322), .Y(n9691) );
  OAI21xp33_ASAP7_75t_SL U51934 ( .A1(n926), .A2(n53448), .B(n77323), .Y(n9689) );
  NAND2x1p5_ASAP7_75t_SL U51935 ( .A(n63497), .B(n63257), .Y(n64743) );
  INVx1_ASAP7_75t_SL U51936 ( .A(n58298), .Y(n74270) );
  NAND2xp33_ASAP7_75t_SL U51937 ( .A(icqmem_adr_qmem[13]), .B(n57136), .Y(
        n77334) );
  NAND2xp33_ASAP7_75t_SL U51938 ( .A(icqmem_adr_qmem[14]), .B(n57136), .Y(
        n77327) );
  NAND2xp33_ASAP7_75t_SL U51939 ( .A(icqmem_adr_qmem[15]), .B(n57136), .Y(
        n77317) );
  NAND2xp33_ASAP7_75t_SL U51940 ( .A(n77315), .B(n57136), .Y(n77316) );
  NAND2xp33_ASAP7_75t_SL U51941 ( .A(icqmem_adr_qmem[16]), .B(n57136), .Y(
        n77332) );
  NAND2xp33_ASAP7_75t_SL U51942 ( .A(icqmem_adr_qmem[17]), .B(n57136), .Y(
        n77335) );
  NAND2xp33_ASAP7_75t_SL U51943 ( .A(icqmem_adr_qmem[19]), .B(n57136), .Y(
        n77321) );
  INVxp67_ASAP7_75t_SL U51944 ( .A(n66607), .Y(n66608) );
  NAND2xp33_ASAP7_75t_SL U51945 ( .A(icqmem_adr_qmem[18]), .B(n57136), .Y(
        n77322) );
  OAI22xp33_ASAP7_75t_SL U51946 ( .A1(or1200_cpu_or1200_except_n208), .A2(
        n77240), .B1(n75781), .B2(n57138), .Y(n63717) );
  OAI22xp33_ASAP7_75t_SL U51947 ( .A1(or1200_cpu_or1200_except_n194), .A2(
        n77240), .B1(n77591), .B2(n57138), .Y(n76573) );
  BUFx3_ASAP7_75t_SL U51948 ( .A(n76931), .Y(n57088) );
  OAI22xp33_ASAP7_75t_SL U51949 ( .A1(or1200_cpu_or1200_except_n188), .A2(
        n77240), .B1(n77583), .B2(n57138), .Y(or1200_cpu_or1200_except_n1784)
         );
  OAI22xp33_ASAP7_75t_SL U51950 ( .A1(or1200_cpu_or1200_except_n206), .A2(
        n77240), .B1(n76508), .B2(n57138), .Y(n76251) );
  OAI22xp33_ASAP7_75t_SL U51951 ( .A1(or1200_cpu_epcr_1_), .A2(n77240), .B1(
        n77585), .B2(n57138), .Y(or1200_cpu_or1200_except_n1783) );
  OAI22xp33_ASAP7_75t_SL U51952 ( .A1(or1200_cpu_or1200_except_n192), .A2(
        n77240), .B1(n76688), .B2(n57138), .Y(n76564) );
  OAI22xp33_ASAP7_75t_SL U51953 ( .A1(or1200_cpu_or1200_except_n216), .A2(
        n77240), .B1(n77019), .B2(n57138), .Y(n63971) );
  OAI22xp33_ASAP7_75t_SL U51954 ( .A1(or1200_cpu_or1200_except_n200), .A2(
        n77240), .B1(n77600), .B2(n57138), .Y(n76597) );
  OAI22xp33_ASAP7_75t_SL U51955 ( .A1(or1200_cpu_or1200_except_n204), .A2(
        n77240), .B1(n76828), .B2(n57138), .Y(n76645) );
  OAI22xp33_ASAP7_75t_SL U51956 ( .A1(or1200_cpu_or1200_except_n214), .A2(
        n77240), .B1(n77637), .B2(n57138), .Y(n63959) );
  OAI22xp33_ASAP7_75t_SL U51957 ( .A1(or1200_cpu_or1200_except_n196), .A2(
        n77240), .B1(n77594), .B2(n57138), .Y(n76583) );
  OAI22xp33_ASAP7_75t_SL U51958 ( .A1(or1200_cpu_or1200_except_n212), .A2(
        n77240), .B1(n77295), .B2(n57138), .Y(n63948) );
  OAI22xp33_ASAP7_75t_SL U51959 ( .A1(or1200_cpu_or1200_except_n198), .A2(
        n77240), .B1(n77597), .B2(n57138), .Y(n76212) );
  OAI22xp33_ASAP7_75t_SL U51960 ( .A1(or1200_cpu_or1200_except_n202), .A2(
        n77240), .B1(n77603), .B2(n57138), .Y(n76702) );
  OAI22xp33_ASAP7_75t_SL U51961 ( .A1(or1200_cpu_or1200_except_n210), .A2(
        n77240), .B1(n77615), .B2(n57138), .Y(n76525) );
  OAI22xp33_ASAP7_75t_SL U51962 ( .A1(or1200_cpu_or1200_except_n224), .A2(
        n77240), .B1(n74984), .B2(n57138), .Y(n74963) );
  OAI22xp33_ASAP7_75t_SL U51963 ( .A1(or1200_cpu_or1200_except_n226), .A2(
        n77240), .B1(n74639), .B2(n57138), .Y(n63922) );
  OAI22xp33_ASAP7_75t_SL U51964 ( .A1(or1200_cpu_or1200_except_n228), .A2(
        n77240), .B1(n74127), .B2(n57138), .Y(n64159) );
  OAI22xp33_ASAP7_75t_SL U51965 ( .A1(or1200_cpu_or1200_except_n230), .A2(
        n77240), .B1(n75431), .B2(n57138), .Y(n75411) );
  OAI22xp33_ASAP7_75t_SL U51966 ( .A1(or1200_cpu_or1200_except_n232), .A2(
        n77240), .B1(n75447), .B2(n57138), .Y(n64261) );
  OAI22xp33_ASAP7_75t_SL U51967 ( .A1(or1200_cpu_or1200_except_n234), .A2(
        n77240), .B1(n75620), .B2(n57138), .Y(n75537) );
  OAI22xp33_ASAP7_75t_SL U51968 ( .A1(or1200_cpu_or1200_except_n236), .A2(
        n77240), .B1(n74045), .B2(n57138), .Y(n65198) );
  OAI22xp33_ASAP7_75t_SL U51969 ( .A1(or1200_cpu_or1200_except_n238), .A2(
        n77240), .B1(n74079), .B2(n57138), .Y(n65215) );
  OAI22xp33_ASAP7_75t_SL U51970 ( .A1(or1200_cpu_or1200_except_n240), .A2(
        n77240), .B1(n69371), .B2(n57138), .Y(n65188) );
  OAI22xp33_ASAP7_75t_SL U51971 ( .A1(or1200_cpu_or1200_except_n242), .A2(
        n77240), .B1(n75796), .B2(n57138), .Y(n75152) );
  OAI22xp33_ASAP7_75t_SL U51972 ( .A1(or1200_cpu_or1200_except_n244), .A2(
        n77240), .B1(n77177), .B2(n57138), .Y(n75166) );
  OAI22xp33_ASAP7_75t_SL U51973 ( .A1(or1200_cpu_or1200_except_n246), .A2(
        n77240), .B1(n75198), .B2(n57138), .Y(n75177) );
  OAI22xp33_ASAP7_75t_SL U51974 ( .A1(or1200_cpu_or1200_except_n248), .A2(
        n77240), .B1(n75675), .B2(n57138), .Y(n75634) );
  OAI22xp33_ASAP7_75t_SL U51975 ( .A1(or1200_cpu_epcr_31_), .A2(n77240), .B1(
        n77673), .B2(n57138), .Y(n76924) );
  OAI22xp33_ASAP7_75t_SL U51976 ( .A1(or1200_cpu_or1200_except_n222), .A2(
        n77240), .B1(n75302), .B2(n57138), .Y(n63927) );
  OAI22xp33_ASAP7_75t_SL U51977 ( .A1(or1200_cpu_or1200_except_n220), .A2(
        n77240), .B1(n76235), .B2(n57138), .Y(n63932) );
  OAI22xp33_ASAP7_75t_SL U51978 ( .A1(or1200_cpu_or1200_except_n218), .A2(
        n77240), .B1(n77646), .B2(n57138), .Y(n63990) );
  NAND2xp5_ASAP7_75t_SL U51979 ( .A(n57650), .B(n62781), .Y(n63242) );
  BUFx6f_ASAP7_75t_SL U51980 ( .A(n77296), .Y(n57070) );
  AOI22xp33_ASAP7_75t_SL U51981 ( .A1(n77237), .A2(n77922), .B1(n77236), .B2(
        n77235), .Y(n77238) );
  NOR2x1p5_ASAP7_75t_SL U51982 ( .A(n69349), .B(n77235), .Y(n77290) );
  AOI22xp33_ASAP7_75t_SL U51983 ( .A1(n57090), .A2(n76584), .B1(n61575), .B2(
        n57137), .Y(n61576) );
  AOI22xp33_ASAP7_75t_SL U51984 ( .A1(n57090), .A2(n76607), .B1(n76606), .B2(
        n57137), .Y(n76608) );
  AOI22xp33_ASAP7_75t_SL U51985 ( .A1(n57090), .A2(n63954), .B1(n63698), .B2(
        n57137), .Y(n63699) );
  AOI22xp33_ASAP7_75t_SL U51986 ( .A1(n57090), .A2(n76252), .B1(n61278), .B2(
        n57137), .Y(n61279) );
  AOI22xp33_ASAP7_75t_SL U51987 ( .A1(n57090), .A2(n76703), .B1(n63739), .B2(
        n57137), .Y(n63740) );
  AOI22xp33_ASAP7_75t_SL U51988 ( .A1(n57090), .A2(n76565), .B1(n63748), .B2(
        n57137), .Y(n63749) );
  AOI22xp33_ASAP7_75t_SL U51989 ( .A1(n57090), .A2(n76574), .B1(n61587), .B2(
        n57137), .Y(n61588) );
  AOI22xp33_ASAP7_75t_SL U51990 ( .A1(n57090), .A2(n63998), .B1(n63997), .B2(
        n57137), .Y(n63999) );
  AOI22xp33_ASAP7_75t_SL U51991 ( .A1(n57090), .A2(n64006), .B1(n64005), .B2(
        n57137), .Y(n64007) );
  AOI22xp33_ASAP7_75t_SL U51992 ( .A1(n57090), .A2(n75186), .B1(n75185), .B2(
        n57137), .Y(n75187) );
  INVx2_ASAP7_75t_SL U51993 ( .A(n63713), .Y(n77240) );
  AOI22xp33_ASAP7_75t_SL U51994 ( .A1(n57090), .A2(n75167), .B1(n75163), .B2(
        n57137), .Y(n75164) );
  AOI22xp33_ASAP7_75t_SL U51995 ( .A1(n57090), .A2(n74970), .B1(n74969), .B2(
        n57137), .Y(n74971) );
  AOI22xp33_ASAP7_75t_SL U51996 ( .A1(n57090), .A2(n64015), .B1(n64014), .B2(
        n57137), .Y(n64016) );
  AOI22xp33_ASAP7_75t_SL U51997 ( .A1(n57090), .A2(n75153), .B1(n75149), .B2(
        n57137), .Y(n75150) );
  AOI22xp33_ASAP7_75t_SL U51998 ( .A1(n57090), .A2(n64165), .B1(n64164), .B2(
        n57137), .Y(n64166) );
  AOI22xp33_ASAP7_75t_SL U51999 ( .A1(n57090), .A2(n75421), .B1(n75420), .B2(
        n57137), .Y(n75422) );
  HB1xp67_ASAP7_75t_SL U52000 ( .A(n76225), .Y(n57245) );
  AOI22xp33_ASAP7_75t_SL U52001 ( .A1(n57090), .A2(n64267), .B1(n64266), .B2(
        n57137), .Y(n64268) );
  AOI22xp33_ASAP7_75t_SL U52002 ( .A1(n57090), .A2(n65234), .B1(n65233), .B2(
        n57137), .Y(n65235) );
  AOI22xp33_ASAP7_75t_SL U52003 ( .A1(n57090), .A2(n75546), .B1(n75545), .B2(
        n57137), .Y(n75547) );
  AOI22xp33_ASAP7_75t_SL U52004 ( .A1(n57090), .A2(n65222), .B1(n65221), .B2(
        n57137), .Y(n65223) );
  AOI22xp33_ASAP7_75t_SL U52005 ( .A1(n57090), .A2(n65218), .B1(n65195), .B2(
        n57137), .Y(n65196) );
  AOI22xp33_ASAP7_75t_SL U52006 ( .A1(n57090), .A2(n76534), .B1(n76533), .B2(
        n57137), .Y(n76535) );
  INVx1_ASAP7_75t_SL U52007 ( .A(n76659), .Y(n77220) );
  INVx1_ASAP7_75t_SL U52008 ( .A(n76507), .Y(n77215) );
  AOI22xp33_ASAP7_75t_SL U52009 ( .A1(n57090), .A2(n63949), .B1(n63945), .B2(
        n57137), .Y(n63946) );
  AOI22xp33_ASAP7_75t_SL U52010 ( .A1(n57090), .A2(n76925), .B1(n76917), .B2(
        n57137), .Y(n76918) );
  BUFx2_ASAP7_75t_SL U52011 ( .A(n77239), .Y(n57138) );
  NAND2xp5_ASAP7_75t_SL U52012 ( .A(n75613), .B(n75612), .Y(n77874) );
  INVxp67_ASAP7_75t_SL U52013 ( .A(n77374), .Y(n61042) );
  OR2x4_ASAP7_75t_SL U52014 ( .A(n59703), .B(n76846), .Y(n58524) );
  INVxp67_ASAP7_75t_SL U52015 ( .A(n74227), .Y(n73859) );
  NAND2xp33_ASAP7_75t_SL U52016 ( .A(n78010), .B(n57092), .Y(n7615) );
  INVxp67_ASAP7_75t_SL U52017 ( .A(n78006), .Y(n78020) );
  NAND2xp33_ASAP7_75t_SL U52018 ( .A(n78016), .B(n57092), .Y(n7625) );
  NAND2xp33_ASAP7_75t_SL U52019 ( .A(n78013), .B(n57092), .Y(n7620) );
  NAND2xp33_ASAP7_75t_SL U52020 ( .A(n78025), .B(n57092), .Y(n7635) );
  XNOR2xp5_ASAP7_75t_SL U52021 ( .A(n66822), .B(n66773), .Y(n66906) );
  INVx1_ASAP7_75t_SL U52022 ( .A(n63609), .Y(n63610) );
  NAND2xp5_ASAP7_75t_SL U52023 ( .A(n67757), .B(n53472), .Y(n58118) );
  NAND2xp33_ASAP7_75t_SL U52024 ( .A(or1200_cpu_rf_datab[3]), .B(n57091), .Y(
        n76872) );
  NAND2xp33_ASAP7_75t_SL U52025 ( .A(or1200_cpu_rf_datab[1]), .B(n57091), .Y(
        n61016) );
  NAND2xp33_ASAP7_75t_SL U52026 ( .A(or1200_cpu_rf_datab[4]), .B(n57091), .Y(
        n77008) );
  INVx1_ASAP7_75t_SL U52027 ( .A(n67757), .Y(n59319) );
  INVx3_ASAP7_75t_SL U52028 ( .A(n77566), .Y(n57093) );
  NAND2xp33_ASAP7_75t_SL U52029 ( .A(or1200_cpu_rf_datab[7]), .B(n57091), .Y(
        n76812) );
  INVx1_ASAP7_75t_SL U52030 ( .A(n78009), .Y(n57092) );
  INVx5_ASAP7_75t_SL U52031 ( .A(n77456), .Y(n57090) );
  NAND2xp33_ASAP7_75t_SL U52032 ( .A(or1200_cpu_rf_datab[2]), .B(n57091), .Y(
        n61266) );
  NAND2xp33_ASAP7_75t_SL U52033 ( .A(or1200_cpu_rf_datab[0]), .B(n57091), .Y(
        n61020) );
  INVxp33_ASAP7_75t_SL U52034 ( .A(n68025), .Y(n67997) );
  INVxp67_ASAP7_75t_SL U52035 ( .A(n71051), .Y(n71035) );
  NOR2xp33_ASAP7_75t_SL U52036 ( .A(n63050), .B(n63051), .Y(n58184) );
  NOR2xp67_ASAP7_75t_SL U52037 ( .A(n63368), .B(n63367), .Y(n62947) );
  O2A1O1Ixp5_ASAP7_75t_SL U52038 ( .A1(n2009), .A2(n65402), .B(n65287), .C(
        n65286), .Y(n65288) );
  BUFx2_ASAP7_75t_SL U52039 ( .A(n77185), .Y(n57091) );
  OAI21xp33_ASAP7_75t_SL U52040 ( .A1(n59671), .A2(n69186), .B(n69185), .Y(
        or1200_cpu_or1200_mult_mac_n1608) );
  INVx5_ASAP7_75t_SL U52041 ( .A(n77566), .Y(n57072) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U52042 ( .A1(n62491), .A2(n75648), .B(n62492), .C(
        n62489), .Y(n62490) );
  OAI21xp33_ASAP7_75t_SL U52043 ( .A1(n66739), .A2(n66737), .B(n66691), .Y(
        n66695) );
  AOI21xp33_ASAP7_75t_SRAM U52044 ( .A1(n74312), .A2(n74311), .B(n74416), .Y(
        n74419) );
  INVx2_ASAP7_75t_SL U52045 ( .A(n58399), .Y(n57142) );
  OAI21xp33_ASAP7_75t_SL U52046 ( .A1(n63003), .A2(n63002), .B(n59226), .Y(
        n59225) );
  XNOR2xp5_ASAP7_75t_SL U52047 ( .A(n63152), .B(n63151), .Y(n63167) );
  NAND2xp33_ASAP7_75t_SL U52048 ( .A(n77381), .B(n59691), .Y(n77553) );
  INVx1_ASAP7_75t_SL U52049 ( .A(n67575), .Y(n67526) );
  OAI21xp5_ASAP7_75t_SL U52050 ( .A1(n64274), .A2(n64273), .B(n64272), .Y(
        n76305) );
  INVx3_ASAP7_75t_SL U52051 ( .A(n57144), .Y(n59693) );
  INVx2_ASAP7_75t_SL U52052 ( .A(n57144), .Y(n59694) );
  NAND2xp33_ASAP7_75t_SRAM U52053 ( .A(n65344), .B(n65343), .Y(n1634) );
  NOR2xp33_ASAP7_75t_SL U52054 ( .A(n66553), .B(n66575), .Y(n66576) );
  INVxp67_ASAP7_75t_SL U52055 ( .A(n70834), .Y(n70820) );
  AOI21xp33_ASAP7_75t_SL U52056 ( .A1(n75213), .A2(
        or1200_cpu_or1200_except_n546), .B(n76791), .Y(n75259) );
  INVxp67_ASAP7_75t_SL U52057 ( .A(n61322), .Y(n62464) );
  NAND2x1p5_ASAP7_75t_SL U52058 ( .A(n62729), .B(n62730), .Y(n63058) );
  INVx4_ASAP7_75t_SL U52059 ( .A(n59695), .Y(n59691) );
  INVx1_ASAP7_75t_SL U52060 ( .A(n70969), .Y(n70922) );
  INVx5_ASAP7_75t_SL U52061 ( .A(n57144), .Y(n57073) );
  OAI21xp33_ASAP7_75t_SL U52062 ( .A1(n64321), .A2(n64145), .B(n64144), .Y(
        n64153) );
  INVx5_ASAP7_75t_SL U52063 ( .A(n59695), .Y(n57074) );
  NOR2xp33_ASAP7_75t_SL U52064 ( .A(n71113), .B(n71112), .Y(n71132) );
  NOR2xp33_ASAP7_75t_SL U52065 ( .A(n64469), .B(n64468), .Y(n64472) );
  NOR2xp33_ASAP7_75t_SL U52066 ( .A(or1200_cpu_or1200_except_n544), .B(n75884), 
        .Y(n75883) );
  INVxp67_ASAP7_75t_SL U52067 ( .A(n70971), .Y(n70960) );
  AOI21xp33_ASAP7_75t_SL U52068 ( .A1(n77662), .A2(n77128), .B(n64797), .Y(
        n64798) );
  AOI21xp5_ASAP7_75t_SL U52069 ( .A1(n70861), .A2(n70860), .B(n70859), .Y(
        n70872) );
  INVxp67_ASAP7_75t_SL U52070 ( .A(n68607), .Y(n68597) );
  INVx1_ASAP7_75t_SL U52071 ( .A(n66407), .Y(n66362) );
  INVxp67_ASAP7_75t_SL U52072 ( .A(n70919), .Y(n70920) );
  INVxp67_ASAP7_75t_SL U52073 ( .A(n61294), .Y(n61290) );
  NOR2xp33_ASAP7_75t_SL U52074 ( .A(n58003), .B(n67063), .Y(n67152) );
  INVxp67_ASAP7_75t_SL U52075 ( .A(n71271), .Y(n71182) );
  NOR2xp33_ASAP7_75t_SL U52076 ( .A(n66569), .B(n68605), .Y(n68607) );
  INVxp67_ASAP7_75t_SL U52077 ( .A(n67592), .Y(n57676) );
  OAI21xp33_ASAP7_75t_SL U52078 ( .A1(n57190), .A2(n72856), .B(n72854), .Y(
        n1968) );
  INVxp67_ASAP7_75t_SL U52079 ( .A(n70816), .Y(n70805) );
  NOR2x1_ASAP7_75t_SL U52080 ( .A(n59637), .B(n67298), .Y(n75467) );
  INVxp33_ASAP7_75t_SL U52081 ( .A(n78076), .Y(n78075) );
  AOI21xp33_ASAP7_75t_SRAM U52082 ( .A1(n76503), .A2(n76502), .B(n76501), .Y(
        n76504) );
  NAND2xp33_ASAP7_75t_SL U52083 ( .A(n66364), .B(n66482), .Y(n66295) );
  NOR2xp33_ASAP7_75t_SL U52084 ( .A(n60059), .B(n64259), .Y(n78252) );
  NOR2x1_ASAP7_75t_SL U52085 ( .A(n59012), .B(n58473), .Y(n57734) );
  AOI21xp33_ASAP7_75t_SL U52086 ( .A1(n71357), .A2(n71365), .B(n71319), .Y(
        n71322) );
  INVxp67_ASAP7_75t_SL U52087 ( .A(n57687), .Y(n57686) );
  OAI22xp33_ASAP7_75t_SL U52088 ( .A1(or1200_cpu_or1200_except_n670), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n550), .B2(n77032), .Y(n61841)
         );
  AOI22xp33_ASAP7_75t_SL U52089 ( .A1(n57126), .A2(n61552), .B1(n62292), .B2(
        n73933), .Y(n61563) );
  NOR2xp33_ASAP7_75t_SL U52090 ( .A(n56983), .B(n66353), .Y(n66467) );
  AOI21xp33_ASAP7_75t_SRAM U52091 ( .A1(n74340), .A2(n74339), .B(n74350), .Y(
        n74352) );
  NAND2xp5_ASAP7_75t_SL U52092 ( .A(n77451), .B(n57160), .Y(n60301) );
  INVxp67_ASAP7_75t_SL U52093 ( .A(n62940), .Y(n62977) );
  OAI21xp33_ASAP7_75t_SL U52094 ( .A1(n59526), .A2(n71212), .B(n71177), .Y(
        n71183) );
  INVxp67_ASAP7_75t_SL U52095 ( .A(n61917), .Y(n60785) );
  NAND2xp5_ASAP7_75t_SL U52096 ( .A(n75947), .B(n75953), .Y(n75951) );
  NAND2xp33_ASAP7_75t_SL U52097 ( .A(n71396), .B(n71117), .Y(n71093) );
  OAI22xp33_ASAP7_75t_SL U52098 ( .A1(or1200_cpu_or1200_except_n206), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n168), .B2(n57102), .Y(n61339)
         );
  OAI21xp33_ASAP7_75t_SL U52099 ( .A1(n57284), .A2(n57109), .B(n63223), .Y(
        n63613) );
  A2O1A1Ixp33_ASAP7_75t_SL U52100 ( .A1(n70028), .A2(n70149), .B(n58583), .C(
        n69848), .Y(n52523) );
  NAND2xp33_ASAP7_75t_SL U52101 ( .A(n67944), .B(n64401), .Y(n64333) );
  NAND2xp5_ASAP7_75t_SL U52102 ( .A(n66054), .B(n66057), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n50) );
  OAI22xp33_ASAP7_75t_SL U52103 ( .A1(or1200_cpu_or1200_except_n210), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n164), .B2(n57102), .Y(n61694)
         );
  OAI22xp33_ASAP7_75t_SL U52104 ( .A1(or1200_cpu_or1200_except_n208), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n166), .B2(n57102), .Y(n61759)
         );
  OAI22xp33_ASAP7_75t_SL U52105 ( .A1(or1200_cpu_or1200_except_n200), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n174), .B2(n57102), .Y(n62247)
         );
  OAI22xp33_ASAP7_75t_SL U52106 ( .A1(or1200_cpu_or1200_except_n202), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n172), .B2(n57102), .Y(n76740)
         );
  INVx3_ASAP7_75t_SL U52107 ( .A(n58554), .Y(n59675) );
  OAI22xp33_ASAP7_75t_SL U52108 ( .A1(or1200_cpu_or1200_except_n216), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n158), .B2(n57102), .Y(n60831)
         );
  NOR2xp33_ASAP7_75t_SL U52109 ( .A(n57284), .B(n59230), .Y(n63822) );
  OAI22xp33_ASAP7_75t_SL U52110 ( .A1(or1200_cpu_or1200_except_n198), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n176), .B2(n57102), .Y(n61615)
         );
  OAI21xp33_ASAP7_75t_SL U52111 ( .A1(n67944), .A2(n57178), .B(n62633), .Y(
        n62940) );
  NOR2xp33_ASAP7_75t_SL U52112 ( .A(n57356), .B(n64083), .Y(n62709) );
  OAI22xp33_ASAP7_75t_SL U52113 ( .A1(n1489), .A2(n74916), .B1(n59543), .B2(
        n74934), .Y(n74811) );
  OAI22xp33_ASAP7_75t_SL U52114 ( .A1(n71149), .A2(n71019), .B1(n71362), .B2(
        n70867), .Y(n70868) );
  OAI22xp33_ASAP7_75t_SL U52115 ( .A1(n71365), .A2(n71364), .B1(n71363), .B2(
        n71362), .Y(n71366) );
  AOI31xp33_ASAP7_75t_SL U52116 ( .A1(n58576), .A2(n66049), .A3(n65993), .B(
        n65879), .Y(n65885) );
  OAI22xp33_ASAP7_75t_SL U52117 ( .A1(or1200_cpu_or1200_except_n220), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n154), .B2(n57102), .Y(n62502)
         );
  INVx5_ASAP7_75t_SL U52118 ( .A(n58401), .Y(n57160) );
  INVxp67_ASAP7_75t_SL U52119 ( .A(n75260), .Y(n75263) );
  AOI21xp33_ASAP7_75t_SL U52120 ( .A1(n57126), .A2(n75251), .B(n75214), .Y(
        n75879) );
  OAI22xp33_ASAP7_75t_SL U52121 ( .A1(or1200_cpu_or1200_except_n196), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n178), .B2(n57102), .Y(n61393)
         );
  OAI22xp33_ASAP7_75t_SL U52122 ( .A1(or1200_cpu_or1200_except_n192), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n182), .B2(n57102), .Y(n61259)
         );
  OAI22xp33_ASAP7_75t_SL U52123 ( .A1(or1200_cpu_or1200_except_n244), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n130), .B2(n57102), .Y(n75816)
         );
  NAND2xp5_ASAP7_75t_SL U52124 ( .A(n57100), .B(n60080), .Y(n4112) );
  OAI22xp33_ASAP7_75t_SL U52125 ( .A1(or1200_cpu_or1200_except_n186), .A2(
        n57102), .B1(or1200_cpu_or1200_except_n188), .B2(n57170), .Y(n60581)
         );
  OAI22xp33_ASAP7_75t_SL U52126 ( .A1(or1200_cpu_or1200_except_n218), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n156), .B2(n57102), .Y(n77053)
         );
  INVxp67_ASAP7_75t_SL U52127 ( .A(n67021), .Y(n67022) );
  OAI22xp33_ASAP7_75t_SL U52128 ( .A1(or1200_cpu_or1200_except_n184), .A2(
        n57102), .B1(or1200_cpu_epcr_1_), .B2(n57170), .Y(n60907) );
  OAI22xp33_ASAP7_75t_SL U52129 ( .A1(or1200_cpu_or1200_except_n204), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n170), .B2(n57102), .Y(n62330)
         );
  INVx3_ASAP7_75t_SL U52130 ( .A(n77269), .Y(n57100) );
  AOI22xp33_ASAP7_75t_SL U52131 ( .A1(n70078), .A2(n69507), .B1(n69512), .B2(
        n69459), .Y(n69517) );
  BUFx3_ASAP7_75t_SL U52132 ( .A(n76172), .Y(n57336) );
  AOI22xp33_ASAP7_75t_SL U52133 ( .A1(n71396), .A2(n70954), .B1(n71394), .B2(
        n70909), .Y(n70917) );
  AOI22xp33_ASAP7_75t_SL U52134 ( .A1(n71209), .A2(n70951), .B1(n59522), .B2(
        n71282), .Y(n70952) );
  INVx3_ASAP7_75t_SL U52135 ( .A(n58416), .Y(n57170) );
  INVx1_ASAP7_75t_SL U52136 ( .A(n74492), .Y(n57103) );
  INVxp67_ASAP7_75t_SL U52137 ( .A(n74224), .Y(n74225) );
  AND2x2_ASAP7_75t_SL U52138 ( .A(n57111), .B(n66332), .Y(n57585) );
  NAND2xp5_ASAP7_75t_SL U52139 ( .A(n63545), .B(n63544), .Y(n63550) );
  NAND2xp33_ASAP7_75t_SL U52140 ( .A(n64181), .B(n64180), .Y(n64182) );
  NOR2xp33_ASAP7_75t_SRAM U52141 ( .A(n78327), .B(n76484), .Y(n76485) );
  AOI22xp33_ASAP7_75t_SL U52142 ( .A1(n70777), .A2(n70725), .B1(n70724), .B2(
        n70931), .Y(n70711) );
  NAND2xp33_ASAP7_75t_SL U52143 ( .A(n65990), .B(n66052), .Y(n65892) );
  INVxp33_ASAP7_75t_SRAM U52144 ( .A(n65250), .Y(n65251) );
  INVxp33_ASAP7_75t_SL U52145 ( .A(n73363), .Y(n73364) );
  AOI21xp33_ASAP7_75t_SL U52146 ( .A1(n73933), .A2(n75876), .B(n73932), .Y(
        n73934) );
  NOR2x1_ASAP7_75t_SL U52147 ( .A(n57111), .B(n75032), .Y(n68133) );
  INVxp67_ASAP7_75t_SL U52148 ( .A(n73279), .Y(n73287) );
  INVx1_ASAP7_75t_SL U52149 ( .A(n66344), .Y(n66372) );
  INVx1_ASAP7_75t_SL U52150 ( .A(n71160), .Y(n71142) );
  INVxp33_ASAP7_75t_SL U52151 ( .A(n71194), .Y(n71045) );
  NAND2x1_ASAP7_75t_SL U52152 ( .A(n66332), .B(n66373), .Y(n67743) );
  NAND2xp33_ASAP7_75t_SL U52153 ( .A(n73363), .B(n73366), .Y(n73317) );
  INVx2_ASAP7_75t_SL U52154 ( .A(n77052), .Y(n57102) );
  OAI21xp33_ASAP7_75t_SL U52155 ( .A1(n61638), .A2(n61637), .B(n61636), .Y(
        n61641) );
  INVxp67_ASAP7_75t_SL U52156 ( .A(n71044), .Y(n71001) );
  NOR2x1_ASAP7_75t_SL U52157 ( .A(n72594), .B(n74276), .Y(n74493) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U52158 ( .A1(n61768), .A2(n62372), .B(n57126), .C(
        n61767), .Y(n61769) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U52159 ( .A1(n73308), .A2(n74502), .B(n73307), 
        .C(n73312), .Y(n73313) );
  OAI21xp5_ASAP7_75t_SL U52160 ( .A1(n71077), .A2(n71076), .B(n71075), .Y(
        n71193) );
  AOI21xp5_ASAP7_75t_SL U52161 ( .A1(n75584), .A2(n75717), .B(n64300), .Y(
        n64312) );
  NAND2xp5_ASAP7_75t_SL U52162 ( .A(n77850), .B(n76735), .Y(n74934) );
  INVxp67_ASAP7_75t_SL U52163 ( .A(n71329), .Y(n71330) );
  INVx1_ASAP7_75t_SL U52164 ( .A(n70882), .Y(n70951) );
  OAI21xp33_ASAP7_75t_SL U52165 ( .A1(n59671), .A2(n65152), .B(n65151), .Y(
        n65153) );
  OAI21xp5_ASAP7_75t_SL U52166 ( .A1(n71281), .A2(n71162), .B(n71161), .Y(
        n71339) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U52167 ( .A1(n71591), .A2(n71590), .B(n71589), .C(
        n71635), .Y(n71592) );
  OAI21xp33_ASAP7_75t_SL U52168 ( .A1(n65872), .A2(n66027), .B(n65968), .Y(
        n65867) );
  INVxp67_ASAP7_75t_SL U52169 ( .A(n71285), .Y(n71243) );
  INVx1_ASAP7_75t_SL U52170 ( .A(n70867), .Y(n70897) );
  INVx3_ASAP7_75t_SL U52171 ( .A(n58600), .Y(n57105) );
  NAND2xp5_ASAP7_75t_SL U52172 ( .A(n62883), .B(n57180), .Y(n62882) );
  INVxp33_ASAP7_75t_SL U52173 ( .A(n66029), .Y(n66030) );
  OAI21xp5_ASAP7_75t_SL U52174 ( .A1(n71076), .A2(n70788), .B(n70787), .Y(
        n70954) );
  INVx6_ASAP7_75t_SL U52175 ( .A(n58440), .Y(n57180) );
  INVxp67_ASAP7_75t_SL U52176 ( .A(n71311), .Y(n71312) );
  AOI22xp5_ASAP7_75t_SL U52177 ( .A1(n73024), .A2(n72966), .B1(n73030), .B2(
        n72965), .Y(n72729) );
  AOI22xp5_ASAP7_75t_SL U52178 ( .A1(n57198), .A2(n62156), .B1(n77920), .B2(
        n77212), .Y(n60232) );
  AOI22xp33_ASAP7_75t_SL U52179 ( .A1(n71087), .A2(n71138), .B1(n70996), .B2(
        n71192), .Y(n71044) );
  INVxp33_ASAP7_75t_SL U52180 ( .A(n78160), .Y(n78159) );
  NAND2xp33_ASAP7_75t_SL U52181 ( .A(n66051), .B(n65955), .Y(n66029) );
  AOI22xp33_ASAP7_75t_SL U52182 ( .A1(n72993), .A2(n72935), .B1(n73030), .B2(
        n72787), .Y(n72791) );
  OAI21xp33_ASAP7_75t_SL U52183 ( .A1(n74196), .A2(n74183), .B(n74182), .Y(
        n74184) );
  INVx3_ASAP7_75t_SL U52184 ( .A(n59503), .Y(n57178) );
  OAI21xp33_ASAP7_75t_SL U52185 ( .A1(n59671), .A2(n68770), .B(n68769), .Y(
        n68771) );
  AOI22xp33_ASAP7_75t_SL U52186 ( .A1(n71209), .A2(n71192), .B1(n71245), .B2(
        n71244), .Y(n71329) );
  OAI21xp33_ASAP7_75t_SL U52187 ( .A1(n1438), .A2(n57114), .B(n74040), .Y(
        n9283) );
  NAND2xp33_ASAP7_75t_SRAM U52188 ( .A(n57128), .B(n62445), .Y(n62446) );
  OAI21xp33_ASAP7_75t_SL U52189 ( .A1(n1450), .A2(n57114), .B(n74980), .Y(
        n9289) );
  OAI21xp33_ASAP7_75t_SL U52190 ( .A1(n1452), .A2(n57114), .B(n75296), .Y(
        n9290) );
  AOI21xp5_ASAP7_75t_SL U52191 ( .A1(n75584), .A2(n77062), .B(n61712), .Y(
        n61713) );
  NAND2xp33_ASAP7_75t_SL U52192 ( .A(n59522), .B(n71138), .Y(n70787) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U52193 ( .A1(n62279), .A2(n62278), .B(n62277), 
        .C(n57126), .Y(n62280) );
  NAND2x1_ASAP7_75t_SL U52194 ( .A(n63246), .B(n63247), .Y(n76633) );
  AOI22xp33_ASAP7_75t_SL U52195 ( .A1(n59522), .A2(n71171), .B1(n71087), .B2(
        n71172), .Y(n70894) );
  BUFx3_ASAP7_75t_SL U52196 ( .A(n76091), .Y(n57310) );
  NAND2xp33_ASAP7_75t_SL U52197 ( .A(n59522), .B(n71244), .Y(n70912) );
  NAND2xp33_ASAP7_75t_SL U52198 ( .A(n66022), .B(n65707), .Y(n65708) );
  AND2x2_ASAP7_75t_SL U52199 ( .A(n63248), .B(n63247), .Y(n58600) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U52200 ( .A1(n77076), .A2(n77075), .B(n77074), 
        .C(n57126), .Y(n77077) );
  OAI211xp5_ASAP7_75t_SRAM U52201 ( .A1(n62353), .A2(n75329), .B(n61355), .C(
        n61354), .Y(n61356) );
  OAI22xp33_ASAP7_75t_SL U52202 ( .A1(n66027), .A2(n65902), .B1(n65929), .B2(
        n65972), .Y(n65903) );
  NAND2x1p5_ASAP7_75t_SL U52203 ( .A(n66375), .B(n66376), .Y(n76172) );
  OAI22xp33_ASAP7_75t_SRAM U52204 ( .A1(n65897), .A2(n66027), .B1(n65972), 
        .B2(n65937), .Y(n65898) );
  AOI22xp33_ASAP7_75t_SL U52205 ( .A1(n71209), .A2(n71074), .B1(n71245), .B2(
        n71138), .Y(n71075) );
  OAI22xp33_ASAP7_75t_SL U52206 ( .A1(n57115), .A2(n70776), .B1(n70767), .B2(
        n70993), .Y(n71040) );
  NOR2xp33_ASAP7_75t_SL U52207 ( .A(or1200_cpu_or1200_except_n498), .B(n76724), 
        .Y(n61603) );
  NAND2xp5_ASAP7_75t_SL U52208 ( .A(n75392), .B(n75387), .Y(n66225) );
  OAI22xp5_ASAP7_75t_SL U52209 ( .A1(n57115), .A2(n70863), .B1(n70850), .B2(
        n70993), .Y(n71192) );
  NAND2xp33_ASAP7_75t_SL U52210 ( .A(n77862), .B(n57114), .Y(n75407) );
  INVxp67_ASAP7_75t_SL U52211 ( .A(n75387), .Y(n75645) );
  INVx3_ASAP7_75t_SL U52212 ( .A(n59672), .Y(n59671) );
  AOI21xp33_ASAP7_75t_SRAM U52213 ( .A1(n76941), .A2(n74887), .B(n76963), .Y(
        n74888) );
  INVxp33_ASAP7_75t_SL U52214 ( .A(n66063), .Y(n65753) );
  OAI21xp5_ASAP7_75t_SL U52215 ( .A1(n64121), .A2(n77749), .B(n61402), .Y(
        n61403) );
  OAI22xp33_ASAP7_75t_SL U52216 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_14_), .A2(n69497), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_15_), .B2(n69496), .Y(
        n69498) );
  INVx1_ASAP7_75t_SL U52217 ( .A(n77107), .Y(n61785) );
  AOI21xp5_ASAP7_75t_SL U52218 ( .A1(n73998), .A2(n61929), .B(n61928), .Y(
        n63545) );
  AOI21xp5_ASAP7_75t_SL U52219 ( .A1(n78359), .A2(n72667), .B(n72656), .Y(
        n72669) );
  OAI21xp33_ASAP7_75t_SRAM U52220 ( .A1(n78429), .A2(n69563), .B(n70078), .Y(
        n69566) );
  INVx4_ASAP7_75t_SL U52221 ( .A(n76631), .Y(n57077) );
  OAI22xp5_ASAP7_75t_SL U52222 ( .A1(n70995), .A2(n57115), .B1(n70994), .B2(
        n59524), .Y(n71331) );
  OAI22xp5_ASAP7_75t_SL U52223 ( .A1(n57115), .A2(n70809), .B1(n70786), .B2(
        n70993), .Y(n71138) );
  OAI22xp5_ASAP7_75t_SL U52224 ( .A1(n57115), .A2(n70983), .B1(n70950), .B2(
        n59524), .Y(n71282) );
  BUFx3_ASAP7_75t_SL U52225 ( .A(n68016), .Y(n59507) );
  NAND2xp5_ASAP7_75t_SL U52226 ( .A(n61750), .B(n61749), .Y(n61751) );
  OAI22xp33_ASAP7_75t_SL U52227 ( .A1(n57115), .A2(n70994), .B1(n70983), .B2(
        n70993), .Y(n71311) );
  OAI22xp33_ASAP7_75t_SL U52228 ( .A1(n75330), .A2(n77103), .B1(n61639), .B2(
        n75587), .Y(n61107) );
  NOR2xp33_ASAP7_75t_SL U52229 ( .A(n62762), .B(n61936), .Y(n76263) );
  OAI21xp5_ASAP7_75t_SL U52230 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[13]), .A2(n58582), 
        .B(n65820), .Y(n66011) );
  AOI22xp33_ASAP7_75t_SL U52231 ( .A1(n66022), .A2(n65887), .B1(n65886), .B2(
        n66051), .Y(n65888) );
  O2A1O1Ixp5_ASAP7_75t_SL U52232 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]), .A2(n65646), 
        .B(n65645), .C(n66160), .Y(n65647) );
  INVxp33_ASAP7_75t_SRAM U52233 ( .A(n65466), .Y(n65467) );
  NAND2xp33_ASAP7_75t_SL U52234 ( .A(n77890), .B(n57114), .Y(n75403) );
  NAND2xp33_ASAP7_75t_SL U52235 ( .A(n77880), .B(n57114), .Y(n64184) );
  NAND2xp33_ASAP7_75t_SL U52236 ( .A(n77873), .B(n57114), .Y(n75404) );
  NAND2xp33_ASAP7_75t_SL U52237 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[10]), .B(
        n59631), .Y(n73160) );
  INVxp67_ASAP7_75t_SL U52238 ( .A(n65958), .Y(n65902) );
  NAND2xp33_ASAP7_75t_SL U52239 ( .A(n77864), .B(n57114), .Y(n75402) );
  NAND2xp33_ASAP7_75t_SL U52240 ( .A(n77866), .B(n57114), .Y(n66223) );
  NAND2xp33_ASAP7_75t_SL U52241 ( .A(n77869), .B(n57114), .Y(n74078) );
  OAI21xp5_ASAP7_75t_SL U52242 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]), .A2(n65500), .B(
        n76977), .Y(n65667) );
  BUFx2_ASAP7_75t_SL U52243 ( .A(n75408), .Y(n57114) );
  INVx2_ASAP7_75t_SL U52244 ( .A(n65974), .Y(n66051) );
  NOR2xp33_ASAP7_75t_SL U52245 ( .A(or1200_cpu_or1200_except_n520), .B(n77081), 
        .Y(n75313) );
  O2A1O1Ixp5_ASAP7_75t_SL U52246 ( .A1(n72169), .A2(n72170), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .C(
        n71903), .Y(n71904) );
  OAI21xp33_ASAP7_75t_SRAM U52247 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n74701), .B(n74700), .Y(n74705) );
  NAND2xp5_ASAP7_75t_SL U52248 ( .A(n70114), .B(n70109), .Y(n70021) );
  O2A1O1Ixp5_ASAP7_75t_SL U52249 ( .A1(n75701), .A2(n75866), .B(n75700), .C(
        n75699), .Y(n75733) );
  AOI21xp33_ASAP7_75t_SL U52250 ( .A1(n74293), .A2(n74292), .B(n74291), .Y(
        n74296) );
  OAI21xp33_ASAP7_75t_SL U52251 ( .A1(n57120), .A2(n57214), .B(n60749), .Y(
        n60759) );
  INVx4_ASAP7_75t_SL U52252 ( .A(n58284), .Y(n57185) );
  OR3x1_ASAP7_75t_SL U52253 ( .A(n60611), .B(n58655), .C(n60612), .Y(n58654)
         );
  INVx3_ASAP7_75t_SL U52254 ( .A(n59485), .Y(n57078) );
  NAND2xp5_ASAP7_75t_SL U52255 ( .A(n57126), .B(n75845), .Y(n75587) );
  INVxp33_ASAP7_75t_SL U52256 ( .A(n61518), .Y(n61520) );
  NAND2xp5_ASAP7_75t_SL U52257 ( .A(n57126), .B(n62374), .Y(n77107) );
  NAND2xp33_ASAP7_75t_SL U52258 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), .B(
        n72920), .Y(n72860) );
  OAI31xp33_ASAP7_75t_SRAM U52259 ( .A1(n1173), .A2(n61746), .A3(n62419), .B(
        n61471), .Y(n61473) );
  NAND2xp5_ASAP7_75t_SL U52260 ( .A(n57126), .B(n77076), .Y(n75574) );
  INVx2_ASAP7_75t_SL U52261 ( .A(n76897), .Y(n59672) );
  AOI22xp33_ASAP7_75t_SL U52262 ( .A1(n73379), .A2(n73119), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[21]), .B2(
        n73382), .Y(n73327) );
  NAND2xp5_ASAP7_75t_SL U52263 ( .A(n57126), .B(n61106), .Y(n77103) );
  INVx3_ASAP7_75t_SL U52264 ( .A(n76897), .Y(n57079) );
  INVx3_ASAP7_75t_SL U52265 ( .A(n76906), .Y(n57080) );
  OAI21xp5_ASAP7_75t_SL U52266 ( .A1(or1200_cpu_or1200_mult_mac_n106), .A2(
        n61826), .B(n61718), .Y(n61832) );
  NAND2xp33_ASAP7_75t_SL U52267 ( .A(n63897), .B(n64167), .Y(n63900) );
  OAI21xp5_ASAP7_75t_SL U52268 ( .A1(n70429), .A2(n70483), .B(n70352), .Y(
        n2344) );
  AOI22xp33_ASAP7_75t_SL U52269 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[39]), .A2(n57187), 
        .B1(n57188), .B2(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[38]), .Y(n65865) );
  NOR2xp33_ASAP7_75t_SL U52270 ( .A(n62254), .B(n61546), .Y(n58285) );
  NAND2xp33_ASAP7_75t_SL U52271 ( .A(n57126), .B(n75322), .Y(n62332) );
  OAI21xp33_ASAP7_75t_SL U52272 ( .A1(n72241), .A2(n72485), .B(n71806), .Y(
        n72305) );
  AND2x2_ASAP7_75t_SL U52273 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[1]), .B(n59628), 
        .Y(n72857) );
  OAI21xp33_ASAP7_75t_SL U52274 ( .A1(n59625), .A2(n72544), .B(n72381), .Y(
        n72172) );
  NAND2xp33_ASAP7_75t_SRAM U52275 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output1_23_), .B(n75625), .Y(n1511)
         );
  INVx1_ASAP7_75t_SL U52276 ( .A(n74255), .Y(n73882) );
  NAND2xp33_ASAP7_75t_SL U52277 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]), .B(n57188), 
        .Y(n65715) );
  INVx1_ASAP7_75t_SL U52278 ( .A(n58420), .Y(n76472) );
  OAI21xp33_ASAP7_75t_SL U52279 ( .A1(or1200_cpu_or1200_mult_mac_n341), .A2(
        n75738), .B(n73922), .Y(n73929) );
  INVxp67_ASAP7_75t_SL U52280 ( .A(n75350), .Y(n75247) );
  NAND2xp33_ASAP7_75t_SL U52281 ( .A(n58203), .B(n62639), .Y(n62642) );
  NAND2xp5_ASAP7_75t_SL U52282 ( .A(n65680), .B(n65827), .Y(n65974) );
  NOR2xp33_ASAP7_75t_SL U52283 ( .A(n57791), .B(n53455), .Y(n60778) );
  OAI21xp33_ASAP7_75t_SL U52284 ( .A1(n57120), .A2(n59443), .B(n60755), .Y(
        n60978) );
  INVx1_ASAP7_75t_SL U52285 ( .A(n66027), .Y(n65978) );
  OAI21xp5_ASAP7_75t_SL U52286 ( .A1(n59627), .A2(n78335), .B(n72831), .Y(
        n72920) );
  NAND2xp33_ASAP7_75t_SL U52287 ( .A(n59539), .B(n57120), .Y(n60734) );
  OAI22xp33_ASAP7_75t_SL U52288 ( .A1(or1200_cpu_or1200_mult_mac_n74), .A2(
        n77058), .B1(n59580), .B2(n75319), .Y(n73938) );
  AOI21xp33_ASAP7_75t_SL U52289 ( .A1(n73921), .A2(n73920), .B(n73919), .Y(
        n73922) );
  INVxp33_ASAP7_75t_SL U52290 ( .A(n71170), .Y(n71168) );
  INVxp33_ASAP7_75t_SL U52291 ( .A(n60142), .Y(n60108) );
  AOI21xp33_ASAP7_75t_SRAM U52292 ( .A1(n73921), .A2(n68814), .B(n61860), .Y(
        n61863) );
  OAI21xp33_ASAP7_75t_SRAM U52293 ( .A1(n1408), .A2(n61599), .B(n61598), .Y(
        n61600) );
  INVxp33_ASAP7_75t_SL U52294 ( .A(n60790), .Y(n60792) );
  NAND2x1_ASAP7_75t_SL U52295 ( .A(n57126), .B(n76753), .Y(n75738) );
  NAND2xp5_ASAP7_75t_SL U52296 ( .A(n57126), .B(n75245), .Y(n75737) );
  INVxp67_ASAP7_75t_SL U52297 ( .A(n69719), .Y(n69722) );
  NAND2xp33_ASAP7_75t_SL U52298 ( .A(n70340), .B(n70370), .Y(n70342) );
  NOR2xp33_ASAP7_75t_SL U52299 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_8_), .B(n65387), .Y(
        n65317) );
  NAND2xp5_ASAP7_75t_SL U52300 ( .A(n63453), .B(n57121), .Y(n61718) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U52301 ( .A1(n61873), .A2(n76768), .B(n62433), .C(
        n61872), .Y(n61874) );
  AOI22xp5_ASAP7_75t_SL U52302 ( .A1(n68789), .A2(n57121), .B1(n61827), .B2(
        n75218), .Y(n75223) );
  NAND2xp5_ASAP7_75t_SL U52303 ( .A(n65146), .B(n57121), .Y(n61819) );
  INVx1_ASAP7_75t_SL U52304 ( .A(n70092), .Y(n69717) );
  INVx4_ASAP7_75t_SL U52305 ( .A(n59629), .Y(n57190) );
  NAND2xp33_ASAP7_75t_SL U52306 ( .A(n69788), .B(n70515), .Y(n69800) );
  AOI22xp5_ASAP7_75t_SL U52307 ( .A1(n68791), .A2(n57121), .B1(n53430), .B2(
        n61815), .Y(n73944) );
  NAND2xp5_ASAP7_75t_SL U52308 ( .A(n65140), .B(n57121), .Y(n61817) );
  OAI21xp33_ASAP7_75t_SL U52309 ( .A1(n62582), .A2(n62556), .B(n57120), .Y(
        n60738) );
  NOR2xp67_ASAP7_75t_SL U52310 ( .A(n64209), .B(n63261), .Y(n77039) );
  AOI22xp33_ASAP7_75t_SL U52311 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[16]), .B2(n57194), .Y(n65839) );
  AOI22xp33_ASAP7_75t_SL U52312 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[18]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]), .B2(n57194), .Y(n65756) );
  NAND2xp5_ASAP7_75t_SL U52313 ( .A(n65078), .B(n57121), .Y(n61821) );
  OAI21xp5_ASAP7_75t_SL U52314 ( .A1(n71946), .A2(n72027), .B(n71860), .Y(
        n71861) );
  NAND2xp33_ASAP7_75t_SL U52315 ( .A(n74956), .B(n74955), .Y(n74958) );
  NAND2xp33_ASAP7_75t_SL U52316 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[10]), .B(n73047), .Y(n72765) );
  INVx4_ASAP7_75t_SL U52317 ( .A(n61828), .Y(n57121) );
  OAI21xp33_ASAP7_75t_SL U52318 ( .A1(n64289), .A2(n75735), .B(n64288), .Y(
        n64290) );
  NAND2xp33_ASAP7_75t_SL U52319 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_44_), .B(n71353), 
        .Y(n71358) );
  NAND2xp5_ASAP7_75t_SL U52320 ( .A(n72544), .B(n57192), .Y(n72278) );
  AOI21xp5_ASAP7_75t_SL U52321 ( .A1(n73781), .A2(n73752), .B(n73738), .Y(
        n73806) );
  INVxp67_ASAP7_75t_SL U52322 ( .A(n75226), .Y(n75230) );
  INVxp67_ASAP7_75t_SL U52323 ( .A(n63248), .Y(n63246) );
  OAI21xp33_ASAP7_75t_SRAM U52324 ( .A1(n72046), .A2(n72147), .B(n71814), .Y(
        n71821) );
  AOI21xp5_ASAP7_75t_SL U52325 ( .A1(n65081), .A2(n65083), .B(n65080), .Y(
        n65170) );
  OAI21xp33_ASAP7_75t_SL U52326 ( .A1(n69787), .A2(n70103), .B(n69616), .Y(
        n70515) );
  OAI21xp5_ASAP7_75t_SL U52327 ( .A1(n69411), .A2(n69446), .B(n69410), .Y(
        n70114) );
  INVxp33_ASAP7_75t_SL U52328 ( .A(n77996), .Y(n61296) );
  NOR2xp33_ASAP7_75t_SRAM U52329 ( .A(n59572), .B(n59584), .Y(n60788) );
  INVx1_ASAP7_75t_SL U52330 ( .A(n76821), .Y(n74956) );
  NOR2xp33_ASAP7_75t_SRAM U52331 ( .A(n59573), .B(n63571), .Y(n60638) );
  AOI22xp33_ASAP7_75t_SL U52332 ( .A1(n57198), .A2(n61567), .B1(n78005), .B2(
        n77253), .Y(n61568) );
  INVx5_ASAP7_75t_SL U52333 ( .A(n58599), .Y(n57192) );
  NAND3xp33_ASAP7_75t_SRAM U52334 ( .A(n74746), .B(n76976), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2), .Y(n66216) );
  INVxp67_ASAP7_75t_SL U52335 ( .A(n70405), .Y(n70427) );
  NAND2xp5_ASAP7_75t_SL U52336 ( .A(n74142), .B(n74143), .Y(n74146) );
  NOR2xp33_ASAP7_75t_SL U52337 ( .A(n61133), .B(n77622), .Y(n60819) );
  AOI21xp5_ASAP7_75t_SL U52338 ( .A1(n73704), .A2(n73752), .B(n73638), .Y(
        n73809) );
  AOI21xp33_ASAP7_75t_SL U52339 ( .A1(n63743), .A2(n77875), .B(n60055), .Y(
        n60056) );
  NOR2xp33_ASAP7_75t_SRAM U52340 ( .A(n59574), .B(n63571), .Y(n60956) );
  AOI22xp33_ASAP7_75t_SL U52341 ( .A1(n71478), .A2(n71477), .B1(n71476), .B2(
        n71475), .Y(n71479) );
  NAND2xp33_ASAP7_75t_SL U52342 ( .A(n62153), .B(n77850), .Y(n76663) );
  NAND2xp33_ASAP7_75t_SL U52343 ( .A(n57126), .B(n75853), .Y(n75723) );
  OAI21xp33_ASAP7_75t_SL U52344 ( .A1(n53311), .A2(n78182), .B(n75486), .Y(
        n77058) );
  OAI211xp5_ASAP7_75t_SRAM U52345 ( .A1(n76435), .A2(n76371), .B(n76370), .C(
        n76369), .Y(n76372) );
  NAND3xp33_ASAP7_75t_SRAM U52346 ( .A(n77996), .B(n77995), .C(n59696), .Y(
        n4306) );
  INVxp33_ASAP7_75t_SL U52347 ( .A(n70241), .Y(n70225) );
  AOI22xp33_ASAP7_75t_SL U52348 ( .A1(n72105), .A2(n72069), .B1(n72126), .B2(
        n72065), .Y(n71999) );
  NOR2xp33_ASAP7_75t_SRAM U52349 ( .A(n59531), .B(n57196), .Y(n61881) );
  NOR2xp33_ASAP7_75t_SRAM U52350 ( .A(n59577), .B(n63571), .Y(n60859) );
  AOI21xp33_ASAP7_75t_SL U52351 ( .A1(n70369), .A2(n74706), .B(n70330), .Y(
        n70548) );
  INVxp67_ASAP7_75t_SL U52352 ( .A(n72087), .Y(n71943) );
  NAND2xp5_ASAP7_75t_SL U52353 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_26_), .B(n70103), 
        .Y(n69718) );
  AOI21xp33_ASAP7_75t_SL U52354 ( .A1(n63743), .A2(n77888), .B(n60110), .Y(
        n60111) );
  OAI21xp33_ASAP7_75t_SL U52355 ( .A1(n76795), .A2(n76794), .B(n76793), .Y(
        n76798) );
  NAND2xp33_ASAP7_75t_SL U52356 ( .A(n77997), .B(n60198), .Y(n60294) );
  NOR2xp33_ASAP7_75t_SL U52357 ( .A(n53473), .B(n70708), .Y(n70695) );
  NOR2xp67_ASAP7_75t_SL U52358 ( .A(n59493), .B(n77965), .Y(n75453) );
  INVxp67_ASAP7_75t_SL U52359 ( .A(n72964), .Y(n72885) );
  INVxp33_ASAP7_75t_SL U52360 ( .A(n60502), .Y(n60492) );
  INVx1_ASAP7_75t_SL U52361 ( .A(n76404), .Y(n59167) );
  INVxp67_ASAP7_75t_SL U52362 ( .A(n78182), .Y(n75507) );
  OAI22xp33_ASAP7_75t_SL U52363 ( .A1(or1200_cpu_or1200_except_n228), .A2(
        n58547), .B1(n1626), .B2(n57124), .Y(n60150) );
  OAI22xp33_ASAP7_75t_SL U52364 ( .A1(n71993), .A2(n57123), .B1(n57203), .B2(
        n71984), .Y(n71986) );
  OAI22xp33_ASAP7_75t_SL U52365 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_), 
        .A2(n57123), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_), 
        .B2(n57203), .Y(n72178) );
  OAI21xp5_ASAP7_75t_SL U52366 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_), .A2(
        n70488), .B(n70265), .Y(n70266) );
  INVxp67_ASAP7_75t_SL U52367 ( .A(n66123), .Y(n65584) );
  OAI21xp33_ASAP7_75t_SL U52368 ( .A1(or1200_cpu_epcr_31_), .A2(n58547), .B(
        n60017), .Y(n59996) );
  NAND2xp5_ASAP7_75t_SL U52369 ( .A(n59493), .B(n77623), .Y(n62419) );
  OAI22xp33_ASAP7_75t_SL U52370 ( .A1(or1200_cpu_or1200_except_n238), .A2(
        n58547), .B1(n74079), .B2(n77254), .Y(n60178) );
  NAND2xp33_ASAP7_75t_SL U52371 ( .A(n57318), .B(n62569), .Y(n60628) );
  AOI22xp33_ASAP7_75t_SL U52372 ( .A1(or1200_cpu_or1200_fpu_result_arith[30]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[30]), 
        .Y(n75721) );
  OAI21xp5_ASAP7_75t_SL U52373 ( .A1(n60226), .A2(n62002), .B(n62476), .Y(
        n77850) );
  INVx1_ASAP7_75t_SL U52374 ( .A(n59587), .Y(n57197) );
  AOI21xp5_ASAP7_75t_SL U52375 ( .A1(n69204), .A2(n69203), .B(n69202), .Y(
        n69205) );
  OAI22xp33_ASAP7_75t_SL U52376 ( .A1(n72080), .A2(n57125), .B1(n57203), .B2(
        n72054), .Y(n72056) );
  NAND2xp5_ASAP7_75t_SL U52377 ( .A(n69522), .B(n78243), .Y(n69977) );
  OAI22xp33_ASAP7_75t_SL U52378 ( .A1(n72162), .A2(n57125), .B1(n57203), .B2(
        n72141), .Y(n72143) );
  INVx2_ASAP7_75t_SL U52379 ( .A(n73379), .Y(n74502) );
  NAND2xp5_ASAP7_75t_SL U52380 ( .A(n74043), .B(n75618), .Y(n78092) );
  NAND2xp5_ASAP7_75t_SL U52381 ( .A(n73381), .B(n59525), .Y(n73386) );
  INVx1_ASAP7_75t_SL U52382 ( .A(n76229), .Y(n59828) );
  INVx1_ASAP7_75t_SL U52383 ( .A(n63427), .Y(n63429) );
  INVx2_ASAP7_75t_SL U52384 ( .A(n72364), .Y(n57123) );
  OAI22xp33_ASAP7_75t_SL U52385 ( .A1(n71936), .A2(n57125), .B1(n71863), .B2(
        n57127), .Y(n71951) );
  OAI22xp33_ASAP7_75t_SL U52386 ( .A1(n71993), .A2(n57127), .B1(n57203), .B2(
        n71952), .Y(n71955) );
  OAI22xp33_ASAP7_75t_SL U52387 ( .A1(n72319), .A2(n57125), .B1(n57203), .B2(
        n72308), .Y(n72252) );
  NOR3xp33_ASAP7_75t_SRAM U52388 ( .A(n66196), .B(n66195), .C(n66194), .Y(
        n66200) );
  OAI22xp33_ASAP7_75t_SL U52389 ( .A1(n72163), .A2(n57125), .B1(n57203), .B2(
        n72154), .Y(n72156) );
  OAI22xp33_ASAP7_75t_SL U52390 ( .A1(n72263), .A2(n57125), .B1(n57203), .B2(
        n72262), .Y(n72265) );
  OR2x2_ASAP7_75t_SL U52391 ( .A(n76657), .B(n75475), .Y(n58547) );
  INVx1_ASAP7_75t_SL U52392 ( .A(n71362), .Y(n71396) );
  AOI21xp33_ASAP7_75t_SL U52393 ( .A1(n70675), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[22]), .B(n71281), 
        .Y(n70673) );
  INVxp67_ASAP7_75t_SL U52394 ( .A(n75849), .Y(n75850) );
  INVxp67_ASAP7_75t_SL U52395 ( .A(n76442), .Y(n76443) );
  NOR2xp33_ASAP7_75t_SL U52396 ( .A(n60855), .B(n60791), .Y(n61855) );
  NAND2xp5_ASAP7_75t_SL U52397 ( .A(n76976), .B(n65670), .Y(n65671) );
  INVx4_ASAP7_75t_SL U52398 ( .A(n77253), .Y(n57124) );
  NAND2xp5_ASAP7_75t_SL U52399 ( .A(n59541), .B(n61212), .Y(n57645) );
  AOI22xp33_ASAP7_75t_SL U52400 ( .A1(n57217), .A2(n73710), .B1(n3331), .B2(
        n57205), .Y(n73636) );
  AOI22xp33_ASAP7_75t_SL U52401 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_17_), 
        .A2(n57207), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_), 
        .B2(n71888), .Y(n71812) );
  INVxp67_ASAP7_75t_SL U52402 ( .A(n77871), .Y(n74045) );
  NAND2xp5_ASAP7_75t_SL U52403 ( .A(n59956), .B(n77210), .Y(n59494) );
  NAND2xp33_ASAP7_75t_SL U52404 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_14_), 
        .B(n57216), .Y(n71778) );
  NOR2xp33_ASAP7_75t_SRAM U52405 ( .A(n59546), .B(n57209), .Y(n74011) );
  INVxp67_ASAP7_75t_SL U52406 ( .A(n69066), .Y(n69071) );
  O2A1O1Ixp5_ASAP7_75t_SL U52407 ( .A1(or1200_cpu_or1200_mult_mac_n235), .A2(
        n69174), .B(n69173), .C(n69172), .Y(n69175) );
  INVxp33_ASAP7_75t_SRAM U52408 ( .A(n77410), .Y(n77411) );
  NAND2xp5_ASAP7_75t_SL U52409 ( .A(n68816), .B(n68815), .Y(n68819) );
  INVx1_ASAP7_75t_SL U52410 ( .A(n75866), .Y(n60635) );
  NAND2x1_ASAP7_75t_SL U52411 ( .A(n59526), .B(n71314), .Y(n71284) );
  OAI21x1_ASAP7_75t_SL U52412 ( .A1(dbg_stb_i), .A2(n77011), .B(n59929), .Y(
        n77623) );
  INVx3_ASAP7_75t_SL U52413 ( .A(n59625), .Y(n59624) );
  NAND2xp5_ASAP7_75t_SL U52414 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]), .B(n74206), .Y(
        n66181) );
  INVxp67_ASAP7_75t_SL U52415 ( .A(n74802), .Y(n74755) );
  INVxp67_ASAP7_75t_SL U52416 ( .A(n3143), .Y(n74828) );
  NAND2x1_ASAP7_75t_SL U52417 ( .A(n58315), .B(n71365), .Y(n71362) );
  INVxp67_ASAP7_75t_SL U52418 ( .A(n74742), .Y(n74743) );
  INVxp67_ASAP7_75t_SL U52419 ( .A(n59881), .Y(n60291) );
  INVx2_ASAP7_75t_SL U52420 ( .A(n71149), .Y(n71263) );
  A2O1A1Ixp33_ASAP7_75t_SL U52421 ( .A1(n62041), .A2(n78438), .B(n62040), .C(
        n62039), .Y(n62043) );
  NOR2xp33_ASAP7_75t_SL U52422 ( .A(n3105), .B(n61289), .Y(n60198) );
  INVxp67_ASAP7_75t_SL U52423 ( .A(n74282), .Y(n74283) );
  OAI21xp5_ASAP7_75t_SL U52424 ( .A1(n75196), .A2(n59867), .B(n59866), .Y(
        n59868) );
  OAI22xp33_ASAP7_75t_SRAM U52425 ( .A1(n73633), .A2(n58400), .B1(n73668), 
        .B2(n58622), .Y(n73634) );
  INVx3_ASAP7_75t_SL U52426 ( .A(n72347), .Y(n57127) );
  OAI21xp33_ASAP7_75t_SL U52427 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[11]), .A2(n71314), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_0_), .Y(n70654) );
  INVxp67_ASAP7_75t_SL U52428 ( .A(n74106), .Y(n74107) );
  INVxp67_ASAP7_75t_SL U52429 ( .A(n73901), .Y(n73902) );
  INVxp33_ASAP7_75t_SRAM U52430 ( .A(n4062), .Y(n61164) );
  INVxp67_ASAP7_75t_SRAM U52431 ( .A(n4058), .Y(n63729) );
  INVxp33_ASAP7_75t_SRAM U52432 ( .A(n4050), .Y(n61275) );
  INVxp67_ASAP7_75t_SL U52433 ( .A(n65225), .Y(n65209) );
  NAND2xp5_ASAP7_75t_SL U52434 ( .A(id_insn_22_), .B(n65218), .Y(n65224) );
  NAND2xp33_ASAP7_75t_SL U52435 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[5]), .B(
        n73221), .Y(n73049) );
  INVx3_ASAP7_75t_SL U52436 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .Y(
        n74706) );
  NAND2xp33_ASAP7_75t_SL U52437 ( .A(or1200_cpu_or1200_except_delayed_tee[1]), 
        .B(n78260), .Y(or1200_cpu_or1200_except_n1694) );
  INVxp33_ASAP7_75t_SRAM U52438 ( .A(n69532), .Y(n69534) );
  INVxp67_ASAP7_75t_SL U52439 ( .A(n59533), .Y(n63668) );
  INVx1_ASAP7_75t_SL U52440 ( .A(n59552), .Y(n57213) );
  INVx2_ASAP7_75t_SL U52441 ( .A(n59573), .Y(n75832) );
  NAND2xp33_ASAP7_75t_SL U52442 ( .A(n72990), .B(n73024), .Y(n72694) );
  INVx4_ASAP7_75t_SL U52443 ( .A(n59577), .Y(n57209) );
  NOR2x1_ASAP7_75t_SL U52444 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .B(
        n59527), .Y(n72347) );
  NAND2xp5_ASAP7_75t_SL U52445 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[3]), .B(
        n70579), .Y(n70581) );
  BUFx2_ASAP7_75t_SL U52446 ( .A(n1621), .Y(n57377) );
  INVx1_ASAP7_75t_SL U52447 ( .A(n59527), .Y(n72517) );
  NAND2xp5_ASAP7_75t_SL U52448 ( .A(n59526), .B(n58315), .Y(n71335) );
  INVx1_ASAP7_75t_SL U52449 ( .A(n71890), .Y(n71888) );
  NAND2x1_ASAP7_75t_SL U52450 ( .A(n1888), .B(n59561), .Y(n69355) );
  NAND2xp5_ASAP7_75t_SL U52451 ( .A(n59562), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]), .Y(n65629) );
  INVx2_ASAP7_75t_SL U52452 ( .A(n59562), .Y(n74206) );
  INVxp33_ASAP7_75t_SL U52453 ( .A(n73522), .Y(n73524) );
  INVx2_ASAP7_75t_SL U52454 ( .A(n59575), .Y(n57215) );
  NAND2xp5_ASAP7_75t_SL U52455 ( .A(n78401), .B(n59699), .Y(n71059) );
  INVxp67_ASAP7_75t_SL U52456 ( .A(n76942), .Y(n74878) );
  NOR2xp33_ASAP7_75t_SL U52457 ( .A(n2814), .B(n61028), .Y(n77427) );
  INVx5_ASAP7_75t_SL U52458 ( .A(ic_en), .Y(n77401) );
  AOI21xp33_ASAP7_75t_SL U52459 ( .A1(or1200_cpu_or1200_mult_mac_n357), .A2(
        or1200_cpu_or1200_mult_mac_n211), .B(n68882), .Y(n68883) );
  INVxp33_ASAP7_75t_SL U52460 ( .A(n68879), .Y(n68880) );
  BUFx2_ASAP7_75t_SL U52461 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[0]), .Y(n59562) );
  INVxp33_ASAP7_75t_SL U52462 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[26]), .Y(n73667) );
  INVx1_ASAP7_75t_SL U52463 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[32]), .Y(n65859) );
  INVx1_ASAP7_75t_SL U52464 ( .A(or1200_cpu_or1200_mult_mac_n309), .Y(n63453)
         );
  INVxp33_ASAP7_75t_SRAM U52465 ( .A(n1832), .Y(n61606) );
  INVxp67_ASAP7_75t_SL U52466 ( .A(or1200_cpu_or1200_genpc_pcreg_default[5]), 
        .Y(n77252) );
  INVxp33_ASAP7_75t_SL U52467 ( .A(or1200_cpu_or1200_mult_mac_n44), .Y(n76038)
         );
  INVxp33_ASAP7_75t_SL U52468 ( .A(n779), .Y(n60172) );
  INVxp33_ASAP7_75t_SRAM U52469 ( .A(n1169), .Y(n62230) );
  INVxp33_ASAP7_75t_SL U52470 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[14]), .Y(n65643) );
  INVxp67_ASAP7_75t_SL U52471 ( .A(n2071), .Y(n60416) );
  INVxp33_ASAP7_75t_SL U52472 ( .A(n2657), .Y(n61152) );
  INVx1_ASAP7_75t_SL U52473 ( .A(or1200_cpu_or1200_mult_mac_n32), .Y(n76085)
         );
  INVxp33_ASAP7_75t_SL U52474 ( .A(ex_insn[26]), .Y(n77522) );
  INVxp67_ASAP7_75t_SL U52475 ( .A(n803), .Y(n59983) );
  INVxp33_ASAP7_75t_SL U52476 ( .A(n2594), .Y(n77524) );
  INVxp67_ASAP7_75t_SL U52477 ( .A(or1200_cpu_or1200_except_n619), .Y(n63972)
         );
  INVxp33_ASAP7_75t_SL U52478 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_0_), .Y(n69377) );
  INVxp33_ASAP7_75t_SL U52479 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_1_), .Y(n74059) );
  INVxp67_ASAP7_75t_SL U52480 ( .A(or1200_cpu_or1200_mult_mac_n76), .Y(n64825)
         );
  INVxp33_ASAP7_75t_SRAM U52481 ( .A(n1129), .Y(n66235) );
  INVxp67_ASAP7_75t_SL U52482 ( .A(or1200_cpu_or1200_mult_mac_n74), .Y(n61815)
         );
  INVxp33_ASAP7_75t_SL U52483 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .Y(n65424) );
  NOR2xp33_ASAP7_75t_SL U52484 ( .A(or1200_cpu_or1200_except_n116), .B(
        or1200_cpu_or1200_except_n120), .Y(n76826) );
  INVxp67_ASAP7_75t_SL U52485 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[47]), .Y(n66089) );
  INVxp67_ASAP7_75t_SL U52486 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_4_), .Y(n65392) );
  INVxp67_ASAP7_75t_SL U52487 ( .A(or1200_cpu_or1200_mult_mac_n72), .Y(n75846)
         );
  INVxp67_ASAP7_75t_SL U52488 ( .A(or1200_cpu_or1200_except_n196), .Y(n61567)
         );
  INVx1_ASAP7_75t_SL U52489 ( .A(n759), .Y(n59987) );
  INVxp33_ASAP7_75t_SRAM U52490 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_14_), .Y(n65303) );
  INVx1_ASAP7_75t_SL U52491 ( .A(or1200_cpu_or1200_mult_mac_n337), .Y(n65160)
         );
  INVxp67_ASAP7_75t_SL U52492 ( .A(or1200_cpu_or1200_mult_mac_n339), .Y(n65159) );
  INVx1_ASAP7_75t_SL U52493 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[5]), .Y(n74367)
         );
  INVx1_ASAP7_75t_SL U52494 ( .A(or1200_cpu_or1200_mult_mac_n167), .Y(n63489)
         );
  INVx1_ASAP7_75t_SL U52495 ( .A(or1200_cpu_or1200_mult_mac_n243), .Y(n74573)
         );
  INVxp67_ASAP7_75t_SL U52496 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_10_), .Y(n65311) );
  INVx4_ASAP7_75t_SL U52497 ( .A(n59540), .Y(n57082) );
  INVxp33_ASAP7_75t_SL U52498 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_), 
        .Y(n72262) );
  INVx1_ASAP7_75t_SL U52499 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[14]), .Y(n74412)
         );
  NAND2xp33_ASAP7_75t_SL U52500 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_1_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_N398), .Y(n66180) );
  INVxp67_ASAP7_75t_SL U52501 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_), .Y(n78371) );
  INVxp33_ASAP7_75t_SL U52502 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_31_), .Y(n78328) );
  INVx6_ASAP7_75t_SL U52503 ( .A(n59706), .Y(n57083) );
  INVx1_ASAP7_75t_SL U52504 ( .A(or1200_cpu_or1200_mult_mac_n171), .Y(n77038)
         );
  INVxp67_ASAP7_75t_SL U52505 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_), 
        .Y(n72319) );
  INVx1_ASAP7_75t_SL U52506 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[13]), .Y(n74407)
         );
  INVx2_ASAP7_75t_SL U52507 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), .Y(
        n72990) );
  INVx1_ASAP7_75t_SL U52508 ( .A(or1200_cpu_or1200_mult_mac_n175), .Y(n75367)
         );
  INVxp67_ASAP7_75t_SL U52509 ( .A(or1200_cpu_or1200_except_n604), .Y(n76252)
         );
  INVx1_ASAP7_75t_SL U52510 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[17]), .Y(n74429)
         );
  INVxp67_ASAP7_75t_SL U52511 ( .A(or1200_cpu_or1200_except_n595), .Y(n76607)
         );
  INVxp67_ASAP7_75t_SL U52512 ( .A(or1200_cpu_or1200_except_n589), .Y(n76584)
         );
  INVxp33_ASAP7_75t_SL U52513 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_16_), .Y(n65301) );
  INVxp33_ASAP7_75t_SRAM U52514 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_17_), .Y(n74865)
         );
  INVx1_ASAP7_75t_SL U52515 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[19]), .Y(n74447)
         );
  INVx1_ASAP7_75t_SL U52516 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[20]), .Y(n74229)
         );
  INVxp67_ASAP7_75t_SL U52517 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .Y(
        n71873) );
  INVxp67_ASAP7_75t_SL U52518 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_11_), .Y(n76953)
         );
  INVxp67_ASAP7_75t_SL U52519 ( .A(or1200_cpu_or1200_except_n646), .Y(n75546)
         );
  INVx1_ASAP7_75t_SL U52520 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[18]), .Y(n74440)
         );
  INVxp67_ASAP7_75t_SL U52521 ( .A(or1200_cpu_or1200_except_n643), .Y(n64267)
         );
  INVx1_ASAP7_75t_SL U52522 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[21]), .Y(n74456)
         );
  INVxp33_ASAP7_75t_SL U52523 ( .A(or1200_cpu_or1200_mult_mac_n183), .Y(n65090) );
  INVxp67_ASAP7_75t_SL U52524 ( .A(or1200_cpu_or1200_except_n210), .Y(n74951)
         );
  INVx1_ASAP7_75t_SL U52525 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[16]), .Y(n74421)
         );
  INVxp33_ASAP7_75t_SL U52526 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[0]), .Y(
        n73868) );
  BUFx3_ASAP7_75t_SL U52527 ( .A(n2006), .Y(n59561) );
  INVxp33_ASAP7_75t_SL U52528 ( .A(or1200_cpu_or1200_mult_mac_n251), .Y(n75558) );
  BUFx5_ASAP7_75t_SL U52529 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_1_), .Y(n59526) );
  INVx1_ASAP7_75t_SL U52530 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[12]), .Y(n74398)
         );
  INVx1_ASAP7_75t_SL U52531 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_2_), .Y(n65238) );
  NAND2x1_ASAP7_75t_SL U52532 ( .A(n53473), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .Y(n71281) );
  INVx1_ASAP7_75t_SL U52533 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_state), .Y(n59697) );
  NAND2xp5_ASAP7_75t_SL U52534 ( .A(or1200_cpu_or1200_mult_mac_n311), .B(
        or1200_cpu_or1200_mult_mac_n165), .Y(n63488) );
  BUFx4f_ASAP7_75t_SL U52535 ( .A(n2856), .Y(n59573) );
  INVx1_ASAP7_75t_SL U52536 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[4]), .Y(n74382)
         );
  INVx1_ASAP7_75t_SL U52537 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[11]), .Y(n74389)
         );
  BUFx3_ASAP7_75t_SL U52538 ( .A(n2867), .Y(n59575) );
  INVxp33_ASAP7_75t_SL U52539 ( .A(or1200_cpu_or1200_mult_mac_n145), .Y(n61249) );
  INVxp33_ASAP7_75t_SRAM U52540 ( .A(or1200_cpu_or1200_except_n266), .Y(n61335) );
  INVxp67_ASAP7_75t_SL U52541 ( .A(n2759), .Y(n59947) );
  INVxp67_ASAP7_75t_SL U52542 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_14_), 
        .Y(n72311) );
  INVxp33_ASAP7_75t_SL U52543 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_27_), .Y(n78227) );
  INVxp33_ASAP7_75t_SL U52544 ( .A(supv), .Y(n76660) );
  INVx3_ASAP7_75t_SL U52545 ( .A(n59700), .Y(n57084) );
  NAND2xp5_ASAP7_75t_SL U52546 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_5_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_4_), .Y(n66207) );
  INVx1_ASAP7_75t_SL U52547 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[7]), .Y(n65823) );
  INVxp33_ASAP7_75t_SL U52548 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_3_), .Y(
        n72531) );
  NAND2xp5_ASAP7_75t_SL U52549 ( .A(dbg_stb_i), .B(dbg_we_i), .Y(n62476) );
  INVx1_ASAP7_75t_SL U52550 ( .A(or1200_ic_top_from_icram[28]), .Y(n60315) );
  INVx1_ASAP7_75t_SL U52551 ( .A(or1200_ic_top_from_icram[26]), .Y(n60323) );
  INVx1_ASAP7_75t_SL U52552 ( .A(or1200_ic_top_from_icram[29]), .Y(n60442) );
  INVx1_ASAP7_75t_SL U52553 ( .A(or1200_dc_top_tag_0_), .Y(n59809) );
  INVxp33_ASAP7_75t_SL U52554 ( .A(or1200_dc_top_dirty), .Y(n61994) );
  OAI21xp33_ASAP7_75t_SL U52555 ( .A1(n68709), .A2(n68714), .B(n68708), .Y(
        n68710) );
  OAI21xp33_ASAP7_75t_SL U52556 ( .A1(n69307), .A2(n59214), .B(n69306), .Y(
        n59213) );
  OAI21xp33_ASAP7_75t_SL U52557 ( .A1(n69155), .A2(n69154), .B(n69153), .Y(
        n69156) );
  AND2x2_ASAP7_75t_SL U52558 ( .A(n74558), .B(n58192), .Y(n58191) );
  INVx1_ASAP7_75t_SL U52559 ( .A(n68958), .Y(n68966) );
  NAND2xp33_ASAP7_75t_SL U52560 ( .A(n69045), .B(n69031), .Y(n69047) );
  INVxp33_ASAP7_75t_SL U52561 ( .A(n69151), .Y(n69122) );
  NAND2xp5_ASAP7_75t_SL U52562 ( .A(n68675), .B(n69295), .Y(n68676) );
  INVxp33_ASAP7_75t_SL U52563 ( .A(n69039), .Y(n69044) );
  INVx1_ASAP7_75t_SL U52564 ( .A(n68919), .Y(n57085) );
  NAND2xp33_ASAP7_75t_SL U52565 ( .A(n68669), .B(n69233), .Y(n68672) );
  NOR2x1_ASAP7_75t_SL U52566 ( .A(n58194), .B(n58193), .Y(n74558) );
  INVxp33_ASAP7_75t_SL U52567 ( .A(n69155), .Y(n69121) );
  NOR2xp33_ASAP7_75t_SL U52568 ( .A(n69032), .B(n69033), .Y(n69039) );
  NAND2xp5_ASAP7_75t_SL U52569 ( .A(n69101), .B(n69102), .Y(n58774) );
  OAI21xp5_ASAP7_75t_SL U52570 ( .A1(n77145), .A2(n77191), .B(n76511), .Y(
        or1200_cpu_or1200_except_n1743) );
  INVxp67_ASAP7_75t_SL U52571 ( .A(n65117), .Y(n65111) );
  NAND2xp5_ASAP7_75t_SL U52572 ( .A(n77192), .B(n77191), .Y(
        or1200_cpu_to_sr[9]) );
  INVxp33_ASAP7_75t_SL U52573 ( .A(n68908), .Y(n68865) );
  INVxp67_ASAP7_75t_SL U52574 ( .A(n59274), .Y(n57901) );
  INVx1_ASAP7_75t_SL U52575 ( .A(n68858), .Y(n68857) );
  INVx1_ASAP7_75t_SL U52576 ( .A(n69102), .Y(n58193) );
  OAI22xp33_ASAP7_75t_SL U52577 ( .A1(n59698), .A2(n71341), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_43_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n232) );
  INVxp67_ASAP7_75t_SL U52578 ( .A(n69040), .Y(n69041) );
  OAI22xp33_ASAP7_75t_SL U52579 ( .A1(n59699), .A2(n71125), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_30_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n193) );
  INVxp67_ASAP7_75t_SL U52580 ( .A(n57376), .Y(n69294) );
  INVx1_ASAP7_75t_SL U52581 ( .A(n67210), .Y(n69119) );
  OAI22xp33_ASAP7_75t_SL U52582 ( .A1(n59698), .A2(n71242), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_38_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n217) );
  NAND2xp33_ASAP7_75t_SL U52583 ( .A(n68685), .B(n68684), .Y(n68691) );
  INVxp67_ASAP7_75t_SL U52584 ( .A(n68709), .Y(n58192) );
  OAI22xp33_ASAP7_75t_SL U52585 ( .A1(n59699), .A2(n71227), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_37_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n214) );
  OAI22xp33_ASAP7_75t_SL U52586 ( .A1(n59698), .A2(n71199), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_35_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n208) );
  INVxp67_ASAP7_75t_SL U52587 ( .A(n68650), .Y(n68670) );
  OAI21xp33_ASAP7_75t_SL U52588 ( .A1(n57211), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_42_), .B(n71328), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n229) );
  INVx1_ASAP7_75t_SL U52589 ( .A(n68685), .Y(n57132) );
  INVx1_ASAP7_75t_SL U52590 ( .A(n68973), .Y(n57086) );
  OAI21xp33_ASAP7_75t_SL U52591 ( .A1(n59677), .A2(n77881), .B(n64157), .Y(
        n9619) );
  OAI21xp33_ASAP7_75t_SL U52592 ( .A1(n57211), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_36_), .B(n71216), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n211) );
  OAI21xp33_ASAP7_75t_SL U52593 ( .A1(n57144), .A2(n75639), .B(n58556), .Y(
        n2980) );
  OAI21xp33_ASAP7_75t_SL U52594 ( .A1(n57144), .A2(n77881), .B(n64155), .Y(
        n1629) );
  OAI22xp33_ASAP7_75t_SL U52595 ( .A1(n59698), .A2(n71361), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_44_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n235) );
  OAI22xp33_ASAP7_75t_SL U52596 ( .A1(n59699), .A2(n70964), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_21_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n166) );
  NOR2xp33_ASAP7_75t_SL U52597 ( .A(n64153), .B(n64152), .Y(n77881) );
  OAI21xp33_ASAP7_75t_SL U52598 ( .A1(n57211), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_23_), .B(n71011), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n172) );
  OAI21xp33_ASAP7_75t_SL U52599 ( .A1(n57211), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_40_), .B(n71280), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n223) );
  NAND2xp5_ASAP7_75t_SL U52600 ( .A(n69375), .B(n69374), .Y(
        or1200_cpu_or1200_except_n1704) );
  OAI21xp33_ASAP7_75t_SL U52601 ( .A1(n57211), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_41_), .B(n71310), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n226) );
  INVx1_ASAP7_75t_SL U52602 ( .A(n69293), .Y(n66602) );
  AOI21xp5_ASAP7_75t_SL U52603 ( .A1(n57135), .A2(n74578), .B(n74577), .Y(
        n74579) );
  AOI21xp5_ASAP7_75t_SL U52604 ( .A1(n57135), .A2(n75312), .B(n75303), .Y(
        n75304) );
  AOI21xp5_ASAP7_75t_SL U52605 ( .A1(n57135), .A2(n74986), .B(n74985), .Y(
        n74987) );
  AOI21xp5_ASAP7_75t_SL U52606 ( .A1(n57135), .A2(n75433), .B(n75432), .Y(
        n75434) );
  AOI21xp5_ASAP7_75t_SL U52607 ( .A1(n57135), .A2(n75622), .B(n75621), .Y(
        n75623) );
  NAND2xp33_ASAP7_75t_SL U52608 ( .A(n57211), .B(n71010), .Y(n71011) );
  NAND2xp5_ASAP7_75t_SL U52609 ( .A(n66609), .B(n66608), .Y(n68633) );
  AOI21xp33_ASAP7_75t_SL U52610 ( .A1(n57135), .A2(n76553), .B(n76552), .Y(
        n76554) );
  AOI21xp33_ASAP7_75t_SL U52611 ( .A1(n57135), .A2(n75783), .B(n75782), .Y(
        n75784) );
  OAI22xp33_ASAP7_75t_SL U52612 ( .A1(n59698), .A2(n71159), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_32_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n199) );
  OAI21xp33_ASAP7_75t_SL U52613 ( .A1(n57211), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_19_), .B(n70927), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n160) );
  OAI22xp33_ASAP7_75t_SL U52614 ( .A1(n59699), .A2(n70946), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_20_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n163) );
  AOI22xp33_ASAP7_75t_SL U52615 ( .A1(n76681), .A2(n57135), .B1(n77290), .B2(
        n76680), .Y(n76686) );
  NAND2xp33_ASAP7_75t_SL U52616 ( .A(n74986), .B(n76927), .Y(n74964) );
  NAND2xp33_ASAP7_75t_SL U52617 ( .A(n75433), .B(n76927), .Y(n75412) );
  NAND2xp33_ASAP7_75t_SL U52618 ( .A(n74047), .B(n76927), .Y(n65199) );
  NAND2xp33_ASAP7_75t_SL U52619 ( .A(n75622), .B(n76927), .Y(n75538) );
  NAND2xp33_ASAP7_75t_SL U52620 ( .A(n76253), .B(n76927), .Y(n76254) );
  AOI22xp33_ASAP7_75t_SL U52621 ( .A1(n76858), .A2(n77290), .B1(n57135), .B2(
        n76857), .Y(n76865) );
  NAND2xp33_ASAP7_75t_SL U52622 ( .A(n76681), .B(n76927), .Y(n76566) );
  INVxp67_ASAP7_75t_SL U52623 ( .A(n77795), .Y(n77801) );
  NAND2xp33_ASAP7_75t_SL U52624 ( .A(n76851), .B(n76927), .Y(n76646) );
  NAND2xp33_ASAP7_75t_SL U52625 ( .A(n77179), .B(n76927), .Y(n75168) );
  NAND2xp33_ASAP7_75t_SL U52626 ( .A(n74578), .B(n76927), .Y(n63923) );
  AOI22xp33_ASAP7_75t_SL U52627 ( .A1(n77291), .A2(n77290), .B1(n57135), .B2(
        n77288), .Y(n77300) );
  NAND2xp33_ASAP7_75t_SL U52628 ( .A(n76857), .B(n76927), .Y(n76575) );
  NAND2xp33_ASAP7_75t_SL U52629 ( .A(n74129), .B(n76927), .Y(n64160) );
  NAND2xp33_ASAP7_75t_SL U52630 ( .A(n77288), .B(n76927), .Y(n63950) );
  AOI22xp33_ASAP7_75t_SL U52631 ( .A1(n76922), .A2(n77290), .B1(n57135), .B2(
        n76928), .Y(n76921) );
  NAND2xp33_ASAP7_75t_SL U52632 ( .A(n76999), .B(n76927), .Y(n76585) );
  NAND2xp33_ASAP7_75t_SL U52633 ( .A(n75312), .B(n76927), .Y(n63928) );
  NAND2xp33_ASAP7_75t_SL U52634 ( .A(n76553), .B(n76927), .Y(n76526) );
  NAND2xp33_ASAP7_75t_SL U52635 ( .A(n77277), .B(n76927), .Y(n76213) );
  NAND2xp33_ASAP7_75t_SL U52636 ( .A(n75783), .B(n76927), .Y(n63727) );
  NAND2xp33_ASAP7_75t_SL U52637 ( .A(n77227), .B(n76927), .Y(n63961) );
  NAND2xp33_ASAP7_75t_SL U52638 ( .A(n76928), .B(n76927), .Y(n76929) );
  NAND2xp33_ASAP7_75t_SL U52639 ( .A(n75686), .B(n76927), .Y(n75635) );
  NAND2xp33_ASAP7_75t_SL U52640 ( .A(n69373), .B(n76927), .Y(n65189) );
  NAND2xp33_ASAP7_75t_SL U52641 ( .A(n75200), .B(n76927), .Y(n75178) );
  NAND2xp33_ASAP7_75t_SL U52642 ( .A(n76232), .B(n76927), .Y(n63933) );
  NAND2xp33_ASAP7_75t_SL U52643 ( .A(n75798), .B(n76927), .Y(n75154) );
  NAND2xp33_ASAP7_75t_SL U52644 ( .A(n76619), .B(n76927), .Y(n76598) );
  NAND2xp33_ASAP7_75t_SL U52645 ( .A(n77021), .B(n76927), .Y(n63973) );
  NAND2xp33_ASAP7_75t_SL U52646 ( .A(n75449), .B(n76927), .Y(n64262) );
  NAND2xp33_ASAP7_75t_SL U52647 ( .A(n76704), .B(n76927), .Y(n76705) );
  INVxp67_ASAP7_75t_SL U52648 ( .A(n70590), .Y(n70591) );
  NAND2xp33_ASAP7_75t_SL U52649 ( .A(n74081), .B(n76927), .Y(n65216) );
  NAND2xp33_ASAP7_75t_SL U52650 ( .A(n77153), .B(n76927), .Y(n63991) );
  INVx2_ASAP7_75t_SL U52651 ( .A(n74503), .Y(n74454) );
  INVx1_ASAP7_75t_SL U52652 ( .A(n69228), .Y(n57087) );
  INVxp67_ASAP7_75t_SL U52653 ( .A(n68629), .Y(n68632) );
  AOI21xp33_ASAP7_75t_SL U52654 ( .A1(n1642), .A2(n57144), .B(n76877), .Y(
        n1643) );
  AOI22xp33_ASAP7_75t_SL U52655 ( .A1(n73610), .A2(n73609), .B1(n73608), .B2(
        n73607), .Y(n1528) );
  NAND2xp33_ASAP7_75t_SL U52656 ( .A(icqmem_adr_qmem[31]), .B(n57136), .Y(
        n77318) );
  NAND2xp33_ASAP7_75t_SL U52657 ( .A(icqmem_adr_qmem[20]), .B(n57136), .Y(
        n77323) );
  NAND2xp33_ASAP7_75t_SL U52658 ( .A(icqmem_adr_qmem[30]), .B(n57136), .Y(
        n77326) );
  NAND2xp33_ASAP7_75t_SL U52659 ( .A(icqmem_adr_qmem[29]), .B(n57136), .Y(
        n77319) );
  AOI21xp33_ASAP7_75t_SL U52660 ( .A1(n2549), .A2(n57144), .B(n73956), .Y(
        n2550) );
  NAND2xp33_ASAP7_75t_SL U52661 ( .A(icqmem_adr_qmem[25]), .B(n57136), .Y(
        n77328) );
  NAND2xp33_ASAP7_75t_SL U52662 ( .A(icqmem_adr_qmem[23]), .B(n57136), .Y(
        n77329) );
  NAND2xp33_ASAP7_75t_SL U52663 ( .A(icqmem_adr_qmem[28]), .B(n57136), .Y(
        n77331) );
  INVxp67_ASAP7_75t_SL U52664 ( .A(n65107), .Y(n65109) );
  NAND2xp33_ASAP7_75t_SL U52665 ( .A(icqmem_adr_qmem[24]), .B(n57136), .Y(
        n77330) );
  NAND2xp33_ASAP7_75t_SL U52666 ( .A(icqmem_adr_qmem[27]), .B(n57136), .Y(
        n77325) );
  NAND2xp33_ASAP7_75t_SL U52667 ( .A(icqmem_adr_qmem[22]), .B(n57136), .Y(
        n77333) );
  NAND2xp33_ASAP7_75t_SL U52668 ( .A(icqmem_adr_qmem[21]), .B(n57136), .Y(
        n77320) );
  NAND2xp33_ASAP7_75t_SL U52669 ( .A(icqmem_adr_qmem[26]), .B(n57136), .Y(
        n77324) );
  NAND2xp33_ASAP7_75t_SL U52670 ( .A(n70609), .B(n70608), .Y(n70611) );
  INVxp67_ASAP7_75t_SL U52671 ( .A(n70601), .Y(n70604) );
  AOI21xp33_ASAP7_75t_SL U52672 ( .A1(n1608), .A2(n57144), .B(n74076), .Y(
        n1609) );
  OAI22xp33_ASAP7_75t_SL U52673 ( .A1(n839), .A2(n58524), .B1(n837), .B2(
        n59683), .Y(n9422) );
  OAI22xp33_ASAP7_75t_SL U52674 ( .A1(n845), .A2(n58524), .B1(n843), .B2(
        n59683), .Y(n9421) );
  INVxp67_ASAP7_75t_SL U52675 ( .A(n77394), .Y(n61048) );
  INVxp67_ASAP7_75t_SL U52676 ( .A(n58812), .Y(n57887) );
  OAI21xp5_ASAP7_75t_SL U52677 ( .A1(n751), .A2(n77385), .B(n77384), .Y(n9165)
         );
  OAI22xp33_ASAP7_75t_SL U52678 ( .A1(n59699), .A2(n70892), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_17_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n154) );
  INVxp67_ASAP7_75t_SL U52679 ( .A(n66603), .Y(n66598) );
  OAI22xp33_ASAP7_75t_SL U52680 ( .A1(n883), .A2(n58524), .B1(n876), .B2(
        n59683), .Y(n9409) );
  OAI22xp33_ASAP7_75t_SL U52681 ( .A1(n1044), .A2(n58524), .B1(n1042), .B2(
        n59682), .Y(n9419) );
  OAI22xp33_ASAP7_75t_SL U52682 ( .A1(n874), .A2(n58524), .B1(n867), .B2(
        n59683), .Y(n9410) );
  OAI22xp33_ASAP7_75t_SL U52683 ( .A1(n892), .A2(n58524), .B1(n885), .B2(
        n59683), .Y(n9408) );
  OAI22xp33_ASAP7_75t_SL U52684 ( .A1(n865), .A2(n58524), .B1(n858), .B2(
        n59683), .Y(n9411) );
  OAI22xp33_ASAP7_75t_SL U52685 ( .A1(n901), .A2(n58524), .B1(n894), .B2(
        n59683), .Y(n9407) );
  OAI22xp33_ASAP7_75t_SL U52686 ( .A1(n1033), .A2(n58524), .B1(n1031), .B2(
        n59683), .Y(n9420) );
  OAI22xp33_ASAP7_75t_SL U52687 ( .A1(n856), .A2(n58524), .B1(n854), .B2(
        n59683), .Y(n9412) );
  OAI22xp33_ASAP7_75t_SL U52688 ( .A1(n910), .A2(n58524), .B1(n903), .B2(
        n59682), .Y(n9406) );
  OAI22xp33_ASAP7_75t_SL U52689 ( .A1(n1027), .A2(n58524), .B1(n1020), .B2(
        n59682), .Y(n9393) );
  OAI22xp33_ASAP7_75t_SL U52690 ( .A1(n1018), .A2(n58524), .B1(n1011), .B2(
        n59682), .Y(n9394) );
  NAND2xp5_ASAP7_75t_SL U52691 ( .A(n74225), .B(n74258), .Y(n74503) );
  OAI22xp33_ASAP7_75t_SL U52692 ( .A1(n1009), .A2(n58524), .B1(n1002), .B2(
        n59682), .Y(n9395) );
  OAI22xp33_ASAP7_75t_SL U52693 ( .A1(n919), .A2(n58524), .B1(n912), .B2(
        n59683), .Y(n9405) );
  OAI22xp33_ASAP7_75t_SL U52694 ( .A1(n1000), .A2(n58524), .B1(n993), .B2(
        n59682), .Y(n9396) );
  OAI22xp33_ASAP7_75t_SL U52695 ( .A1(n1055), .A2(n58524), .B1(n1053), .B2(
        n59682), .Y(n9418) );
  OAI22xp33_ASAP7_75t_SL U52696 ( .A1(n991), .A2(n58524), .B1(n984), .B2(
        n59682), .Y(n9397) );
  OAI22xp33_ASAP7_75t_SL U52697 ( .A1(n1066), .A2(n58524), .B1(n1064), .B2(
        n59683), .Y(n9417) );
  OAI22xp33_ASAP7_75t_SL U52698 ( .A1(n982), .A2(n58524), .B1(n975), .B2(
        n59682), .Y(n9398) );
  OAI22xp33_ASAP7_75t_SL U52699 ( .A1(n973), .A2(n58524), .B1(n966), .B2(
        n59682), .Y(n9399) );
  OAI22xp33_ASAP7_75t_SL U52700 ( .A1(n1110), .A2(n58524), .B1(n1108), .B2(
        n59682), .Y(n9413) );
  OAI22xp33_ASAP7_75t_SL U52701 ( .A1(n928), .A2(n58524), .B1(n921), .B2(
        n59682), .Y(n9404) );
  OAI22xp33_ASAP7_75t_SL U52702 ( .A1(n964), .A2(n58524), .B1(n957), .B2(
        n59682), .Y(n9400) );
  OAI22xp33_ASAP7_75t_SL U52703 ( .A1(n1099), .A2(n58524), .B1(n1097), .B2(
        n59683), .Y(n9414) );
  OAI22xp33_ASAP7_75t_SL U52704 ( .A1(n955), .A2(n58524), .B1(n948), .B2(
        n59682), .Y(n9401) );
  OAI22xp33_ASAP7_75t_SL U52705 ( .A1(n946), .A2(n58524), .B1(n939), .B2(
        n59682), .Y(n9402) );
  INVxp67_ASAP7_75t_SL U52706 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_27_), .Y(n73850)
         );
  OAI22xp33_ASAP7_75t_SL U52707 ( .A1(n937), .A2(n58524), .B1(n930), .B2(
        n59682), .Y(n9403) );
  OAI22xp33_ASAP7_75t_SL U52708 ( .A1(n1088), .A2(n58524), .B1(n1086), .B2(
        n59683), .Y(n9415) );
  NAND2xp5_ASAP7_75t_SL U52709 ( .A(n60353), .B(n60352), .Y(n9451) );
  NAND2xp5_ASAP7_75t_SL U52710 ( .A(n60346), .B(n60345), .Y(n9452) );
  NAND2xp33_ASAP7_75t_SL U52711 ( .A(n66606), .B(n66605), .Y(n66609) );
  XNOR2xp5_ASAP7_75t_SL U52712 ( .A(n66601), .B(n66600), .Y(n66603) );
  NAND2xp5_ASAP7_75t_SL U52713 ( .A(n60374), .B(n60373), .Y(n9453) );
  NAND2xp5_ASAP7_75t_SL U52714 ( .A(n60364), .B(n60363), .Y(n9454) );
  AND3x2_ASAP7_75t_SL U52715 ( .A(n63726), .B(n63725), .C(n63724), .Y(n76927)
         );
  NAND2xp5_ASAP7_75t_SL U52716 ( .A(n60384), .B(n60383), .Y(n9447) );
  NAND2xp5_ASAP7_75t_SL U52717 ( .A(n60390), .B(n60389), .Y(n9446) );
  INVxp33_ASAP7_75t_SL U52718 ( .A(n66441), .Y(n66444) );
  AOI22xp33_ASAP7_75t_SL U52719 ( .A1(n77237), .A2(n77920), .B1(n77168), .B2(
        n77235), .Y(n77169) );
  OAI22xp33_ASAP7_75t_SL U52720 ( .A1(n59698), .A2(n71038), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_24_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n175) );
  OAI21xp5_ASAP7_75t_SL U52721 ( .A1(n1095), .A2(n76523), .B(n74948), .Y(n9186) );
  INVxp67_ASAP7_75t_SL U52722 ( .A(n76256), .Y(n76318) );
  OAI21xp5_ASAP7_75t_SL U52723 ( .A1(n1084), .A2(n76523), .B(n76522), .Y(n9187) );
  OAI21xp5_ASAP7_75t_SL U52724 ( .A1(n59677), .A2(n77886), .B(n63604), .Y(
        n9621) );
  OAI22xp33_ASAP7_75t_SL U52725 ( .A1(n1853), .A2(n59156), .B1(n77348), .B2(
        n77344), .Y(n9164) );
  INVxp67_ASAP7_75t_SL U52726 ( .A(n75098), .Y(n75100) );
  OAI21xp33_ASAP7_75t_SL U52727 ( .A1(n57144), .A2(n77886), .B(n63602), .Y(
        n1659) );
  NAND2xp5_ASAP7_75t_SL U52728 ( .A(or1200_cpu_rf_rdb), .B(n77841), .Y(n77845)
         );
  OAI21xp33_ASAP7_75t_SL U52729 ( .A1(n57144), .A2(n77867), .B(n64866), .Y(
        n1574) );
  OAI21xp33_ASAP7_75t_SL U52730 ( .A1(n74899), .A2(n76941), .B(n77170), .Y(
        n74898) );
  INVxp67_ASAP7_75t_SL U52731 ( .A(n64696), .Y(n64550) );
  OAI21xp33_ASAP7_75t_SL U52732 ( .A1(n76664), .A2(n76663), .B(n76662), .Y(
        n77143) );
  AOI22xp33_ASAP7_75t_SL U52733 ( .A1(n60347), .A2(n57139), .B1(
        or1200_ic_top_from_icram[2]), .B2(n78022), .Y(n60345) );
  XNOR2xp5_ASAP7_75t_SL U52734 ( .A(n57041), .B(n57897), .Y(n63103) );
  AOI22xp33_ASAP7_75t_SL U52735 ( .A1(n60365), .A2(n57139), .B1(
        or1200_ic_top_from_icram[0]), .B2(n78022), .Y(n60363) );
  AOI22xp33_ASAP7_75t_SL U52736 ( .A1(n60375), .A2(n57139), .B1(
        or1200_ic_top_from_icram[1]), .B2(n59497), .Y(n60373) );
  OAI21xp5_ASAP7_75t_SL U52737 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_12_), .A2(n74858), 
        .B(n74857), .Y(n52507) );
  OAI21xp5_ASAP7_75t_SL U52738 ( .A1(n759), .A2(n76523), .B(n75175), .Y(n9167)
         );
  AOI22xp33_ASAP7_75t_SL U52739 ( .A1(n60385), .A2(n57139), .B1(
        or1200_ic_top_from_icram[7]), .B2(n78022), .Y(n60383) );
  OAI21xp5_ASAP7_75t_SL U52740 ( .A1(n767), .A2(n76523), .B(n75162), .Y(n9169)
         );
  AOI22xp33_ASAP7_75t_SL U52741 ( .A1(n60391), .A2(n57139), .B1(
        or1200_ic_top_from_icram[8]), .B2(n59497), .Y(n60389) );
  AOI22xp33_ASAP7_75t_SL U52742 ( .A1(n59701), .A2(n77383), .B1(n77382), .B2(
        n53441), .Y(n77384) );
  INVxp67_ASAP7_75t_SL U52743 ( .A(n66593), .Y(n66594) );
  NAND2xp5_ASAP7_75t_SL U52744 ( .A(n59499), .B(n76311), .Y(n74630) );
  AOI22xp33_ASAP7_75t_SL U52745 ( .A1(n60354), .A2(n57139), .B1(
        or1200_ic_top_from_icram[3]), .B2(n59497), .Y(n60352) );
  OA21x2_ASAP7_75t_SL U52746 ( .A1(n63294), .A2(n63293), .B(n63346), .Y(n63295) );
  INVxp67_ASAP7_75t_SL U52747 ( .A(n68639), .Y(n66580) );
  XNOR2xp5_ASAP7_75t_SL U52748 ( .A(n59007), .B(n66906), .Y(n59006) );
  INVx1_ASAP7_75t_SL U52749 ( .A(n78021), .Y(n77423) );
  INVxp33_ASAP7_75t_SL U52750 ( .A(n60451), .Y(n60452) );
  OAI21xp5_ASAP7_75t_SL U52751 ( .A1(n75310), .A2(n75309), .B(n75308), .Y(
        n76275) );
  OAI21xp5_ASAP7_75t_SL U52752 ( .A1(n59677), .A2(n77897), .B(n77029), .Y(
        n9625) );
  OAI21xp5_ASAP7_75t_SL U52753 ( .A1(n59677), .A2(n77905), .B(n61805), .Y(
        n9629) );
  NOR2xp33_ASAP7_75t_SL U52754 ( .A(n73860), .B(n73859), .Y(n73863) );
  NAND2xp33_ASAP7_75t_SL U52755 ( .A(iwb_dat_i[13]), .B(n78020), .Y(n7627) );
  NAND2xp33_ASAP7_75t_SL U52756 ( .A(iwb_dat_i[12]), .B(n78020), .Y(n7632) );
  INVxp33_ASAP7_75t_SL U52757 ( .A(n63476), .Y(n63479) );
  OAI21xp5_ASAP7_75t_SL U52758 ( .A1(n59677), .A2(n77891), .B(n62548), .Y(
        n9623) );
  AOI21xp33_ASAP7_75t_SL U52759 ( .A1(n1787), .A2(n57144), .B(n76556), .Y(
        n1788) );
  OAI21xp33_ASAP7_75t_SL U52760 ( .A1(n74629), .A2(n74628), .B(n74627), .Y(
        n76311) );
  NAND2xp33_ASAP7_75t_SL U52761 ( .A(iwb_dat_i[11]), .B(n78020), .Y(n7637) );
  NAND2xp33_ASAP7_75t_SL U52762 ( .A(iwb_dat_i[14]), .B(n78020), .Y(n7622) );
  OAI22xp33_ASAP7_75t_SL U52763 ( .A1(n59699), .A2(n70748), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_7_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n124) );
  INVx2_ASAP7_75t_SL U52764 ( .A(n69370), .Y(n77294) );
  NAND2xp33_ASAP7_75t_SL U52765 ( .A(iwb_dat_i[15]), .B(n78020), .Y(n7617) );
  OAI21xp5_ASAP7_75t_SL U52766 ( .A1(n59677), .A2(n77232), .B(n61130), .Y(
        n9626) );
  NAND2xp5_ASAP7_75t_SL U52767 ( .A(n76692), .B(n76691), .Y(n9668) );
  NAND2xp5_ASAP7_75t_SL U52768 ( .A(or1200_ic_top_from_icram[15]), .B(n58387), 
        .Y(n7616) );
  INVx2_ASAP7_75t_SL U52769 ( .A(n77454), .Y(n77376) );
  NAND2xp5_ASAP7_75t_SL U52770 ( .A(n61566), .B(n61565), .Y(n9667) );
  AOI21xp33_ASAP7_75t_SL U52771 ( .A1(n2564), .A2(n57144), .B(n75459), .Y(
        n2565) );
  NAND2xp5_ASAP7_75t_SL U52772 ( .A(n76656), .B(n76655), .Y(n9662) );
  NAND2xp5_ASAP7_75t_SL U52773 ( .A(n77245), .B(n77244), .Y(n9670) );
  XOR2xp5_ASAP7_75t_SL U52774 ( .A(n58946), .B(n58945), .Y(n63164) );
  AOI22xp33_ASAP7_75t_SL U52775 ( .A1(or1200_cpu_or1200_except_n555), .A2(
        n57144), .B1(n61059), .B2(n77567), .Y(or1200_cpu_or1200_except_n1821)
         );
  NAND2xp5_ASAP7_75t_SL U52776 ( .A(or1200_ic_top_from_icram[11]), .B(n58387), 
        .Y(n7636) );
  NAND2xp5_ASAP7_75t_SL U52777 ( .A(n77031), .B(n77030), .Y(n77130) );
  NAND2xp5_ASAP7_75t_SL U52778 ( .A(or1200_ic_top_from_icram[13]), .B(n58387), 
        .Y(n7626) );
  NOR2x1_ASAP7_75t_SL U52779 ( .A(n60317), .B(n77454), .Y(n77359) );
  INVxp67_ASAP7_75t_SL U52780 ( .A(n77362), .Y(n57089) );
  NAND2xp5_ASAP7_75t_SL U52781 ( .A(or1200_ic_top_from_icram[12]), .B(n58387), 
        .Y(n7631) );
  AOI21xp5_ASAP7_75t_SL U52782 ( .A1(n76274), .A2(n77031), .B(n75608), .Y(
        n75612) );
  NAND2xp5_ASAP7_75t_SL U52783 ( .A(or1200_ic_top_from_icram[14]), .B(n58387), 
        .Y(n7621) );
  OAI22xp33_ASAP7_75t_SL U52784 ( .A1(n59698), .A2(n70808), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_11_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n136) );
  INVxp67_ASAP7_75t_SL U52785 ( .A(n66449), .Y(n57435) );
  AOI22xp33_ASAP7_75t_SL U52786 ( .A1(n2045), .A2(n57144), .B1(n2054), .B2(
        n60486), .Y(n9198) );
  XNOR2xp5_ASAP7_75t_SL U52787 ( .A(n63682), .B(n63681), .Y(n63791) );
  AOI22xp33_ASAP7_75t_SL U52788 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[24]), 
        .B1(n74074), .B2(n77279), .Y(n74075) );
  AOI22xp33_ASAP7_75t_SL U52789 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[27]), 
        .B1(n73954), .B2(n77279), .Y(n73955) );
  NAND2xp33_ASAP7_75t_SL U52790 ( .A(n63710), .B(n74940), .Y(n74931) );
  AOI22xp33_ASAP7_75t_SL U52791 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[19]), 
        .B1(n76875), .B2(n77279), .Y(n76876) );
  AOI22xp33_ASAP7_75t_SL U52792 ( .A1(n77280), .A2(n77279), .B1(n77465), .B2(
        or1200_cpu_spr_dat_rf[7]), .Y(n77281) );
  AOI22xp33_ASAP7_75t_SL U52793 ( .A1(n75888), .A2(n77279), .B1(n77465), .B2(
        or1200_cpu_spr_dat_rf[28]), .Y(n75892) );
  OAI21xp5_ASAP7_75t_SL U52794 ( .A1(n70753), .A2(n70746), .B(n70752), .Y(
        n70747) );
  AOI22xp33_ASAP7_75t_SL U52795 ( .A1(or1200_cpu_rf_dataa_0_), .A2(n77465), 
        .B1(n77923), .B2(n77243), .Y(n77244) );
  AOI22xp33_ASAP7_75t_SL U52796 ( .A1(n77156), .A2(n77279), .B1(n77465), .B2(
        or1200_cpu_spr_dat_rf[15]), .Y(n77159) );
  INVxp67_ASAP7_75t_SL U52797 ( .A(n60330), .Y(n61043) );
  NAND2xp5_ASAP7_75t_SL U52798 ( .A(n70641), .B(n74220), .Y(n74271) );
  AOI22xp33_ASAP7_75t_SL U52799 ( .A1(n77242), .A2(n57144), .B1(n77241), .B2(
        n77279), .Y(n77245) );
  AOI21xp33_ASAP7_75t_SL U52800 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[12]), 
        .B(n77302), .Y(n77303) );
  XNOR2xp5_ASAP7_75t_SL U52801 ( .A(n63019), .B(n63020), .Y(n63038) );
  AOI22xp33_ASAP7_75t_SL U52802 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[11]), 
        .B1(n61741), .B2(n77279), .Y(n61742) );
  INVxp67_ASAP7_75t_SL U52803 ( .A(n57832), .Y(n58627) );
  AOI21xp33_ASAP7_75t_SL U52804 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[16]), 
        .B(n76240), .Y(n76241) );
  AOI21xp33_ASAP7_75t_SL U52805 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[13]), 
        .B(n77230), .Y(n77231) );
  INVx1_ASAP7_75t_SL U52806 ( .A(n77537), .Y(n62004) );
  AOI21xp33_ASAP7_75t_SL U52807 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[10]), 
        .B(n75786), .Y(n75787) );
  INVx1_ASAP7_75t_SL U52808 ( .A(n77137), .Y(n59678) );
  AOI22xp33_ASAP7_75t_SL U52809 ( .A1(n2575), .A2(n57144), .B1(n3117), .B2(
        n60486), .Y(n9201) );
  AOI22xp33_ASAP7_75t_SL U52810 ( .A1(n59079), .A2(n57144), .B1(n76870), .B2(
        n77279), .Y(n61566) );
  AOI22xp33_ASAP7_75t_SL U52811 ( .A1(or1200_cpu_spr_dat_rf[3]), .A2(n77465), 
        .B1(n77917), .B2(n77243), .Y(n61565) );
  AOI22xp33_ASAP7_75t_SL U52812 ( .A1(n75376), .A2(n77279), .B1(n77465), .B2(
        or1200_cpu_spr_dat_rf[17]), .Y(n75380) );
  NOR2xp33_ASAP7_75t_SL U52813 ( .A(n68615), .B(n68614), .Y(n75057) );
  AOI21xp33_ASAP7_75t_SL U52814 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[25]), 
        .B(n74108), .Y(n74109) );
  AOI21xp33_ASAP7_75t_SL U52815 ( .A1(n3068), .A2(n57144), .B(n77282), .Y(
        n3069) );
  AOI21xp33_ASAP7_75t_SL U52816 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[18]), 
        .B(n74989), .Y(n74990) );
  OAI21xp33_ASAP7_75t_SL U52817 ( .A1(n75554), .A2(n75553), .B(n75552), .Y(
        n76274) );
  AOI21xp33_ASAP7_75t_SL U52818 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[26]), 
        .B(n73903), .Y(n73904) );
  INVxp67_ASAP7_75t_SL U52819 ( .A(n75261), .Y(n75262) );
  INVxp33_ASAP7_75t_SL U52820 ( .A(n75306), .Y(n75309) );
  NOR2x1_ASAP7_75t_SL U52821 ( .A(n74221), .B(n74220), .Y(n74464) );
  AOI22xp33_ASAP7_75t_SL U52822 ( .A1(n76627), .A2(n57144), .B1(n76626), .B2(
        n77279), .Y(n76630) );
  AOI22xp33_ASAP7_75t_SL U52823 ( .A1(or1200_cpu_spr_dat_rf[6]), .A2(n77465), 
        .B1(n77912), .B2(n77243), .Y(n76629) );
  AOI22xp33_ASAP7_75t_SL U52824 ( .A1(n76220), .A2(n77279), .B1(n77465), .B2(
        or1200_cpu_spr_dat_rf[5]), .Y(n76223) );
  AO21x1_ASAP7_75t_SL U52825 ( .A1(n57144), .A2(n58084), .B(n77243), .Y(n58083) );
  INVxp33_ASAP7_75t_SL U52826 ( .A(n66446), .Y(n66447) );
  OAI21xp33_ASAP7_75t_SL U52827 ( .A1(n77206), .A2(n77205), .B(n77204), .Y(
        or1200_du_N108) );
  AOI22xp33_ASAP7_75t_SL U52828 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[14]), 
        .B1(n60730), .B2(n77279), .Y(n60890) );
  AOI22xp33_ASAP7_75t_SL U52829 ( .A1(or1200_cpu_spr_dat_rf[4]), .A2(n77465), 
        .B1(n77915), .B2(n77243), .Y(n61462) );
  AOI22xp33_ASAP7_75t_SL U52830 ( .A1(n59182), .A2(n57144), .B1(n77006), .B2(
        n77279), .Y(n61463) );
  AOI22xp33_ASAP7_75t_SL U52831 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[22]), 
        .B1(n75457), .B2(n77279), .Y(n75458) );
  AOI22xp33_ASAP7_75t_SL U52832 ( .A1(or1200_cpu_spr_dat_rf[8]), .A2(n77465), 
        .B1(n77909), .B2(n77243), .Y(n76655) );
  OAI22xp33_ASAP7_75t_SL U52833 ( .A1(n75260), .A2(n75261), .B1(n61985), .B2(
        n57215), .Y(n75680) );
  AOI22xp33_ASAP7_75t_SL U52834 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[23]), 
        .B1(n75626), .B2(n77279), .Y(n75630) );
  OAI21xp33_ASAP7_75t_SL U52835 ( .A1(n57144), .A2(n77907), .B(n76512), .Y(
        n1822) );
  AOI22xp33_ASAP7_75t_SL U52836 ( .A1(n53316), .A2(n57144), .B1(n76689), .B2(
        n77279), .Y(n76692) );
  AOI21xp33_ASAP7_75t_SL U52837 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[9]), 
        .B(n61377), .Y(n61378) );
  AOI22xp33_ASAP7_75t_SL U52838 ( .A1(or1200_cpu_spr_dat_rf[2]), .A2(n77465), 
        .B1(n77919), .B2(n77243), .Y(n76691) );
  AOI21xp33_ASAP7_75t_SL U52839 ( .A1(n77465), .A2(or1200_cpu_spr_dat_rf[20]), 
        .B(n74552), .Y(n74553) );
  OAI21xp33_ASAP7_75t_SL U52840 ( .A1(or1200_cpu_or1200_mult_mac_n187), .A2(
        n76889), .B(n65139), .Y(or1200_cpu_or1200_mult_mac_n1570) );
  INVxp67_ASAP7_75t_SL U52841 ( .A(n68616), .Y(n68618) );
  OAI21xp33_ASAP7_75t_SL U52842 ( .A1(or1200_cpu_or1200_mult_mac_n179), .A2(
        n76889), .B(n63906), .Y(or1200_cpu_or1200_mult_mac_n1574) );
  AOI21xp33_ASAP7_75t_SL U52843 ( .A1(n69184), .A2(n57080), .B(n69183), .Y(
        n69185) );
  AOI22xp5_ASAP7_75t_SL U52844 ( .A1(n57198), .A2(n73959), .B1(n73958), .B2(
        n73961), .Y(n74037) );
  OAI21xp33_ASAP7_75t_SL U52845 ( .A1(or1200_cpu_or1200_mult_mac_n177), .A2(
        n76889), .B(n63789), .Y(or1200_cpu_or1200_mult_mac_n1575) );
  INVxp67_ASAP7_75t_SL U52846 ( .A(n68637), .Y(n66564) );
  NAND2xp5_ASAP7_75t_SL U52847 ( .A(n62905), .B(n62904), .Y(n63311) );
  AOI21xp33_ASAP7_75t_SL U52848 ( .A1(n68969), .A2(n57080), .B(n68952), .Y(
        n68953) );
  AOI21xp33_ASAP7_75t_SL U52849 ( .A1(n73427), .A2(n73426), .B(n73425), .Y(
        n78214) );
  OAI22xp33_ASAP7_75t_SL U52850 ( .A1(n1804), .A2(n77463), .B1(n59541), .B2(
        n57073), .Y(n75786) );
  XNOR2xp5_ASAP7_75t_SL U52851 ( .A(n66837), .B(n66836), .Y(n66838) );
  OAI21xp33_ASAP7_75t_SL U52852 ( .A1(or1200_cpu_or1200_mult_mac_n193), .A2(
        n76889), .B(n65186), .Y(or1200_cpu_or1200_mult_mac_n1567) );
  OAI21xp33_ASAP7_75t_SL U52853 ( .A1(or1200_cpu_or1200_mult_mac_n195), .A2(
        n76889), .B(n68776), .Y(or1200_cpu_or1200_mult_mac_n1566) );
  OAI21xp33_ASAP7_75t_SL U52854 ( .A1(or1200_cpu_or1200_mult_mac_n191), .A2(
        n76889), .B(n65158), .Y(or1200_cpu_or1200_mult_mac_n1568) );
  OAI21xp33_ASAP7_75t_SL U52855 ( .A1(or1200_cpu_or1200_mult_mac_n197), .A2(
        n76889), .B(n75005), .Y(or1200_cpu_or1200_mult_mac_n1565) );
  AOI21xp33_ASAP7_75t_SL U52856 ( .A1(n69263), .A2(n57080), .B(n69262), .Y(
        n69269) );
  XNOR2xp5_ASAP7_75t_SL U52857 ( .A(n67577), .B(n67576), .Y(n67764) );
  OAI21xp33_ASAP7_75t_SL U52858 ( .A1(or1200_cpu_or1200_mult_mac_n201), .A2(
        n76889), .B(n68802), .Y(or1200_cpu_or1200_mult_mac_n1563) );
  OAI21xp33_ASAP7_75t_SL U52859 ( .A1(or1200_cpu_or1200_mult_mac_n159), .A2(
        n76889), .B(n63421), .Y(or1200_cpu_or1200_mult_mac_n1584) );
  OAI22xp33_ASAP7_75t_SL U52860 ( .A1(n2196), .A2(n77463), .B1(n59570), .B2(
        n57074), .Y(n77302) );
  AOI21xp5_ASAP7_75t_SL U52861 ( .A1(n63703), .A2(n77445), .B(
        or1200_cpu_or1200_except_n565), .Y(n63705) );
  OAI21xp33_ASAP7_75t_SL U52862 ( .A1(or1200_cpu_or1200_mult_mac_n165), .A2(
        n76889), .B(n63466), .Y(or1200_cpu_or1200_mult_mac_n1581) );
  INVx1_ASAP7_75t_SL U52863 ( .A(n71201), .Y(n71181) );
  OAI21xp33_ASAP7_75t_SL U52864 ( .A1(or1200_cpu_or1200_mult_mac_n151), .A2(
        n76889), .B(n63333), .Y(or1200_cpu_or1200_mult_mac_n1588) );
  INVx2_ASAP7_75t_SL U52865 ( .A(n77463), .Y(n77279) );
  INVx2_ASAP7_75t_SL U52866 ( .A(n77467), .Y(n77243) );
  OAI21xp33_ASAP7_75t_SL U52867 ( .A1(or1200_cpu_or1200_mult_mac_n167), .A2(
        n76889), .B(n63474), .Y(or1200_cpu_or1200_mult_mac_n1580) );
  INVxp67_ASAP7_75t_SL U52868 ( .A(n66428), .Y(n57712) );
  OAI21xp33_ASAP7_75t_SL U52869 ( .A1(or1200_cpu_or1200_mult_mac_n147), .A2(
        n76889), .B(n63291), .Y(or1200_cpu_or1200_mult_mac_n1590) );
  OAI21xp33_ASAP7_75t_SL U52870 ( .A1(or1200_cpu_or1200_mult_mac_n169), .A2(
        n76889), .B(n63496), .Y(or1200_cpu_or1200_mult_mac_n1579) );
  NAND2xp5_ASAP7_75t_SL U52871 ( .A(n57954), .B(n57953), .Y(n68025) );
  NOR2x1p5_ASAP7_75t_SL U52872 ( .A(n60312), .B(or1200_cpu_or1200_if_if_bypass), .Y(n60330) );
  NAND2x1p5_ASAP7_75t_SL U52873 ( .A(n77834), .B(n77459), .Y(n77454) );
  OAI21xp33_ASAP7_75t_SL U52874 ( .A1(or1200_cpu_or1200_mult_mac_n157), .A2(
        n76889), .B(n63408), .Y(or1200_cpu_or1200_mult_mac_n1585) );
  OAI21xp33_ASAP7_75t_SL U52875 ( .A1(or1200_cpu_or1200_mult_mac_n155), .A2(
        n76889), .B(n63360), .Y(or1200_cpu_or1200_mult_mac_n1586) );
  AOI21xp33_ASAP7_75t_SL U52876 ( .A1(n69217), .A2(n57080), .B(n69216), .Y(
        n69224) );
  INVxp67_ASAP7_75t_SL U52877 ( .A(n75058), .Y(n57846) );
  AOI22xp33_ASAP7_75t_SL U52878 ( .A1(or1200_dc_top_tag_17_), .A2(n59501), 
        .B1(n78073), .B2(n57142), .Y(n78074) );
  AND3x2_ASAP7_75t_SL U52879 ( .A(n57073), .B(n60728), .C(n61056), .Y(n77465)
         );
  NAND2x1_ASAP7_75t_SL U52880 ( .A(n60729), .B(n59691), .Y(n77463) );
  INVxp67_ASAP7_75t_SL U52881 ( .A(n63718), .Y(n77445) );
  AOI22xp5_ASAP7_75t_SL U52882 ( .A1(n71744), .A2(n71789), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_0_), .B2(
        n71749), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n114) );
  AOI22xp33_ASAP7_75t_SL U52883 ( .A1(or1200_dc_top_tag_19_), .A2(n59501), 
        .B1(n78065), .B2(n57142), .Y(n78066) );
  AOI22xp33_ASAP7_75t_SL U52884 ( .A1(or1200_dc_top_tag_18_), .A2(n59500), 
        .B1(n78069), .B2(n57142), .Y(n78070) );
  INVxp67_ASAP7_75t_SL U52885 ( .A(n63139), .Y(n63142) );
  NAND2xp5_ASAP7_75t_SL U52886 ( .A(or1200_cpu_or1200_except_n563), .B(n63718), 
        .Y(n63722) );
  INVxp33_ASAP7_75t_SL U52887 ( .A(n71406), .Y(n71398) );
  AOI22xp33_ASAP7_75t_SL U52888 ( .A1(or1200_dc_top_tag_9_), .A2(n59500), .B1(
        n78114), .B2(n57142), .Y(n78115) );
  AOI22xp33_ASAP7_75t_SL U52889 ( .A1(or1200_dc_top_tag_5_), .A2(n59501), .B1(
        n78130), .B2(n57142), .Y(n78131) );
  AOI22xp33_ASAP7_75t_SL U52890 ( .A1(or1200_dc_top_tag_14_), .A2(n59501), 
        .B1(n78085), .B2(n57142), .Y(n78086) );
  AOI22xp33_ASAP7_75t_SL U52891 ( .A1(or1200_dc_top_tag_2_), .A2(n59501), .B1(
        n78145), .B2(n57142), .Y(n78146) );
  AOI22xp33_ASAP7_75t_SL U52892 ( .A1(or1200_dc_top_tag_12_), .A2(n59500), 
        .B1(n78102), .B2(n57142), .Y(n78103) );
  INVx1_ASAP7_75t_SL U52893 ( .A(n65345), .Y(n65352) );
  AOI22xp33_ASAP7_75t_SL U52894 ( .A1(or1200_dc_top_tag_6_), .A2(n59500), .B1(
        n78126), .B2(n57142), .Y(n78127) );
  AOI22xp33_ASAP7_75t_SL U52895 ( .A1(or1200_dc_top_tag_13_), .A2(n78157), 
        .B1(n78097), .B2(n57142), .Y(n78098) );
  NAND2xp5_ASAP7_75t_SL U52896 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_21_), .B(
        n74430), .Y(n74443) );
  AOI22xp33_ASAP7_75t_SL U52897 ( .A1(or1200_dc_top_tag_1_), .A2(n78157), .B1(
        n78151), .B2(n57142), .Y(n78152) );
  AOI22xp33_ASAP7_75t_SL U52898 ( .A1(or1200_dc_top_tag_7_), .A2(n78157), .B1(
        n78122), .B2(n57142), .Y(n78123) );
  AOI22xp33_ASAP7_75t_SL U52899 ( .A1(or1200_dc_top_tag_8_), .A2(n59501), .B1(
        n78118), .B2(n57142), .Y(n78119) );
  AOI22xp33_ASAP7_75t_SL U52900 ( .A1(or1200_dc_top_tag_10_), .A2(n78157), 
        .B1(n78110), .B2(n57142), .Y(n78111) );
  AOI22xp33_ASAP7_75t_SL U52901 ( .A1(or1200_dc_top_tag_16_), .A2(n78157), 
        .B1(n78077), .B2(n57142), .Y(n78078) );
  AOI22xp33_ASAP7_75t_SL U52902 ( .A1(or1200_dc_top_tag_3_), .A2(n59500), .B1(
        n78141), .B2(n57142), .Y(n78142) );
  AOI22xp33_ASAP7_75t_SL U52903 ( .A1(or1200_dc_top_tag_0_), .A2(n59500), .B1(
        n78156), .B2(n57142), .Y(n78158) );
  NOR2xp33_ASAP7_75t_SL U52904 ( .A(n73456), .B(n73461), .Y(n73464) );
  AOI22xp33_ASAP7_75t_SL U52905 ( .A1(or1200_dc_top_tag_4_), .A2(n78157), .B1(
        n78135), .B2(n57142), .Y(n78136) );
  AOI22xp33_ASAP7_75t_SL U52906 ( .A1(or1200_dc_top_tag_11_), .A2(n59501), 
        .B1(n78106), .B2(n57142), .Y(n78107) );
  AOI22xp33_ASAP7_75t_SL U52907 ( .A1(or1200_dc_top_tag_15_), .A2(n59500), 
        .B1(n78081), .B2(n57142), .Y(n78082) );
  XNOR2xp5_ASAP7_75t_SL U52908 ( .A(n63651), .B(n63239), .Y(n63240) );
  XNOR2xp5_ASAP7_75t_SL U52909 ( .A(n63158), .B(n63071), .Y(n63139) );
  INVx1_ASAP7_75t_SL U52910 ( .A(n71788), .Y(n71749) );
  OAI21xp5_ASAP7_75t_SL U52911 ( .A1(n75882), .A2(n75881), .B(n58548), .Y(
        n75886) );
  NAND2x1_ASAP7_75t_SL U52912 ( .A(n68787), .B(n68813), .Y(n76889) );
  INVxp67_ASAP7_75t_SL U52913 ( .A(n71032), .Y(n70981) );
  NAND2xp33_ASAP7_75t_SL U52914 ( .A(n76514), .B(n57144), .Y(n76512) );
  AOI21xp33_ASAP7_75t_SL U52915 ( .A1(n74219), .A2(n76956), .B(n77171), .Y(
        n58821) );
  INVxp67_ASAP7_75t_SL U52916 ( .A(n70939), .Y(n70923) );
  NAND2xp33_ASAP7_75t_SL U52917 ( .A(n63601), .B(n57144), .Y(n63602) );
  NAND2xp5_ASAP7_75t_SL U52918 ( .A(n67730), .B(n58136), .Y(n67732) );
  XOR2xp5_ASAP7_75t_SL U52919 ( .A(n64449), .B(n64688), .Y(n57770) );
  OAI21xp5_ASAP7_75t_SL U52920 ( .A1(n62799), .A2(n62856), .B(n62798), .Y(
        n62811) );
  AOI21xp5_ASAP7_75t_SL U52921 ( .A1(n62464), .A2(n62463), .B(n62462), .Y(
        n62465) );
  NAND2xp33_ASAP7_75t_SL U52922 ( .A(n64154), .B(n57144), .Y(n64155) );
  NAND2xp33_ASAP7_75t_SL U52923 ( .A(n64865), .B(n57144), .Y(n64866) );
  OAI21xp33_ASAP7_75t_SL U52924 ( .A1(n66586), .A2(n66567), .B(n66566), .Y(
        n57967) );
  NAND2xp33_ASAP7_75t_SL U52925 ( .A(n71400), .B(n71399), .Y(n71403) );
  INVxp67_ASAP7_75t_SL U52926 ( .A(n66592), .Y(n66595) );
  INVx1_ASAP7_75t_SL U52927 ( .A(n66437), .Y(n66393) );
  AOI21xp33_ASAP7_75t_SL U52928 ( .A1(n69213), .A2(n69212), .B(n69279), .Y(
        n69214) );
  INVx1_ASAP7_75t_SL U52929 ( .A(n59313), .Y(n58796) );
  INVxp67_ASAP7_75t_SL U52930 ( .A(n69338), .Y(n69336) );
  NAND2xp33_ASAP7_75t_SL U52931 ( .A(n73571), .B(n73559), .Y(n73566) );
  INVx1_ASAP7_75t_SL U52932 ( .A(n62148), .Y(n62151) );
  INVx6_ASAP7_75t_SL U52933 ( .A(n78173), .Y(n59695) );
  INVx8_ASAP7_75t_SL U52934 ( .A(n78173), .Y(n57144) );
  NAND2xp5_ASAP7_75t_SL U52935 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_33_), .B(
        n74338), .Y(n74348) );
  INVxp67_ASAP7_75t_SL U52936 ( .A(n67178), .Y(n67188) );
  NAND2xp5_ASAP7_75t_SL U52937 ( .A(n66760), .B(n66759), .Y(n66815) );
  XNOR2xp5_ASAP7_75t_SL U52938 ( .A(n57146), .B(n57622), .Y(n57621) );
  INVx1_ASAP7_75t_SL U52939 ( .A(n63852), .Y(n63619) );
  NOR2xp33_ASAP7_75t_SL U52940 ( .A(n75815), .B(n75814), .Y(n75222) );
  NAND2xp5_ASAP7_75t_SL U52941 ( .A(n70922), .B(n70978), .Y(n70939) );
  OAI21xp33_ASAP7_75t_SL U52942 ( .A1(or1200_cpu_or1200_except_n548), .A2(
        n75685), .B(n76928), .Y(n61900) );
  INVxp33_ASAP7_75t_SL U52943 ( .A(n75685), .Y(n61840) );
  INVx2_ASAP7_75t_SL U52944 ( .A(n67767), .Y(n57095) );
  XNOR2xp5_ASAP7_75t_SL U52945 ( .A(n68358), .B(n68359), .Y(n68458) );
  OAI22xp33_ASAP7_75t_SL U52946 ( .A1(n59700), .A2(n77807), .B1(n57084), .B2(
        n1035), .Y(n1036) );
  OAI22xp33_ASAP7_75t_SL U52947 ( .A1(n59700), .A2(n77815), .B1(n57084), .B2(
        n849), .Y(n850) );
  OAI21xp33_ASAP7_75t_SL U52948 ( .A1(n62315), .A2(n62314), .B(n53470), .Y(
        n76298) );
  NAND2xp33_ASAP7_75t_SL U52949 ( .A(n63003), .B(n63002), .Y(n59224) );
  NOR2xp33_ASAP7_75t_SL U52950 ( .A(n64598), .B(n64597), .Y(n58028) );
  INVxp67_ASAP7_75t_SL U52951 ( .A(n61961), .Y(n64270) );
  NAND2xp5_ASAP7_75t_SL U52952 ( .A(n66642), .B(n66970), .Y(n66643) );
  NOR2xp33_ASAP7_75t_SL U52953 ( .A(n71799), .B(n71686), .Y(n71796) );
  NAND2xp5_ASAP7_75t_SL U52954 ( .A(n75200), .B(n75883), .Y(n75685) );
  XNOR2xp5_ASAP7_75t_SL U52955 ( .A(n58333), .B(n67098), .Y(n67178) );
  INVx1_ASAP7_75t_SL U52956 ( .A(n67132), .Y(n67135) );
  OAI22xp33_ASAP7_75t_SL U52957 ( .A1(n59700), .A2(n77811), .B1(n57084), .B2(
        n1079), .Y(n1080) );
  INVxp67_ASAP7_75t_SL U52958 ( .A(n67138), .Y(n67139) );
  NAND2xp5_ASAP7_75t_SL U52959 ( .A(n58528), .B(n59052), .Y(n62998) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U52960 ( .A1(n77998), .A2(n3105), .B(n61319), .C(
        n59889), .Y(n59892) );
  INVxp67_ASAP7_75t_SL U52961 ( .A(n70975), .Y(n70942) );
  OAI22xp33_ASAP7_75t_SL U52962 ( .A1(n59700), .A2(n77813), .B1(n57084), .B2(
        n1101), .Y(n1102) );
  OAI22xp33_ASAP7_75t_SL U52963 ( .A1(n59700), .A2(n77808), .B1(n57084), .B2(
        n1046), .Y(n1047) );
  NAND2xp5_ASAP7_75t_SL U52964 ( .A(n57676), .B(n57675), .Y(n57674) );
  OAI21xp33_ASAP7_75t_SL U52965 ( .A1(n68597), .A2(n68596), .B(n68595), .Y(
        n68598) );
  INVxp67_ASAP7_75t_SL U52966 ( .A(n67546), .Y(n67549) );
  MAJx2_ASAP7_75t_SL U52967 ( .A(n57868), .B(n59076), .C(n57867), .Y(n68447)
         );
  OAI22xp33_ASAP7_75t_SL U52968 ( .A1(n59700), .A2(n77822), .B1(n57084), .B2(
        n914), .Y(n915) );
  INVx2_ASAP7_75t_SL U52969 ( .A(n57467), .Y(n64879) );
  AOI21xp5_ASAP7_75t_SL U52970 ( .A1(n62077), .A2(n60785), .B(n60784), .Y(
        n61120) );
  INVx1_ASAP7_75t_SL U52971 ( .A(n59439), .Y(n57151) );
  NAND2xp5_ASAP7_75t_SL U52972 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_17_), .B(
        n74409), .Y(n74408) );
  INVx1_ASAP7_75t_SL U52973 ( .A(n70860), .Y(n70849) );
  XOR2xp5_ASAP7_75t_SL U52974 ( .A(n62771), .B(n62652), .Y(n58510) );
  INVx1_ASAP7_75t_SL U52975 ( .A(n67133), .Y(n67134) );
  OAI22xp33_ASAP7_75t_SL U52976 ( .A1(n59700), .A2(n77814), .B1(n57084), .B2(
        n2769), .Y(n2770) );
  INVx1_ASAP7_75t_SL U52977 ( .A(n71130), .Y(n71100) );
  NOR2xp33_ASAP7_75t_SRAM U52978 ( .A(n2796), .B(n76541), .Y(n77679) );
  NOR2xp33_ASAP7_75t_SL U52979 ( .A(n74059), .B(n74179), .Y(n74060) );
  OAI22xp33_ASAP7_75t_SL U52980 ( .A1(n59700), .A2(n77809), .B1(n57084), .B2(
        n1057), .Y(n1058) );
  NOR2xp33_ASAP7_75t_SL U52981 ( .A(n62089), .B(n61949), .Y(n61961) );
  OAI21xp5_ASAP7_75t_SL U52982 ( .A1(n67444), .A2(n67232), .B(n58493), .Y(
        n59052) );
  OAI22xp33_ASAP7_75t_SL U52983 ( .A1(n59700), .A2(n77810), .B1(n57084), .B2(
        n1068), .Y(n1069) );
  INVxp67_ASAP7_75t_SL U52984 ( .A(n65364), .Y(n65370) );
  NOR2x1_ASAP7_75t_SL U52985 ( .A(n58446), .B(n59077), .Y(n59076) );
  NOR2xp33_ASAP7_75t_SL U52986 ( .A(n64856), .B(n64857), .Y(n73937) );
  NAND2xp33_ASAP7_75t_SL U52987 ( .A(n57321), .B(n66352), .Y(n66325) );
  NOR2xp33_ASAP7_75t_SL U52988 ( .A(n70921), .B(n70920), .Y(n58303) );
  AOI21xp5_ASAP7_75t_SL U52989 ( .A1(n67464), .A2(n64936), .B(n64935), .Y(
        n65014) );
  INVxp67_ASAP7_75t_SL U52990 ( .A(n64470), .Y(n64468) );
  INVxp67_ASAP7_75t_SL U52991 ( .A(n53470), .Y(n61320) );
  XNOR2xp5_ASAP7_75t_SL U52992 ( .A(n57313), .B(n67618), .Y(n57634) );
  OAI22xp33_ASAP7_75t_SL U52993 ( .A1(n59700), .A2(n77812), .B1(n57084), .B2(
        n1090), .Y(n1091) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U52994 ( .A1(n61119), .A2(n77641), .B(n77128), .C(
        n61118), .Y(n61122) );
  AOI22xp5_ASAP7_75t_SL U52995 ( .A1(n77672), .A2(n77869), .B1(n77671), .B2(
        n77664), .Y(n52474) );
  INVxp33_ASAP7_75t_SL U52996 ( .A(n66557), .Y(n66321) );
  INVxp67_ASAP7_75t_SL U52997 ( .A(n67024), .Y(n67025) );
  NAND2xp5_ASAP7_75t_SL U52998 ( .A(or1200_dc_top_dirty), .B(n59890), .Y(
        n77470) );
  NOR2xp33_ASAP7_75t_SL U52999 ( .A(n75037), .B(n75039), .Y(n75064) );
  NOR2xp33_ASAP7_75t_SL U53000 ( .A(n67544), .B(n67543), .Y(n67546) );
  OAI21xp33_ASAP7_75t_SL U53001 ( .A1(n64339), .A2(n64336), .B(n64340), .Y(
        n58127) );
  NAND2xp5_ASAP7_75t_SL U53002 ( .A(n60215), .B(n76538), .Y(n76542) );
  OAI21xp33_ASAP7_75t_SL U53003 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[1]), .A2(n57190), .B(n72869), .Y(n1986) );
  NOR2xp33_ASAP7_75t_SL U53004 ( .A(n58011), .B(n66921), .Y(n66922) );
  NOR2xp33_ASAP7_75t_SL U53005 ( .A(n62796), .B(n62795), .Y(n62797) );
  INVxp67_ASAP7_75t_SL U53006 ( .A(n64559), .Y(n64560) );
  INVxp33_ASAP7_75t_SL U53007 ( .A(n64471), .Y(n64469) );
  INVxp67_ASAP7_75t_SL U53008 ( .A(n64558), .Y(n64561) );
  NAND2xp5_ASAP7_75t_SL U53009 ( .A(n59123), .B(n67304), .Y(n67800) );
  NAND2xp5_ASAP7_75t_SL U53010 ( .A(n68606), .B(n68605), .Y(n68609) );
  OAI21xp33_ASAP7_75t_SL U53011 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[9]), .A2(n57190), .B(n72802), .Y(n1816) );
  NAND2xp5_ASAP7_75t_SL U53012 ( .A(n4114), .B(n78252), .Y(icqmem_adr_qmem[22]) );
  INVxp67_ASAP7_75t_SL U53013 ( .A(n64571), .Y(n64508) );
  NAND2xp5_ASAP7_75t_SL U53014 ( .A(n64251), .B(n64755), .Y(n64857) );
  INVxp67_ASAP7_75t_SL U53015 ( .A(n62785), .Y(n62792) );
  INVxp67_ASAP7_75t_SL U53016 ( .A(n70712), .Y(n70730) );
  INVxp33_ASAP7_75t_SL U53017 ( .A(n61957), .Y(n61958) );
  AOI21xp33_ASAP7_75t_SL U53018 ( .A1(n69085), .A2(n57080), .B(n69075), .Y(
        n69081) );
  INVx1_ASAP7_75t_SL U53019 ( .A(n64598), .Y(n57154) );
  OA21x2_ASAP7_75t_SL U53020 ( .A1(n75076), .A2(n66540), .B(n66539), .Y(n57762) );
  NAND2xp5_ASAP7_75t_SL U53021 ( .A(n58498), .B(n59613), .Y(n58750) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U53022 ( .A1(n75030), .A2(n62404), .B(n62403), 
        .C(n62407), .Y(n62405) );
  INVx1_ASAP7_75t_SL U53023 ( .A(n68402), .Y(n68400) );
  INVxp33_ASAP7_75t_SL U53024 ( .A(n62309), .Y(n62311) );
  OAI21xp33_ASAP7_75t_SL U53025 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[17]), .A2(
        n57190), .B(n72737), .Y(n1669) );
  OAI21xp33_ASAP7_75t_SL U53026 ( .A1(n70986), .A2(n71149), .B(n70934), .Y(
        n70936) );
  NOR2xp33_ASAP7_75t_SL U53027 ( .A(n75648), .B(n62403), .Y(n62398) );
  INVxp33_ASAP7_75t_SL U53028 ( .A(n62888), .Y(n62891) );
  INVxp67_ASAP7_75t_SL U53029 ( .A(n63853), .Y(n63618) );
  INVxp67_ASAP7_75t_SL U53030 ( .A(n62824), .Y(n62825) );
  INVxp67_ASAP7_75t_SL U53031 ( .A(n62829), .Y(n62826) );
  INVxp67_ASAP7_75t_SL U53032 ( .A(n67282), .Y(n58011) );
  OAI21xp5_ASAP7_75t_SL U53033 ( .A1(n59163), .A2(n53612), .B(n59162), .Y(
        n68402) );
  AOI21xp33_ASAP7_75t_SL U53034 ( .A1(n71090), .A2(n71315), .B(n70933), .Y(
        n70934) );
  INVxp67_ASAP7_75t_SL U53035 ( .A(n62788), .Y(n62790) );
  INVxp33_ASAP7_75t_SL U53036 ( .A(n70698), .Y(n70696) );
  OAI22xp33_ASAP7_75t_SL U53037 ( .A1(n72763), .A2(n72762), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[12]), .B2(
        n57190), .Y(n1939) );
  OAI21xp33_ASAP7_75t_SL U53038 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[8]), .A2(n57190), .B(n72794), .Y(n1946) );
  NOR2xp33_ASAP7_75t_SL U53039 ( .A(n57911), .B(n57686), .Y(n66764) );
  OAI22xp33_ASAP7_75t_SL U53040 ( .A1(n71285), .A2(n71149), .B1(n71284), .B2(
        n71139), .Y(n71144) );
  OAI21xp33_ASAP7_75t_SL U53041 ( .A1(n72963), .A2(n72969), .B(n72962), .Y(
        n72983) );
  OAI22xp33_ASAP7_75t_SL U53042 ( .A1(n72721), .A2(n72720), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]), .B2(
        n57190), .Y(n1926) );
  OAI21xp33_ASAP7_75t_SL U53043 ( .A1(n77600), .A2(n76890), .B(n62304), .Y(
        n9269) );
  AOI21xp5_ASAP7_75t_SL U53044 ( .A1(n63473), .A2(n59674), .B(n63472), .Y(
        n63474) );
  OAI21xp33_ASAP7_75t_SL U53045 ( .A1(n74079), .A2(n76890), .B(n66234), .Y(
        n9250) );
  NOR2xp33_ASAP7_75t_SL U53046 ( .A(n60082), .B(n65191), .Y(n78263) );
  INVxp67_ASAP7_75t_SL U53047 ( .A(n62966), .Y(n62926) );
  NOR2xp33_ASAP7_75t_SL U53048 ( .A(n60070), .B(n64258), .Y(n78259) );
  INVx1_ASAP7_75t_SL U53049 ( .A(n71359), .Y(n71381) );
  NAND3xp33_ASAP7_75t_SRAM U53050 ( .A(n75770), .B(n75769), .C(n76719), .Y(
        n75771) );
  OAI21xp33_ASAP7_75t_SL U53051 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[18]), .A2(
        n57190), .B(n72705), .Y(n1653) );
  AOI21xp33_ASAP7_75t_SL U53052 ( .A1(n71117), .A2(n71315), .B(n70988), .Y(
        n70989) );
  INVxp33_ASAP7_75t_SL U53053 ( .A(n62308), .Y(n62312) );
  BUFx3_ASAP7_75t_SL U53054 ( .A(n59650), .Y(n57325) );
  AOI22xp33_ASAP7_75t_SL U53055 ( .A1(n71396), .A2(n71001), .B1(n71394), .B2(
        n71000), .Y(n71002) );
  OAI22xp33_ASAP7_75t_SL U53056 ( .A1(or1200_cpu_spr_dat_ppc[22]), .A2(n59676), 
        .B1(or1200_cpu_or1200_except_n232), .B2(n57170), .Y(n64287) );
  OAI21xp33_ASAP7_75t_SL U53057 ( .A1(or1200_cpu_or1200_except_n230), .A2(
        n57170), .B(n62100), .Y(n62101) );
  AOI22xp33_ASAP7_75t_SL U53058 ( .A1(n59526), .A2(n70813), .B1(n71365), .B2(
        n70846), .Y(n70814) );
  OAI22xp33_ASAP7_75t_SL U53059 ( .A1(or1200_cpu_or1200_except_n646), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n534), .B2(n77032), .Y(n75566)
         );
  OAI22xp33_ASAP7_75t_SL U53060 ( .A1(or1200_cpu_or1200_except_n461), .A2(
        n59676), .B1(or1200_cpu_or1200_except_n234), .B2(n57170), .Y(n75565)
         );
  OAI21xp5_ASAP7_75t_SL U53061 ( .A1(n75644), .A2(n75927), .B(n67280), .Y(
        n67747) );
  INVxp67_ASAP7_75t_SL U53062 ( .A(n75358), .Y(n64216) );
  NAND2xp33_ASAP7_75t_SL U53063 ( .A(n69902), .B(n70001), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[4]) );
  INVxp33_ASAP7_75t_SL U53064 ( .A(n66537), .Y(n66540) );
  NAND2xp5_ASAP7_75t_SL U53065 ( .A(n72806), .B(n72868), .Y(n72801) );
  NAND2xp33_ASAP7_75t_SL U53066 ( .A(n58549), .B(n75358), .Y(n75359) );
  OAI22xp33_ASAP7_75t_SL U53067 ( .A1(n65354), .A2(n65304), .B1(n65322), .B2(
        n65303), .Y(n65305) );
  OAI22xp33_ASAP7_75t_SL U53068 ( .A1(or1200_cpu_or1200_except_n607), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n508), .B2(n77032), .Y(n61760)
         );
  OAI22xp33_ASAP7_75t_SL U53069 ( .A1(or1200_cpu_or1200_except_n401), .A2(
        n59676), .B1(or1200_cpu_or1200_except_n194), .B2(n57170), .Y(n61466)
         );
  AOI22xp33_ASAP7_75t_SL U53070 ( .A1(n71263), .A2(n71001), .B1(n71315), .B2(
        n71000), .Y(n70854) );
  AOI21xp5_ASAP7_75t_SL U53071 ( .A1(n67444), .A2(n57485), .B(n59211), .Y(
        n63113) );
  OAI22xp33_ASAP7_75t_SL U53072 ( .A1(or1200_cpu_spr_dat_ppc[27]), .A2(n59676), 
        .B1(or1200_cpu_or1200_except_n242), .B2(n57170), .Y(n73913) );
  OAI21xp33_ASAP7_75t_SL U53073 ( .A1(n856), .A2(n57168), .B(n63943), .Y(
        n63944) );
  AOI21xp33_ASAP7_75t_SL U53074 ( .A1(n72897), .A2(n72947), .B(n72940), .Y(
        n72927) );
  OAI21xp33_ASAP7_75t_SL U53075 ( .A1(or1200_cpu_or1200_except_n228), .A2(
        n57170), .B(n64103), .Y(n64104) );
  NAND2xp33_ASAP7_75t_SL U53076 ( .A(n67148), .B(n57336), .Y(n67149) );
  INVx2_ASAP7_75t_SL U53077 ( .A(n57567), .Y(n67975) );
  OAI21xp5_ASAP7_75t_SL U53078 ( .A1(n72879), .A2(n72868), .B(n72867), .Y(
        n72870) );
  AOI21xp5_ASAP7_75t_SL U53079 ( .A1(n63465), .A2(n59674), .B(n63464), .Y(
        n63466) );
  INVx1_ASAP7_75t_SL U53080 ( .A(n71210), .Y(n71230) );
  AOI22xp33_ASAP7_75t_SL U53081 ( .A1(n71263), .A2(n71248), .B1(n71315), .B2(
        n71193), .Y(n71107) );
  INVxp67_ASAP7_75t_SL U53082 ( .A(n71140), .Y(n71141) );
  AOI21xp5_ASAP7_75t_SL U53083 ( .A1(n73005), .A2(n72987), .B(n72778), .Y(
        n72779) );
  AOI22xp33_ASAP7_75t_SL U53084 ( .A1(n58861), .A2(n67948), .B1(n67276), .B2(
        n67431), .Y(n67277) );
  NAND2xp33_ASAP7_75t_SL U53085 ( .A(n57321), .B(n68101), .Y(n67372) );
  INVx1_ASAP7_75t_SL U53086 ( .A(n57067), .Y(n57096) );
  NAND2xp5_ASAP7_75t_SL U53087 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_14_), 
        .B(n74350), .Y(n74387) );
  NAND2xp5_ASAP7_75t_SL U53088 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[3]), .B(n65416), .Y(
        n65559) );
  OAI22xp33_ASAP7_75t_SL U53089 ( .A1(or1200_cpu_or1200_except_n667), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n548), .B2(n77032), .Y(n75698)
         );
  INVxp67_ASAP7_75t_SL U53090 ( .A(n63800), .Y(n57874) );
  INVxp33_ASAP7_75t_SL U53091 ( .A(n60210), .Y(n59884) );
  NOR2xp33_ASAP7_75t_SL U53092 ( .A(n63909), .B(n62397), .Y(n62403) );
  OAI21xp33_ASAP7_75t_SL U53093 ( .A1(or1200_cpu_or1200_except_n226), .A2(
        n57170), .B(n74589), .Y(n74590) );
  INVxp67_ASAP7_75t_SL U53094 ( .A(n78133), .Y(n78132) );
  INVx1_ASAP7_75t_SL U53095 ( .A(n67327), .Y(n58642) );
  INVxp67_ASAP7_75t_SL U53096 ( .A(n64441), .Y(n64443) );
  XNOR2xp5_ASAP7_75t_SL U53097 ( .A(n57109), .B(n75947), .Y(n67411) );
  INVxp67_ASAP7_75t_SL U53098 ( .A(n62750), .Y(n62751) );
  NAND2xp5_ASAP7_75t_SL U53099 ( .A(n58701), .B(n57180), .Y(n58700) );
  OAI21xp33_ASAP7_75t_SL U53100 ( .A1(n59604), .A2(n58431), .B(n63079), .Y(
        n63110) );
  INVxp67_ASAP7_75t_SL U53101 ( .A(n67473), .Y(n67476) );
  INVxp67_ASAP7_75t_SL U53102 ( .A(n67557), .Y(n67558) );
  NOR2x1_ASAP7_75t_SL U53103 ( .A(n67341), .B(n58449), .Y(n67844) );
  INVxp67_ASAP7_75t_SL U53104 ( .A(n65060), .Y(n67952) );
  INVx2_ASAP7_75t_SL U53105 ( .A(n67329), .Y(n57098) );
  INVxp33_ASAP7_75t_SL U53106 ( .A(n58849), .Y(n64480) );
  AOI21xp33_ASAP7_75t_SL U53107 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[19]), 
        .B(n74588), .Y(n74589) );
  NOR2xp33_ASAP7_75t_SRAM U53108 ( .A(n77943), .B(n76739), .Y(n76741) );
  NAND2xp33_ASAP7_75t_SL U53109 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_0_), .B(
        n76477), .Y(n76489) );
  OAI21xp5_ASAP7_75t_SL U53110 ( .A1(n69899), .A2(n69904), .B(n69572), .Y(
        n70001) );
  INVxp67_ASAP7_75t_SL U53111 ( .A(n60767), .Y(n60768) );
  INVx2_ASAP7_75t_SL U53112 ( .A(n77051), .Y(n59676) );
  OAI22xp33_ASAP7_75t_SL U53113 ( .A1(n71284), .A2(n70880), .B1(n71362), .B2(
        n70768), .Y(n70769) );
  AOI21xp33_ASAP7_75t_SL U53114 ( .A1(n75019), .A2(n57080), .B(n75001), .Y(
        n75002) );
  AOI21xp5_ASAP7_75t_SL U53115 ( .A1(n65185), .A2(n57080), .B(n65184), .Y(
        n65186) );
  OAI21xp33_ASAP7_75t_SL U53116 ( .A1(n1066), .A2(n57168), .B(n76816), .Y(
        n63738) );
  AOI21xp5_ASAP7_75t_SL U53117 ( .A1(n65138), .A2(n59674), .B(n65137), .Y(
        n65139) );
  OAI21xp33_ASAP7_75t_SL U53118 ( .A1(n1055), .A2(n57168), .B(n76603), .Y(
        n76605) );
  NAND2xp5_ASAP7_75t_SL U53119 ( .A(n73404), .B(n73408), .Y(n73349) );
  OAI22xp33_ASAP7_75t_SL U53120 ( .A1(n71149), .A2(n71046), .B1(n70885), .B2(
        n71362), .Y(n70886) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U53121 ( .A1(n76906), .A2(n63903), .B(n63902), .C(
        n63901), .Y(n63904) );
  INVx1_ASAP7_75t_SL U53122 ( .A(n71046), .Y(n71073) );
  INVx1_ASAP7_75t_SL U53123 ( .A(n73367), .Y(n73371) );
  INVx1_ASAP7_75t_SL U53124 ( .A(n73359), .Y(n73361) );
  OAI22xp33_ASAP7_75t_SL U53125 ( .A1(n71284), .A2(n71142), .B1(n71362), .B2(
        n71046), .Y(n71047) );
  OAI22xp33_ASAP7_75t_SL U53126 ( .A1(n71149), .A2(n71045), .B1(n71044), .B2(
        n71335), .Y(n71048) );
  OAI22xp33_ASAP7_75t_SL U53127 ( .A1(n71334), .A2(n71362), .B1(n71335), .B2(
        n71285), .Y(n71286) );
  AOI22xp33_ASAP7_75t_SL U53128 ( .A1(or1200_cpu_esr[0]), .A2(n77048), .B1(
        n59686), .B2(or1200_cpu_rf_dataa_0_), .Y(n60578) );
  AOI21xp33_ASAP7_75t_SL U53129 ( .A1(n77587), .A2(supv), .B(n60571), .Y(
        n60579) );
  NAND2xp5_ASAP7_75t_SL U53130 ( .A(n76009), .B(n76008), .Y(n76014) );
  NOR2xp33_ASAP7_75t_SL U53131 ( .A(n62135), .B(n75214), .Y(n75358) );
  NOR2xp33_ASAP7_75t_SL U53132 ( .A(n71413), .B(n70711), .Y(n70716) );
  OR2x2_ASAP7_75t_SL U53133 ( .A(n57317), .B(n70723), .Y(n58328) );
  OAI21xp33_ASAP7_75t_SL U53134 ( .A1(n1088), .A2(n57168), .B(n61276), .Y(
        n61277) );
  INVxp33_ASAP7_75t_SL U53135 ( .A(n68970), .Y(n68949) );
  NOR2xp33_ASAP7_75t_SL U53136 ( .A(n771), .B(n60173), .Y(n60031) );
  AOI21xp33_ASAP7_75t_SL U53137 ( .A1(n73963), .A2(n78253), .B(
        or1200_cpu_to_sr[2]), .Y(n60263) );
  OAI22xp33_ASAP7_75t_SL U53138 ( .A1(n1110), .A2(n57168), .B1(n4042), .B2(
        n76837), .Y(n76531) );
  OAI22xp33_ASAP7_75t_SL U53139 ( .A1(n1536), .A2(n74916), .B1(n59556), .B2(
        n74934), .Y(n74758) );
  NAND2xp33_ASAP7_75t_SL U53140 ( .A(or1200_cpu_spr_dat_rf[18]), .B(n59686), 
        .Y(n63559) );
  INVxp67_ASAP7_75t_SL U53141 ( .A(n75812), .Y(n61980) );
  NAND2xp5_ASAP7_75t_SL U53142 ( .A(n57260), .B(n75043), .Y(n75075) );
  NAND2xp33_ASAP7_75t_SL U53143 ( .A(n60174), .B(n60173), .Y(n60181) );
  INVx1_ASAP7_75t_SL U53144 ( .A(n71231), .Y(n71356) );
  OAI21xp5_ASAP7_75t_SL U53145 ( .A1(n73178), .A2(n73177), .B(n73175), .Y(
        n73433) );
  NAND2xp33_ASAP7_75t_SL U53146 ( .A(n64932), .B(n57180), .Y(n63812) );
  NOR2xp33_ASAP7_75t_SL U53147 ( .A(n68994), .B(n53432), .Y(n68970) );
  NAND2xp33_ASAP7_75t_SL U53148 ( .A(n70149), .B(n69825), .Y(n69483) );
  AOI21xp5_ASAP7_75t_SL U53149 ( .A1(n73294), .A2(n73293), .B(n73292), .Y(
        n73441) );
  INVx1_ASAP7_75t_SL U53150 ( .A(n73267), .Y(n73266) );
  OAI21xp5_ASAP7_75t_SL U53151 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), 
        .A2(n72711), .B(n72704), .Y(n72878) );
  INVx1_ASAP7_75t_SL U53152 ( .A(n62074), .Y(n74629) );
  OAI21xp5_ASAP7_75t_SL U53153 ( .A1(n1768), .A2(n77214), .B(n77213), .Y(
        or1200_cpu_to_sr[13]) );
  INVx2_ASAP7_75t_SL U53154 ( .A(n75958), .Y(n76176) );
  INVxp67_ASAP7_75t_SL U53155 ( .A(n67248), .Y(n62678) );
  OAI21xp33_ASAP7_75t_SL U53156 ( .A1(n1733), .A2(n61755), .B(n61255), .Y(
        n61256) );
  AOI21xp5_ASAP7_75t_SL U53157 ( .A1(n73282), .A2(n73281), .B(n73280), .Y(
        n73439) );
  INVxp67_ASAP7_75t_SL U53158 ( .A(n62767), .Y(n62727) );
  NAND2x1_ASAP7_75t_SL U53159 ( .A(n66332), .B(n66373), .Y(n64569) );
  INVxp67_ASAP7_75t_SL U53160 ( .A(n62725), .Y(n62726) );
  OAI21xp5_ASAP7_75t_SL U53161 ( .A1(n74123), .A2(n75298), .B(n74122), .Y(
        n74575) );
  NAND2xp5_ASAP7_75t_SL U53162 ( .A(n76675), .B(n61060), .Y(n77032) );
  BUFx2_ASAP7_75t_SL U53163 ( .A(n77848), .Y(n59686) );
  OAI22xp33_ASAP7_75t_SL U53164 ( .A1(n71231), .A2(n71284), .B1(n71362), .B2(
        n71262), .Y(n71232) );
  NAND2xp5_ASAP7_75t_SL U53165 ( .A(n61065), .B(n61480), .Y(n76739) );
  AOI21xp5_ASAP7_75t_SL U53166 ( .A1(n73274), .A2(n73273), .B(n73272), .Y(
        n73424) );
  NAND2xp33_ASAP7_75t_SL U53167 ( .A(n74043), .B(n74042), .Y(n78096) );
  OAI22xp33_ASAP7_75t_SL U53168 ( .A1(n66000), .A2(n66078), .B1(n65999), .B2(
        n65998), .Y(n66004) );
  OAI21xp33_ASAP7_75t_SL U53169 ( .A1(n70078), .A2(n69507), .B(n69506), .Y(
        n69562) );
  INVxp67_ASAP7_75t_SL U53170 ( .A(n71395), .Y(n71283) );
  OAI21xp33_ASAP7_75t_SL U53171 ( .A1(n73578), .A2(n73577), .B(n73576), .Y(
        n73653) );
  A2O1A1Ixp33_ASAP7_75t_SL U53172 ( .A1(n59168), .A2(n61523), .B(n61522), .C(
        n61521), .Y(n61541) );
  NOR2xp33_ASAP7_75t_SRAM U53173 ( .A(n76530), .B(n77269), .Y(n76532) );
  INVxp67_ASAP7_75t_SL U53174 ( .A(n73201), .Y(n73199) );
  NAND2xp5_ASAP7_75t_SL U53175 ( .A(n59985), .B(n60171), .Y(n60173) );
  AOI21xp33_ASAP7_75t_SL U53176 ( .A1(n65156), .A2(n57080), .B(n65153), .Y(
        n65154) );
  NAND2xp5_ASAP7_75t_SL U53177 ( .A(n73201), .B(n73200), .Y(n73460) );
  NOR2xp33_ASAP7_75t_SRAM U53178 ( .A(n76818), .B(n77269), .Y(n63737) );
  AOI21xp5_ASAP7_75t_SL U53179 ( .A1(n70954), .A2(n71314), .B(n70790), .Y(
        n70828) );
  INVx1_ASAP7_75t_SL U53180 ( .A(n66782), .Y(n63218) );
  INVx1_ASAP7_75t_SL U53181 ( .A(n65990), .Y(n66067) );
  AOI21xp5_ASAP7_75t_SL U53182 ( .A1(n73327), .A2(n73326), .B(n73325), .Y(
        n73328) );
  AOI21xp5_ASAP7_75t_SL U53183 ( .A1(n72864), .A2(n72876), .B(n72863), .Y(
        n72865) );
  NAND2xp33_ASAP7_75t_SL U53184 ( .A(n57221), .B(n59668), .Y(n66251) );
  AOI21xp5_ASAP7_75t_SL U53185 ( .A1(n73348), .A2(n73347), .B(n73346), .Y(
        n73404) );
  NAND2xp33_ASAP7_75t_SRAM U53186 ( .A(n75208), .B(n58416), .Y(n75209) );
  NOR2xp33_ASAP7_75t_SL U53187 ( .A(n60291), .B(n75673), .Y(n60292) );
  OAI22xp33_ASAP7_75t_SL U53188 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n72975), .B1(n72990), .B2(n72797), .Y(n72866) );
  AOI21xp5_ASAP7_75t_SL U53189 ( .A1(n73324), .A2(n73323), .B(n73322), .Y(
        n73369) );
  AOI22xp33_ASAP7_75t_SL U53190 ( .A1(n70777), .A2(n70812), .B1(n71314), .B2(
        n70898), .Y(n70813) );
  AOI22xp33_ASAP7_75t_SL U53191 ( .A1(n76216), .A2(n77587), .B1(n76217), .B2(
        n62508), .Y(n61613) );
  INVxp67_ASAP7_75t_SL U53192 ( .A(n61943), .Y(n61942) );
  NOR2xp33_ASAP7_75t_SL U53193 ( .A(n63543), .B(n61935), .Y(n62084) );
  OAI21xp33_ASAP7_75t_SL U53194 ( .A1(n60196), .A2(n75673), .B(n60195), .Y(
        n60206) );
  NAND2xp33_ASAP7_75t_SL U53195 ( .A(n57078), .B(n59668), .Y(n75054) );
  AOI22xp33_ASAP7_75t_SL U53196 ( .A1(n67960), .A2(n59508), .B1(n67962), .B2(
        n67961), .Y(n59155) );
  AND2x2_ASAP7_75t_SL U53197 ( .A(n62477), .B(n77250), .Y(n58401) );
  OAI21xp5_ASAP7_75t_SL U53198 ( .A1(n59630), .A2(n73115), .B(n73114), .Y(
        n73389) );
  NAND2xp33_ASAP7_75t_SL U53199 ( .A(n70118), .B(n69743), .Y(n69744) );
  NAND2xp33_ASAP7_75t_SL U53200 ( .A(n71314), .B(n71313), .Y(n71173) );
  INVxp33_ASAP7_75t_SL U53201 ( .A(n62228), .Y(n62227) );
  INVxp67_ASAP7_75t_SL U53202 ( .A(n71162), .Y(n71101) );
  INVxp67_ASAP7_75t_SL U53203 ( .A(n70778), .Y(n70779) );
  OAI22xp33_ASAP7_75t_SL U53204 ( .A1(n76897), .A2(n68788), .B1(n75675), .B2(
        n68787), .Y(n68801) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U53205 ( .A1(n62447), .A2(n57196), .B(n62446), .C(
        n75872), .Y(n62449) );
  OAI21xp33_ASAP7_75t_SL U53206 ( .A1(or1200_pic_picmr_19_), .A2(n74641), .B(
        n74640), .Y(n1353) );
  AOI21xp33_ASAP7_75t_SL U53207 ( .A1(n72738), .A2(n73028), .B(n72990), .Y(
        n72739) );
  NAND2xp5_ASAP7_75t_SL U53208 ( .A(n75903), .B(n57180), .Y(n62925) );
  NOR2xp33_ASAP7_75t_SRAM U53209 ( .A(n69890), .B(n69657), .Y(n69658) );
  INVx3_ASAP7_75t_SL U53210 ( .A(n75044), .Y(n75032) );
  OAI21xp5_ASAP7_75t_SL U53211 ( .A1(n72993), .A2(n72728), .B(n72703), .Y(
        n72711) );
  AOI21xp5_ASAP7_75t_SL U53212 ( .A1(n59674), .A2(n63290), .B(n63289), .Y(
        n63291) );
  OR2x2_ASAP7_75t_SL U53213 ( .A(n67288), .B(n57178), .Y(n58040) );
  INVxp67_ASAP7_75t_SL U53214 ( .A(n73200), .Y(n73198) );
  NAND2x1_ASAP7_75t_SL U53215 ( .A(n77210), .B(n73960), .Y(n77214) );
  O2A1O1Ixp33_ASAP7_75t_SL U53216 ( .A1(n61753), .A2(n61254), .B(n77589), .C(
        n61253), .Y(n61255) );
  NAND2xp33_ASAP7_75t_SRAM U53217 ( .A(n74578), .B(n74593), .Y(n64142) );
  OAI21xp33_ASAP7_75t_SL U53218 ( .A1(n70896), .A2(n70895), .B(n70894), .Y(
        n71090) );
  INVxp67_ASAP7_75t_SL U53219 ( .A(n61396), .Y(n61398) );
  AOI22xp5_ASAP7_75t_SL U53220 ( .A1(n73024), .A2(n72728), .B1(n72990), .B2(
        n72699), .Y(n72847) );
  AOI211xp5_ASAP7_75t_SL U53221 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[21]), .B(n70037), .C(n70036), .Y(n70039) );
  OAI21xp33_ASAP7_75t_SL U53222 ( .A1(n78342), .A2(n70054), .B(n69797), .Y(
        n70030) );
  INVx2_ASAP7_75t_SL U53223 ( .A(n59659), .Y(n57101) );
  INVxp67_ASAP7_75t_SL U53224 ( .A(n74276), .Y(n74239) );
  NAND2xp33_ASAP7_75t_SL U53225 ( .A(n65237), .B(n76735), .Y(n60906) );
  NAND2xp33_ASAP7_75t_SL U53226 ( .A(n70078), .B(n69505), .Y(n69506) );
  AOI22xp33_ASAP7_75t_SL U53227 ( .A1(n66024), .A2(n65916), .B1(n66051), .B2(
        n65915), .Y(n65919) );
  AOI21xp33_ASAP7_75t_SL U53228 ( .A1(n72768), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_), .B(
        n72877), .Y(n72777) );
  AOI21xp33_ASAP7_75t_SL U53229 ( .A1(n65610), .A2(n66092), .B(n65609), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n1) );
  INVxp67_ASAP7_75t_SL U53230 ( .A(n76750), .Y(n76757) );
  AOI22xp33_ASAP7_75t_SL U53231 ( .A1(n71209), .A2(n71208), .B1(n71245), .B2(
        n71207), .Y(n71231) );
  AND2x2_ASAP7_75t_SL U53232 ( .A(n53473), .B(n70896), .Y(n70723) );
  NOR2xp33_ASAP7_75t_SRAM U53233 ( .A(or1200_cpu_or1200_except_n276), .B(
        n76731), .Y(n61388) );
  NOR2xp67_ASAP7_75t_SL U53234 ( .A(n60818), .B(n60833), .Y(n77587) );
  OAI22xp5_ASAP7_75t_SL U53235 ( .A1(n71314), .A2(n71313), .B1(n71312), .B2(
        n71355), .Y(n71357) );
  AOI22xp33_ASAP7_75t_SL U53236 ( .A1(n66022), .A2(n65967), .B1(n65978), .B2(
        n65917), .Y(n65918) );
  O2A1O1Ixp33_ASAP7_75t_SL U53237 ( .A1(n61753), .A2(n61332), .B(n77610), .C(
        n61331), .Y(n61333) );
  AOI22xp33_ASAP7_75t_SL U53238 ( .A1(n57198), .A2(n75145), .B1(n77896), .B2(
        n58296), .Y(n75142) );
  NAND2xp5_ASAP7_75t_SL U53239 ( .A(n77125), .B(n62544), .Y(n60698) );
  INVx5_ASAP7_75t_SL U53240 ( .A(n75897), .Y(n57104) );
  NAND2xp33_ASAP7_75t_SRAM U53241 ( .A(n65653), .B(n65651), .Y(n65652) );
  INVxp33_ASAP7_75t_SL U53242 ( .A(n73170), .Y(n73174) );
  INVx2_ASAP7_75t_SL U53243 ( .A(n76091), .Y(n75912) );
  OAI21xp5_ASAP7_75t_SL U53244 ( .A1(n59630), .A2(n73193), .B(n73192), .Y(
        n73204) );
  BUFx3_ASAP7_75t_SL U53245 ( .A(n59644), .Y(n57322) );
  OAI22xp5_ASAP7_75t_SL U53246 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n72898), .B1(n72885), .B2(n72990), .Y(n72728) );
  O2A1O1Ixp33_ASAP7_75t_SL U53247 ( .A1(n60904), .A2(n61753), .B(n60977), .C(
        n60903), .Y(n60905) );
  AOI22xp33_ASAP7_75t_SL U53248 ( .A1(n66024), .A2(n65952), .B1(n66022), .B2(
        n65951), .Y(n65930) );
  NOR2x1_ASAP7_75t_SL U53249 ( .A(n58938), .B(n57554), .Y(n57553) );
  AOI22xp33_ASAP7_75t_SL U53250 ( .A1(n71209), .A2(n71172), .B1(n71245), .B2(
        n71171), .Y(n71313) );
  AOI21xp5_ASAP7_75t_SL U53251 ( .A1(n74249), .A2(n73891), .B(n74240), .Y(
        n74247) );
  NAND2xp33_ASAP7_75t_SL U53252 ( .A(n71245), .B(n71219), .Y(n71161) );
  NAND2xp33_ASAP7_75t_SL U53253 ( .A(n71245), .B(n70997), .Y(n70913) );
  NAND2xp33_ASAP7_75t_SL U53254 ( .A(n71087), .B(n71192), .Y(n70914) );
  NAND2xp33_ASAP7_75t_SL U53255 ( .A(n71245), .B(n71208), .Y(n71147) );
  OAI21xp5_ASAP7_75t_SL U53256 ( .A1(n59631), .A2(n73219), .B(n73218), .Y(
        n73254) );
  AOI21xp5_ASAP7_75t_SL U53257 ( .A1(n63420), .A2(n59674), .B(n63419), .Y(
        n63421) );
  AOI22xp33_ASAP7_75t_SL U53258 ( .A1(n71245), .A2(n71039), .B1(n71087), .B2(
        n71219), .Y(n70953) );
  INVxp67_ASAP7_75t_SL U53259 ( .A(n71085), .Y(n71089) );
  AOI22xp33_ASAP7_75t_SL U53260 ( .A1(n57198), .A2(n76217), .B1(n77977), .B2(
        n77212), .Y(n76215) );
  OAI22xp33_ASAP7_75t_SL U53261 ( .A1(n53473), .A2(n71311), .B1(n71015), .B2(
        n71171), .Y(n71228) );
  NAND2xp33_ASAP7_75t_SL U53262 ( .A(n71015), .B(n58301), .Y(n71014) );
  INVx1_ASAP7_75t_SL U53263 ( .A(n71012), .Y(n71207) );
  NAND2xp33_ASAP7_75t_SL U53264 ( .A(n71245), .B(n71040), .Y(n71041) );
  INVxp67_ASAP7_75t_SL U53265 ( .A(n73539), .Y(n73578) );
  INVxp67_ASAP7_75t_SL U53266 ( .A(n75869), .Y(n64237) );
  AOI22xp33_ASAP7_75t_SL U53267 ( .A1(n77089), .A2(n75577), .B1(n76761), .B2(
        n75576), .Y(n75581) );
  AOI21xp33_ASAP7_75t_SL U53268 ( .A1(n70706), .A2(n70695), .B(n70693), .Y(
        n70702) );
  NAND2xp33_ASAP7_75t_SL U53269 ( .A(n71332), .B(n71282), .Y(n71333) );
  NAND2xp5_ASAP7_75t_SL U53270 ( .A(n76065), .B(n75906), .Y(n76074) );
  INVxp33_ASAP7_75t_SL U53271 ( .A(n71244), .Y(n71247) );
  INVxp33_ASAP7_75t_SL U53272 ( .A(n71219), .Y(n71221) );
  NAND2xp33_ASAP7_75t_SL U53273 ( .A(n71245), .B(n71282), .Y(n71220) );
  AOI211xp5_ASAP7_75t_SRAM U53274 ( .A1(n77623), .A2(n61609), .B(n61604), .C(
        n61603), .Y(n61612) );
  AOI22xp33_ASAP7_75t_SL U53275 ( .A1(n71087), .A2(n71039), .B1(n70996), .B2(
        n71040), .Y(n70885) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U53276 ( .A1(n76749), .A2(n76748), .B(n76747), .C(
        n76746), .Y(n76758) );
  OAI21xp5_ASAP7_75t_SL U53277 ( .A1(n74196), .A2(n74195), .B(n74194), .Y(
        n74197) );
  INVx11_ASAP7_75t_SL U53278 ( .A(n59652), .Y(n57107) );
  AOI21xp33_ASAP7_75t_SL U53279 ( .A1(n71465), .A2(n71464), .B(n71463), .Y(
        n71466) );
  NAND2xp33_ASAP7_75t_SL U53280 ( .A(n69364), .B(n69363), .Y(n75194) );
  BUFx12f_ASAP7_75t_SL U53281 ( .A(n75761), .Y(n57108) );
  INVx3_ASAP7_75t_SL U53282 ( .A(n59608), .Y(n57109) );
  INVxp67_ASAP7_75t_SL U53283 ( .A(n61673), .Y(n61675) );
  OAI21xp33_ASAP7_75t_SL U53284 ( .A1(n72415), .A2(n72414), .B(n72413), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n74) );
  NAND2xp5_ASAP7_75t_SL U53285 ( .A(n74730), .B(n74727), .Y(n74276) );
  AOI22xp33_ASAP7_75t_SL U53286 ( .A1(n66024), .A2(n66007), .B1(n66022), .B2(
        n66006), .Y(n66010) );
  NAND2xp33_ASAP7_75t_SL U53287 ( .A(n74639), .B(n74641), .Y(n74640) );
  NAND2xp5_ASAP7_75t_SL U53288 ( .A(n66063), .B(n66076), .Y(n66052) );
  NAND2x1p5_ASAP7_75t_SL U53289 ( .A(n56854), .B(n58057), .Y(n75908) );
  AOI22xp33_ASAP7_75t_SL U53290 ( .A1(n73030), .A2(n72908), .B1(n73028), .B2(
        n72889), .Y(n72742) );
  NAND2xp5_ASAP7_75t_SL U53291 ( .A(n75618), .B(n78089), .Y(n75617) );
  O2A1O1Ixp5_ASAP7_75t_SL U53292 ( .A1(n76784), .A2(n76783), .B(n76782), .C(
        n76781), .Y(n76785) );
  INVxp67_ASAP7_75t_SL U53293 ( .A(n63545), .Y(n61934) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U53294 ( .A1(n61753), .A2(n61752), .B(n77613), .C(
        n61751), .Y(n61754) );
  OAI21xp33_ASAP7_75t_SL U53295 ( .A1(n72996), .A2(n72995), .B(n72994), .Y(
        n72997) );
  INVxp67_ASAP7_75t_SL U53296 ( .A(n60745), .Y(n60746) );
  AOI22xp33_ASAP7_75t_SL U53297 ( .A1(n57198), .A2(n63764), .B1(n77918), .B2(
        n77212), .Y(n60262) );
  NAND2xp33_ASAP7_75t_SL U53298 ( .A(n72886), .B(n72898), .Y(n72928) );
  NAND2xp5_ASAP7_75t_SL U53299 ( .A(n63545), .B(n75310), .Y(n62085) );
  INVx1_ASAP7_75t_SL U53300 ( .A(n67749), .Y(n57177) );
  INVx1_ASAP7_75t_SL U53301 ( .A(n72890), .Y(n72908) );
  INVxp67_ASAP7_75t_SL U53302 ( .A(n72916), .Y(n72787) );
  INVxp67_ASAP7_75t_SL U53303 ( .A(n65928), .Y(n65952) );
  INVxp33_ASAP7_75t_SL U53304 ( .A(n77101), .Y(n61109) );
  NAND2xp33_ASAP7_75t_SL U53305 ( .A(n66022), .B(n65934), .Y(n65801) );
  INVx1_ASAP7_75t_SL U53306 ( .A(n65920), .Y(n65977) );
  OAI22xp33_ASAP7_75t_SL U53307 ( .A1(n73217), .A2(n57185), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[4]), .B2(
        n73379), .Y(n73218) );
  INVxp67_ASAP7_75t_SL U53308 ( .A(n72912), .Y(n72788) );
  BUFx4f_ASAP7_75t_SL U53309 ( .A(n59507), .Y(n57110) );
  OAI22xp33_ASAP7_75t_SL U53310 ( .A1(n73009), .A2(n72830), .B1(n73008), .B2(
        n72915), .Y(n72834) );
  INVxp67_ASAP7_75t_SL U53311 ( .A(n71716), .Y(n71722) );
  AOI21x1_ASAP7_75t_SL U53312 ( .A1(n62645), .A2(n62646), .B(n58220), .Y(
        n59470) );
  OAI22xp33_ASAP7_75t_SL U53313 ( .A1(n73191), .A2(n57185), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[7]), .B2(
        n59525), .Y(n73192) );
  AOI22xp33_ASAP7_75t_SL U53314 ( .A1(n73030), .A2(n72915), .B1(n73028), .B2(
        n72935), .Y(n72774) );
  OAI22xp33_ASAP7_75t_SL U53315 ( .A1(n73227), .A2(n57185), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[1]), .B2(
        n59525), .Y(n73228) );
  INVxp67_ASAP7_75t_SL U53316 ( .A(n65921), .Y(n65707) );
  NAND2xp5_ASAP7_75t_SL U53317 ( .A(n76229), .B(n76228), .Y(n78139) );
  NAND2xp5_ASAP7_75t_SL U53318 ( .A(n75428), .B(n75429), .Y(n75445) );
  OAI21xp33_ASAP7_75t_SRAM U53319 ( .A1(or1200_cpu_or1200_except_n540), .A2(
        n76724), .B(n75687), .Y(n64816) );
  AOI21xp33_ASAP7_75t_SL U53320 ( .A1(n74193), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .B(n74752), .Y(
        n74182) );
  INVxp33_ASAP7_75t_SL U53321 ( .A(n63191), .Y(n63094) );
  NAND2xp33_ASAP7_75t_SL U53322 ( .A(n69355), .B(n75442), .Y(n78089) );
  AOI21xp33_ASAP7_75t_SL U53323 ( .A1(n74193), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]), .B(n74752), .Y(
        n74194) );
  O2A1O1Ixp5_ASAP7_75t_SL U53324 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .A2(n72319), .B(n71570), .C(n71569), .Y(n71571) );
  BUFx2_ASAP7_75t_SL U53325 ( .A(n75916), .Y(n59657) );
  XNOR2xp5_ASAP7_75t_SL U53326 ( .A(n59182), .B(n60762), .Y(n61400) );
  INVxp67_ASAP7_75t_SL U53327 ( .A(n60758), .Y(n60751) );
  INVx8_ASAP7_75t_SL U53328 ( .A(n59656), .Y(n57111) );
  OA21x2_ASAP7_75t_SL U53329 ( .A1(n74373), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_7_), 
        .B(n74372), .Y(n74374) );
  AOI21xp33_ASAP7_75t_SL U53330 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_17_), .A2(n70109), .B(
        n69475), .Y(n69499) );
  NOR2xp33_ASAP7_75t_SRAM U53331 ( .A(or1200_cpu_or1200_except_n500), .B(
        n76724), .Y(n62240) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U53332 ( .A1(n62604), .A2(n58206), .B(n61500), .C(
        n60967), .Y(n60968) );
  NAND2xp33_ASAP7_75t_SL U53333 ( .A(n73027), .B(n73029), .Y(n72940) );
  AOI21xp33_ASAP7_75t_SL U53334 ( .A1(n72131), .A2(n72389), .B(n72053), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n93) );
  AOI211xp5_ASAP7_75t_SRAM U53335 ( .A1(n68812), .A2(n69256), .B(n64277), .C(
        n64276), .Y(n64278) );
  NOR2xp33_ASAP7_75t_SRAM U53336 ( .A(or1200_cpu_or1200_except_n502), .B(
        n76724), .Y(n76725) );
  INVxp33_ASAP7_75t_SL U53337 ( .A(n71419), .Y(n71465) );
  AOI21xp33_ASAP7_75t_SL U53338 ( .A1(n76422), .A2(n76421), .B(n76469), .Y(
        n76424) );
  AOI21xp5_ASAP7_75t_SL U53339 ( .A1(n69859), .A2(n69864), .B(n69863), .Y(
        n69860) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U53340 ( .A1(n75735), .A2(n75595), .B(n75594), .C(
        n59547), .Y(n75596) );
  NAND2xp5_ASAP7_75t_SL U53341 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[23]), .B(
        n57185), .Y(n73351) );
  NAND2xp5_ASAP7_75t_SL U53342 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[22]), .B(
        n57185), .Y(n73347) );
  NAND2xp5_ASAP7_75t_SL U53343 ( .A(n73341), .B(n57185), .Y(n73342) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U53344 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), 
        .A2(n73025), .B(n72860), .C(n72999), .Y(n72861) );
  NAND2xp5_ASAP7_75t_SL U53345 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[21]), .B(
        n57185), .Y(n73326) );
  NAND2xp5_ASAP7_75t_SL U53346 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[12]), .B(
        n57185), .Y(n73273) );
  NAND2xp5_ASAP7_75t_SL U53347 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[20]), .B(
        n57185), .Y(n73323) );
  XNOR2xp5_ASAP7_75t_SL U53348 ( .A(n62762), .B(n61936), .Y(n76258) );
  NAND2xp33_ASAP7_75t_SL U53349 ( .A(or1200_cpu_sr_15_), .B(n77040), .Y(n77045) );
  NAND2xp5_ASAP7_75t_SL U53350 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[19]), .B(
        n57185), .Y(n73319) );
  AND2x2_ASAP7_75t_SL U53351 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[23]), .B(n71013), 
        .Y(n71354) );
  INVx1_ASAP7_75t_SL U53352 ( .A(n61938), .Y(n76259) );
  NAND2xp33_ASAP7_75t_SL U53353 ( .A(n59535), .B(n61940), .Y(n63546) );
  NAND2xp33_ASAP7_75t_SL U53354 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[13]), .B(
        n57185), .Y(n73277) );
  INVx1_ASAP7_75t_SL U53355 ( .A(n58058), .Y(n57554) );
  NAND2xp5_ASAP7_75t_SL U53356 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[17]), .B(
        n57185), .Y(n73298) );
  INVxp67_ASAP7_75t_SL U53357 ( .A(n72889), .Y(n72909) );
  NAND2xp5_ASAP7_75t_SL U53358 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[14]), .B(
        n57185), .Y(n73281) );
  BUFx3_ASAP7_75t_SL U53359 ( .A(n68005), .Y(n59503) );
  NAND2xp5_ASAP7_75t_SL U53360 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[16]), .B(
        n57185), .Y(n73293) );
  NAND2xp33_ASAP7_75t_SL U53361 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[15]), .B(
        n57185), .Y(n73286) );
  OAI22xp33_ASAP7_75t_SL U53362 ( .A1(n75316), .A2(n75314), .B1(n61369), .B2(
        n76796), .Y(n61370) );
  AOI22xp33_ASAP7_75t_SL U53363 ( .A1(n73030), .A2(n72830), .B1(n73028), .B2(
        n72915), .Y(n72821) );
  NAND2xp33_ASAP7_75t_SL U53364 ( .A(n58206), .B(n60741), .Y(n61672) );
  NAND2xp5_ASAP7_75t_SL U53365 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[25]), .B(
        n57185), .Y(n73392) );
  OAI22xp33_ASAP7_75t_SL U53366 ( .A1(n73161), .A2(n57185), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[10]), .B2(
        n73379), .Y(n73162) );
  INVxp67_ASAP7_75t_SL U53367 ( .A(n61410), .Y(n61413) );
  OAI21xp5_ASAP7_75t_SL U53368 ( .A1(n78353), .A2(n57190), .B(n72714), .Y(
        n72889) );
  INVxp67_ASAP7_75t_SL U53369 ( .A(n72891), .Y(n72913) );
  OAI22xp33_ASAP7_75t_SL U53370 ( .A1(n78354), .A2(n70035), .B1(n78356), .B2(
        n70034), .Y(n70037) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U53371 ( .A1(n57506), .A2(n61214), .B(n61213), 
        .C(n61521), .Y(n61220) );
  AOI22xp33_ASAP7_75t_SRAM U53372 ( .A1(n57424), .A2(n61215), .B1(n61630), 
        .B2(n62274), .Y(n61219) );
  NOR2xp33_ASAP7_75t_SRAM U53373 ( .A(or1200_cpu_or1200_mult_mac_n185), .B(
        n64275), .Y(n64276) );
  NOR2x1_ASAP7_75t_SL U53374 ( .A(n61226), .B(n75766), .Y(n77246) );
  INVxp67_ASAP7_75t_SL U53375 ( .A(n75865), .Y(n61439) );
  INVxp33_ASAP7_75t_SL U53376 ( .A(n64316), .Y(n64320) );
  AOI22xp33_ASAP7_75t_SL U53377 ( .A1(n75570), .A2(
        or1200_dc_top_from_dcram_20_), .B1(dwb_dat_i[20]), .B2(n75569), .Y(
        n64108) );
  NOR2xp33_ASAP7_75t_SL U53378 ( .A(n61810), .B(n78170), .Y(n75760) );
  INVx1_ASAP7_75t_SL U53379 ( .A(n70018), .Y(n69563) );
  INVxp67_ASAP7_75t_SL U53380 ( .A(n64136), .Y(n61448) );
  INVxp67_ASAP7_75t_SL U53381 ( .A(n63564), .Y(n61227) );
  NAND2xp5_ASAP7_75t_SL U53382 ( .A(or1200_dc_top_tag_0_), .B(n77293), .Y(
        n59727) );
  INVx1_ASAP7_75t_SL U53383 ( .A(n66162), .Y(n66105) );
  AOI21xp33_ASAP7_75t_SL U53384 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_), .A2(n57190), .B(n72618), 
        .Y(n72625) );
  AOI211xp5_ASAP7_75t_SRAM U53385 ( .A1(n69884), .A2(n69912), .B(n69891), .C(
        n69908), .Y(n69676) );
  NAND2xp5_ASAP7_75t_SL U53386 ( .A(n64775), .B(n64774), .Y(n64778) );
  AOI22xp33_ASAP7_75t_SRAM U53387 ( .A1(n76772), .A2(n58084), .B1(n61631), 
        .B2(n61630), .Y(n61632) );
  INVxp33_ASAP7_75t_SL U53388 ( .A(n77598), .Y(n61608) );
  INVxp33_ASAP7_75t_SL U53389 ( .A(n77610), .Y(n61369) );
  INVx1_ASAP7_75t_SL U53390 ( .A(n72893), .Y(n72911) );
  NAND2xp5_ASAP7_75t_SL U53391 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[0]), .B(n58291), 
        .Y(n70864) );
  OAI21xp5_ASAP7_75t_SL U53392 ( .A1(n78347), .A2(n57190), .B(n72764), .Y(
        n72912) );
  INVxp67_ASAP7_75t_SL U53393 ( .A(n76771), .Y(n76780) );
  OAI21xp5_ASAP7_75t_SL U53394 ( .A1(n71714), .A2(n71724), .B(n71654), .Y(
        n71716) );
  NAND2xp33_ASAP7_75t_SRAM U53395 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        n72203), .Y(n72204) );
  OAI22xp33_ASAP7_75t_SL U53396 ( .A1(n59708), .A2(n77056), .B1(n59709), .B2(
        n77089), .Y(n74608) );
  OAI21xp33_ASAP7_75t_SL U53397 ( .A1(or1200_cpu_or1200_mult_mac_n299), .A2(
        n75738), .B(n62261), .Y(n62272) );
  AOI21xp33_ASAP7_75t_SL U53398 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_27_), .A2(n57190), .B(n72668), 
        .Y(n72679) );
  INVxp67_ASAP7_75t_SL U53399 ( .A(n72923), .Y(n73025) );
  AOI21xp33_ASAP7_75t_SL U53400 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_29_), .A2(n57190), .B(n72647), 
        .Y(n72672) );
  INVxp33_ASAP7_75t_SL U53401 ( .A(n66637), .Y(n57183) );
  NOR2x1_ASAP7_75t_SL U53402 ( .A(n68810), .B(n77035), .Y(n74641) );
  NAND2xp5_ASAP7_75t_SL U53403 ( .A(n59984), .B(n60149), .Y(n60147) );
  NAND2xp33_ASAP7_75t_SL U53404 ( .A(n77713), .B(n61929), .Y(n61926) );
  NOR2x1p5_ASAP7_75t_SL U53405 ( .A(n68810), .B(n63254), .Y(n77287) );
  AOI21xp33_ASAP7_75t_SL U53406 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_), .A2(n57190), .B(n72653), 
        .Y(n72670) );
  INVx1_ASAP7_75t_SL U53407 ( .A(n66024), .Y(n65972) );
  INVx1_ASAP7_75t_SL U53408 ( .A(n77663), .Y(n59973) );
  INVxp67_ASAP7_75t_SL U53409 ( .A(n65929), .Y(n65951) );
  INVx1_ASAP7_75t_SL U53410 ( .A(n72966), .Y(n72900) );
  OAI21xp33_ASAP7_75t_SL U53411 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[38]), .A2(n58582), 
        .B(n65744), .Y(n65748) );
  INVx1_ASAP7_75t_SL U53412 ( .A(n72937), .Y(n72830) );
  AOI22xp33_ASAP7_75t_SL U53413 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_12_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_11_), .B2(n70018), .Y(
        n69422) );
  NOR2xp33_ASAP7_75t_SL U53414 ( .A(n62200), .B(n62199), .Y(n75387) );
  NAND2xp33_ASAP7_75t_SL U53415 ( .A(n65853), .B(n57187), .Y(n65746) );
  NAND2xp33_ASAP7_75t_SL U53416 ( .A(n78053), .B(n57189), .Y(n596) );
  NAND2xp33_ASAP7_75t_SL U53417 ( .A(n78043), .B(n57189), .Y(n636) );
  NAND2xp33_ASAP7_75t_SL U53418 ( .A(n78047), .B(n57189), .Y(n617) );
  NAND2xp33_ASAP7_75t_SL U53419 ( .A(n65743), .B(n57188), .Y(n65744) );
  AOI21xp33_ASAP7_75t_SL U53420 ( .A1(n63350), .A2(n63396), .B(n63394), .Y(
        n63351) );
  INVxp33_ASAP7_75t_SL U53421 ( .A(n72010), .Y(n71996) );
  NAND2xp5_ASAP7_75t_SL U53422 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_7_), .B(
        n74379), .Y(n74378) );
  OAI21xp33_ASAP7_75t_SL U53423 ( .A1(n72495), .A2(n72484), .B(n57192), .Y(
        n71987) );
  AOI22xp33_ASAP7_75t_SL U53424 ( .A1(n57194), .A2(n65804), .B1(n65853), .B2(
        n57188), .Y(n65706) );
  NAND2xp33_ASAP7_75t_SL U53425 ( .A(n78042), .B(n57189), .Y(n643) );
  NAND2xp33_ASAP7_75t_SL U53426 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[32]), .B(n57188), 
        .Y(n65713) );
  NAND2xp33_ASAP7_75t_SL U53427 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[33]), .B(n57187), 
        .Y(n65712) );
  NAND2xp33_ASAP7_75t_SL U53428 ( .A(n78045), .B(n57189), .Y(n626) );
  NAND2xp33_ASAP7_75t_SL U53429 ( .A(n72474), .B(n72421), .Y(n72152) );
  NAND2xp33_ASAP7_75t_SL U53430 ( .A(n78049), .B(n57189), .Y(n610) );
  NAND2xp33_ASAP7_75t_SL U53431 ( .A(n78051), .B(n57189), .Y(n603) );
  NAND2xp33_ASAP7_75t_SL U53432 ( .A(n72474), .B(n72404), .Y(n72405) );
  NAND2xp33_ASAP7_75t_SL U53433 ( .A(n78044), .B(n57189), .Y(n631) );
  NAND2xp33_ASAP7_75t_SL U53434 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[16]), .B(n57187), 
        .Y(n65755) );
  NAND2xp33_ASAP7_75t_SL U53435 ( .A(n78432), .B(n57190), .Y(n72724) );
  NAND2xp33_ASAP7_75t_SL U53436 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[15]), .B(n57188), 
        .Y(n65754) );
  NAND2xp5_ASAP7_75t_SL U53437 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_7_), .B(
        n71673), .Y(n71675) );
  NAND2xp5_ASAP7_75t_SL U53438 ( .A(n70049), .B(n70048), .Y(n70050) );
  NAND2xp33_ASAP7_75t_SL U53439 ( .A(n70092), .B(n70091), .Y(n70093) );
  INVxp67_ASAP7_75t_SL U53440 ( .A(n76759), .Y(n76762) );
  OAI22xp33_ASAP7_75t_SL U53441 ( .A1(n76765), .A2(n77100), .B1(n76764), .B2(
        n77102), .Y(n76784) );
  AOI21xp5_ASAP7_75t_SL U53442 ( .A1(n75736), .A2(n59443), .B(n60982), .Y(
        n60983) );
  NOR2xp33_ASAP7_75t_SL U53443 ( .A(n59709), .B(n64218), .Y(n75845) );
  AOI21xp33_ASAP7_75t_SL U53444 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[14]), .A2(n70502), .B(
        n70495), .Y(n69867) );
  NAND2xp33_ASAP7_75t_SL U53445 ( .A(n78064), .B(n57189), .Y(n572) );
  NAND2xp33_ASAP7_75t_SL U53446 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .B(n57187), 
        .Y(n65716) );
  NAND2xp33_ASAP7_75t_SL U53447 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]), .B(n57187), 
        .Y(n65740) );
  NAND2xp33_ASAP7_75t_SL U53448 ( .A(n78062), .B(n57189), .Y(n579) );
  OAI22xp33_ASAP7_75t_SL U53449 ( .A1(n75350), .A2(n75702), .B1(n76764), .B2(
        n75324), .Y(n62109) );
  NAND2xp33_ASAP7_75t_SL U53450 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[39]), .B(n57188), 
        .Y(n65739) );
  NAND2xp33_ASAP7_75t_SL U53451 ( .A(n78060), .B(n57189), .Y(n589) );
  NAND2xp5_ASAP7_75t_SL U53452 ( .A(n65383), .B(n65317), .Y(n65385) );
  NOR2xp33_ASAP7_75t_SL U53453 ( .A(n66081), .B(n66060), .Y(n66058) );
  INVxp33_ASAP7_75t_SL U53454 ( .A(n74290), .Y(n74291) );
  AOI22xp33_ASAP7_75t_SL U53455 ( .A1(n75220), .A2(n63485), .B1(n60811), .B2(
        n57191), .Y(n60812) );
  OAI21xp33_ASAP7_75t_SL U53456 ( .A1(n73942), .A2(n75702), .B(n61874), .Y(
        n61890) );
  OAI22xp33_ASAP7_75t_SL U53457 ( .A1(n75590), .A2(n76764), .B1(n75325), .B2(
        n77104), .Y(n61888) );
  INVx1_ASAP7_75t_SL U53458 ( .A(n63583), .Y(n64293) );
  NAND2xp33_ASAP7_75t_SL U53459 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[15]), .B(n57187), 
        .Y(n65838) );
  OAI22xp33_ASAP7_75t_SL U53460 ( .A1(n76764), .A2(n77104), .B1(n75702), .B2(
        n75586), .Y(n73924) );
  NAND2xp33_ASAP7_75t_SL U53461 ( .A(n65833), .B(n57188), .Y(n65834) );
  NAND2xp33_ASAP7_75t_SL U53462 ( .A(n78037), .B(n57189), .Y(n668) );
  NAND2xp33_ASAP7_75t_SL U53463 ( .A(n78028), .B(n57189), .Y(n713) );
  NAND2xp33_ASAP7_75t_SL U53464 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[11]), .B(n57190), .Y(n72764) );
  OAI21xp5_ASAP7_75t_SL U53465 ( .A1(n78351), .A2(n57190), .B(n72752), .Y(
        n72891) );
  INVxp33_ASAP7_75t_SL U53466 ( .A(n65317), .Y(n65384) );
  NAND2xp33_ASAP7_75t_SL U53467 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[10]), .B(n57188), 
        .Y(n65817) );
  NAND2xp33_ASAP7_75t_SL U53468 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]), .B(n57187), 
        .Y(n65779) );
  NAND2xp33_ASAP7_75t_SL U53469 ( .A(n78032), .B(n57189), .Y(n693) );
  NAND2xp33_ASAP7_75t_SL U53470 ( .A(n78038), .B(n57189), .Y(n663) );
  AOI22xp33_ASAP7_75t_SL U53471 ( .A1(n57193), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[7]), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[5]), .B2(n57187), 
        .Y(n65693) );
  AOI22xp33_ASAP7_75t_SL U53472 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[4]), .A2(n57194), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[2]), .B2(n57188), 
        .Y(n65813) );
  NAND2xp33_ASAP7_75t_SL U53473 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[25]), .B(n57188), 
        .Y(n65780) );
  AOI22xp33_ASAP7_75t_SL U53474 ( .A1(n57194), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[6]), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[4]), .B2(n57188), 
        .Y(n65692) );
  AOI22xp33_ASAP7_75t_SL U53475 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[5]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[3]), .B2(n57187), 
        .Y(n65814) );
  OAI21xp5_ASAP7_75t_SL U53476 ( .A1(n78349), .A2(n57190), .B(n72765), .Y(
        n72893) );
  INVx1_ASAP7_75t_SL U53477 ( .A(n70117), .Y(n70119) );
  NAND2xp33_ASAP7_75t_SL U53478 ( .A(n78034), .B(n57189), .Y(n683) );
  AOI21x1_ASAP7_75t_SL U53479 ( .A1(n69557), .A2(n78364), .B(n71512), .Y(
        n70104) );
  NAND2xp33_ASAP7_75t_SL U53480 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]), .B(n57188), 
        .Y(n65843) );
  NAND2xp33_ASAP7_75t_SL U53481 ( .A(n78035), .B(n57189), .Y(n678) );
  NAND2xp33_ASAP7_75t_SL U53482 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]), .B(n57187), 
        .Y(n65678) );
  NAND2xp33_ASAP7_75t_SL U53483 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[16]), .B(n57188), 
        .Y(n65677) );
  NAND2xp33_ASAP7_75t_SL U53484 ( .A(n78027), .B(n57189), .Y(n720) );
  AOI22xp33_ASAP7_75t_SL U53485 ( .A1(n76767), .A2(n64839), .B1(n76766), .B2(
        n75705), .Y(n64842) );
  NAND2xp5_ASAP7_75t_SL U53486 ( .A(n70124), .B(n69557), .Y(n70034) );
  NAND2xp33_ASAP7_75t_SL U53487 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .B(n57187), 
        .Y(n65844) );
  OR2x4_ASAP7_75t_SL U53488 ( .A(n63262), .B(n63266), .Y(n76906) );
  NAND2xp33_ASAP7_75t_SL U53489 ( .A(n78036), .B(n57189), .Y(n673) );
  NAND2xp33_ASAP7_75t_SL U53490 ( .A(n78026), .B(n57189), .Y(n727) );
  NAND2xp33_ASAP7_75t_SL U53491 ( .A(n78033), .B(n57189), .Y(n688) );
  INVxp67_ASAP7_75t_SL U53492 ( .A(n73552), .Y(n73546) );
  NAND2xp33_ASAP7_75t_SL U53493 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[14]), .B(n57188), 
        .Y(n65837) );
  NAND2xp33_ASAP7_75t_SL U53494 ( .A(n78162), .B(n57189), .Y(n235) );
  OAI21xp5_ASAP7_75t_SL U53495 ( .A1(n78367), .A2(n57190), .B(n72682), .Y(
        n72966) );
  NAND2xp33_ASAP7_75t_SL U53496 ( .A(n78040), .B(n57189), .Y(n653) );
  AOI21xp33_ASAP7_75t_SL U53497 ( .A1(n57122), .A2(n59443), .B(
        or1200_cpu_or1200_mult_mac_n62), .Y(n75918) );
  INVxp67_ASAP7_75t_SL U53498 ( .A(n77043), .Y(n75364) );
  NAND2xp33_ASAP7_75t_SL U53499 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[3]), .B(n57188), .Y(
        n65730) );
  NAND2xp33_ASAP7_75t_SL U53500 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[4]), .B(n57187), .Y(
        n65731) );
  NAND2xp33_ASAP7_75t_SL U53501 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[18]), .B(n57187), 
        .Y(n65773) );
  NAND2xp33_ASAP7_75t_SL U53502 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[1]), .B(n57187), .Y(
        n65695) );
  OAI21xp33_ASAP7_75t_SL U53503 ( .A1(n78333), .A2(n57190), .B(n72843), .Y(
        n72923) );
  AOI22xp33_ASAP7_75t_SL U53504 ( .A1(n57193), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[2]), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[0]), .B2(n57187), 
        .Y(n65733) );
  INVxp33_ASAP7_75t_SL U53505 ( .A(n67307), .Y(n67310) );
  NAND2xp33_ASAP7_75t_SL U53506 ( .A(n78029), .B(n57189), .Y(n708) );
  NAND2xp33_ASAP7_75t_SL U53507 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]), .B(n57190), .Y(n72714) );
  NAND2xp33_ASAP7_75t_SL U53508 ( .A(n78369), .B(n57190), .Y(n72688) );
  INVx1_ASAP7_75t_SL U53509 ( .A(n75860), .Y(n62525) );
  NAND2xp33_ASAP7_75t_SL U53510 ( .A(n78031), .B(n57189), .Y(n698) );
  NAND2xp33_ASAP7_75t_SL U53511 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[12]), .B(n57187), 
        .Y(n65726) );
  NAND2xp33_ASAP7_75t_SL U53512 ( .A(n78030), .B(n57189), .Y(n703) );
  NAND2xp33_ASAP7_75t_SL U53513 ( .A(n78041), .B(n57189), .Y(n648) );
  NAND2xp33_ASAP7_75t_SL U53514 ( .A(n69850), .B(n69858), .Y(n69659) );
  AOI21xp33_ASAP7_75t_SL U53515 ( .A1(n57191), .A2(n62365), .B(n62364), .Y(
        n62369) );
  NAND2xp33_ASAP7_75t_SL U53516 ( .A(n65832), .B(n57187), .Y(n65762) );
  NAND2xp33_ASAP7_75t_SL U53517 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[0]), .B(n57188), .Y(
        n65694) );
  NAND2xp33_ASAP7_75t_SL U53518 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[7]), .B(n57188), .Y(
        n65734) );
  NAND2xp33_ASAP7_75t_SL U53519 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]), .B(n57188), 
        .Y(n65772) );
  NAND2xp33_ASAP7_75t_SL U53520 ( .A(n77802), .B(n57189), .Y(n7192) );
  INVxp33_ASAP7_75t_SL U53521 ( .A(n70754), .Y(n70757) );
  OAI21xp5_ASAP7_75t_SL U53522 ( .A1(n78430), .A2(n57190), .B(n72710), .Y(
        n72904) );
  AND2x2_ASAP7_75t_SL U53523 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[19]), .B(n57190), .Y(n72697) );
  OAI21xp5_ASAP7_75t_SL U53524 ( .A1(n73806), .A2(n73770), .B(n73750), .Y(
        n3303) );
  NAND2xp33_ASAP7_75t_SL U53525 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[8]), .B(n57187), .Y(
        n65735) );
  OAI21xp5_ASAP7_75t_SL U53526 ( .A1(n73803), .A2(n73770), .B(n73735), .Y(
        n3304) );
  OAI21xp5_ASAP7_75t_SL U53527 ( .A1(n78355), .A2(n57190), .B(n72701), .Y(
        n72901) );
  NAND2xp33_ASAP7_75t_SL U53528 ( .A(n78039), .B(n57189), .Y(n658) );
  NAND2xp5_ASAP7_75t_SL U53529 ( .A(n57209), .B(n66271), .Y(n58209) );
  OAI22xp5_ASAP7_75t_SL U53530 ( .A1(n70448), .A2(n70447), .B1(n70446), .B2(
        n70471), .Y(n70449) );
  AOI21xp33_ASAP7_75t_SL U53531 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]), .A2(n57193), 
        .B(n65759), .Y(n65760) );
  NAND2xp33_ASAP7_75t_SL U53532 ( .A(n65725), .B(n57194), .Y(n65729) );
  INVx1_ASAP7_75t_SL U53533 ( .A(n77058), .Y(n57191) );
  INVxp67_ASAP7_75t_SL U53534 ( .A(n73555), .Y(n73575) );
  NOR2xp67_ASAP7_75t_SL U53535 ( .A(n75872), .B(n77058), .Y(n75727) );
  AOI22xp33_ASAP7_75t_SL U53536 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[6]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[5]), .B2(n57194), 
        .Y(n65732) );
  NOR2xp33_ASAP7_75t_SL U53537 ( .A(n62319), .B(n76716), .Y(n77043) );
  INVx2_ASAP7_75t_SL U53538 ( .A(n64026), .Y(n57116) );
  NAND2xp33_ASAP7_75t_SL U53539 ( .A(n57219), .B(n53455), .Y(n60742) );
  NAND2xp33_ASAP7_75t_SL U53540 ( .A(n57213), .B(n53455), .Y(n60733) );
  AOI21xp33_ASAP7_75t_SL U53541 ( .A1(n76996), .A2(n76615), .B(n76614), .Y(
        n76637) );
  NAND2x1_ASAP7_75t_SL U53542 ( .A(n60584), .B(n61999), .Y(n61546) );
  INVxp67_ASAP7_75t_SL U53543 ( .A(n75835), .Y(n64235) );
  OAI21xp5_ASAP7_75t_SL U53544 ( .A1(n73816), .A2(n73806), .B(n73805), .Y(
        n3295) );
  INVx1_ASAP7_75t_SL U53545 ( .A(n77097), .Y(n75734) );
  INVxp33_ASAP7_75t_SL U53546 ( .A(n71323), .Y(n71321) );
  INVxp33_ASAP7_75t_SL U53547 ( .A(n75233), .Y(n61631) );
  NAND2xp33_ASAP7_75t_SL U53548 ( .A(n77730), .B(n53455), .Y(n61967) );
  OAI21xp5_ASAP7_75t_SL U53549 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[4]), .A2(n73872), 
        .B(n73545), .Y(n73552) );
  NAND2xp33_ASAP7_75t_SL U53550 ( .A(n63300), .B(n76753), .Y(n61497) );
  INVxp67_ASAP7_75t_SL U53551 ( .A(n70641), .Y(n74272) );
  NAND2xp33_ASAP7_75t_SL U53552 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[14]), .B(n57194), 
        .Y(n65702) );
  NAND2xp33_ASAP7_75t_SL U53553 ( .A(n70118), .B(n70114), .Y(n69578) );
  AOI21xp5_ASAP7_75t_SL U53554 ( .A1(n74163), .A2(n74055), .B(n74164), .Y(
        n66219) );
  INVxp33_ASAP7_75t_SL U53555 ( .A(n65387), .Y(n65328) );
  AOI22xp33_ASAP7_75t_SL U53556 ( .A1(n65831), .A2(n57193), .B1(n65833), .B2(
        n57194), .Y(n65687) );
  INVxp33_ASAP7_75t_SL U53557 ( .A(n72467), .Y(n72191) );
  AOI21xp5_ASAP7_75t_SL U53558 ( .A1(n65666), .A2(n74169), .B(n74751), .Y(
        n65668) );
  NAND2xp5_ASAP7_75t_SL U53559 ( .A(n65816), .B(n65827), .Y(n66027) );
  AND2x2_ASAP7_75t_SL U53560 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[11]), .B(n57193), 
        .Y(n65699) );
  NOR2xp33_ASAP7_75t_SL U53561 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_4_), .B(n69751), .Y(
        n69758) );
  OAI22xp33_ASAP7_75t_SRAM U53562 ( .A1(n72355), .A2(n71819), .B1(n72085), 
        .B2(n71818), .Y(n71820) );
  INVx2_ASAP7_75t_SL U53563 ( .A(n58418), .Y(n57187) );
  INVx1_ASAP7_75t_SL U53564 ( .A(n58571), .Y(n57188) );
  AOI211xp5_ASAP7_75t_SL U53565 ( .A1(n72072), .A2(n72105), .B(n72071), .C(
        n72070), .Y(n72074) );
  NAND2xp5_ASAP7_75t_SL U53566 ( .A(n57211), .B(n71413), .Y(n71186) );
  AOI22xp33_ASAP7_75t_SL U53567 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[10]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[9]), .B2(n57194), 
        .Y(n65736) );
  INVxp33_ASAP7_75t_SL U53568 ( .A(n65625), .Y(n65597) );
  NAND2xp33_ASAP7_75t_SL U53569 ( .A(n65832), .B(n57194), .Y(n65835) );
  INVx1_ASAP7_75t_SL U53570 ( .A(n72278), .Y(n72474) );
  INVxp67_ASAP7_75t_SL U53571 ( .A(n70145), .Y(n70151) );
  NAND2xp5_ASAP7_75t_SL U53572 ( .A(n59983), .B(n60142), .Y(n60140) );
  NAND2xp5_ASAP7_75t_SL U53573 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_5_), 
        .B(n74333), .Y(n74345) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U53574 ( .A1(n61774), .A2(n76253), .B(n75783), 
        .C(n61773), .Y(n61779) );
  AOI22xp33_ASAP7_75t_SL U53575 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .B2(n57194), .Y(n65774) );
  OAI22xp33_ASAP7_75t_SL U53576 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]), .A2(n58418), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .B2(n58571), .Y(n65776) );
  OAI21xp33_ASAP7_75t_SL U53577 ( .A1(n72064), .A2(n72147), .B(n72063), .Y(
        n72282) );
  BUFx6f_ASAP7_75t_SL U53578 ( .A(n59589), .Y(n57117) );
  O2A1O1Ixp5_ASAP7_75t_SL U53579 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]), .B(n65423), 
        .C(n65422), .Y(n65427) );
  NAND2xp5_ASAP7_75t_SL U53580 ( .A(n60635), .B(n76782), .Y(n61531) );
  NOR2xp33_ASAP7_75t_SL U53581 ( .A(n71637), .B(n71694), .Y(n71673) );
  INVxp33_ASAP7_75t_SL U53582 ( .A(n76469), .Y(n76419) );
  NAND2xp33_ASAP7_75t_SL U53583 ( .A(n57214), .B(n62362), .Y(n60846) );
  BUFx4f_ASAP7_75t_SL U53584 ( .A(n59588), .Y(n57118) );
  INVx3_ASAP7_75t_SL U53585 ( .A(n66256), .Y(n57119) );
  NOR2xp33_ASAP7_75t_SRAM U53586 ( .A(n1424), .B(n60897), .Y(n60555) );
  NAND2xp5_ASAP7_75t_SL U53587 ( .A(n62433), .B(n76782), .Y(n76779) );
  INVx1_ASAP7_75t_SL U53588 ( .A(n59629), .Y(n59626) );
  AOI21xp33_ASAP7_75t_SRAM U53589 ( .A1(n74603), .A2(n78003), .B(n64290), .Y(
        n64291) );
  AOI22xp33_ASAP7_75t_SL U53590 ( .A1(n75689), .A2(n1119), .B1(
        or1200_cpu_or1200_mult_mac_n267), .B2(n75823), .Y(n61846) );
  NOR2xp33_ASAP7_75t_SL U53591 ( .A(n62319), .B(n61599), .Y(n74582) );
  INVx1_ASAP7_75t_SL U53592 ( .A(n70135), .Y(n69899) );
  INVxp67_ASAP7_75t_SL U53593 ( .A(n75722), .Y(n74603) );
  NOR2xp33_ASAP7_75t_SL U53594 ( .A(n72147), .B(n72086), .Y(n72004) );
  AOI21xp33_ASAP7_75t_SL U53595 ( .A1(n72109), .A2(n72116), .B(n57192), .Y(
        n71880) );
  NOR2x1_ASAP7_75t_SL U53596 ( .A(n71512), .B(n69766), .Y(n70124) );
  INVxp67_ASAP7_75t_SL U53597 ( .A(n75723), .Y(n73921) );
  NOR2x1p5_ASAP7_75t_SL U53598 ( .A(n57218), .B(n61918), .Y(n66451) );
  NAND2xp5_ASAP7_75t_SL U53599 ( .A(n65350), .B(n65349), .Y(n65351) );
  NAND2xp5_ASAP7_75t_SL U53600 ( .A(n60834), .B(n60819), .Y(n76716) );
  AOI21xp5_ASAP7_75t_SL U53601 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_48_), .A2(n70103), 
        .B(n69705), .Y(n70068) );
  O2A1O1Ixp5_ASAP7_75t_SL U53602 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[4]), 
        .A2(n73888), .B(n73879), .C(n73878), .Y(n73880) );
  OAI21xp33_ASAP7_75t_SL U53603 ( .A1(n72441), .A2(n72422), .B(n57192), .Y(
        n72423) );
  NAND2xp33_ASAP7_75t_SL U53604 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_41_), .B(n59523), 
        .Y(n71291) );
  OAI22xp33_ASAP7_75t_SL U53605 ( .A1(n72085), .A2(n72084), .B1(n72112), .B2(
        n72083), .Y(n72089) );
  NOR2xp33_ASAP7_75t_SL U53606 ( .A(n61289), .B(n60582), .Y(n60584) );
  AOI22xp33_ASAP7_75t_SL U53607 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_15_), .A2(
        n70476), .B1(n70485), .B2(n70354), .Y(n70340) );
  OAI22xp33_ASAP7_75t_SL U53608 ( .A1(n72434), .A2(n72418), .B1(n72465), .B2(
        n59623), .Y(n72419) );
  OAI22xp33_ASAP7_75t_SL U53609 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[24]), .A2(n58582), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .B2(n58419), .Y(n65775) );
  INVx2_ASAP7_75t_SL U53610 ( .A(n71353), .Y(n71413) );
  NAND2xp5_ASAP7_75t_SL U53611 ( .A(n75453), .B(n60819), .Y(n61599) );
  NAND2xp5_ASAP7_75t_SL U53612 ( .A(n62205), .B(n61242), .Y(n77621) );
  NAND2xp5_ASAP7_75t_SL U53613 ( .A(n75507), .B(n57504), .Y(n64858) );
  OAI21xp5_ASAP7_75t_SL U53614 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]), .A2(n74145), .B(
        n74153), .Y(n74150) );
  OAI21xp33_ASAP7_75t_SL U53615 ( .A1(n3036), .A2(n74953), .B(n74952), .Y(
        n74960) );
  AOI22xp33_ASAP7_75t_SL U53616 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_6_), .A2(
        n70476), .B1(n70485), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_5_), .Y(
        n70428) );
  NAND2xp5_ASAP7_75t_SL U53617 ( .A(n76942), .B(n76949), .Y(n76954) );
  AOI22xp33_ASAP7_75t_SL U53618 ( .A1(n72095), .A2(n71992), .B1(n72093), .B2(
        n72072), .Y(n71998) );
  NAND2xp33_ASAP7_75t_SL U53619 ( .A(n60560), .B(n76711), .Y(n60561) );
  NAND2xp5_ASAP7_75t_SL U53620 ( .A(n65327), .B(n65326), .Y(n65387) );
  OAI21xp33_ASAP7_75t_SL U53621 ( .A1(n72355), .A2(n72146), .B(n71938), .Y(
        n72467) );
  OAI21xp33_ASAP7_75t_SL U53622 ( .A1(n69724), .A2(n70103), .B(n69593), .Y(
        n69730) );
  AOI21xp33_ASAP7_75t_SL U53623 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_38_), .A2(n70103), 
        .B(n69639), .Y(n69853) );
  OAI31xp33_ASAP7_75t_SL U53624 ( .A1(n76985), .A2(n1502), .A3(n76984), .B(
        n2944), .Y(n76986) );
  AOI21xp33_ASAP7_75t_SL U53625 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_39_), .A2(n70103), 
        .B(n69645), .Y(n69866) );
  OR2x2_ASAP7_75t_SL U53626 ( .A(n57195), .B(n75915), .Y(n62575) );
  INVx1_ASAP7_75t_SL U53627 ( .A(n58419), .Y(n57194) );
  O2A1O1Ixp5_ASAP7_75t_SL U53628 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .A2(n65684), 
        .B(n65681), .C(n65660), .Y(n65453) );
  OAI21xp5_ASAP7_75t_SL U53629 ( .A1(n76449), .A2(n75735), .B(n75335), .Y(
        n75336) );
  AOI22xp33_ASAP7_75t_SL U53630 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .A2(
        n70476), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_12_), .B2(
        n70485), .Y(n70358) );
  INVx1_ASAP7_75t_SL U53631 ( .A(n58582), .Y(n57193) );
  INVxp33_ASAP7_75t_SL U53632 ( .A(n72044), .Y(n71819) );
  NAND2xp5_ASAP7_75t_SL U53633 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_49_), .B(n70103), 
        .Y(n69712) );
  INVxp33_ASAP7_75t_SL U53634 ( .A(n76378), .Y(n76379) );
  INVxp33_ASAP7_75t_SL U53635 ( .A(n74798), .Y(n76409) );
  NOR2xp67_ASAP7_75t_SL U53636 ( .A(n77994), .B(n60552), .Y(n61242) );
  NAND2xp5_ASAP7_75t_SL U53637 ( .A(n59494), .B(n76821), .Y(n77370) );
  INVx1_ASAP7_75t_SL U53638 ( .A(n77257), .Y(n74953) );
  NOR2xp33_ASAP7_75t_SRAM U53639 ( .A(n59574), .B(n57196), .Y(n60636) );
  NOR2xp33_ASAP7_75t_SRAM U53640 ( .A(n59559), .B(n57196), .Y(n61434) );
  NOR2xp33_ASAP7_75t_SL U53641 ( .A(n60842), .B(n62333), .Y(n61772) );
  AOI21xp33_ASAP7_75t_SL U53642 ( .A1(n2761), .A2(n77793), .B(n60276), .Y(
        n9482) );
  NAND2xp5_ASAP7_75t_SL U53643 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]), .B(n74145), .Y(
        n74153) );
  NAND2xp33_ASAP7_75t_SL U53644 ( .A(n64780), .B(n57197), .Y(n64782) );
  NAND2xp33_ASAP7_75t_SL U53645 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_27_), .B(n70103), 
        .Y(n69591) );
  NAND2xp5_ASAP7_75t_SL U53646 ( .A(n60799), .B(n61855), .Y(n75863) );
  NAND2xp33_ASAP7_75t_SL U53647 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_28_), .B(n70103), 
        .Y(n69593) );
  NOR2xp33_ASAP7_75t_SRAM U53648 ( .A(n59538), .B(n59584), .Y(n60796) );
  NOR2xp33_ASAP7_75t_SRAM U53649 ( .A(n59560), .B(n57196), .Y(n60797) );
  NAND2xp33_ASAP7_75t_SL U53650 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_34_), .B(n70103), 
        .Y(n69616) );
  NAND2xp33_ASAP7_75t_SL U53651 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_32_), .B(n70103), 
        .Y(n69612) );
  NAND2xp5_ASAP7_75t_SL U53652 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_47_), .B(n70103), 
        .Y(n69703) );
  NOR2xp33_ASAP7_75t_SRAM U53653 ( .A(n73976), .B(n76351), .Y(n73978) );
  INVxp67_ASAP7_75t_SL U53654 ( .A(n62419), .Y(n76711) );
  AOI21xp33_ASAP7_75t_SL U53655 ( .A1(n63743), .A2(n77880), .B(n60150), .Y(
        n60151) );
  NAND2xp5_ASAP7_75t_SL U53656 ( .A(n77850), .B(n61131), .Y(n68810) );
  INVxp67_ASAP7_75t_SL U53657 ( .A(n76764), .Y(n64840) );
  INVx1_ASAP7_75t_SL U53658 ( .A(n75876), .Y(n75602) );
  INVxp67_ASAP7_75t_SL U53659 ( .A(n70429), .Y(n70430) );
  INVxp33_ASAP7_75t_SL U53660 ( .A(n75326), .Y(n61357) );
  NAND2xp5_ASAP7_75t_SL U53661 ( .A(n75579), .B(n53430), .Y(n61820) );
  AOI22xp33_ASAP7_75t_SL U53662 ( .A1(n57198), .A2(n64758), .B1(n77871), .B2(
        n63743), .Y(n60037) );
  NOR2xp33_ASAP7_75t_SRAM U53663 ( .A(n59579), .B(n59584), .Y(n60858) );
  AOI22xp33_ASAP7_75t_SL U53664 ( .A1(n57198), .A2(n61165), .B1(n77980), .B2(
        n63743), .Y(n61166) );
  INVx1_ASAP7_75t_SL U53665 ( .A(n65830), .Y(n65841) );
  OR3x1_ASAP7_75t_SL U53666 ( .A(n74780), .B(n2410), .C(n74771), .Y(n74772) );
  INVx1_ASAP7_75t_SL U53667 ( .A(n75862), .Y(n64769) );
  AOI22xp33_ASAP7_75t_SL U53668 ( .A1(n75475), .A2(n75531), .B1(n75474), .B2(
        n57198), .Y(n75530) );
  NAND2xp5_ASAP7_75t_SL U53669 ( .A(n70686), .B(n70695), .Y(n71353) );
  NOR2xp33_ASAP7_75t_SL U53670 ( .A(n72321), .B(n72320), .Y(n72506) );
  OAI21xp5_ASAP7_75t_SL U53671 ( .A1(n69191), .A2(n69190), .B(n69189), .Y(
        n69192) );
  AOI22xp33_ASAP7_75t_SL U53672 ( .A1(n57198), .A2(n63731), .B1(n78002), .B2(
        n77253), .Y(n63732) );
  NAND2xp33_ASAP7_75t_SL U53673 ( .A(n72286), .B(n72045), .Y(n72222) );
  INVxp67_ASAP7_75t_SL U53674 ( .A(n71747), .Y(n71743) );
  OAI22xp33_ASAP7_75t_SL U53675 ( .A1(n72146), .A2(n72112), .B1(n72085), .B2(
        n72064), .Y(n71991) );
  INVxp33_ASAP7_75t_SL U53676 ( .A(n76765), .Y(n64771) );
  NAND2xp5_ASAP7_75t_SL U53677 ( .A(n70686), .B(n70695), .Y(n59523) );
  INVxp67_ASAP7_75t_SL U53678 ( .A(n72069), .Y(n71765) );
  NAND2xp5_ASAP7_75t_SL U53679 ( .A(n59990), .B(n59991), .Y(n76821) );
  NAND2xp33_ASAP7_75t_SL U53680 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), .B(n65621), 
        .Y(n65623) );
  NAND2xp33_ASAP7_75t_SL U53681 ( .A(n66181), .B(n65636), .Y(n66161) );
  INVxp67_ASAP7_75t_SL U53682 ( .A(n73070), .Y(n73073) );
  OAI21xp5_ASAP7_75t_SL U53683 ( .A1(n74447), .A2(n57202), .B(n74446), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N102) );
  AOI22xp33_ASAP7_75t_SL U53684 ( .A1(or1200_cpu_or1200_except_n494), .A2(
        n77082), .B1(or1200_cpu_or1200_fpu_result_arith[3]), .B2(n77091), .Y(
        n61555) );
  NAND2xp33_ASAP7_75t_SL U53685 ( .A(n74026), .B(n76416), .Y(n74023) );
  NOR2xp33_ASAP7_75t_SL U53686 ( .A(n57640), .B(n57639), .Y(n59127) );
  OAI21xp5_ASAP7_75t_SL U53687 ( .A1(n74440), .A2(n57202), .B(n74439), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N101) );
  OAI21xp33_ASAP7_75t_SL U53688 ( .A1(n58422), .A2(n72317), .B(n71844), .Y(
        n71845) );
  OAI21xp5_ASAP7_75t_SL U53689 ( .A1(n74398), .A2(n57202), .B(n74397), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N95) );
  NAND2xp5_ASAP7_75t_SL U53690 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_6_), .B(n74846), 
        .Y(n76950) );
  NAND2xp5_ASAP7_75t_SL U53691 ( .A(n57407), .B(n60645), .Y(n77066) );
  OAI21xp5_ASAP7_75t_SL U53692 ( .A1(n74389), .A2(n57202), .B(n74388), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N94) );
  OAI21xp5_ASAP7_75t_SL U53693 ( .A1(n74382), .A2(n57202), .B(n74381), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N87) );
  AOI22xp33_ASAP7_75t_SL U53694 ( .A1(or1200_cpu_or1200_fpu_result_arith[15]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[15]), 
        .Y(n77092) );
  INVxp33_ASAP7_75t_SL U53695 ( .A(n72582), .Y(n72562) );
  INVxp67_ASAP7_75t_SL U53696 ( .A(n61134), .Y(n61135) );
  AND2x2_ASAP7_75t_SL U53697 ( .A(n71768), .B(n72502), .Y(n58599) );
  NAND3xp33_ASAP7_75t_SL U53698 ( .A(n69276), .B(n69284), .C(n69275), .Y(
        n69289) );
  AOI22xp5_ASAP7_75t_SL U53699 ( .A1(n65205), .A2(n75541), .B1(n65204), .B2(
        n65203), .Y(n65206) );
  NAND2xp33_ASAP7_75t_SL U53700 ( .A(n71229), .B(n71315), .Y(n70758) );
  OAI21xp5_ASAP7_75t_SL U53701 ( .A1(n74412), .A2(n57202), .B(n74411), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N97) );
  NOR2xp33_ASAP7_75t_SL U53702 ( .A(n60669), .B(n60622), .Y(n60799) );
  OAI21xp5_ASAP7_75t_SL U53703 ( .A1(n74407), .A2(n57202), .B(n74406), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N96) );
  INVxp67_ASAP7_75t_SL U53704 ( .A(n71648), .Y(n71649) );
  AOI22xp5_ASAP7_75t_SL U53705 ( .A1(or1200_cpu_or1200_fpu_result_arith[0]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[0]), 
        .Y(n60693) );
  AOI22xp33_ASAP7_75t_SL U53706 ( .A1(or1200_cpu_or1200_fpu_result_arith[28]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[28]), 
        .Y(n75870) );
  AOI22xp33_ASAP7_75t_SL U53707 ( .A1(n77082), .A2(n61452), .B1(
        or1200_cpu_or1200_fpu_result_arith[4]), .B2(n77091), .Y(n61454) );
  OAI21xp5_ASAP7_75t_SL U53708 ( .A1(n74429), .A2(n57202), .B(n74428), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N100) );
  INVx1_ASAP7_75t_SL U53709 ( .A(n74136), .Y(n74143) );
  INVxp67_ASAP7_75t_SL U53710 ( .A(n65483), .Y(n65482) );
  AOI22xp33_ASAP7_75t_SL U53711 ( .A1(or1200_cpu_or1200_fpu_result_arith[29]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[29]), 
        .Y(n75215) );
  NAND2xp5_ASAP7_75t_SL U53712 ( .A(n64209), .B(n77623), .Y(n62418) );
  AOI22xp33_ASAP7_75t_SL U53713 ( .A1(or1200_cpu_or1200_fpu_result_conv[17]), 
        .A2(n77090), .B1(n77091), .B2(or1200_cpu_or1200_fpu_result_arith[17]), 
        .Y(n75335) );
  NAND2xp5_ASAP7_75t_SL U53714 ( .A(n65348), .B(n65391), .Y(n65347) );
  OAI21xp5_ASAP7_75t_SL U53715 ( .A1(n74421), .A2(n57202), .B(n74420), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N99) );
  AOI22xp33_ASAP7_75t_SL U53716 ( .A1(or1200_cpu_or1200_fpu_result_arith[7]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[7]), 
        .Y(n76793) );
  INVxp67_ASAP7_75t_SL U53717 ( .A(n74132), .Y(n74156) );
  OAI21xp5_ASAP7_75t_SL U53718 ( .A1(n74367), .A2(n57202), .B(n74366), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N88) );
  INVx1_ASAP7_75t_SL U53719 ( .A(n71728), .Y(n71792) );
  NAND2xp33_ASAP7_75t_SL U53720 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .B(n71315), .Y(
        n71317) );
  NAND2xp33_ASAP7_75t_SRAM U53721 ( .A(n73613), .B(n73612), .Y(n73615) );
  OAI21xp5_ASAP7_75t_SL U53722 ( .A1(n74229), .A2(n57202), .B(n74228), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N103) );
  OAI21xp33_ASAP7_75t_SL U53723 ( .A1(n57208), .A2(n72348), .B(n71836), .Y(
        n71837) );
  NOR2x1_ASAP7_75t_SL U53724 ( .A(n60554), .B(n64208), .Y(n75687) );
  INVxp33_ASAP7_75t_SRAM U53725 ( .A(n76405), .Y(n76408) );
  OAI21xp5_ASAP7_75t_SL U53726 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_ine), .A2(n57202), .B(
        n74743), .Y(n1561) );
  OAI21xp5_ASAP7_75t_SL U53727 ( .A1(n74456), .A2(n57202), .B(n74455), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N104) );
  NOR2xp33_ASAP7_75t_SRAM U53728 ( .A(n76394), .B(n76399), .Y(n76402) );
  AOI22xp33_ASAP7_75t_SL U53729 ( .A1(or1200_cpu_or1200_fpu_result_arith[1]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[1]), 
        .Y(n60981) );
  AOI22xp33_ASAP7_75t_SL U53730 ( .A1(or1200_cpu_or1200_fpu_result_arith[9]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[9]), 
        .Y(n61363) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U53731 ( .A1(n2561), .A2(n61056), .B(n61055), .C(
        n61058), .Y(n61057) );
  OAI21xp5_ASAP7_75t_SL U53732 ( .A1(n59871), .A2(n75193), .B(n59870), .Y(
        n59872) );
  AOI22xp33_ASAP7_75t_SL U53733 ( .A1(or1200_cpu_or1200_fpu_result_arith[24]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[24]), 
        .Y(n64786) );
  AOI22xp33_ASAP7_75t_SL U53734 ( .A1(or1200_cpu_or1200_fpu_result_arith[22]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[22]), 
        .Y(n64288) );
  NAND3xp33_ASAP7_75t_SL U53735 ( .A(n74757), .B(n74759), .C(n75455), .Y(n1537) );
  NAND2xp5_ASAP7_75t_SL U53736 ( .A(n77757), .B(n77125), .Y(n61628) );
  OAI21xp5_ASAP7_75t_SL U53737 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[26]), .A2(n57202), 
        .B(n73902), .Y(n1576) );
  INVxp33_ASAP7_75t_SL U53738 ( .A(n74708), .Y(n74709) );
  OAI21xp5_ASAP7_75t_SL U53739 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[30]), .A2(n57202), 
        .B(n74283), .Y(n1539) );
  INVxp33_ASAP7_75t_SRAM U53740 ( .A(n76367), .Y(n76371) );
  NAND2xp33_ASAP7_75t_SL U53741 ( .A(n61289), .B(n78166), .Y(n59879) );
  AOI22xp33_ASAP7_75t_SL U53742 ( .A1(or1200_cpu_or1200_fpu_result_arith[25]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[25]), 
        .Y(n64238) );
  OAI21xp5_ASAP7_75t_SL U53743 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[25]), .A2(n57202), 
        .B(n74107), .Y(n1593) );
  INVx2_ASAP7_75t_SL U53744 ( .A(n77623), .Y(n62319) );
  NAND2xp33_ASAP7_75t_SL U53745 ( .A(n57208), .B(n71895), .Y(n71897) );
  OAI21xp33_ASAP7_75t_SL U53746 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_), 
        .A2(n57203), .B(n72363), .Y(n72504) );
  OAI21xp33_ASAP7_75t_SL U53747 ( .A1(n72219), .A2(n57208), .B(n71808), .Y(
        n71809) );
  AOI22xp33_ASAP7_75t_SL U53748 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[3]), .A2(n57204), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[2]), .B2(n59632), .Y(
        n73740) );
  OAI21xp33_ASAP7_75t_SL U53749 ( .A1(n58423), .A2(n73739), .B(n3309), .Y(
        n73742) );
  NAND2xp33_ASAP7_75t_SL U53750 ( .A(n72079), .B(n57207), .Y(n71759) );
  AOI22xp33_ASAP7_75t_SL U53751 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_), 
        .A2(n57216), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_), 
        .B2(n57207), .Y(n71804) );
  AOI22xp33_ASAP7_75t_SL U53752 ( .A1(n57216), .A2(n72351), .B1(n72350), .B2(
        n57207), .Y(n71833) );
  NOR2xp33_ASAP7_75t_SL U53753 ( .A(n59703), .B(n60041), .Y(n76822) );
  AOI22xp33_ASAP7_75t_SL U53754 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_), 
        .A2(n57207), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_), 
        .B2(n71888), .Y(n71817) );
  NAND2xp5_ASAP7_75t_SL U53755 ( .A(n66179), .B(n66186), .Y(n74136) );
  AOI22xp33_ASAP7_75t_SL U53756 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_), 
        .A2(n57216), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_), 
        .B2(n57207), .Y(n71774) );
  AOI22xp33_ASAP7_75t_SL U53757 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[3]), .A2(n57205), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[1]), .B2(n59632), .Y(
        n73756) );
  OAI22xp33_ASAP7_75t_SL U53758 ( .A1(n72163), .A2(n57208), .B1(n72197), .B2(
        n71890), .Y(n71815) );
  NAND2xp5_ASAP7_75t_SL U53759 ( .A(n60572), .B(n60573), .Y(n59936) );
  OAI21xp33_ASAP7_75t_SL U53760 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_24_), 
        .A2(n57208), .B(n71847), .Y(n71848) );
  NAND2xp33_ASAP7_75t_SL U53761 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_), 
        .B(n57207), .Y(n71844) );
  INVxp67_ASAP7_75t_SL U53762 ( .A(n70132), .Y(n70136) );
  NAND2xp5_ASAP7_75t_SL U53763 ( .A(n72005), .B(n71542), .Y(n71584) );
  AOI22xp33_ASAP7_75t_SL U53764 ( .A1(n72262), .A2(n57207), .B1(n72346), .B2(
        n71888), .Y(n71771) );
  NAND2xp33_ASAP7_75t_SL U53765 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_2_), 
        .B(n57207), .Y(n71870) );
  NAND2xp33_ASAP7_75t_SL U53766 ( .A(n59255), .B(n61911), .Y(n59265) );
  AOI22xp33_ASAP7_75t_SL U53767 ( .A1(n70666), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[1]), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[9]), .B2(n70665), 
        .Y(n70671) );
  AOI22xp33_ASAP7_75t_SL U53768 ( .A1(n70666), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[0]), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[8]), .B2(n70665), 
        .Y(n70664) );
  OAI22xp33_ASAP7_75t_SL U53769 ( .A1(n72250), .A2(n57208), .B1(n71869), .B2(
        n71890), .Y(n71872) );
  AOI22xp33_ASAP7_75t_SL U53770 ( .A1(n70666), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[2]), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[10]), .B2(n70665), 
        .Y(n70659) );
  OAI21xp33_ASAP7_75t_SL U53771 ( .A1(n70654), .A2(n70653), .B(n71229), .Y(
        n70655) );
  O2A1O1Ixp5_ASAP7_75t_SL U53772 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_), 
        .A2(n71607), .B(n71863), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_), 
        .Y(n71608) );
  NOR2xp33_ASAP7_75t_SL U53773 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .B(
        n59622), .Y(n72490) );
  AOI22xp33_ASAP7_75t_SL U53774 ( .A1(n57216), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_), 
        .B2(n57207), .Y(n71879) );
  INVxp67_ASAP7_75t_SL U53775 ( .A(n65322), .Y(n65357) );
  NAND2xp33_ASAP7_75t_SL U53776 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_), 
        .B(n57207), .Y(n71753) );
  NAND2xp33_ASAP7_75t_SL U53777 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .B(n57207), .Y(n71836) );
  INVx1_ASAP7_75t_SL U53778 ( .A(n71438), .Y(n71460) );
  OAI22xp33_ASAP7_75t_SL U53779 ( .A1(n72317), .A2(n57208), .B1(n72310), .B2(
        n71890), .Y(n71752) );
  NAND2xp33_ASAP7_75t_SL U53780 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_), 
        .B(n57207), .Y(n71750) );
  NAND2xp5_ASAP7_75t_SL U53781 ( .A(n2616), .B(n60720), .Y(n60502) );
  NAND2xp33_ASAP7_75t_SL U53782 ( .A(n72080), .B(n57207), .Y(n71857) );
  NAND2xp33_ASAP7_75t_SL U53783 ( .A(n72351), .B(n72364), .Y(n72352) );
  INVx1_ASAP7_75t_SL U53784 ( .A(n59493), .Y(n64209) );
  AOI21xp33_ASAP7_75t_SL U53785 ( .A1(n70646), .A2(n71314), .B(n70666), .Y(
        n70647) );
  NAND2x1_ASAP7_75t_SL U53786 ( .A(n59876), .B(n77773), .Y(n78166) );
  INVxp33_ASAP7_75t_SL U53787 ( .A(n73923), .Y(n73927) );
  AOI21xp33_ASAP7_75t_SL U53788 ( .A1(n70646), .A2(n71229), .B(n59522), .Y(
        n70645) );
  INVxp33_ASAP7_75t_SRAM U53789 ( .A(n74018), .Y(n73918) );
  INVx1_ASAP7_75t_SL U53790 ( .A(n68884), .Y(n68881) );
  NOR2xp33_ASAP7_75t_SRAM U53791 ( .A(n73968), .B(n73990), .Y(n76377) );
  NAND2xp33_ASAP7_75t_SL U53792 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[22]), .B(n57205), .Y(
        n73716) );
  AOI22xp33_ASAP7_75t_SL U53793 ( .A1(n73708), .A2(n57204), .B1(n73680), .B2(
        n59632), .Y(n73637) );
  AOI21xp33_ASAP7_75t_SL U53794 ( .A1(n68823), .A2(n75008), .B(n68822), .Y(
        n68824) );
  AOI22xp33_ASAP7_75t_SL U53795 ( .A1(n73680), .A2(n57204), .B1(n59632), .B2(
        n73828), .Y(n73624) );
  AOI22xp33_ASAP7_75t_SL U53796 ( .A1(n3331), .A2(n57217), .B1(n73708), .B2(
        n57205), .Y(n73625) );
  INVxp33_ASAP7_75t_SL U53797 ( .A(n66181), .Y(n65621) );
  INVxp67_ASAP7_75t_SL U53798 ( .A(n75672), .Y(n59749) );
  NOR2xp33_ASAP7_75t_SL U53799 ( .A(n74093), .B(n66146), .Y(n65483) );
  AOI21xp5_ASAP7_75t_SL U53800 ( .A1(n59854), .A2(n59817), .B(n59793), .Y(
        n59796) );
  NOR2xp33_ASAP7_75t_SRAM U53801 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[14]), .B(
        n73379), .Y(n73138) );
  NAND2xp5_ASAP7_75t_SL U53802 ( .A(n59865), .B(n59869), .Y(n75195) );
  NAND2xp33_ASAP7_75t_SL U53803 ( .A(n74121), .B(n59854), .Y(n59857) );
  AOI21xp33_ASAP7_75t_SL U53804 ( .A1(n69169), .A2(n69168), .B(n69167), .Y(
        n69178) );
  NAND2xp5_ASAP7_75t_SL U53805 ( .A(n76639), .B(n76636), .Y(n76696) );
  NAND2xp33_ASAP7_75t_SL U53806 ( .A(n63125), .B(n57753), .Y(n61408) );
  NAND2xp33_ASAP7_75t_SL U53807 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[29]), .B(n66182), 
        .Y(n65574) );
  NAND2xp33_ASAP7_75t_SL U53808 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[20]), .B(n57205), .Y(
        n73744) );
  AOI22xp33_ASAP7_75t_SL U53809 ( .A1(n73833), .A2(n57204), .B1(n73679), .B2(
        n59632), .Y(n73682) );
  NAND2xp5_ASAP7_75t_SL U53810 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[1]), .B(
        n73889), .Y(n73896) );
  INVx1_ASAP7_75t_SL U53811 ( .A(n74066), .Y(n73895) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U53812 ( .A1(n59573), .A2(n75890), .B(n57212), 
        .C(n60604), .Y(n60605) );
  AOI22xp33_ASAP7_75t_SL U53813 ( .A1(n57217), .A2(n73680), .B1(n73828), .B2(
        n57205), .Y(n73681) );
  INVxp33_ASAP7_75t_SL U53814 ( .A(n74016), .Y(n76336) );
  NAND2xp33_ASAP7_75t_SL U53815 ( .A(n73685), .B(n57205), .Y(n73672) );
  AOI21xp33_ASAP7_75t_SL U53816 ( .A1(n57205), .A2(n73680), .B(n73752), .Y(
        n73670) );
  AOI22xp33_ASAP7_75t_SL U53817 ( .A1(n57217), .A2(n73708), .B1(n73828), .B2(
        n57204), .Y(n73671) );
  INVxp67_ASAP7_75t_SL U53818 ( .A(n64779), .Y(n59587) );
  INVx1_ASAP7_75t_SL U53819 ( .A(n77859), .Y(n75198) );
  INVxp67_ASAP7_75t_SL U53820 ( .A(n77875), .Y(n75447) );
  INVx1_ASAP7_75t_SL U53821 ( .A(n77856), .Y(n75675) );
  NAND2xp33_ASAP7_75t_SL U53822 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_), 
        .B(n72516), .Y(n71972) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U53823 ( .A1(n59527), .A2(n72362), .B(n72361), 
        .C(n72367), .Y(n72363) );
  INVx2_ASAP7_75t_SL U53824 ( .A(n72417), .Y(n59622) );
  INVxp33_ASAP7_75t_SL U53825 ( .A(n60668), .Y(n60622) );
  INVx2_ASAP7_75t_SL U53826 ( .A(n58611), .Y(n57208) );
  HB1xp67_ASAP7_75t_SL U53827 ( .A(n59079), .Y(n58175) );
  INVx1_ASAP7_75t_SL U53828 ( .A(n72507), .Y(n72494) );
  INVx1_ASAP7_75t_SL U53829 ( .A(n63531), .Y(n63440) );
  NAND2xp5_ASAP7_75t_SL U53830 ( .A(n65225), .B(n65224), .Y(n65231) );
  INVxp67_ASAP7_75t_SL U53831 ( .A(n65142), .Y(n65125) );
  INVx1_ASAP7_75t_SL U53832 ( .A(n74062), .Y(n74097) );
  NAND2xp33_ASAP7_75t_SL U53833 ( .A(n72313), .B(n57216), .Y(n71875) );
  NAND2xp5_ASAP7_75t_SL U53834 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_0_), 
        .B(n57216), .Y(n72411) );
  NAND2xp5_ASAP7_75t_SL U53835 ( .A(n59956), .B(n77210), .Y(n77254) );
  NAND2xp33_ASAP7_75t_SL U53836 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .B(n57216), .Y(n71811) );
  NAND2xp5_ASAP7_75t_SL U53837 ( .A(n74265), .B(n74064), .Y(n74065) );
  NOR2xp33_ASAP7_75t_SL U53838 ( .A(n59544), .B(n58084), .Y(n76363) );
  INVxp67_ASAP7_75t_SL U53839 ( .A(n61156), .Y(n76675) );
  BUFx2_ASAP7_75t_SL U53840 ( .A(n77953), .Y(n59493) );
  NAND4xp25_ASAP7_75t_SRAM U53841 ( .A(n60290), .B(n3080), .C(n1494), .D(n1492), .Y(n60200) );
  NOR2x1_ASAP7_75t_SL U53842 ( .A(n74802), .B(n60690), .Y(n77091) );
  INVx1_ASAP7_75t_SL U53843 ( .A(n57377), .Y(n64114) );
  NAND2xp33_ASAP7_75t_SL U53844 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[22]), .B(n57217), .Y(
        n73729) );
  NAND2xp5_ASAP7_75t_SL U53845 ( .A(n72141), .B(n71497), .Y(n71437) );
  NOR2xp33_ASAP7_75t_SL U53846 ( .A(n74093), .B(n65629), .Y(n74137) );
  NAND2xp5_ASAP7_75t_SL U53847 ( .A(n70229), .B(n70371), .Y(n59521) );
  OAI22xp5_ASAP7_75t_SL U53848 ( .A1(dbg_stb_i), .A2(n59945), .B1(
        dbg_adr_i[12]), .B2(n78439), .Y(n77994) );
  INVxp33_ASAP7_75t_SL U53849 ( .A(n70535), .Y(n70491) );
  INVx1_ASAP7_75t_SL U53850 ( .A(n70844), .Y(n70812) );
  AOI31xp33_ASAP7_75t_SL U53851 ( .A1(n71588), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .A3(n72351), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_), 
        .Y(n71589) );
  NAND2xp33_ASAP7_75t_SL U53852 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[11]), .B(n57217), .Y(
        n73632) );
  INVx1_ASAP7_75t_SL U53853 ( .A(n65629), .Y(n66182) );
  INVx1_ASAP7_75t_SL U53854 ( .A(n65653), .Y(n66146) );
  NAND2xp5_ASAP7_75t_SL U53855 ( .A(n57217), .B(n73685), .Y(n73831) );
  NAND2xp5_ASAP7_75t_SL U53856 ( .A(n65629), .B(n65653), .Y(n65670) );
  INVxp67_ASAP7_75t_SL U53857 ( .A(n65646), .Y(n65634) );
  INVx1_ASAP7_75t_SL U53858 ( .A(n74122), .Y(n59793) );
  INVxp33_ASAP7_75t_SL U53859 ( .A(n76202), .Y(n76203) );
  OAI21xp33_ASAP7_75t_SL U53860 ( .A1(n58423), .A2(n73755), .B(n3309), .Y(
        n73758) );
  NOR2xp33_ASAP7_75t_SL U53861 ( .A(n74672), .B(n74671), .Y(n74673) );
  INVxp67_ASAP7_75t_SL U53862 ( .A(n74121), .Y(n59818) );
  NAND2xp33_ASAP7_75t_SL U53863 ( .A(n77752), .B(n77756), .Y(n77753) );
  INVx1_ASAP7_75t_SL U53864 ( .A(n71335), .Y(n71394) );
  INVxp67_ASAP7_75t_SL U53865 ( .A(n66136), .Y(n65523) );
  NOR2xp33_ASAP7_75t_SL U53866 ( .A(dbg_stb_i), .B(n59926), .Y(n59927) );
  INVx1_ASAP7_75t_SL U53867 ( .A(n70674), .Y(n70669) );
  AOI22xp5_ASAP7_75t_SL U53868 ( .A1(n70676), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[20]), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[21]), .B2(n70674), 
        .Y(n70672) );
  INVxp33_ASAP7_75t_SL U53869 ( .A(n59799), .Y(n59760) );
  NAND2xp33_ASAP7_75t_SL U53870 ( .A(n72234), .B(n57216), .Y(n71847) );
  INVxp67_ASAP7_75t_SL U53871 ( .A(n59839), .Y(n75441) );
  AOI21xp33_ASAP7_75t_SL U53872 ( .A1(n70542), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_24_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .Y(
        n70275) );
  INVx1_ASAP7_75t_SL U53873 ( .A(n72877), .Y(n73031) );
  NAND2xp33_ASAP7_75t_SL U53874 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_), 
        .B(n57216), .Y(n71808) );
  OAI22xp33_ASAP7_75t_SL U53875 ( .A1(n73679), .A2(n58400), .B1(n3337), .B2(
        n58622), .Y(n73640) );
  INVxp33_ASAP7_75t_SL U53876 ( .A(n74495), .Y(n69525) );
  OAI22xp33_ASAP7_75t_SL U53877 ( .A1(n73833), .A2(n58619), .B1(n73828), .B2(
        n58423), .Y(n73639) );
  INVx1_ASAP7_75t_SL U53878 ( .A(n70540), .Y(n70543) );
  INVx1_ASAP7_75t_SL U53879 ( .A(n70676), .Y(n70662) );
  INVxp33_ASAP7_75t_SL U53880 ( .A(n69526), .Y(n69531) );
  O2A1O1Ixp5_ASAP7_75t_SL U53881 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .A2(n71502), .B(n72365), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_1_), 
        .Y(n71503) );
  NAND2xp33_ASAP7_75t_SL U53882 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[15]), .B(n58315), 
        .Y(n70651) );
  INVxp33_ASAP7_75t_SL U53883 ( .A(n65658), .Y(n65455) );
  A2O1A1Ixp33_ASAP7_75t_SL U53884 ( .A1(n65804), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[37]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[39]), .C(n65805), 
        .Y(n65430) );
  INVx1_ASAP7_75t_SL U53885 ( .A(n72437), .Y(n59625) );
  INVxp67_ASAP7_75t_SL U53886 ( .A(n59106), .Y(n59105) );
  INVx1_ASAP7_75t_SL U53887 ( .A(n70686), .Y(n58302) );
  INVxp67_ASAP7_75t_SL U53888 ( .A(n63751), .Y(n63754) );
  INVx1_ASAP7_75t_SL U53889 ( .A(n69385), .Y(n69411) );
  INVxp67_ASAP7_75t_SL U53890 ( .A(n59550), .Y(n76429) );
  NAND2xp33_ASAP7_75t_SL U53891 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .B(n78372), .Y(
        n72599) );
  INVxp33_ASAP7_75t_SL U53892 ( .A(n72266), .Y(n72267) );
  INVx1_ASAP7_75t_SL U53893 ( .A(n68821), .Y(n68822) );
  NAND2xp33_ASAP7_75t_SL U53894 ( .A(n78344), .B(n78342), .Y(n69537) );
  INVx1_ASAP7_75t_SL U53895 ( .A(n72994), .Y(n72963) );
  NAND2xp5_ASAP7_75t_SL U53896 ( .A(n72996), .B(n72994), .Y(n72877) );
  NAND2xp33_ASAP7_75t_SL U53897 ( .A(n65745), .B(n65544), .Y(n65379) );
  INVxp33_ASAP7_75t_SL U53898 ( .A(n69386), .Y(n69402) );
  NAND2xp33_ASAP7_75t_SL U53899 ( .A(n74751), .B(n66197), .Y(n66198) );
  INVxp67_ASAP7_75t_SL U53900 ( .A(n65495), .Y(n65506) );
  NOR3x1_ASAP7_75t_SL U53901 ( .A(n65487), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_1_), .C(n2491), .Y(
        n76976) );
  INVx3_ASAP7_75t_SL U53902 ( .A(n59526), .Y(n71365) );
  NAND2xp5_ASAP7_75t_SL U53903 ( .A(n69532), .B(n69535), .Y(n69530) );
  INVxp67_ASAP7_75t_SL U53904 ( .A(n74731), .Y(n74732) );
  NAND2xp5_ASAP7_75t_SL U53905 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[23]), .B(
        n73333), .Y(n73088) );
  NAND2xp5_ASAP7_75t_SL U53906 ( .A(n2450), .B(n69583), .Y(n70478) );
  INVx1_ASAP7_75t_SL U53907 ( .A(n74133), .Y(n65528) );
  AOI21xp5_ASAP7_75t_SL U53908 ( .A1(n70530), .A2(n69377), .B(n2451), .Y(
        n70289) );
  NAND2xp33_ASAP7_75t_SL U53909 ( .A(n76253), .B(n75783), .Y(n60842) );
  NAND2xp5_ASAP7_75t_SL U53910 ( .A(n72132), .B(n72080), .Y(n71484) );
  INVx1_ASAP7_75t_SL U53911 ( .A(n59546), .Y(n57218) );
  NAND2xp5_ASAP7_75t_SL U53912 ( .A(n1894), .B(n59533), .Y(n59854) );
  NAND2xp33_ASAP7_75t_SL U53913 ( .A(n74644), .B(n74686), .Y(n70336) );
  INVx3_ASAP7_75t_SL U53914 ( .A(n59580), .Y(n57219) );
  NAND2xp5_ASAP7_75t_SL U53915 ( .A(n1876), .B(n59576), .Y(n59881) );
  NAND2xp33_ASAP7_75t_SL U53916 ( .A(n58315), .B(n71229), .Y(n70844) );
  NAND2xp33_ASAP7_75t_SL U53917 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_9_), .B(
        n74686), .Y(n70423) );
  NOR2x1_ASAP7_75t_SL U53918 ( .A(n1915), .B(n59573), .Y(n75189) );
  INVx1_ASAP7_75t_SL U53919 ( .A(n71281), .Y(n71209) );
  NAND2xp5_ASAP7_75t_SL U53920 ( .A(n70183), .B(n70184), .Y(n70169) );
  NAND2xp5_ASAP7_75t_SL U53921 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_), .B(
        n74682), .Y(n70540) );
  NAND2xp5_ASAP7_75t_SL U53922 ( .A(n72309), .B(n71629), .Y(n71418) );
  INVx1_ASAP7_75t_SL U53923 ( .A(n59924), .Y(n77581) );
  NAND2xp5_ASAP7_75t_SL U53924 ( .A(n62477), .B(dbg_dat_i[11]), .Y(n4042) );
  NAND2xp33_ASAP7_75t_SL U53925 ( .A(n62477), .B(dbg_dat_i[5]), .Y(n4067) );
  NAND2xp33_ASAP7_75t_SL U53926 ( .A(n62477), .B(dbg_dat_i[8]), .Y(n4054) );
  NOR2xp33_ASAP7_75t_SL U53927 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .Y(n71579) );
  INVxp33_ASAP7_75t_SRAM U53928 ( .A(n1519), .Y(n61390) );
  INVxp67_ASAP7_75t_SL U53929 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_1_), .Y(
        n74682) );
  INVxp67_ASAP7_75t_SL U53930 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .Y(n72250) );
  INVxp67_ASAP7_75t_SL U53931 ( .A(n3024), .Y(n60095) );
  INVxp67_ASAP7_75t_SL U53932 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_5_), .Y(
        n70486) );
  NAND2xp5_ASAP7_75t_SL U53933 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .Y(
        n71890) );
  INVx1_ASAP7_75t_SL U53934 ( .A(n2600), .Y(n60304) );
  INVx1_ASAP7_75t_SL U53935 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[1]), .Y(
        n73864) );
  NOR2xp33_ASAP7_75t_SL U53936 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[37]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[38]), .Y(n65462) );
  INVxp67_ASAP7_75t_SL U53937 ( .A(n3054), .Y(n77258) );
  INVxp67_ASAP7_75t_SL U53938 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_10_), 
        .Y(n72341) );
  INVx2_ASAP7_75t_SL U53939 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .Y(
        n72544) );
  NOR2xp33_ASAP7_75t_SL U53940 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[24]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[27]), .Y(n74761) );
  INVx1_ASAP7_75t_SL U53941 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_4_), .Y(n69583) );
  NOR2xp33_ASAP7_75t_SL U53942 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[26]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[25]), .Y(n74762) );
  NOR2xp33_ASAP7_75t_SL U53943 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output1_23_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[30]), .Y(n74763) );
  INVx1_ASAP7_75t_SL U53944 ( .A(n3105), .Y(n78184) );
  INVx1_ASAP7_75t_SL U53945 ( .A(n3074), .Y(n61995) );
  INVx1_ASAP7_75t_SL U53946 ( .A(or1200_cpu_or1200_mult_mac_n24), .Y(n58850)
         );
  INVxp67_ASAP7_75t_SL U53947 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[0]), .Y(n65405) );
  NOR2xp33_ASAP7_75t_SL U53948 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_3_), .Y(
        n74483) );
  INVxp67_ASAP7_75t_SL U53949 ( .A(n2860), .Y(n65264) );
  INVx1_ASAP7_75t_SL U53950 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_22_), .Y(n69708) );
  BUFx3_ASAP7_75t_SL U53951 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_0_), .Y(
        n59527) );
  INVxp67_ASAP7_75t_SL U53952 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]), .Y(n65507) );
  NOR2xp33_ASAP7_75t_SL U53953 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[28]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[29]), .Y(n74760) );
  INVx1_ASAP7_75t_SL U53954 ( .A(or1200_cpu_or1200_except_n561), .Y(n60217) );
  INVxp67_ASAP7_75t_SL U53955 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_0_), .Y(
        n78438) );
  INVxp33_ASAP7_75t_SL U53956 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_0_), .Y(n74202) );
  INVxp67_ASAP7_75t_SL U53957 ( .A(or1200_cpu_or1200_mult_mac_n48), .Y(n76023)
         );
  INVxp67_ASAP7_75t_SL U53958 ( .A(n2807), .Y(n60590) );
  INVxp67_ASAP7_75t_SL U53959 ( .A(n3033), .Y(n63938) );
  INVxp67_ASAP7_75t_SL U53960 ( .A(n3060), .Y(n61583) );
  INVxp67_ASAP7_75t_SL U53961 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_), 
        .Y(n72306) );
  INVxp67_ASAP7_75t_SL U53962 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_), 
        .Y(n72308) );
  INVxp67_ASAP7_75t_SL U53963 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_), 
        .Y(n72197) );
  INVx1_ASAP7_75t_SL U53964 ( .A(n767), .Y(n59986) );
  INVxp67_ASAP7_75t_SL U53965 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_), 
        .Y(n72162) );
  INVxp67_ASAP7_75t_SL U53966 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_6_), .Y(n69613) );
  INVxp67_ASAP7_75t_SL U53967 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_), 
        .Y(n72164) );
  INVxp67_ASAP7_75t_SL U53968 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_), .Y(n78360) );
  INVx1_ASAP7_75t_SL U53969 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_7_), .Y(n69601) );
  INVxp67_ASAP7_75t_SL U53970 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .Y(n72219) );
  INVx1_ASAP7_75t_SL U53971 ( .A(n2585), .Y(n59921) );
  INVx1_ASAP7_75t_SL U53972 ( .A(n1830), .Y(n76216) );
  INVxp67_ASAP7_75t_SL U53973 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_), 
        .Y(n72307) );
  INVx3_ASAP7_75t_SL U53974 ( .A(n3374), .Y(n59700) );
  INVxp67_ASAP7_75t_SL U53975 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_), 
        .Y(n72310) );
  INVxp67_ASAP7_75t_SL U53976 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_13_), .Y(n69655) );
  INVx1_ASAP7_75t_SL U53977 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_1_), .Y(n65672) );
  INVxp67_ASAP7_75t_SL U53978 ( .A(or1200_cpu_or1200_mult_mac_n327), .Y(n65078) );
  INVxp67_ASAP7_75t_SL U53979 ( .A(or1200_cpu_or1200_mult_mac_n90), .Y(n74609)
         );
  INVx1_ASAP7_75t_SL U53980 ( .A(n1943), .Y(n76648) );
  INVx1_ASAP7_75t_SL U53981 ( .A(or1200_cpu_or1200_mult_mac_n317), .Y(n63501)
         );
  INVxp67_ASAP7_75t_SL U53982 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_30_), .Y(n78383) );
  INVxp67_ASAP7_75t_SL U53983 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_20_), .Y(n69702) );
  INVx1_ASAP7_75t_SL U53984 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_14_), .Y(n78432) );
  INVxp67_ASAP7_75t_SL U53985 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_), .Y(n78378) );
  INVxp67_ASAP7_75t_SL U53986 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_), 
        .Y(n72360) );
  INVxp67_ASAP7_75t_SL U53987 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_), .Y(n78375) );
  INVxp33_ASAP7_75t_SL U53988 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_), 
        .Y(n72362) );
  INVx1_ASAP7_75t_SL U53989 ( .A(or1200_cpu_or1200_mult_mac_n345), .Y(n68789)
         );
  INVxp67_ASAP7_75t_SL U53990 ( .A(or1200_cpu_or1200_mult_mac_n70), .Y(n75218)
         );
  INVx1_ASAP7_75t_SL U53991 ( .A(n1951), .Y(n76622) );
  INVxp67_ASAP7_75t_SL U53992 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_12_), .Y(n69641) );
  INVxp67_ASAP7_75t_SL U53993 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .Y(
        n72400) );
  INVxp67_ASAP7_75t_SL U53994 ( .A(or1200_cpu_or1200_mult_mac_n78), .Y(n64240)
         );
  INVxp33_ASAP7_75t_SL U53995 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[12]), .Y(
        n73064) );
  INVx2_ASAP7_75t_SL U53996 ( .A(n53473), .Y(n71015) );
  INVxp67_ASAP7_75t_SL U53997 ( .A(n1237), .Y(dwb_adr_o[21]) );
  INVxp67_ASAP7_75t_SL U53998 ( .A(or1200_cpu_or1200_except_n661), .Y(n75167)
         );
  NAND2xp5_ASAP7_75t_SL U53999 ( .A(or1200_cpu_or1200_mult_mac_n225), .B(
        or1200_cpu_or1200_mult_mac_n371), .Y(n69108) );
  INVxp67_ASAP7_75t_SL U54000 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[24]), .Y(
        n73111) );
  INVx1_ASAP7_75t_SL U54001 ( .A(or1200_cpu_or1200_mult_mac_n247), .Y(n69220)
         );
  INVx1_ASAP7_75t_SL U54002 ( .A(n1588), .Y(n77732) );
  NAND2xp5_ASAP7_75t_SL U54003 ( .A(or1200_cpu_or1200_mult_mac_n243), .B(
        or1200_cpu_or1200_mult_mac_n389), .Y(n69210) );
  INVxp33_ASAP7_75t_SL U54004 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[20]), .Y(n73767) );
  NAND2xp5_ASAP7_75t_SL U54005 ( .A(or1200_cpu_or1200_mult_mac_n213), .B(
        or1200_cpu_or1200_mult_mac_n359), .Y(n68931) );
  NAND2xp5_ASAP7_75t_SL U54006 ( .A(or1200_cpu_or1200_except_n592), .B(n2464), 
        .Y(n63750) );
  NAND2xp5_ASAP7_75t_SL U54007 ( .A(or1200_cpu_or1200_except_n589), .B(n2499), 
        .Y(n63751) );
  INVxp33_ASAP7_75t_SL U54008 ( .A(n1626), .Y(n77717) );
  INVxp67_ASAP7_75t_SL U54009 ( .A(or1200_cpu_or1200_except_n598), .Y(n76703)
         );
  INVxp33_ASAP7_75t_SL U54010 ( .A(n2569), .Y(n77708) );
  INVxp67_ASAP7_75t_SL U54011 ( .A(n3331), .Y(n73823) );
  BUFx2_ASAP7_75t_SL U54012 ( .A(n1929), .Y(n59551) );
  INVx1_ASAP7_75t_SL U54013 ( .A(or1200_cpu_or1200_mult_mac_n207), .Y(n68846)
         );
  INVx1_ASAP7_75t_SL U54014 ( .A(n1171), .Y(n62229) );
  INVx1_ASAP7_75t_SL U54015 ( .A(n3313), .Y(n73706) );
  INVx1_ASAP7_75t_SL U54016 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_8_), .Y(
        n70633) );
  BUFx2_ASAP7_75t_SL U54017 ( .A(n1774), .Y(n59539) );
  BUFx2_ASAP7_75t_SL U54018 ( .A(n1934), .Y(n59552) );
  INVx1_ASAP7_75t_SL U54019 ( .A(n1768), .Y(n77219) );
  INVxp33_ASAP7_75t_SL U54020 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_6_), .Y(n65321) );
  INVxp33_ASAP7_75t_SL U54021 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[17]), .Y(n73687) );
  INVxp67_ASAP7_75t_SL U54022 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_output_o_31_), .Y(
        n27324) );
  NAND2xp5_ASAP7_75t_SL U54023 ( .A(n3090), .B(n3086), .Y(n77473) );
  INVxp33_ASAP7_75t_SRAM U54024 ( .A(n2450), .Y(n69382) );
  INVxp33_ASAP7_75t_SL U54025 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[4]), .Y(n73680) );
  INVxp33_ASAP7_75t_SL U54026 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[11]), .Y(n73810) );
  INVxp33_ASAP7_75t_SL U54027 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[8]), .Y(n73668) );
  INVxp67_ASAP7_75t_SL U54028 ( .A(n3071), .Y(n77241) );
  INVxp33_ASAP7_75t_SL U54029 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[15]), .Y(n73696) );
  NAND2xp33_ASAP7_75t_SL U54030 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .B(
        n3309), .Y(n73791) );
  INVxp33_ASAP7_75t_SL U54031 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[18]), .Y(n73688) );
  INVxp67_ASAP7_75t_SL U54032 ( .A(or1200_cpu_or1200_except_n601), .Y(n76849)
         );
  INVxp33_ASAP7_75t_SL U54033 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_19_), .Y(n74868)
         );
  INVx2_ASAP7_75t_SL U54034 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_0_), .Y(n70686) );
  INVxp33_ASAP7_75t_SL U54035 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_18_), .Y(n74863)
         );
  INVxp67_ASAP7_75t_SL U54036 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_31_), .Y(n78226) );
  INVx1_ASAP7_75t_SL U54037 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[0]), .Y(n78329)
         );
  INVx1_ASAP7_75t_SL U54038 ( .A(or1200_dc_top_tag_5_), .Y(n59815) );
  INVxp67_ASAP7_75t_SL U54039 ( .A(n59421), .Y(n59420) );
  AOI21xp33_ASAP7_75t_SL U54040 ( .A1(n65071), .A2(n68757), .B(n68765), .Y(
        n52057) );
  NAND2xp5_ASAP7_75t_SL U54041 ( .A(n58866), .B(n58339), .Y(n68921) );
  INVxp67_ASAP7_75t_SL U54042 ( .A(n58772), .Y(n58769) );
  INVxp67_ASAP7_75t_SL U54043 ( .A(n75279), .Y(n68713) );
  NAND2xp33_ASAP7_75t_SL U54044 ( .A(n59295), .B(n58881), .Y(n69105) );
  AND2x4_ASAP7_75t_SL U54045 ( .A(n58190), .B(n58830), .Y(n75109) );
  NAND2xp33_ASAP7_75t_SL U54046 ( .A(n69297), .B(n59214), .Y(n58827) );
  INVxp67_ASAP7_75t_SL U54047 ( .A(n68976), .Y(n68977) );
  INVxp67_ASAP7_75t_SL U54048 ( .A(n69123), .Y(n58869) );
  INVxp67_ASAP7_75t_SL U54049 ( .A(n69236), .Y(n59251) );
  INVxp67_ASAP7_75t_SL U54050 ( .A(n65123), .Y(n52053) );
  NAND2xp5_ASAP7_75t_SL U54051 ( .A(n74565), .B(n74564), .Y(n74566) );
  NAND2xp5_ASAP7_75t_SL U54052 ( .A(n69041), .B(n69043), .Y(n69042) );
  O2A1O1Ixp33_ASAP7_75t_SL U54053 ( .A1(n65122), .A2(n75790), .B(n65121), .C(
        n65120), .Y(n65123) );
  NAND2xp33_ASAP7_75t_SL U54054 ( .A(n68644), .B(n68645), .Y(n59422) );
  AOI21xp33_ASAP7_75t_SL U54055 ( .A1(n69100), .A2(n69101), .B(n69099), .Y(
        n69104) );
  INVxp33_ASAP7_75t_SL U54056 ( .A(n75114), .Y(n75108) );
  AOI21xp33_ASAP7_75t_SL U54057 ( .A1(n75790), .A2(n75789), .B(n75788), .Y(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N22) );
  OAI21xp33_ASAP7_75t_SL U54058 ( .A1(n75091), .A2(n75085), .B(n75461), .Y(
        n75086) );
  INVxp67_ASAP7_75t_SL U54059 ( .A(n69157), .Y(n69154) );
  INVxp33_ASAP7_75t_SL U54060 ( .A(n57085), .Y(n58339) );
  NAND2xp33_ASAP7_75t_SL U54061 ( .A(n69115), .B(n69151), .Y(n69120) );
  AND2x2_ASAP7_75t_SL U54062 ( .A(n68701), .B(n68652), .Y(n69298) );
  NAND2xp33_ASAP7_75t_SL U54063 ( .A(n69239), .B(n69241), .Y(n69237) );
  INVx1_ASAP7_75t_SL U54064 ( .A(n58442), .Y(n58637) );
  INVxp67_ASAP7_75t_SL U54065 ( .A(n74558), .Y(n68716) );
  AOI21xp5_ASAP7_75t_SL U54066 ( .A1(n68964), .A2(n58345), .B(n68960), .Y(
        n68927) );
  INVxp33_ASAP7_75t_SL U54067 ( .A(n68686), .Y(n58745) );
  NAND2xp33_ASAP7_75t_SL U54068 ( .A(n74111), .B(n68686), .Y(n68690) );
  NAND2xp5_ASAP7_75t_SL U54069 ( .A(n70617), .B(n70615), .Y(n12856) );
  NAND2xp33_ASAP7_75t_SL U54070 ( .A(n68902), .B(n76881), .Y(n68903) );
  INVxp67_ASAP7_75t_SL U54071 ( .A(n68681), .Y(n68683) );
  INVx1_ASAP7_75t_SL U54072 ( .A(n68869), .Y(n57129) );
  INVxp67_ASAP7_75t_SL U54073 ( .A(n75110), .Y(n67222) );
  NAND2xp33_ASAP7_75t_SL U54074 ( .A(n69155), .B(n69152), .Y(n69159) );
  NOR2xp33_ASAP7_75t_SL U54075 ( .A(n71416), .B(n71415), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n244) );
  INVxp67_ASAP7_75t_SL U54076 ( .A(n68854), .Y(n58867) );
  INVxp67_ASAP7_75t_SL U54077 ( .A(n69229), .Y(n69240) );
  INVxp67_ASAP7_75t_SL U54078 ( .A(n69032), .Y(n68731) );
  INVxp33_ASAP7_75t_SL U54079 ( .A(n68651), .Y(n68653) );
  INVxp67_ASAP7_75t_SL U54080 ( .A(n58958), .Y(n58956) );
  INVx1_ASAP7_75t_SL U54081 ( .A(n68675), .Y(n68671) );
  INVxp33_ASAP7_75t_SL U54082 ( .A(n69235), .Y(n68679) );
  INVxp33_ASAP7_75t_SL U54083 ( .A(n68868), .Y(n68866) );
  NAND2x1_ASAP7_75t_SL U54084 ( .A(n58329), .B(n68749), .Y(n68808) );
  INVxp33_ASAP7_75t_SL U54085 ( .A(n69303), .Y(n69297) );
  INVxp33_ASAP7_75t_SL U54086 ( .A(n68961), .Y(n58345) );
  AOI21xp33_ASAP7_75t_SL U54087 ( .A1(n68707), .A2(n74561), .B(n68706), .Y(
        n68708) );
  INVxp67_ASAP7_75t_SL U54088 ( .A(n69307), .Y(n69308) );
  INVx2_ASAP7_75t_SL U54089 ( .A(n68916), .Y(n58686) );
  INVxp33_ASAP7_75t_SL U54090 ( .A(n70607), .Y(n70614) );
  INVxp33_ASAP7_75t_SL U54091 ( .A(n68807), .Y(n68745) );
  O2A1O1Ixp33_ASAP7_75t_SL U54092 ( .A1(n53482), .A2(n57341), .B(n59434), .C(
        n68739), .Y(n68741) );
  INVxp67_ASAP7_75t_SL U54093 ( .A(n71414), .Y(n71412) );
  NAND2xp5_ASAP7_75t_SL U54094 ( .A(n69305), .B(n69302), .Y(n69307) );
  INVx2_ASAP7_75t_SL U54095 ( .A(n69116), .Y(n57130) );
  INVxp33_ASAP7_75t_SL U54096 ( .A(n68654), .Y(n68656) );
  INVxp67_ASAP7_75t_SL U54097 ( .A(n76880), .Y(n58349) );
  INVxp67_ASAP7_75t_SL U54098 ( .A(n76195), .Y(n76196) );
  OAI21xp33_ASAP7_75t_SL U54099 ( .A1(n2972), .A2(n77454), .B(n77366), .Y(
        n9456) );
  INVx3_ASAP7_75t_SL U54100 ( .A(n58377), .Y(n76881) );
  OAI21xp33_ASAP7_75t_SL U54101 ( .A1(n57074), .A2(n2976), .B(n77393), .Y(
        n2977) );
  AOI22xp33_ASAP7_75t_SL U54102 ( .A1(n58600), .A2(n76112), .B1(n76111), .B2(
        n76195), .Y(n76113) );
  AOI22xp33_ASAP7_75t_SL U54103 ( .A1(n58600), .A2(n76106), .B1(n76105), .B2(
        n76195), .Y(n76107) );
  INVxp33_ASAP7_75t_SL U54104 ( .A(n68732), .Y(n68729) );
  AOI22xp33_ASAP7_75t_SL U54105 ( .A1(n58600), .A2(n76085), .B1(n76084), .B2(
        n76195), .Y(n76086) );
  OAI21xp33_ASAP7_75t_SL U54106 ( .A1(n2982), .A2(n57073), .B(n75184), .Y(
        n2983) );
  INVxp33_ASAP7_75t_SL U54107 ( .A(n69230), .Y(n69234) );
  AOI22xp33_ASAP7_75t_SL U54108 ( .A1(n58600), .A2(n76065), .B1(n76064), .B2(
        n76195), .Y(n76066) );
  INVx1_ASAP7_75t_SL U54109 ( .A(n68837), .Y(n68826) );
  AOI22xp33_ASAP7_75t_SL U54110 ( .A1(n58600), .A2(n76045), .B1(n76044), .B2(
        n76195), .Y(n76046) );
  AOI22xp33_ASAP7_75t_SL U54111 ( .A1(n58600), .A2(n75980), .B1(n75979), .B2(
        n76195), .Y(n75981) );
  AOI22xp33_ASAP7_75t_SL U54112 ( .A1(n58600), .A2(n76038), .B1(n76037), .B2(
        n76195), .Y(n76039) );
  AOI22xp33_ASAP7_75t_SL U54113 ( .A1(n58600), .A2(n76005), .B1(n75999), .B2(
        n76195), .Y(n76000) );
  AOI22xp33_ASAP7_75t_SL U54114 ( .A1(n58600), .A2(n76023), .B1(n76022), .B2(
        n76195), .Y(n76024) );
  NAND2xp33_ASAP7_75t_SL U54115 ( .A(n57421), .B(n68907), .Y(n68868) );
  NAND2xp33_ASAP7_75t_SL U54116 ( .A(n76005), .B(n76004), .Y(n76006) );
  AOI22xp33_ASAP7_75t_SL U54117 ( .A1(n74454), .A2(n74329), .B1(n74352), .B2(
        n74444), .Y(n2889) );
  AOI22xp33_ASAP7_75t_SL U54118 ( .A1(n74454), .A2(n74352), .B1(n74351), .B2(
        n74437), .Y(n2888) );
  AOI22xp33_ASAP7_75t_SL U54119 ( .A1(n74454), .A2(n74351), .B1(n74396), .B2(
        n74444), .Y(n2887) );
  AOI22xp33_ASAP7_75t_SL U54120 ( .A1(n74454), .A2(n74323), .B1(n74330), .B2(
        n74444), .Y(n2891) );
  AOI22xp33_ASAP7_75t_SL U54121 ( .A1(n74454), .A2(n74365), .B1(n74323), .B2(
        n74437), .Y(n2892) );
  AOI22xp33_ASAP7_75t_SL U54122 ( .A1(n74454), .A2(n74330), .B1(n74329), .B2(
        n74437), .Y(n2890) );
  NAND2xp5_ASAP7_75t_SL U54123 ( .A(n74086), .B(n74085), .Y(
        or1200_cpu_or1200_except_n1705) );
  NOR2xp67_ASAP7_75t_SL U54124 ( .A(n58818), .B(n64744), .Y(n57890) );
  NAND2xp5_ASAP7_75t_SL U54125 ( .A(n76865), .B(n76864), .Y(
        or1200_cpu_or1200_except_n1727) );
  NAND2xp5_ASAP7_75t_SL U54126 ( .A(n76686), .B(n76685), .Y(
        or1200_cpu_or1200_except_n1728) );
  NAND2xp5_ASAP7_75t_SL U54127 ( .A(n77155), .B(n77154), .Y(
        or1200_cpu_or1200_except_n1715) );
  NAND2xp5_ASAP7_75t_SL U54128 ( .A(n77001), .B(n77000), .Y(
        or1200_cpu_or1200_except_n1726) );
  INVxp33_ASAP7_75t_SL U54129 ( .A(n68703), .Y(n68704) );
  INVxp33_ASAP7_75t_SL U54130 ( .A(n68702), .Y(n68705) );
  INVxp67_ASAP7_75t_SL U54131 ( .A(n70610), .Y(n70605) );
  OAI21xp5_ASAP7_75t_SL U54132 ( .A1(n59677), .A2(n77878), .B(n62141), .Y(
        n9618) );
  OAI21xp33_ASAP7_75t_SL U54133 ( .A1(n77960), .A2(n77936), .B(n77935), .Y(
        or1200_cpu_or1200_rf_n7) );
  OAI21xp33_ASAP7_75t_SL U54134 ( .A1(n77960), .A2(n77946), .B(n77945), .Y(
        or1200_cpu_or1200_rf_n9) );
  OAI21xp33_ASAP7_75t_SL U54135 ( .A1(n77960), .A2(n77942), .B(n77941), .Y(
        or1200_cpu_or1200_rf_n8) );
  AOI22xp33_ASAP7_75t_SL U54136 ( .A1(n74454), .A2(n74374), .B1(n74380), .B2(
        n74444), .Y(n2894) );
  NAND2xp5_ASAP7_75t_SL U54137 ( .A(n77181), .B(n77180), .Y(
        or1200_cpu_or1200_except_n1702) );
  OAI21xp33_ASAP7_75t_SL U54138 ( .A1(n77960), .A2(n77951), .B(n77950), .Y(
        or1200_cpu_or1200_rf_n10) );
  OAI21xp33_ASAP7_75t_SL U54139 ( .A1(n74450), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_45_), .B(
        n74466), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n46) );
  NAND2xp5_ASAP7_75t_SL U54140 ( .A(n76921), .B(n76920), .Y(
        or1200_cpu_or1200_except_n1699) );
  AOI22xp33_ASAP7_75t_SL U54141 ( .A1(n74454), .A2(n74375), .B1(n74374), .B2(
        n74437), .Y(n2895) );
  OAI21xp33_ASAP7_75t_SL U54142 ( .A1(n77467), .A2(n77878), .B(n75437), .Y(
        n9649) );
  NAND2xp5_ASAP7_75t_SL U54143 ( .A(n74131), .B(n74130), .Y(
        or1200_cpu_or1200_except_n1710) );
  INVxp33_ASAP7_75t_SL U54144 ( .A(n69100), .Y(n69094) );
  NAND2xp5_ASAP7_75t_SL U54145 ( .A(n76642), .B(n76641), .Y(
        or1200_cpu_or1200_except_n1722) );
  NAND2xp5_ASAP7_75t_SL U54146 ( .A(n76555), .B(n76554), .Y(
        or1200_cpu_or1200_except_n1719) );
  INVxp67_ASAP7_75t_SL U54147 ( .A(n69299), .Y(n69305) );
  NAND2xp5_ASAP7_75t_SL U54148 ( .A(n76699), .B(n76698), .Y(
        or1200_cpu_or1200_except_n1723) );
  AOI22xp33_ASAP7_75t_SL U54149 ( .A1(n74454), .A2(n74445), .B1(n74453), .B2(
        n74437), .Y(n2878) );
  AOI22xp33_ASAP7_75t_SL U54150 ( .A1(n74454), .A2(n74436), .B1(n74445), .B2(
        n74444), .Y(n2879) );
  NAND2xp33_ASAP7_75t_SL U54151 ( .A(n59694), .B(n77392), .Y(n77393) );
  AOI22xp33_ASAP7_75t_SL U54152 ( .A1(n74454), .A2(n74438), .B1(n74436), .B2(
        n74437), .Y(n2880) );
  AOI22xp33_ASAP7_75t_SL U54153 ( .A1(n74438), .A2(n74437), .B1(n74454), .B2(
        n74427), .Y(n2881) );
  NAND2xp5_ASAP7_75t_SL U54154 ( .A(n77300), .B(n77299), .Y(
        or1200_cpu_or1200_except_n1718) );
  AOI22xp33_ASAP7_75t_SL U54155 ( .A1(n74454), .A2(n74419), .B1(n53460), .B2(
        n74427), .Y(n2882) );
  AOI21xp5_ASAP7_75t_SL U54156 ( .A1(n74281), .A2(n74280), .B(n74279), .Y(
        n1540) );
  NAND2xp5_ASAP7_75t_SL U54157 ( .A(n76621), .B(n76620), .Y(
        or1200_cpu_or1200_except_n1724) );
  AOI22xp33_ASAP7_75t_SL U54158 ( .A1(n74454), .A2(n74310), .B1(n74419), .B2(
        n74444), .Y(n2883) );
  AOI22xp33_ASAP7_75t_SL U54159 ( .A1(n74454), .A2(n74410), .B1(n74310), .B2(
        n74437), .Y(n2884) );
  AOI22xp33_ASAP7_75t_SL U54160 ( .A1(n74454), .A2(n74395), .B1(n74410), .B2(
        n74444), .Y(n2885) );
  OAI21xp33_ASAP7_75t_SL U54161 ( .A1(n77467), .A2(n77881), .B(n74553), .Y(
        n9650) );
  OAI21xp33_ASAP7_75t_SL U54162 ( .A1(n77961), .A2(n77960), .B(n77959), .Y(
        or1200_cpu_or1200_rf_n11) );
  NAND2xp33_ASAP7_75t_SL U54163 ( .A(n59694), .B(n75183), .Y(n75184) );
  OA21x2_ASAP7_75t_SRAM U54164 ( .A1(n57332), .A2(n65106), .B(n65101), .Y(
        n65103) );
  AOI22xp33_ASAP7_75t_SL U54165 ( .A1(n74454), .A2(n74396), .B1(n74395), .B2(
        n74437), .Y(n2886) );
  INVx1_ASAP7_75t_SL U54166 ( .A(n68828), .Y(n68570) );
  AOI22xp33_ASAP7_75t_SL U54167 ( .A1(n74454), .A2(n74334), .B1(n74375), .B2(
        n74444), .Y(n2896) );
  AOI22xp33_ASAP7_75t_SL U54168 ( .A1(n74454), .A2(n74335), .B1(n74334), .B2(
        n74444), .Y(n2897) );
  INVxp33_ASAP7_75t_SL U54169 ( .A(n57369), .Y(n69144) );
  AOI21xp33_ASAP7_75t_SL U54170 ( .A1(n74437), .A2(n74335), .B(n74306), .Y(
        n2898) );
  AOI21xp33_ASAP7_75t_SL U54171 ( .A1(n59681), .A2(n78160), .B(n77297), .Y(
        n77299) );
  NAND2xp5_ASAP7_75t_SL U54172 ( .A(n70602), .B(n70594), .Y(n70595) );
  INVxp67_ASAP7_75t_SL U54173 ( .A(n75042), .Y(n68641) );
  OAI21xp33_ASAP7_75t_SL U54174 ( .A1(n74242), .A2(n74313), .B(n74503), .Y(
        n74281) );
  AOI22xp33_ASAP7_75t_SL U54175 ( .A1(n77987), .A2(n59681), .B1(n77290), .B2(
        n76249), .Y(n76248) );
  AOI22xp33_ASAP7_75t_SL U54176 ( .A1(n74576), .A2(n77290), .B1(n59681), .B2(
        n78125), .Y(n74580) );
  INVxp67_ASAP7_75t_SL U54177 ( .A(n71388), .Y(n71410) );
  AOI22xp33_ASAP7_75t_SL U54178 ( .A1(n77151), .A2(n77290), .B1(n59681), .B2(
        n78144), .Y(n77155) );
  INVx1_ASAP7_75t_SL U54179 ( .A(n68972), .Y(n57131) );
  AOI22xp33_ASAP7_75t_SL U54180 ( .A1(n77225), .A2(n59681), .B1(n77290), .B2(
        n77224), .Y(n77229) );
  AOI22xp33_ASAP7_75t_SL U54181 ( .A1(n76551), .A2(n77290), .B1(n59681), .B2(
        n77970), .Y(n76555) );
  AOI22xp33_ASAP7_75t_SL U54182 ( .A1(n75780), .A2(n77290), .B1(n59681), .B2(
        n77964), .Y(n75785) );
  AOI21xp33_ASAP7_75t_SL U54183 ( .A1(n71407), .A2(n71406), .B(n71405), .Y(
        n71408) );
  AOI22xp33_ASAP7_75t_SL U54184 ( .A1(n74126), .A2(n77290), .B1(n59681), .B2(
        n78121), .Y(n74131) );
  AOI22xp33_ASAP7_75t_SL U54185 ( .A1(n75301), .A2(n77290), .B1(n59681), .B2(
        n78133), .Y(n75305) );
  AOI22xp33_ASAP7_75t_SL U54186 ( .A1(n78134), .A2(n59681), .B1(n77290), .B2(
        n76230), .Y(n76234) );
  AOI22xp33_ASAP7_75t_SL U54187 ( .A1(n78129), .A2(n59681), .B1(n77290), .B2(
        n74983), .Y(n74988) );
  AOI22xp33_ASAP7_75t_SL U54188 ( .A1(n77985), .A2(n59681), .B1(n77290), .B2(
        n76643), .Y(n76642) );
  AOI22xp33_ASAP7_75t_SL U54189 ( .A1(n77018), .A2(n77290), .B1(n59681), .B2(
        n78148), .Y(n77023) );
  AOI21xp33_ASAP7_75t_SL U54190 ( .A1(n70586), .A2(n70592), .B(n70603), .Y(
        n51979) );
  AOI22xp33_ASAP7_75t_SL U54191 ( .A1(n78084), .A2(n59681), .B1(n77290), .B2(
        n75795), .Y(n75800) );
  AOI22xp33_ASAP7_75t_SL U54192 ( .A1(n69367), .A2(n77290), .B1(n59681), .B2(
        n78088), .Y(n69375) );
  AOI22xp33_ASAP7_75t_SL U54193 ( .A1(n74084), .A2(n59681), .B1(n77290), .B2(
        n74083), .Y(n74085) );
  NAND2xp5_ASAP7_75t_SL U54194 ( .A(n68693), .B(n74565), .Y(n68702) );
  AOI22xp33_ASAP7_75t_SL U54195 ( .A1(n74044), .A2(n77290), .B1(n59681), .B2(
        n78105), .Y(n74049) );
  AOI21xp33_ASAP7_75t_SL U54196 ( .A1(n59681), .A2(n77495), .B(n76684), .Y(
        n76685) );
  NAND2xp5_ASAP7_75t_SL U54197 ( .A(n77934), .B(n77960), .Y(n77935) );
  INVxp67_ASAP7_75t_SL U54198 ( .A(n53296), .Y(n59098) );
  AOI22xp33_ASAP7_75t_SL U54199 ( .A1(n75619), .A2(n77290), .B1(n59681), .B2(
        n78109), .Y(n75624) );
  NAND2xp5_ASAP7_75t_SL U54200 ( .A(n77944), .B(n77960), .Y(n77945) );
  NAND2xp33_ASAP7_75t_SL U54201 ( .A(n71184), .B(n71188), .Y(n71191) );
  NAND2xp5_ASAP7_75t_SL U54202 ( .A(n77940), .B(n77960), .Y(n77941) );
  NAND2xp5_ASAP7_75t_SL U54203 ( .A(n77949), .B(n77960), .Y(n77950) );
  INVxp67_ASAP7_75t_SL U54204 ( .A(n65116), .Y(n65112) );
  AOI22xp33_ASAP7_75t_SL U54205 ( .A1(n75446), .A2(n77290), .B1(n59681), .B2(
        n78113), .Y(n75451) );
  AOI21xp33_ASAP7_75t_SL U54206 ( .A1(n59681), .A2(n77494), .B(n76863), .Y(
        n76864) );
  AOI22xp33_ASAP7_75t_SL U54207 ( .A1(n78080), .A2(n59681), .B1(n77290), .B2(
        n77176), .Y(n77181) );
  OAI21xp33_ASAP7_75t_SL U54208 ( .A1(n59698), .A2(n71195), .B(n71186), .Y(
        n71187) );
  INVxp33_ASAP7_75t_SL U54209 ( .A(n68668), .Y(n68669) );
  AOI22xp33_ASAP7_75t_SL U54210 ( .A1(n76997), .A2(n77290), .B1(n59681), .B2(
        n77973), .Y(n77001) );
  AOI22xp33_ASAP7_75t_SL U54211 ( .A1(n77982), .A2(n59681), .B1(n77290), .B2(
        n76700), .Y(n76699) );
  INVxp67_ASAP7_75t_SL U54212 ( .A(n58546), .Y(n58834) );
  AOI21xp33_ASAP7_75t_SL U54213 ( .A1(n78068), .A2(n59681), .B(n76919), .Y(
        n76920) );
  AOI22xp33_ASAP7_75t_SL U54214 ( .A1(n77976), .A2(n59681), .B1(n77290), .B2(
        n76210), .Y(n76209) );
  AOI22xp33_ASAP7_75t_SL U54215 ( .A1(n78076), .A2(n59681), .B1(n77290), .B2(
        n75197), .Y(n75202) );
  AOI22xp33_ASAP7_75t_SL U54216 ( .A1(n78117), .A2(n59681), .B1(n77290), .B2(
        n75430), .Y(n75435) );
  NAND2xp5_ASAP7_75t_SL U54217 ( .A(n69293), .B(n75042), .Y(n69299) );
  AOI22xp33_ASAP7_75t_SL U54218 ( .A1(n76617), .A2(n77290), .B1(n59681), .B2(
        n77979), .Y(n76621) );
  AOI22xp33_ASAP7_75t_SL U54219 ( .A1(n75674), .A2(n77290), .B1(n59681), .B2(
        n78072), .Y(n75678) );
  NAND2xp5_ASAP7_75t_SL U54220 ( .A(n75892), .B(n75891), .Y(n9642) );
  INVxp67_ASAP7_75t_SL U54221 ( .A(n75284), .Y(n68712) );
  OAI21xp33_ASAP7_75t_SL U54222 ( .A1(n74278), .A2(n58298), .B(n74362), .Y(
        n74279) );
  INVxp33_ASAP7_75t_SL U54223 ( .A(n68338), .Y(n64752) );
  INVxp33_ASAP7_75t_SL U54224 ( .A(n71185), .Y(n71188) );
  O2A1O1Ixp33_ASAP7_75t_SL U54225 ( .A1(n70970), .A2(n70963), .B(n70962), .C(
        n70961), .Y(n70964) );
  OAI21xp33_ASAP7_75t_SL U54226 ( .A1(n3419), .A2(n77298), .B(n77238), .Y(
        or1200_cpu_or1200_except_n1730) );
  INVx1_ASAP7_75t_SL U54227 ( .A(n74505), .Y(n57134) );
  OAI21xp5_ASAP7_75t_SL U54228 ( .A1(n59677), .A2(n74638), .B(n74637), .Y(
        n9620) );
  OAI21xp33_ASAP7_75t_SL U54229 ( .A1(n2843), .A2(n77298), .B(n77169), .Y(
        or1200_cpu_or1200_except_n1729) );
  NAND2xp5_ASAP7_75t_SL U54230 ( .A(n77189), .B(n77188), .Y(n9611) );
  NAND2x1p5_ASAP7_75t_SL U54231 ( .A(n77933), .B(or1200_cpu_or1200_rf_rf_ena), 
        .Y(n77960) );
  OAI21xp5_ASAP7_75t_SL U54232 ( .A1(n59677), .A2(n76989), .B(n61992), .Y(
        n9676) );
  AOI22xp33_ASAP7_75t_SL U54233 ( .A1(n74068), .A2(n74270), .B1(n74067), .B2(
        n74258), .Y(n74073) );
  OAI21xp33_ASAP7_75t_SL U54234 ( .A1(n74431), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_43_), .B(
        n74223), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n42) );
  OAI21xp33_ASAP7_75t_SL U54235 ( .A1(n77137), .A2(n75805), .B(n75804), .Y(
        n9612) );
  INVxp67_ASAP7_75t_SL U54236 ( .A(n74250), .Y(n74267) );
  OAI21xp33_ASAP7_75t_SL U54237 ( .A1(n3136), .A2(n77399), .B(n58280), .Y(
        n9474) );
  INVx1_ASAP7_75t_SL U54238 ( .A(n74362), .Y(n74260) );
  INVxp67_ASAP7_75t_SL U54239 ( .A(n68591), .Y(n68593) );
  OAI21xp33_ASAP7_75t_SL U54240 ( .A1(n77467), .A2(n76989), .B(n76988), .Y(
        n9673) );
  NAND2x1p5_ASAP7_75t_SL U54241 ( .A(n75278), .B(n57962), .Y(n68694) );
  OAI21xp33_ASAP7_75t_SL U54242 ( .A1(n58316), .A2(n4134), .B(n78161), .Y(
        n9698) );
  OAI21xp33_ASAP7_75t_SL U54243 ( .A1(n58316), .A2(n4135), .B(n78063), .Y(
        n9699) );
  NAND2xp5_ASAP7_75t_SL U54244 ( .A(n74269), .B(n74266), .Y(n74268) );
  AOI22xp33_ASAP7_75t_SL U54245 ( .A1(n77376), .A2(n61041), .B1(n61040), .B2(
        n61039), .Y(n61054) );
  NAND2xp5_ASAP7_75t_SL U54246 ( .A(n75380), .B(n75379), .Y(n9653) );
  NAND2xp5_ASAP7_75t_SL U54247 ( .A(n75385), .B(n75384), .Y(n9622) );
  NAND2x1_ASAP7_75t_SL U54248 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_43_), .B(
        n74431), .Y(n74223) );
  NAND2xp5_ASAP7_75t_SL U54249 ( .A(n75530), .B(n75529), .Y(
        or1200_cpu_to_sr[11]) );
  OAI22xp33_ASAP7_75t_SL U54250 ( .A1(n77397), .A2(n77396), .B1(n2600), .B2(
        n77454), .Y(n9457) );
  OAI21xp33_ASAP7_75t_SL U54251 ( .A1(n74740), .A2(n74739), .B(n74738), .Y(
        n2899) );
  INVxp67_ASAP7_75t_SL U54252 ( .A(n68587), .Y(n68590) );
  OAI21xp33_ASAP7_75t_SL U54253 ( .A1(n58316), .A2(n4091), .B(n78046), .Y(
        n9705) );
  OA21x2_ASAP7_75t_SL U54254 ( .A1(n59688), .A2(n75888), .B(n75889), .Y(n75887) );
  OAI21xp33_ASAP7_75t_SL U54255 ( .A1(n58316), .A2(n4090), .B(n78048), .Y(
        n9704) );
  OAI21xp33_ASAP7_75t_SL U54256 ( .A1(n58316), .A2(n4089), .B(n78050), .Y(
        n9703) );
  OAI21xp33_ASAP7_75t_SL U54257 ( .A1(n58316), .A2(n4138), .B(n78052), .Y(
        n9702) );
  NAND2xp5_ASAP7_75t_SL U54258 ( .A(n77507), .B(n77795), .Y(n77508) );
  INVxp33_ASAP7_75t_SL U54259 ( .A(n77363), .Y(n60446) );
  AOI22xp5_ASAP7_75t_SL U54260 ( .A1(n77799), .A2(n77802), .B1(n77798), .B2(
        n77797), .Y(n77800) );
  OAI21xp5_ASAP7_75t_SL U54261 ( .A1(n815), .A2(n77385), .B(n63988), .Y(n9181)
         );
  OAI21xp33_ASAP7_75t_SL U54262 ( .A1(n58316), .A2(n4136), .B(n78061), .Y(
        n9700) );
  OAI21xp5_ASAP7_75t_SL U54263 ( .A1(n775), .A2(n77385), .B(n65194), .Y(n9171)
         );
  OAI21xp5_ASAP7_75t_SL U54264 ( .A1(n763), .A2(n77385), .B(n75172), .Y(n9168)
         );
  OAI21xp5_ASAP7_75t_SL U54265 ( .A1(n819), .A2(n77385), .B(n63985), .Y(n9182)
         );
  AOI21xp33_ASAP7_75t_SL U54266 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[25]), .A2(n70502), .B(
        n70100), .Y(n2265) );
  AOI22xp33_ASAP7_75t_SL U54267 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[26]), .A2(n70502), .B1(
        n59621), .B2(n70102), .Y(n2263) );
  NAND2x1p5_ASAP7_75t_SL U54268 ( .A(n64987), .B(n64986), .Y(n68758) );
  NAND2xp33_ASAP7_75t_SL U54269 ( .A(n77386), .B(n77388), .Y(n75637) );
  NAND2xp33_ASAP7_75t_SL U54270 ( .A(n59678), .B(n77863), .Y(n77188) );
  AO21x1_ASAP7_75t_SL U54271 ( .A1(n63348), .A2(n63347), .B(n63369), .Y(n63349) );
  NAND2xp5_ASAP7_75t_SL U54272 ( .A(n66581), .B(n66580), .Y(n69293) );
  AOI22xp33_ASAP7_75t_SL U54273 ( .A1(n73610), .A2(n73592), .B1(n73591), .B2(
        n73607), .Y(n1525) );
  OAI22xp33_ASAP7_75t_SL U54274 ( .A1(n74249), .A2(n74503), .B1(n74248), .B2(
        n58298), .Y(n74251) );
  INVx1_ASAP7_75t_SL U54275 ( .A(n77884), .Y(n74638) );
  OAI21xp5_ASAP7_75t_SL U54276 ( .A1(n77796), .A2(n60285), .B(n60284), .Y(
        n9475) );
  OAI21xp33_ASAP7_75t_SL U54277 ( .A1(n77467), .A2(n74110), .B(n74109), .Y(
        n9645) );
  INVx1_ASAP7_75t_SL U54278 ( .A(n77865), .Y(n75805) );
  AOI21xp33_ASAP7_75t_SL U54279 ( .A1(n68638), .A2(n68637), .B(n68636), .Y(
        n68640) );
  NAND2x1p5_ASAP7_75t_SL U54280 ( .A(n57043), .B(n63160), .Y(n63257) );
  OAI21xp33_ASAP7_75t_SL U54281 ( .A1(n2585), .A2(n77567), .B(n61160), .Y(
        n9608) );
  NAND2xp5_ASAP7_75t_SL U54282 ( .A(n76239), .B(n76238), .Y(
        or1200_cpu_or1200_except_n1736) );
  OAI22xp33_ASAP7_75t_SL U54283 ( .A1(n2688), .A2(n77145), .B1(n77144), .B2(
        n77143), .Y(n77146) );
  NAND2xp33_ASAP7_75t_SL U54284 ( .A(n59678), .B(n77889), .Y(n75384) );
  INVxp67_ASAP7_75t_SL U54285 ( .A(n70210), .Y(n51958) );
  OAI21xp33_ASAP7_75t_SL U54286 ( .A1(n845), .A2(n77276), .B(n61588), .Y(
        or1200_cpu_or1200_except_n587) );
  OAI21xp33_ASAP7_75t_SL U54287 ( .A1(n964), .A2(n77276), .B(n65196), .Y(
        or1200_cpu_or1200_except_n650) );
  OAI21xp33_ASAP7_75t_SL U54288 ( .A1(n937), .A2(n77276), .B(n75422), .Y(
        or1200_cpu_or1200_except_n641) );
  OAI21xp33_ASAP7_75t_SL U54289 ( .A1(n1099), .A2(n77276), .B(n63699), .Y(
        or1200_cpu_or1200_except_n608) );
  INVxp67_ASAP7_75t_SL U54290 ( .A(n68624), .Y(n66534) );
  OAI21xp33_ASAP7_75t_SL U54291 ( .A1(n1110), .A2(n77276), .B(n76535), .Y(
        or1200_cpu_or1200_except_n611) );
  OAI21xp33_ASAP7_75t_SL U54292 ( .A1(n1009), .A2(n77276), .B(n75187), .Y(
        or1200_cpu_or1200_except_n665) );
  INVxp33_ASAP7_75t_SL U54293 ( .A(n61038), .Y(n60447) );
  NAND2xp5_ASAP7_75t_SL U54294 ( .A(n62158), .B(n62157), .Y(
        or1200_cpu_or1200_except_n1751) );
  NAND2xp5_ASAP7_75t_SL U54295 ( .A(n75147), .B(n75146), .Y(
        or1200_cpu_or1200_except_n1738) );
  NAND2xp5_ASAP7_75t_SL U54296 ( .A(n63766), .B(n63765), .Y(
        or1200_cpu_or1200_except_n1750) );
  NAND2xp33_ASAP7_75t_SL U54297 ( .A(n78060), .B(n58434), .Y(n78057) );
  OAI21xp33_ASAP7_75t_SL U54298 ( .A1(n1033), .A2(n77276), .B(n61576), .Y(
        or1200_cpu_or1200_except_n590) );
  INVxp33_ASAP7_75t_SL U54299 ( .A(n68635), .Y(n68638) );
  NAND2xp5_ASAP7_75t_SL U54300 ( .A(n77222), .B(n77221), .Y(
        or1200_cpu_or1200_except_n1739) );
  OAI21xp33_ASAP7_75t_SL U54301 ( .A1(n1027), .A2(n77276), .B(n76918), .Y(
        or1200_cpu_or1200_except_n671) );
  OAI21xp33_ASAP7_75t_SL U54302 ( .A1(n955), .A2(n77276), .B(n75547), .Y(
        or1200_cpu_or1200_except_n647) );
  OAI21xp33_ASAP7_75t_SL U54303 ( .A1(n1088), .A2(n77276), .B(n61279), .Y(
        or1200_cpu_or1200_except_n605) );
  NAND2xp5_ASAP7_75t_SL U54304 ( .A(n75535), .B(n75534), .Y(
        or1200_cpu_or1200_except_n1740) );
  NAND2xp5_ASAP7_75t_SL U54305 ( .A(n76868), .B(n76867), .Y(
        or1200_cpu_or1200_except_n1749) );
  OAI21xp33_ASAP7_75t_SL U54306 ( .A1(n946), .A2(n77276), .B(n64268), .Y(
        or1200_cpu_or1200_except_n644) );
  OAI21xp33_ASAP7_75t_SL U54307 ( .A1(n1066), .A2(n77276), .B(n63740), .Y(
        or1200_cpu_or1200_except_n599) );
  NAND2xp5_ASAP7_75t_SL U54308 ( .A(n77004), .B(n77003), .Y(
        or1200_cpu_or1200_except_n1748) );
  NAND2xp5_ASAP7_75t_SL U54309 ( .A(n76651), .B(n76650), .Y(
        or1200_cpu_or1200_except_n1744) );
  OAI21xp33_ASAP7_75t_SL U54310 ( .A1(n1055), .A2(n77276), .B(n76608), .Y(
        or1200_cpu_or1200_except_n596) );
  NAND2xp5_ASAP7_75t_SL U54311 ( .A(n76710), .B(n76709), .Y(
        or1200_cpu_or1200_except_n1745) );
  NAND2xp5_ASAP7_75t_SL U54312 ( .A(n76625), .B(n76624), .Y(
        or1200_cpu_or1200_except_n1746) );
  NAND2xp5_ASAP7_75t_SL U54313 ( .A(n76219), .B(n76218), .Y(
        or1200_cpu_or1200_except_n1747) );
  NAND2xp33_ASAP7_75t_SL U54314 ( .A(n78053), .B(n58434), .Y(n78052) );
  NAND2xp5_ASAP7_75t_SL U54315 ( .A(n64806), .B(n64805), .Y(n77872) );
  OAI21xp33_ASAP7_75t_SL U54316 ( .A1(n910), .A2(n77276), .B(n74971), .Y(
        or1200_cpu_or1200_except_n632) );
  AOI21xp33_ASAP7_75t_SL U54317 ( .A1(n66565), .A2(n68635), .B(n66564), .Y(
        n66581) );
  OAI21xp33_ASAP7_75t_SL U54318 ( .A1(n77467), .A2(n77857), .B(n77466), .Y(
        n9640) );
  NAND2xp33_ASAP7_75t_SL U54319 ( .A(n78064), .B(n58434), .Y(n78063) );
  OAI21xp33_ASAP7_75t_SL U54320 ( .A1(n919), .A2(n77276), .B(n64016), .Y(
        or1200_cpu_or1200_except_n635) );
  NAND2xp33_ASAP7_75t_SL U54321 ( .A(n78047), .B(n58434), .Y(n78046) );
  NAND2xp5_ASAP7_75t_SL U54322 ( .A(n61989), .B(n61988), .Y(n77855) );
  NAND2xp33_ASAP7_75t_SL U54323 ( .A(n78049), .B(n58434), .Y(n78048) );
  OAI21xp33_ASAP7_75t_SL U54324 ( .A1(n892), .A2(n77276), .B(n64007), .Y(
        or1200_cpu_or1200_except_n626) );
  OAI21xp33_ASAP7_75t_SL U54325 ( .A1(n74424), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_41_), .B(
        n74433), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n38) );
  AOI21xp5_ASAP7_75t_SL U54326 ( .A1(n76820), .A2(
        or1200_cpu_or1200_genpc_pcreg_default[6]), .B(n61177), .Y(n1050) );
  OAI21xp33_ASAP7_75t_SL U54327 ( .A1(n973), .A2(n77276), .B(n65223), .Y(
        or1200_cpu_or1200_except_n653) );
  INVxp67_ASAP7_75t_SL U54328 ( .A(n66604), .Y(n66599) );
  OAI21xp33_ASAP7_75t_SL U54329 ( .A1(n982), .A2(n77276), .B(n65235), .Y(
        or1200_cpu_or1200_except_n656) );
  OAI21xp33_ASAP7_75t_SL U54330 ( .A1(n883), .A2(n77276), .B(n63999), .Y(
        or1200_cpu_or1200_except_n623) );
  AOI21xp5_ASAP7_75t_SL U54331 ( .A1(n76820), .A2(
        or1200_cpu_or1200_genpc_pcreg_default[4]), .B(n76595), .Y(n1028) );
  NAND2xp33_ASAP7_75t_SL U54332 ( .A(n78062), .B(n58434), .Y(n78061) );
  INVxp67_ASAP7_75t_SL U54333 ( .A(n73652), .Y(n73607) );
  NAND2xp5_ASAP7_75t_SL U54334 ( .A(n60362), .B(n60361), .Y(n9236) );
  NOR2x1_ASAP7_75t_SL U54335 ( .A(n58618), .B(n75180), .Y(n77388) );
  NAND2xp5_ASAP7_75t_SL U54336 ( .A(n60342), .B(n61160), .Y(n9464) );
  OAI21xp33_ASAP7_75t_SL U54337 ( .A1(n839), .A2(n77276), .B(n63749), .Y(
        or1200_cpu_or1200_except_n584) );
  NAND2xp33_ASAP7_75t_SL U54338 ( .A(n52493), .B(n52492), .Y(n74912) );
  OAI21xp33_ASAP7_75t_SL U54339 ( .A1(n991), .A2(n77276), .B(n75150), .Y(
        or1200_cpu_or1200_except_n659) );
  OAI21xp33_ASAP7_75t_SL U54340 ( .A1(n928), .A2(n77276), .B(n64166), .Y(
        or1200_cpu_or1200_except_n638) );
  NAND2xp33_ASAP7_75t_SL U54341 ( .A(n78051), .B(n58434), .Y(n78050) );
  OAI21xp33_ASAP7_75t_SL U54342 ( .A1(n856), .A2(n77276), .B(n63946), .Y(
        or1200_cpu_or1200_except_n614) );
  AOI21xp5_ASAP7_75t_SL U54343 ( .A1(n76820), .A2(
        or1200_cpu_or1200_genpc_pcreg_default[7]), .B(n76819), .Y(n1061) );
  OAI21xp33_ASAP7_75t_SL U54344 ( .A1(n1000), .A2(n77276), .B(n75164), .Y(
        or1200_cpu_or1200_except_n662) );
  OA21x2_ASAP7_75t_SL U54345 ( .A1(n59688), .A2(n75376), .B(n75377), .Y(n75375) );
  INVxp67_ASAP7_75t_SL U54346 ( .A(n77870), .Y(n74110) );
  NAND2xp33_ASAP7_75t_SL U54347 ( .A(n78162), .B(n58434), .Y(n78161) );
  NAND2xp5_ASAP7_75t_SL U54348 ( .A(n60288), .B(n77796), .Y(n60284) );
  INVxp67_ASAP7_75t_SL U54349 ( .A(n60289), .Y(n9476) );
  NAND2xp33_ASAP7_75t_SL U54350 ( .A(n77187), .B(n77186), .Y(n77863) );
  NAND2xp5_ASAP7_75t_SL U54351 ( .A(n75273), .B(n75272), .Y(n9610) );
  INVx1_ASAP7_75t_SL U54352 ( .A(n68643), .Y(n68644) );
  INVxp67_ASAP7_75t_SL U54353 ( .A(n61046), .Y(n61047) );
  OAI21xp33_ASAP7_75t_SL U54354 ( .A1(n77137), .A2(n77857), .B(n75758), .Y(
        n9609) );
  OAI21xp33_ASAP7_75t_SL U54355 ( .A1(n847), .A2(n76523), .B(n63957), .Y(n9184) );
  INVxp67_ASAP7_75t_SL U54356 ( .A(n74258), .Y(n74266) );
  AOI21xp5_ASAP7_75t_SL U54357 ( .A1(n76820), .A2(
        or1200_cpu_or1200_genpc_pcreg_default[3]), .B(n58545), .Y(n840) );
  INVxp67_ASAP7_75t_SL U54358 ( .A(n64150), .Y(n62095) );
  NAND2xp5_ASAP7_75t_SL U54359 ( .A(n74028), .B(n74027), .Y(n76323) );
  NAND2xp33_ASAP7_75t_SL U54360 ( .A(n77395), .B(n77394), .Y(n77396) );
  AOI21xp5_ASAP7_75t_SL U54361 ( .A1(n76820), .A2(
        or1200_cpu_or1200_genpc_pcreg_default[2]), .B(n76571), .Y(n826) );
  OAI22xp33_ASAP7_75t_SL U54362 ( .A1(n69334), .A2(n69333), .B1(
        or1200_cpu_or1200_except_n677), .B2(n77454), .Y(
        or1200_cpu_or1200_except_n1830) );
  OAI21xp33_ASAP7_75t_SL U54363 ( .A1(n2596), .A2(n77454), .B(n60332), .Y(
        n9574) );
  OAI21xp33_ASAP7_75t_SL U54364 ( .A1(n77467), .A2(n77860), .B(n76854), .Y(
        n9641) );
  OR2x2_ASAP7_75t_SL U54365 ( .A(n69354), .B(n77235), .Y(n77298) );
  INVx1_ASAP7_75t_SL U54366 ( .A(n77235), .Y(n77296) );
  INVxp67_ASAP7_75t_SL U54367 ( .A(n77796), .Y(n77797) );
  INVxp33_ASAP7_75t_SL U54368 ( .A(n75111), .Y(n75089) );
  AOI22xp33_ASAP7_75t_SL U54369 ( .A1(n77220), .A2(n78260), .B1(n77920), .B2(
        n76707), .Y(n62158) );
  INVxp33_ASAP7_75t_SL U54370 ( .A(n77249), .Y(n77265) );
  AOI22xp33_ASAP7_75t_SL U54371 ( .A1(n77220), .A2(n78253), .B1(n77918), .B2(
        n76707), .Y(n63766) );
  INVxp67_ASAP7_75t_SL U54372 ( .A(n75041), .Y(n68642) );
  AOI22xp33_ASAP7_75t_SL U54373 ( .A1(dc_en), .A2(n77220), .B1(n77916), .B2(
        n77218), .Y(n76868) );
  AOI22xp33_ASAP7_75t_SL U54374 ( .A1(n77217), .A2(or1200_cpu_to_sr[3]), .B1(
        n76866), .B2(n77215), .Y(n76867) );
  NAND2xp5_ASAP7_75t_SL U54375 ( .A(n75615), .B(n75614), .Y(n9616) );
  AOI22xp33_ASAP7_75t_SL U54376 ( .A1(ic_en), .A2(n77220), .B1(n77974), .B2(
        n77218), .Y(n77004) );
  OAI22xp33_ASAP7_75t_SL U54377 ( .A1(n76537), .A2(n76536), .B1(n2033), .B2(
        n77567), .Y(n9569) );
  AOI22xp33_ASAP7_75t_SL U54378 ( .A1(n77217), .A2(or1200_cpu_to_sr[4]), .B1(
        n77002), .B2(n77215), .Y(n77003) );
  NAND2xp5_ASAP7_75t_SL U54379 ( .A(n74631), .B(n74630), .Y(n74634) );
  AOI22xp33_ASAP7_75t_SL U54380 ( .A1(n77220), .A2(n76216), .B1(n77977), .B2(
        n76707), .Y(n76219) );
  AOI22xp33_ASAP7_75t_SL U54381 ( .A1(n77217), .A2(or1200_cpu_to_sr[5]), .B1(
        n76217), .B2(n77215), .Y(n76218) );
  OAI21xp33_ASAP7_75t_SL U54382 ( .A1(or1200_cpu_or1200_if_insn_saved[26]), 
        .A2(n59683), .B(n60319), .Y(n2696) );
  NAND2xp33_ASAP7_75t_SL U54383 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[6]), .B(
        n70600), .Y(n70606) );
  AOI22xp33_ASAP7_75t_SL U54384 ( .A1(n77220), .A2(n76622), .B1(n77980), .B2(
        n76707), .Y(n76625) );
  OAI21xp33_ASAP7_75t_SL U54385 ( .A1(n77467), .A2(n77886), .B(n74990), .Y(
        n9652) );
  AOI22xp33_ASAP7_75t_SL U54386 ( .A1(n77217), .A2(or1200_cpu_to_sr[6]), .B1(
        n76623), .B2(n77215), .Y(n76624) );
  AOI22xp33_ASAP7_75t_SL U54387 ( .A1(n77220), .A2(n76736), .B1(n77983), .B2(
        n76707), .Y(n76710) );
  AOI22xp33_ASAP7_75t_SL U54388 ( .A1(n77217), .A2(or1200_cpu_to_sr[7]), .B1(
        n76708), .B2(n77215), .Y(n76709) );
  AOI22xp33_ASAP7_75t_SL U54389 ( .A1(n77220), .A2(n76648), .B1(n77986), .B2(
        n76707), .Y(n76651) );
  AOI22xp33_ASAP7_75t_SL U54390 ( .A1(n77217), .A2(or1200_cpu_to_sr[8]), .B1(
        n76649), .B2(n77215), .Y(n76650) );
  OAI21xp33_ASAP7_75t_SL U54391 ( .A1(n1075), .A2(n53428), .B(n76850), .Y(
        or1200_cpu_or1200_except_n602) );
  AOI21xp33_ASAP7_75t_SL U54392 ( .A1(n77220), .A2(n74034), .B(n74033), .Y(
        n74035) );
  INVxp67_ASAP7_75t_SL U54393 ( .A(n61050), .Y(n60332) );
  AOI22xp33_ASAP7_75t_SL U54394 ( .A1(n77220), .A2(n75532), .B1(n77901), .B2(
        n76707), .Y(n75535) );
  AOI22xp33_ASAP7_75t_SL U54395 ( .A1(n77217), .A2(or1200_cpu_to_sr[12]), .B1(
        n75533), .B2(n77215), .Y(n75534) );
  AOI22xp33_ASAP7_75t_SL U54396 ( .A1(n77217), .A2(or1200_cpu_to_sr[13]), .B1(
        n77216), .B2(n77215), .Y(n77222) );
  AOI21xp33_ASAP7_75t_SL U54397 ( .A1(n77843), .A2(n78440), .B(n77952), .Y(
        n77844) );
  AOI22xp33_ASAP7_75t_SL U54398 ( .A1(n77220), .A2(n77219), .B1(n77899), .B2(
        n77218), .Y(n77221) );
  AOI22xp33_ASAP7_75t_SL U54399 ( .A1(n75144), .A2(n77220), .B1(n77217), .B2(
        n75148), .Y(n75147) );
  AOI22xp33_ASAP7_75t_SL U54400 ( .A1(n77896), .A2(n76707), .B1(n75145), .B2(
        n77215), .Y(n75146) );
  NAND2xp5_ASAP7_75t_SL U54401 ( .A(n73356), .B(n73355), .Y(n51957) );
  NAND2xp33_ASAP7_75t_SL U54402 ( .A(n71082), .B(n71057), .Y(n71060) );
  OAI21xp33_ASAP7_75t_SL U54403 ( .A1(n77467), .A2(n77867), .B(n73904), .Y(
        n9644) );
  OAI21xp33_ASAP7_75t_SL U54404 ( .A1(n77137), .A2(n77867), .B(n64868), .Y(
        n9613) );
  NAND2xp5_ASAP7_75t_SL U54405 ( .A(n60499), .B(n60498), .Y(n9466) );
  INVxp33_ASAP7_75t_SL U54406 ( .A(n68556), .Y(n68557) );
  NAND2xp5_ASAP7_75t_SL U54407 ( .A(n77159), .B(n77158), .Y(n9655) );
  NAND2xp5_ASAP7_75t_SL U54408 ( .A(n60892), .B(n60891), .Y(n9450) );
  NAND2xp5_ASAP7_75t_SL U54409 ( .A(n61590), .B(n61589), .Y(n9449) );
  OAI22xp33_ASAP7_75t_SL U54410 ( .A1(n2054), .A2(n76536), .B1(n2035), .B2(
        n77567), .Y(n9570) );
  NAND2xp5_ASAP7_75t_SL U54411 ( .A(n61023), .B(n61022), .Y(n9448) );
  OAI21xp33_ASAP7_75t_SL U54412 ( .A1(n60434), .A2(n77423), .B(n60433), .Y(
        n9424) );
  INVx1_ASAP7_75t_SL U54413 ( .A(n70600), .Y(n70608) );
  NAND2xp5_ASAP7_75t_SL U54414 ( .A(n60396), .B(n60395), .Y(n9445) );
  NAND2xp5_ASAP7_75t_SL U54415 ( .A(n77372), .B(n77371), .Y(n9444) );
  NAND2xp5_ASAP7_75t_SL U54416 ( .A(n78024), .B(n78023), .Y(n9443) );
  NAND2xp5_ASAP7_75t_SL U54417 ( .A(n78018), .B(n78017), .Y(n9442) );
  OAI21xp33_ASAP7_75t_SL U54418 ( .A1(n3423), .A2(n77567), .B(n77461), .Y(
        n9460) );
  NAND2xp5_ASAP7_75t_SL U54419 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[0]), .B(
        n70600), .Y(n70575) );
  NAND2xp5_ASAP7_75t_SL U54420 ( .A(n78015), .B(n78014), .Y(n9441) );
  NAND2xp5_ASAP7_75t_SL U54421 ( .A(n78012), .B(n78011), .Y(n9440) );
  AO21x1_ASAP7_75t_SL U54422 ( .A1(n77354), .A2(n77353), .B(n77352), .Y(n77355) );
  NAND2xp5_ASAP7_75t_SL U54423 ( .A(n78008), .B(n78007), .Y(n9439) );
  OAI21xp33_ASAP7_75t_SL U54424 ( .A1(n60513), .A2(n77423), .B(n60512), .Y(
        n9437) );
  OAI21xp33_ASAP7_75t_SL U54425 ( .A1(n60533), .A2(n77423), .B(n60532), .Y(
        n9436) );
  OAI21xp33_ASAP7_75t_SL U54426 ( .A1(n60520), .A2(n77423), .B(n60519), .Y(
        n9435) );
  INVxp33_ASAP7_75t_SL U54427 ( .A(n64147), .Y(n64148) );
  OAI21xp33_ASAP7_75t_SL U54428 ( .A1(n60528), .A2(n77423), .B(n60527), .Y(
        n9434) );
  NAND2xp5_ASAP7_75t_SL U54429 ( .A(n60419), .B(n60418), .Y(n9433) );
  NAND2xp5_ASAP7_75t_SL U54430 ( .A(n60411), .B(n60410), .Y(n9431) );
  INVxp67_ASAP7_75t_SL U54431 ( .A(n68625), .Y(n66523) );
  NAND2xp5_ASAP7_75t_SL U54432 ( .A(n60481), .B(n60480), .Y(n9430) );
  NAND2xp5_ASAP7_75t_SL U54433 ( .A(n60472), .B(n60471), .Y(n9429) );
  INVxp33_ASAP7_75t_SL U54434 ( .A(n64804), .Y(n64805) );
  OAI21xp33_ASAP7_75t_SL U54435 ( .A1(n60331), .A2(n77423), .B(n60329), .Y(
        n9427) );
  OAI21xp33_ASAP7_75t_SL U54436 ( .A1(n77406), .A2(n77423), .B(n77405), .Y(
        n9425) );
  AOI22xp33_ASAP7_75t_SL U54437 ( .A1(n77376), .A2(n2609), .B1(n60456), .B2(
        n77456), .Y(n9575) );
  NOR2x1_ASAP7_75t_SL U54438 ( .A(n75158), .B(n75159), .Y(n75180) );
  INVxp67_ASAP7_75t_SL U54439 ( .A(n75975), .Y(n75973) );
  NAND2xp5_ASAP7_75t_SL U54440 ( .A(n71131), .B(n71137), .Y(n71099) );
  INVxp67_ASAP7_75t_SL U54441 ( .A(n68626), .Y(n66524) );
  INVxp33_ASAP7_75t_SL U54442 ( .A(n60462), .Y(n60463) );
  INVxp67_ASAP7_75t_SL U54443 ( .A(n77217), .Y(n77145) );
  BUFx2_ASAP7_75t_SL U54444 ( .A(n68329), .Y(n57420) );
  AOI22xp33_ASAP7_75t_SL U54445 ( .A1(n59701), .A2(n65193), .B1(n65192), .B2(
        n53441), .Y(n65194) );
  AND2x2_ASAP7_75t_SL U54446 ( .A(n74868), .B(n74867), .Y(n74869) );
  OAI21xp33_ASAP7_75t_SL U54447 ( .A1(n77947), .A2(n57090), .B(n60517), .Y(
        n9588) );
  OAI21xp5_ASAP7_75t_SL U54448 ( .A1(n70942), .A2(n70941), .B(n70940), .Y(
        n70948) );
  NAND2xp5_ASAP7_75t_SL U54449 ( .A(n74842), .B(n74841), .Y(n52498) );
  OAI21xp33_ASAP7_75t_SL U54450 ( .A1(or1200_cpu_or1200_if_insn_saved[28]), 
        .A2(n59683), .B(n77361), .Y(n2694) );
  OAI21xp33_ASAP7_75t_SL U54451 ( .A1(n77424), .A2(n77423), .B(n77422), .Y(
        n9423) );
  AOI22xp33_ASAP7_75t_SL U54452 ( .A1(dbg_dat_i[10]), .A2(n76521), .B1(n74947), 
        .B2(n53441), .Y(n74948) );
  INVxp67_ASAP7_75t_SL U54453 ( .A(n59156), .Y(n58280) );
  OAI22xp33_ASAP7_75t_SL U54454 ( .A1(n57090), .A2(n60535), .B1(n2671), .B2(
        n77454), .Y(n9587) );
  AND2x2_ASAP7_75t_SL U54455 ( .A(n76953), .B(n74858), .Y(n74853) );
  OAI21xp33_ASAP7_75t_SL U54456 ( .A1(n77938), .A2(n57090), .B(n60525), .Y(
        n9586) );
  NAND2xp5_ASAP7_75t_SL U54457 ( .A(n75630), .B(n75629), .Y(n9647) );
  INVxp67_ASAP7_75t_SL U54458 ( .A(n64720), .Y(n59154) );
  OAI22xp33_ASAP7_75t_SL U54459 ( .A1(n78055), .A2(n76846), .B1(n1075), .B2(
        n59682), .Y(n9416) );
  OAI21xp33_ASAP7_75t_SL U54460 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_16_), .A2(n77171), 
        .B(n74860), .Y(n74864) );
  OAI22xp33_ASAP7_75t_SL U54461 ( .A1(n57090), .A2(n60530), .B1(n2685), .B2(
        n77454), .Y(n9585) );
  NAND2xp5_ASAP7_75t_SL U54462 ( .A(n75521), .B(n75520), .Y(n75527) );
  NAND2xp5_ASAP7_75t_SL U54463 ( .A(n61151), .B(n61150), .Y(n51982) );
  NAND2xp5_ASAP7_75t_SL U54464 ( .A(n59499), .B(n76314), .Y(n77186) );
  OAI21xp33_ASAP7_75t_SL U54465 ( .A1(n1073), .A2(n76839), .B(n76838), .Y(
        n9188) );
  NAND2xp5_ASAP7_75t_SL U54466 ( .A(n76223), .B(n76222), .Y(n9665) );
  INVxp33_ASAP7_75t_SL U54467 ( .A(n77350), .Y(n77342) );
  OAI21xp5_ASAP7_75t_SL U54468 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_21_), .A2(n74876), 
        .B(n74874), .Y(n52497) );
  AOI22xp33_ASAP7_75t_SL U54469 ( .A1(n59701), .A2(n63956), .B1(n63955), .B2(
        n53441), .Y(n63957) );
  NAND2xp33_ASAP7_75t_SL U54470 ( .A(n75383), .B(n75382), .Y(n77889) );
  AOI22xp33_ASAP7_75t_SL U54471 ( .A1(n77217), .A2(n78187), .B1(n76236), .B2(
        n77215), .Y(n76239) );
  AOI21xp5_ASAP7_75t_SL U54472 ( .A1(n70941), .A2(n70923), .B(n70938), .Y(
        n70925) );
  AOI22xp33_ASAP7_75t_SL U54473 ( .A1(dbg_dat_i[9]), .A2(n76521), .B1(n76520), 
        .B2(n53441), .Y(n76522) );
  AOI22xp33_ASAP7_75t_SL U54474 ( .A1(n77220), .A2(n76237), .B1(n77890), .B2(
        n77218), .Y(n76238) );
  AOI21xp33_ASAP7_75t_SL U54475 ( .A1(n77376), .A2(n2814), .B(n77395), .Y(
        n51945) );
  OAI21xp33_ASAP7_75t_SL U54476 ( .A1(n74458), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_25_), .B(
        n74457), .Y(n2953) );
  NAND2xp5_ASAP7_75t_SL U54477 ( .A(n70203), .B(n70209), .Y(n3254) );
  AND3x1_ASAP7_75t_SL U54478 ( .A(n74494), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_27_), 
        .C(n74507), .Y(n74452) );
  OA21x2_ASAP7_75t_SL U54479 ( .A1(n75469), .A2(n75462), .B(n75461), .Y(n75463) );
  INVxp67_ASAP7_75t_SL U54480 ( .A(n66525), .Y(n66528) );
  OAI21xp33_ASAP7_75t_SL U54481 ( .A1(n70199), .A2(n70198), .B(n70209), .Y(
        n3256) );
  NOR2x1_ASAP7_75t_SL U54482 ( .A(n73863), .B(n73862), .Y(n74418) );
  AOI21xp33_ASAP7_75t_SL U54483 ( .A1(n74899), .A2(n76933), .B(n74885), .Y(
        n74874) );
  NAND2xp5_ASAP7_75t_SL U54484 ( .A(n75060), .B(n57842), .Y(n75102) );
  INVx1_ASAP7_75t_SL U54485 ( .A(n57842), .Y(n75061) );
  AOI22xp33_ASAP7_75t_SL U54486 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_8_), .A2(n74905), 
        .B1(n76944), .B2(n74904), .Y(n74906) );
  OAI21xp33_ASAP7_75t_SL U54487 ( .A1(n74308), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_39_), .B(
        n74415), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n34) );
  INVxp33_ASAP7_75t_SL U54488 ( .A(n74872), .Y(n74849) );
  NOR2x1_ASAP7_75t_SL U54489 ( .A(n68324), .B(n68323), .Y(n68332) );
  NAND2xp5_ASAP7_75t_SL U54490 ( .A(n76934), .B(n74899), .Y(n74870) );
  AOI22xp33_ASAP7_75t_SL U54491 ( .A1(n60432), .A2(n57089), .B1(
        or1200_ic_top_from_icram[30]), .B2(n59497), .Y(n60433) );
  OAI21xp5_ASAP7_75t_SL U54492 ( .A1(n59677), .A2(n76562), .B(n76561), .Y(
        n9628) );
  NAND2xp5_ASAP7_75t_SL U54493 ( .A(n74851), .B(n74899), .Y(n74854) );
  INVxp67_ASAP7_75t_SL U54494 ( .A(n63104), .Y(n63102) );
  OA21x2_ASAP7_75t_SL U54495 ( .A1(n57074), .A2(n77156), .B(n77157), .Y(n77129) );
  NAND2xp5_ASAP7_75t_SL U54496 ( .A(n64332), .B(n64331), .Y(n9617) );
  XNOR2xp5_ASAP7_75t_SL U54497 ( .A(n64696), .B(n64695), .Y(n64697) );
  XNOR2xp5_ASAP7_75t_SL U54498 ( .A(n68193), .B(n68192), .Y(n68334) );
  INVxp67_ASAP7_75t_SL U54499 ( .A(n68323), .Y(n68226) );
  AOI21xp33_ASAP7_75t_SL U54500 ( .A1(n74899), .A2(n74902), .B(n74885), .Y(
        n74842) );
  INVxp67_ASAP7_75t_SL U54501 ( .A(n68324), .Y(n68225) );
  AOI22xp33_ASAP7_75t_SL U54502 ( .A1(n57090), .A2(n76849), .B1(n76848), .B2(
        n76847), .Y(n76850) );
  AOI22xp33_ASAP7_75t_SL U54503 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_1_), .A2(n74882), 
        .B1(n74901), .B2(n74881), .Y(n77170) );
  OAI22xp33_ASAP7_75t_SL U54504 ( .A1(n77583), .A2(n76661), .B1(n76660), .B2(
        n76659), .Y(n76667) );
  NAND2xp33_ASAP7_75t_SL U54505 ( .A(n74929), .B(n77442), .Y(n74930) );
  OAI21xp33_ASAP7_75t_SL U54506 ( .A1(n77954), .A2(n60448), .B(n60441), .Y(
        n60462) );
  AOI22xp33_ASAP7_75t_SL U54507 ( .A1(n77376), .A2(n60516), .B1(
        or1200_ic_top_from_icram[17]), .B2(n53436), .Y(n60517) );
  INVxp67_ASAP7_75t_SL U54508 ( .A(n77946), .Y(n60535) );
  AOI22xp33_ASAP7_75t_SL U54509 ( .A1(n77376), .A2(n60524), .B1(
        or1200_ic_top_from_icram[19]), .B2(n53436), .Y(n60525) );
  INVxp67_ASAP7_75t_SL U54510 ( .A(n76191), .Y(n76186) );
  AOI21xp5_ASAP7_75t_SL U54511 ( .A1(n76313), .A2(n59499), .B(n63600), .Y(
        n77886) );
  INVxp67_ASAP7_75t_SL U54512 ( .A(n77936), .Y(n60530) );
  NAND2xp33_ASAP7_75t_SL U54513 ( .A(n58083), .B(n76221), .Y(n76222) );
  NAND2xp33_ASAP7_75t_SL U54514 ( .A(n74944), .B(n77442), .Y(n74945) );
  OAI21xp33_ASAP7_75t_SL U54515 ( .A1(n77954), .A2(n77948), .B(n77947), .Y(
        n77951) );
  OAI21xp33_ASAP7_75t_SL U54516 ( .A1(n77954), .A2(n77939), .B(n77938), .Y(
        n77942) );
  AOI22xp33_ASAP7_75t_SL U54517 ( .A1(n77421), .A2(n59685), .B1(
        or1200_ic_top_from_icram[31]), .B2(n59497), .Y(n77422) );
  AOI21xp33_ASAP7_75t_SL U54518 ( .A1(n65277), .A2(n65308), .B(n2900), .Y(
        n65276) );
  INVxp67_ASAP7_75t_SL U54519 ( .A(n71301), .Y(n71257) );
  AOI22xp33_ASAP7_75t_SL U54520 ( .A1(n77376), .A2(n69335), .B1(n60354), .B2(
        n77374), .Y(n60355) );
  NAND2xp33_ASAP7_75t_SL U54521 ( .A(iwb_dat_i[3]), .B(n77373), .Y(n60356) );
  NAND2xp33_ASAP7_75t_SL U54522 ( .A(or1200_cpu_or1200_if_insn_saved[22]), .B(
        n77374), .Y(n60407) );
  INVx2_ASAP7_75t_SL U54523 ( .A(n59685), .Y(n59683) );
  NAND2xp33_ASAP7_75t_SL U54524 ( .A(iwb_dat_i[10]), .B(n77373), .Y(n77378) );
  AOI22xp33_ASAP7_75t_SL U54525 ( .A1(n77376), .A2(n77381), .B1(n77375), .B2(
        n77374), .Y(n77377) );
  NAND2xp33_ASAP7_75t_SL U54526 ( .A(iwb_dat_i[9]), .B(n77373), .Y(n60399) );
  NAND2xp33_ASAP7_75t_SL U54527 ( .A(n59678), .B(n77874), .Y(n75614) );
  AOI22xp33_ASAP7_75t_SL U54528 ( .A1(n77376), .A2(n61161), .B1(n60397), .B2(
        n77374), .Y(n60398) );
  INVx2_ASAP7_75t_SL U54529 ( .A(n59685), .Y(n59682) );
  AOI22xp33_ASAP7_75t_SL U54530 ( .A1(n77404), .A2(n59684), .B1(
        or1200_ic_top_from_icram[29]), .B2(n78022), .Y(n77405) );
  NAND2xp33_ASAP7_75t_SL U54531 ( .A(iwb_dat_i[8]), .B(n77373), .Y(n60393) );
  AOI22xp33_ASAP7_75t_SL U54532 ( .A1(n77376), .A2(n63953), .B1(n60391), .B2(
        n77374), .Y(n60392) );
  AOI22xp33_ASAP7_75t_SL U54533 ( .A1(n60328), .A2(n59684), .B1(
        or1200_ic_top_from_icram[27]), .B2(n59497), .Y(n60329) );
  AOI22xp33_ASAP7_75t_SL U54534 ( .A1(n77376), .A2(n61314), .B1(n60473), .B2(
        n77374), .Y(n60474) );
  OAI21xp33_ASAP7_75t_SL U54535 ( .A1(n76603), .A2(n59703), .B(n61176), .Y(
        n61177) );
  AOI22xp33_ASAP7_75t_SL U54536 ( .A1(n77376), .A2(n62052), .B1(n60365), .B2(
        n77374), .Y(n60366) );
  INVx1_ASAP7_75t_SL U54537 ( .A(n58357), .Y(n58358) );
  OAI21xp33_ASAP7_75t_SL U54538 ( .A1(n70906), .A2(n70982), .B(n70967), .Y(
        n70890) );
  NAND2xp33_ASAP7_75t_SL U54539 ( .A(iwb_dat_i[25]), .B(n77373), .Y(n60475) );
  OAI22xp33_ASAP7_75t_SL U54540 ( .A1(n76594), .A2(n76593), .B1(n76592), .B2(
        n76591), .Y(n76595) );
  INVxp33_ASAP7_75t_SL U54541 ( .A(n73398), .Y(n73355) );
  NAND2xp5_ASAP7_75t_SL U54542 ( .A(n62147), .B(n62146), .Y(n76536) );
  NAND2xp33_ASAP7_75t_SL U54543 ( .A(iwb_dat_i[0]), .B(n77373), .Y(n60367) );
  INVxp33_ASAP7_75t_SL U54544 ( .A(n65211), .Y(n76839) );
  AOI22xp33_ASAP7_75t_SL U54545 ( .A1(n60370), .A2(n62146), .B1(n60725), .B2(
        n61155), .Y(n60372) );
  NAND2xp33_ASAP7_75t_SL U54546 ( .A(n60491), .B(n61153), .Y(n60382) );
  AOI22xp33_ASAP7_75t_SL U54547 ( .A1(n77376), .A2(n69337), .B1(n60375), .B2(
        n77374), .Y(n60376) );
  NAND2xp33_ASAP7_75t_SL U54548 ( .A(iwb_dat_i[1]), .B(n77373), .Y(n60377) );
  NAND2xp5_ASAP7_75t_SL U54549 ( .A(n60440), .B(n60439), .Y(n77841) );
  NAND2x1_ASAP7_75t_SL U54550 ( .A(n59702), .B(n65211), .Y(n76523) );
  NAND2xp5_ASAP7_75t_SL U54551 ( .A(n69320), .B(n69319), .Y(
        or1200_cpu_or1200_mult_mac_n1599) );
  OAI22xp33_ASAP7_75t_SL U54552 ( .A1(or1200_cpu_or1200_except_n264), .A2(
        n76507), .B1(n75781), .B2(n76661), .Y(n74033) );
  NAND2xp33_ASAP7_75t_SL U54553 ( .A(iwb_dat_i[24]), .B(n77373), .Y(n60484) );
  AOI22xp33_ASAP7_75t_SL U54554 ( .A1(n77376), .A2(n76537), .B1(n60482), .B2(
        n77374), .Y(n60483) );
  INVxp33_ASAP7_75t_SL U54555 ( .A(n71154), .Y(n71057) );
  NAND2xp5_ASAP7_75t_SL U54556 ( .A(n77837), .B(n60443), .Y(n60454) );
  OAI22xp33_ASAP7_75t_SL U54557 ( .A1(n76508), .A2(n76661), .B1(n3123), .B2(
        n76659), .Y(n76509) );
  AOI22xp33_ASAP7_75t_SL U54558 ( .A1(n77376), .A2(n69343), .B1(n60347), .B2(
        n77374), .Y(n60348) );
  NAND2xp33_ASAP7_75t_SL U54559 ( .A(iwb_dat_i[2]), .B(n77373), .Y(n60349) );
  OAI21xp33_ASAP7_75t_SL U54560 ( .A1(n76592), .A2(n76570), .B(n76569), .Y(
        n76571) );
  NAND2xp33_ASAP7_75t_SL U54561 ( .A(iwb_dat_i[23]), .B(n77373), .Y(n60414) );
  AOI22xp33_ASAP7_75t_SL U54562 ( .A1(n77376), .A2(n60416), .B1(n60412), .B2(
        n77374), .Y(n60413) );
  AOI22xp33_ASAP7_75t_SL U54563 ( .A1(n60518), .A2(n57071), .B1(
        or1200_ic_top_from_icram[19]), .B2(n59497), .Y(n60519) );
  AOI22xp33_ASAP7_75t_SL U54564 ( .A1(n60526), .A2(n57071), .B1(
        or1200_ic_top_from_icram[20]), .B2(n78022), .Y(n60527) );
  OAI21xp33_ASAP7_75t_SL U54565 ( .A1(n74508), .A2(n74507), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_27_), 
        .Y(n74506) );
  OAI21xp33_ASAP7_75t_SL U54566 ( .A1(or1200_cpu_or1200_except_n601), .A2(
        n57093), .B(n76852), .Y(or1200_cpu_or1200_except_n1797) );
  AOI22xp33_ASAP7_75t_SL U54567 ( .A1(n60531), .A2(n57071), .B1(
        or1200_ic_top_from_icram[18]), .B2(n59497), .Y(n60532) );
  NAND2xp33_ASAP7_75t_SL U54568 ( .A(iwb_dat_i[5]), .B(n77373), .Y(n61593) );
  AOI22xp33_ASAP7_75t_SL U54569 ( .A1(n60417), .A2(n57089), .B1(
        or1200_ic_top_from_icram[21]), .B2(n78022), .Y(n60418) );
  AOI22xp33_ASAP7_75t_SL U54570 ( .A1(n77375), .A2(n59684), .B1(
        or1200_ic_top_from_icram[10]), .B2(n59497), .Y(n77371) );
  AOI22xp33_ASAP7_75t_SL U54571 ( .A1(n61024), .A2(n57071), .B1(
        or1200_ic_top_from_icram[6]), .B2(n59497), .Y(n61022) );
  AOI22xp33_ASAP7_75t_SL U54572 ( .A1(n78016), .A2(n57071), .B1(
        or1200_ic_top_from_icram[13]), .B2(n78022), .Y(n78014) );
  INVx1_ASAP7_75t_SL U54573 ( .A(n65281), .Y(n1560) );
  AOI22xp33_ASAP7_75t_SL U54574 ( .A1(n77376), .A2(n74796), .B1(n61024), .B2(
        n77374), .Y(n61025) );
  AOI22xp33_ASAP7_75t_SL U54575 ( .A1(n77376), .A2(n76809), .B1(n60385), .B2(
        n77374), .Y(n60386) );
  NAND2xp33_ASAP7_75t_SL U54576 ( .A(iwb_dat_i[7]), .B(n77373), .Y(n60387) );
  AOI22xp33_ASAP7_75t_SL U54577 ( .A1(n60412), .A2(n57089), .B1(
        or1200_ic_top_from_icram[23]), .B2(n59497), .Y(n60410) );
  AOI22xp33_ASAP7_75t_SL U54578 ( .A1(n60511), .A2(n57071), .B1(
        or1200_ic_top_from_icram[17]), .B2(n78022), .Y(n60512) );
  AOI22xp33_ASAP7_75t_SL U54579 ( .A1(n77376), .A2(n74793), .B1(n61591), .B2(
        n77374), .Y(n61592) );
  NAND2xp5_ASAP7_75t_SL U54580 ( .A(n63294), .B(n63293), .Y(n63346) );
  INVxp67_ASAP7_75t_SL U54581 ( .A(n57986), .Y(n57985) );
  NAND2xp33_ASAP7_75t_SL U54582 ( .A(iwb_dat_i[6]), .B(n77373), .Y(n61026) );
  NAND2xp33_ASAP7_75t_SL U54583 ( .A(iwb_dat_i[4]), .B(n77373), .Y(n60895) );
  OAI21xp33_ASAP7_75t_SL U54584 ( .A1(n77902), .A2(n77137), .B(n62475), .Y(
        n9627) );
  NAND2xp33_ASAP7_75t_SL U54585 ( .A(iwb_dat_i[15]), .B(n59496), .Y(n78008) );
  NAND2xp33_ASAP7_75t_SL U54586 ( .A(iwb_dat_i[12]), .B(n59496), .Y(n78018) );
  AOI22xp33_ASAP7_75t_SL U54587 ( .A1(n77376), .A2(n74790), .B1(n60893), .B2(
        n77374), .Y(n60894) );
  AOI22xp33_ASAP7_75t_SL U54588 ( .A1(n60482), .A2(n57089), .B1(
        or1200_ic_top_from_icram[24]), .B2(n59497), .Y(n60480) );
  AOI22xp33_ASAP7_75t_SL U54589 ( .A1(n78013), .A2(n59685), .B1(
        or1200_ic_top_from_icram[14]), .B2(n59497), .Y(n78011) );
  AOI22xp33_ASAP7_75t_SL U54590 ( .A1(n78025), .A2(n59684), .B1(
        or1200_ic_top_from_icram[11]), .B2(n78022), .Y(n78023) );
  NAND2xp33_ASAP7_75t_SL U54591 ( .A(iwb_dat_i[23]), .B(n78021), .Y(n60411) );
  AOI22xp33_ASAP7_75t_SL U54592 ( .A1(n78010), .A2(n59685), .B1(
        or1200_ic_top_from_icram[15]), .B2(n78022), .Y(n78007) );
  NAND2xp33_ASAP7_75t_SL U54593 ( .A(n77443), .B(n77442), .Y(n77444) );
  NAND2xp33_ASAP7_75t_SL U54594 ( .A(iwb_dat_i[24]), .B(n78021), .Y(n60481) );
  NAND2xp33_ASAP7_75t_SL U54595 ( .A(iwb_dat_i[25]), .B(n59496), .Y(n60472) );
  NAND2xp33_ASAP7_75t_SL U54596 ( .A(iwb_dat_i[14]), .B(n78021), .Y(n78012) );
  AOI22xp33_ASAP7_75t_SL U54597 ( .A1(n60893), .A2(n57071), .B1(
        or1200_ic_top_from_icram[4]), .B2(n78022), .Y(n60891) );
  OAI21xp5_ASAP7_75t_SL U54598 ( .A1(n59677), .A2(n77894), .B(n77136), .Y(
        n9624) );
  AOI22xp33_ASAP7_75t_SL U54599 ( .A1(n60397), .A2(n57089), .B1(
        or1200_ic_top_from_icram[9]), .B2(n78022), .Y(n60395) );
  XOR2xp5_ASAP7_75t_SL U54600 ( .A(n68235), .B(n68234), .Y(n68236) );
  AOI22xp33_ASAP7_75t_SL U54601 ( .A1(n78019), .A2(n57071), .B1(
        or1200_ic_top_from_icram[12]), .B2(n59497), .Y(n78017) );
  AOI22xp33_ASAP7_75t_SL U54602 ( .A1(n60473), .A2(n57089), .B1(
        or1200_ic_top_from_icram[25]), .B2(n78022), .Y(n60471) );
  AOI22xp33_ASAP7_75t_SL U54603 ( .A1(n61591), .A2(n59684), .B1(
        or1200_ic_top_from_icram[5]), .B2(n78022), .Y(n61589) );
  NAND2xp33_ASAP7_75t_SL U54604 ( .A(n74507), .B(n74494), .Y(n74504) );
  NAND2xp33_ASAP7_75t_SL U54605 ( .A(iwb_dat_i[11]), .B(n78021), .Y(n78024) );
  OAI22xp33_ASAP7_75t_SL U54606 ( .A1(n2628), .A2(n77567), .B1(n2630), .B2(
        n57072), .Y(n9221) );
  AOI21xp33_ASAP7_75t_SL U54607 ( .A1(n76810), .A2(n69337), .B(n61014), .Y(
        n61015) );
  OAI21xp33_ASAP7_75t_SL U54608 ( .A1(n2129), .A2(n77567), .B(n77543), .Y(
        n9242) );
  OAI21xp33_ASAP7_75t_SL U54609 ( .A1(n2127), .A2(n77567), .B(n77543), .Y(
        n9226) );
  NAND2xp5_ASAP7_75t_SL U54610 ( .A(n75609), .B(n75612), .Y(n75627) );
  NAND2x1_ASAP7_75t_SL U54611 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_39_), .B(
        n74308), .Y(n74415) );
  NAND2xp5_ASAP7_75t_SL U54612 ( .A(n65201), .B(n75419), .Y(n75542) );
  OAI21xp33_ASAP7_75t_SL U54613 ( .A1(n76791), .A2(n75755), .B(n75754), .Y(
        n75756) );
  INVxp67_ASAP7_75t_SL U54614 ( .A(n66529), .Y(n66532) );
  OAI22xp33_ASAP7_75t_SL U54615 ( .A1(n2524), .A2(n77567), .B1(n3390), .B2(
        n57072), .Y(n9233) );
  NAND2xp5_ASAP7_75t_SL U54616 ( .A(n77272), .B(n77263), .Y(n77264) );
  OAI22xp33_ASAP7_75t_SL U54617 ( .A1(ex_insn[22]), .A2(n77567), .B1(
        id_insn_22_), .B2(n57072), .Y(n2083) );
  NAND2xp5_ASAP7_75t_SL U54618 ( .A(n68618), .B(n68617), .Y(n68619) );
  OAI22xp33_ASAP7_75t_SL U54619 ( .A1(n2621), .A2(n77567), .B1(n2623), .B2(
        n57072), .Y(n9222) );
  NAND2xp5_ASAP7_75t_SL U54620 ( .A(n59499), .B(n76265), .Y(n75264) );
  OAI21xp33_ASAP7_75t_SL U54621 ( .A1(n2139), .A2(n77567), .B(n77540), .Y(
        n9227) );
  OAI21xp33_ASAP7_75t_SL U54622 ( .A1(n2141), .A2(n77567), .B(n77540), .Y(
        n9243) );
  AND4x1_ASAP7_75t_SL U54623 ( .A(n78211), .B(n53190), .C(n78216), .D(n73836), 
        .Y(n73837) );
  NAND2xp33_ASAP7_75t_SL U54624 ( .A(n73354), .B(n73396), .Y(n73356) );
  OAI21xp33_ASAP7_75t_SL U54625 ( .A1(n65283), .A2(n65270), .B(n65269), .Y(
        n1581) );
  AOI21xp33_ASAP7_75t_SL U54626 ( .A1(n76810), .A2(n62052), .B(n61018), .Y(
        n61019) );
  XNOR2xp5_ASAP7_75t_SL U54627 ( .A(n58359), .B(n64547), .Y(n64696) );
  OAI22xp33_ASAP7_75t_SL U54628 ( .A1(n2031), .A2(n77567), .B1(n2037), .B2(
        n57072), .Y(n9208) );
  OAI22xp33_ASAP7_75t_SL U54629 ( .A1(ex_insn[26]), .A2(n77567), .B1(n57072), 
        .B2(n61154), .Y(n2604) );
  OAI22xp33_ASAP7_75t_SL U54630 ( .A1(n2598), .A2(n77567), .B1(n2600), .B2(
        n57072), .Y(n9607) );
  OAI21xp33_ASAP7_75t_SL U54631 ( .A1(n65307), .A2(n65331), .B(n65330), .Y(
        n1763) );
  OAI22xp33_ASAP7_75t_SL U54632 ( .A1(n2153), .A2(n77567), .B1(n2160), .B2(
        n77537), .Y(n9228) );
  OAI21xp33_ASAP7_75t_SL U54633 ( .A1(n65312), .A2(n65331), .B(n65330), .Y(
        n52484) );
  OAI22xp33_ASAP7_75t_SL U54634 ( .A1(n2594), .A2(n77567), .B1(n2596), .B2(
        n57072), .Y(n9206) );
  XOR2xp5_ASAP7_75t_SL U54635 ( .A(n67206), .B(n67205), .Y(n67207) );
  OAI22xp33_ASAP7_75t_SL U54636 ( .A1(n2569), .A2(n77567), .B1(n77457), .B2(
        n57072), .Y(n9461) );
  OAI22xp33_ASAP7_75t_SL U54637 ( .A1(n2184), .A2(n77567), .B1(n2464), .B2(
        n77537), .Y(n9230) );
  OAI22xp33_ASAP7_75t_SL U54638 ( .A1(n2970), .A2(n77567), .B1(n2972), .B2(
        n57072), .Y(n9606) );
  NAND2xp5_ASAP7_75t_SL U54639 ( .A(n76630), .B(n76629), .Y(n9664) );
  NAND3xp33_ASAP7_75t_SL U54640 ( .A(n63365), .B(n63364), .C(n58477), .Y(
        n58816) );
  OAI22xp33_ASAP7_75t_SL U54641 ( .A1(n2662), .A2(n77567), .B1(n2664), .B2(
        n57072), .Y(n9216) );
  OAI22xp33_ASAP7_75t_SL U54642 ( .A1(n2086), .A2(n77567), .B1(n62469), .B2(
        n57072), .Y(n9579) );
  NAND2xp5_ASAP7_75t_SL U54643 ( .A(n70199), .B(n70198), .Y(n70209) );
  OAI21xp33_ASAP7_75t_SL U54644 ( .A1(n65388), .A2(n65331), .B(n65330), .Y(
        n2489) );
  OAI21xp33_ASAP7_75t_SL U54645 ( .A1(n65302), .A2(n65331), .B(n65330), .Y(
        n52485) );
  OAI22xp33_ASAP7_75t_SL U54646 ( .A1(n2676), .A2(n77567), .B1(n2678), .B2(
        n57072), .Y(n9214) );
  OAI21xp33_ASAP7_75t_SL U54647 ( .A1(n76906), .A2(n76893), .B(n75666), .Y(
        n75667) );
  OAI22xp33_ASAP7_75t_SL U54648 ( .A1(n2683), .A2(n77567), .B1(n2685), .B2(
        n57072), .Y(n9213) );
  OAI21xp33_ASAP7_75t_SL U54649 ( .A1(n2069), .A2(n77567), .B(n77556), .Y(
        n9578) );
  OA211x2_ASAP7_75t_SL U54650 ( .A1(n74902), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_3_), .B(n74901), 
        .C(n74900), .Y(n74903) );
  NAND2xp5_ASAP7_75t_SL U54651 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_25_), 
        .B(n74451), .Y(n74507) );
  OAI21xp33_ASAP7_75t_SL U54652 ( .A1(n2067), .A2(n77567), .B(n77556), .Y(
        n9210) );
  OAI22xp33_ASAP7_75t_SL U54653 ( .A1(ex_insn[16]), .A2(n77567), .B1(n61152), 
        .B2(n57072), .Y(n2654) );
  NAND2xp33_ASAP7_75t_SL U54654 ( .A(n76568), .B(n53440), .Y(n76569) );
  OAI22xp33_ASAP7_75t_SL U54655 ( .A1(n2691), .A2(n77567), .B1(n2693), .B2(
        n57072), .Y(n9674) );
  INVxp33_ASAP7_75t_SL U54656 ( .A(n77500), .Y(n77502) );
  INVxp67_ASAP7_75t_SL U54657 ( .A(n77839), .Y(n61051) );
  INVxp67_ASAP7_75t_SL U54658 ( .A(n61036), .Y(n60408) );
  INVxp67_ASAP7_75t_SL U54659 ( .A(n76269), .Y(n64201) );
  OAI22xp33_ASAP7_75t_SL U54660 ( .A1(n2469), .A2(n77567), .B1(n2499), .B2(
        n77537), .Y(n9231) );
  OAI22xp33_ASAP7_75t_SL U54661 ( .A1(n2649), .A2(n77567), .B1(n3392), .B2(
        n57072), .Y(n9218) );
  NAND2xp33_ASAP7_75t_SL U54662 ( .A(n77360), .B(n77359), .Y(n77361) );
  NAND2xp5_ASAP7_75t_SL U54663 ( .A(n59280), .B(n75084), .Y(n75461) );
  OAI21xp33_ASAP7_75t_SL U54664 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_3_), .A2(
        n62035), .B(n62034), .Y(n2458) );
  OAI22xp33_ASAP7_75t_SL U54665 ( .A1(n2506), .A2(n77567), .B1(n2517), .B2(
        n77537), .Y(n9232) );
  NAND2xp5_ASAP7_75t_SL U54666 ( .A(n74888), .B(n74901), .Y(n77138) );
  OAI21xp33_ASAP7_75t_SL U54667 ( .A1(n2103), .A2(n77567), .B(n77549), .Y(
        n9224) );
  NAND2xp33_ASAP7_75t_SL U54668 ( .A(n60318), .B(n77359), .Y(n60319) );
  NAND2xp5_ASAP7_75t_SL U54669 ( .A(n60890), .B(n60889), .Y(n9656) );
  OAI22xp33_ASAP7_75t_SL U54670 ( .A1(n2642), .A2(n77567), .B1(n2644), .B2(
        n57072), .Y(n9219) );
  OAI21xp33_ASAP7_75t_SL U54671 ( .A1(n2105), .A2(n77567), .B(n77549), .Y(
        n9240) );
  NAND2xp5_ASAP7_75t_SL U54672 ( .A(n60404), .B(n77376), .Y(n60405) );
  INVxp67_ASAP7_75t_SL U54673 ( .A(n76160), .Y(n76156) );
  OAI21xp33_ASAP7_75t_SL U54674 ( .A1(n53457), .A2(n64812), .B(n64811), .Y(
        n76273) );
  OAI21xp33_ASAP7_75t_SL U54675 ( .A1(n2052), .A2(n77567), .B(n77561), .Y(
        n9577) );
  OAI21xp33_ASAP7_75t_SL U54676 ( .A1(n2050), .A2(n77567), .B(n77561), .Y(
        n9209) );
  OAI22xp33_ASAP7_75t_SL U54677 ( .A1(n2635), .A2(n77567), .B1(n2637), .B2(
        n57072), .Y(n9220) );
  OAI21xp33_ASAP7_75t_SL U54678 ( .A1(n2115), .A2(n77567), .B(n77546), .Y(
        n9225) );
  NAND2xp5_ASAP7_75t_SL U54679 ( .A(n61463), .B(n61462), .Y(n9666) );
  OAI21xp33_ASAP7_75t_SL U54680 ( .A1(n2117), .A2(n77567), .B(n77546), .Y(
        n9241) );
  OAI22xp33_ASAP7_75t_SL U54681 ( .A1(n2669), .A2(n77567), .B1(n2671), .B2(
        n57072), .Y(n9215) );
  OAI21xp33_ASAP7_75t_SL U54682 ( .A1(n2826), .A2(n77567), .B(n77511), .Y(
        n9580) );
  OAI21xp33_ASAP7_75t_SL U54683 ( .A1(n2824), .A2(n77567), .B(n77511), .Y(
        n9212) );
  OA21x2_ASAP7_75t_SL U54684 ( .A1(n69352), .A2(n69347), .B(n77209), .Y(n69348) );
  OAI22xp33_ASAP7_75t_SL U54685 ( .A1(n2819), .A2(n77567), .B1(n3078), .B2(
        n57072), .Y(n9202) );
  AOI21xp33_ASAP7_75t_SL U54686 ( .A1(n76810), .A2(n76809), .B(n76808), .Y(
        n76811) );
  INVxp67_ASAP7_75t_SL U54687 ( .A(n60320), .Y(n60324) );
  INVx1_ASAP7_75t_SL U54688 ( .A(n68343), .Y(n57488) );
  OAI21xp33_ASAP7_75t_SL U54689 ( .A1(n67756), .A2(n67757), .B(n53472), .Y(
        n58074) );
  NAND2xp33_ASAP7_75t_SL U54690 ( .A(n76851), .B(n57093), .Y(n76852) );
  OAI21xp5_ASAP7_75t_SL U54691 ( .A1(n71056), .A2(n71055), .B(n71054), .Y(
        n71154) );
  OAI22xp33_ASAP7_75t_SL U54692 ( .A1(or1200_cpu_or1200_except_n567), .A2(
        n77567), .B1(n77370), .B2(n57072), .Y(or1200_cpu_or1200_except_n1827)
         );
  OAI22xp33_ASAP7_75t_SL U54693 ( .A1(or1200_cpu_or1200_except_n563), .A2(
        n77567), .B1(or1200_cpu_or1200_except_n565), .B2(n57072), .Y(
        or1200_cpu_or1200_except_n1825) );
  OAI22xp33_ASAP7_75t_SL U54694 ( .A1(or1200_cpu_or1200_except_n561), .A2(
        n77567), .B1(or1200_cpu_or1200_except_n677), .B2(n57072), .Y(
        or1200_cpu_or1200_except_n1824) );
  NAND2xp33_ASAP7_75t_SL U54695 ( .A(n57090), .B(n61059), .Y(
        or1200_cpu_or1200_except_n1831) );
  INVxp67_ASAP7_75t_SL U54696 ( .A(n77209), .Y(n76662) );
  NAND2xp5_ASAP7_75t_SL U54697 ( .A(n60271), .B(n60270), .Y(n77402) );
  NAND2xp5_ASAP7_75t_SL U54698 ( .A(n73963), .B(n77209), .Y(n76659) );
  NAND2xp33_ASAP7_75t_SL U54699 ( .A(n74037), .B(n74039), .Y(n73964) );
  NAND2xp33_ASAP7_75t_SL U54700 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[5]), .B(
        n74464), .Y(n5508) );
  NAND2xp33_ASAP7_75t_SL U54701 ( .A(n61161), .B(n77566), .Y(n77549) );
  OAI22xp33_ASAP7_75t_SL U54702 ( .A1(or1200_cpu_or1200_except_n565), .A2(
        n77567), .B1(or1200_cpu_or1200_except_n567), .B2(n77537), .Y(
        or1200_cpu_or1200_except_n1826) );
  OAI21xp33_ASAP7_75t_SL U54703 ( .A1(n77467), .A2(n77902), .B(n77303), .Y(
        n9658) );
  NAND2xp33_ASAP7_75t_SL U54704 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[10]), .B(
        n74464), .Y(n5549) );
  OAI22xp33_ASAP7_75t_SL U54705 ( .A1(n1692), .A2(n59679), .B1(n57312), .B2(
        n57074), .Y(n62547) );
  OAI21xp33_ASAP7_75t_SL U54706 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_1_), .A2(
        n74272), .B(n74271), .Y(n1612) );
  OAI21xp33_ASAP7_75t_SL U54707 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_0_), .A2(
        n74272), .B(n74271), .Y(n1614) );
  NAND2xp33_ASAP7_75t_SL U54708 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[21]), .B(
        n74464), .Y(n5537) );
  NAND2xp5_ASAP7_75t_SL U54709 ( .A(n68898), .B(n68897), .Y(
        or1200_cpu_or1200_mult_mac_n1620) );
  AOI21xp5_ASAP7_75t_SL U54710 ( .A1(n65324), .A2(n65395), .B(n65323), .Y(
        n1563) );
  NAND2xp33_ASAP7_75t_SL U54711 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[16]), .B(
        n74464), .Y(n5543) );
  NAND2xp33_ASAP7_75t_SL U54712 ( .A(n76537), .B(n77566), .Y(n77561) );
  NAND2xp33_ASAP7_75t_SL U54713 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[3]), .B(
        n74464), .Y(n5510) );
  NAND2xp33_ASAP7_75t_SL U54714 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[4]), .B(
        n74464), .Y(n5509) );
  NAND2xp33_ASAP7_75t_SL U54715 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[11]), .B(
        n74464), .Y(n5548) );
  NAND2xp5_ASAP7_75t_SL U54716 ( .A(n69136), .B(n69135), .Y(
        or1200_cpu_or1200_mult_mac_n1610) );
  XNOR2xp5_ASAP7_75t_SL U54717 ( .A(n63790), .B(n63791), .Y(n58823) );
  NAND2xp33_ASAP7_75t_SL U54718 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[12]), .B(
        n74464), .Y(n5547) );
  NAND2xp5_ASAP7_75t_SL U54719 ( .A(n76153), .B(n76152), .Y(n76160) );
  NAND2xp5_ASAP7_75t_SL U54720 ( .A(n64264), .B(n65207), .Y(n75417) );
  NAND2xp33_ASAP7_75t_SL U54721 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[20]), .B(
        n74464), .Y(n5538) );
  OAI21xp33_ASAP7_75t_SL U54722 ( .A1(n74441), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_23_), .B(
        n74449), .Y(n2331) );
  INVxp33_ASAP7_75t_SL U54723 ( .A(n62069), .Y(n62034) );
  NAND2xp33_ASAP7_75t_SL U54724 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[13]), .B(
        n74464), .Y(n5546) );
  OAI21xp33_ASAP7_75t_SL U54725 ( .A1(n74402), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_37_), .B(
        n74401), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n30) );
  NAND2xp33_ASAP7_75t_SL U54726 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[14]), .B(
        n74464), .Y(n5545) );
  OR2x2_ASAP7_75t_SL U54727 ( .A(n57966), .B(n57965), .Y(n57964) );
  INVxp67_ASAP7_75t_SL U54728 ( .A(n75970), .Y(n75956) );
  AOI21xp33_ASAP7_75t_SL U54729 ( .A1(n65313), .A2(n65334), .B(n65361), .Y(
        n65294) );
  NAND2xp33_ASAP7_75t_SL U54730 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[7]), .B(
        n74464), .Y(n5506) );
  NAND2xp33_ASAP7_75t_SL U54731 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[6]), .B(
        n74464), .Y(n5507) );
  NAND2xp33_ASAP7_75t_SL U54732 ( .A(n74796), .B(n77566), .Y(n77540) );
  OAI21xp33_ASAP7_75t_SL U54733 ( .A1(n74797), .A2(n74796), .B(n74795), .Y(
        n2142) );
  NAND2xp33_ASAP7_75t_SL U54734 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[18]), .B(
        n74464), .Y(n5541) );
  OAI22xp33_ASAP7_75t_SL U54735 ( .A1(n1658), .A2(n59679), .B1(n59534), .B2(
        n59688), .Y(n63603) );
  AOI21xp33_ASAP7_75t_SL U54736 ( .A1(n65313), .A2(n65374), .B(n65371), .Y(
        n65290) );
  OAI22xp33_ASAP7_75t_SL U54737 ( .A1(n1573), .A2(n59679), .B1(n1571), .B2(
        n57074), .Y(n64867) );
  OAI21xp33_ASAP7_75t_SL U54738 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_3_), .A2(
        n74272), .B(n74271), .Y(n1577) );
  OAI21xp33_ASAP7_75t_SL U54739 ( .A1(n74797), .A2(n74793), .B(n74792), .Y(
        n2154) );
  NAND2xp5_ASAP7_75t_SL U54740 ( .A(n76809), .B(n62004), .Y(n77543) );
  INVx2_ASAP7_75t_SL U54741 ( .A(n77195), .Y(n74885) );
  NAND2xp33_ASAP7_75t_SL U54742 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[0]), .B(
        n74464), .Y(n5550) );
  OAI21xp33_ASAP7_75t_SL U54743 ( .A1(n74797), .A2(n74790), .B(n74789), .Y(
        n2166) );
  OAI21xp33_ASAP7_75t_SL U54744 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_5_), .A2(
        n74272), .B(n74271), .Y(n1553) );
  OAI22xp33_ASAP7_75t_SL U54745 ( .A1(n1674), .A2(n59679), .B1(n59536), .B2(
        n57073), .Y(n75381) );
  INVx1_ASAP7_75t_SL U54746 ( .A(n65313), .Y(n65262) );
  INVxp67_ASAP7_75t_SL U54747 ( .A(n75060), .Y(n75062) );
  OAI21xp33_ASAP7_75t_SL U54748 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_6_), .A2(
        n74272), .B(n74271), .Y(n1552) );
  OAI21xp33_ASAP7_75t_SL U54749 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_7_), .A2(
        n74272), .B(n74271), .Y(n1551) );
  OAI22xp33_ASAP7_75t_SL U54750 ( .A1(n1590), .A2(n59679), .B1(n1588), .B2(
        n57074), .Y(n64257) );
  NAND2xp33_ASAP7_75t_SL U54751 ( .A(n69343), .B(n62069), .Y(n2179) );
  NAND2xp33_ASAP7_75t_SL U54752 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[8]), .B(
        n74464), .Y(n5505) );
  NAND2xp33_ASAP7_75t_SL U54753 ( .A(n60416), .B(n77566), .Y(n77556) );
  AOI21xp33_ASAP7_75t_SL U54754 ( .A1(n62000), .A2(n57333), .B(n60359), .Y(
        n60362) );
  NAND2xp33_ASAP7_75t_SL U54755 ( .A(n63953), .B(n77566), .Y(n77546) );
  OAI21xp33_ASAP7_75t_SL U54756 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_2_), .A2(
        n74272), .B(n74271), .Y(n1594) );
  NAND2xp33_ASAP7_75t_SL U54757 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[19]), .B(
        n74464), .Y(n5540) );
  OR2x2_ASAP7_75t_SL U54758 ( .A(n57846), .B(n75057), .Y(n57842) );
  NAND2xp33_ASAP7_75t_SL U54759 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[1]), .B(
        n74464), .Y(n5539) );
  NAND2xp33_ASAP7_75t_SL U54760 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[17]), .B(
        n74464), .Y(n5542) );
  NAND2xp33_ASAP7_75t_SL U54761 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[9]), .B(
        n74464), .Y(n5503) );
  OAI21xp33_ASAP7_75t_SL U54762 ( .A1(n74797), .A2(n62052), .B(n62051), .Y(
        n2529) );
  OAI21xp33_ASAP7_75t_SL U54763 ( .A1(n76104), .A2(n76108), .B(n76103), .Y(
        n76105) );
  INVxp67_ASAP7_75t_SL U54764 ( .A(n75969), .Y(n75964) );
  OAI21xp33_ASAP7_75t_SL U54765 ( .A1(n74797), .A2(n69337), .B(n62050), .Y(
        n2511) );
  OAI21xp33_ASAP7_75t_SL U54766 ( .A1(n74878), .A2(n74877), .B(n77195), .Y(
        n74879) );
  AOI21xp33_ASAP7_75t_SL U54767 ( .A1(n65313), .A2(n65298), .B(n65301), .Y(
        n65299) );
  NAND2xp33_ASAP7_75t_SL U54768 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[2]), .B(
        n74464), .Y(n5513) );
  OAI21xp33_ASAP7_75t_SL U54769 ( .A1(n77467), .A2(n77891), .B(n76241), .Y(
        n9654) );
  OAI22xp33_ASAP7_75t_SL U54770 ( .A1(n1642), .A2(n59679), .B1(n59532), .B2(
        n57074), .Y(n74636) );
  INVxp67_ASAP7_75t_SL U54771 ( .A(n70015), .Y(n2273) );
  OAI21xp33_ASAP7_75t_SL U54772 ( .A1(n77467), .A2(n77232), .B(n77231), .Y(
        n9657) );
  OAI22xp33_ASAP7_75t_SL U54773 ( .A1(n2558), .A2(n59679), .B1(n59550), .B2(
        n57073), .Y(n75757) );
  INVx2_ASAP7_75t_SL U54774 ( .A(n59678), .Y(n59677) );
  AOI21xp33_ASAP7_75t_SL U54775 ( .A1(n74434), .A2(n74226), .B(n74227), .Y(
        n74445) );
  NAND2xp5_ASAP7_75t_SL U54776 ( .A(n77270), .B(n77262), .Y(n77263) );
  INVxp67_ASAP7_75t_SL U54777 ( .A(n75307), .Y(n75308) );
  OAI22xp33_ASAP7_75t_SL U54778 ( .A1(n2555), .A2(n59679), .B1(n59549), .B2(
        n57073), .Y(n75267) );
  OAI22xp33_ASAP7_75t_SL U54779 ( .A1(n2552), .A2(n59679), .B1(n1868), .B2(
        n57074), .Y(n77183) );
  INVxp33_ASAP7_75t_SL U54780 ( .A(n75808), .Y(n64811) );
  OAI22xp33_ASAP7_75t_SL U54781 ( .A1(n2581), .A2(n77567), .B1(n77552), .B2(
        n74797), .Y(n9463) );
  OAI22xp33_ASAP7_75t_SL U54782 ( .A1(n2963), .A2(n59679), .B1(n59547), .B2(
        n57073), .Y(n75610) );
  OAI22xp33_ASAP7_75t_SL U54783 ( .A1(n2941), .A2(n59679), .B1(n59546), .B2(
        n57074), .Y(n62140) );
  NAND2xp33_ASAP7_75t_SL U54784 ( .A(or1200_cpu_rf_datab[5]), .B(n57091), .Y(
        n61670) );
  OAI21xp33_ASAP7_75t_SL U54785 ( .A1(n75809), .A2(n75808), .B(n75807), .Y(
        n75810) );
  INVxp33_ASAP7_75t_SL U54786 ( .A(n75680), .Y(n75681) );
  NAND2xp33_ASAP7_75t_SL U54787 ( .A(n59672), .B(n69261), .Y(n69268) );
  OAI21xp33_ASAP7_75t_SL U54788 ( .A1(n77467), .A2(n77905), .B(n75787), .Y(
        n9660) );
  NAND2xp33_ASAP7_75t_SL U54789 ( .A(n78019), .B(n57092), .Y(n7630) );
  OAI21xp33_ASAP7_75t_SL U54790 ( .A1(n76906), .A2(n69318), .B(n69315), .Y(
        n69316) );
  INVxp67_ASAP7_75t_SL U54791 ( .A(n77362), .Y(n57139) );
  AOI21xp33_ASAP7_75t_SL U54792 ( .A1(n65313), .A2(n65385), .B(n65311), .Y(
        n65310) );
  AOI21xp33_ASAP7_75t_SL U54793 ( .A1(n65313), .A2(n65384), .B(n65383), .Y(
        n65315) );
  NAND2xp33_ASAP7_75t_SL U54794 ( .A(n77401), .B(n77307), .Y(n60270) );
  NAND2xp33_ASAP7_75t_SL U54795 ( .A(or1200_cpu_rf_datab[8]), .B(n57091), .Y(
        n62393) );
  NAND2xp33_ASAP7_75t_SL U54796 ( .A(or1200_cpu_rf_datab[9]), .B(n57091), .Y(
        n76516) );
  OAI21xp33_ASAP7_75t_SL U54797 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_4_), .A2(
        n74272), .B(n74271), .Y(n2859) );
  OAI21xp33_ASAP7_75t_SL U54798 ( .A1(n77907), .A2(n77467), .B(n61378), .Y(
        n9661) );
  INVxp33_ASAP7_75t_SL U54799 ( .A(n77904), .Y(n76562) );
  NAND2xp33_ASAP7_75t_SL U54800 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco2[15]), .B(
        n74464), .Y(n5544) );
  NAND2xp33_ASAP7_75t_SL U54801 ( .A(or1200_cpu_rf_datab[6]), .B(n57091), .Y(
        n62301) );
  OAI22xp33_ASAP7_75t_SL U54802 ( .A1(n3071), .A2(n59679), .B1(n59711), .B2(
        n57074), .Y(n61018) );
  NAND2xp33_ASAP7_75t_SL U54803 ( .A(n76558), .B(n77566), .Y(n77511) );
  INVx1_ASAP7_75t_SL U54804 ( .A(n67756), .Y(n58117) );
  NAND2xp5_ASAP7_75t_SL U54805 ( .A(n70878), .B(n58288), .Y(n70862) );
  AOI22xp33_ASAP7_75t_SL U54806 ( .A1(n59673), .A2(n77974), .B1(n68892), .B2(
        n75650), .Y(n68898) );
  AOI22xp33_ASAP7_75t_SL U54807 ( .A1(n59673), .A2(n77971), .B1(n69084), .B2(
        n75650), .Y(n69078) );
  INVxp67_ASAP7_75t_SL U54808 ( .A(n69970), .Y(n2277) );
  INVx1_ASAP7_75t_SL U54809 ( .A(n66340), .Y(n66339) );
  AOI22xp33_ASAP7_75t_SL U54810 ( .A1(n59673), .A2(n77869), .B1(n69324), .B2(
        n75650), .Y(n69320) );
  INVxp33_ASAP7_75t_SL U54811 ( .A(n65271), .Y(n65272) );
  INVxp67_ASAP7_75t_SL U54812 ( .A(n76181), .Y(n75954) );
  INVxp67_ASAP7_75t_SL U54813 ( .A(n75078), .Y(n75083) );
  AO21x1_ASAP7_75t_SL U54814 ( .A1(n74392), .A2(n74391), .B(n74402), .Y(n74393) );
  INVxp33_ASAP7_75t_SL U54815 ( .A(n74797), .Y(n62035) );
  NAND2xp5_ASAP7_75t_SL U54816 ( .A(n68954), .B(n68953), .Y(
        or1200_cpu_or1200_mult_mac_n1618) );
  OAI21xp33_ASAP7_75t_SL U54817 ( .A1(n69323), .A2(n69310), .B(n69322), .Y(
        n69318) );
  NAND2xp33_ASAP7_75t_SL U54818 ( .A(n57079), .B(n69215), .Y(n69223) );
  NAND2xp33_ASAP7_75t_SL U54819 ( .A(n74809), .B(n74797), .Y(n74789) );
  AOI22xp33_ASAP7_75t_SL U54820 ( .A1(n59673), .A2(n77877), .B1(n69220), .B2(
        n75650), .Y(n69221) );
  INVxp67_ASAP7_75t_SL U54821 ( .A(n66843), .Y(n66844) );
  OAI21xp33_ASAP7_75t_SL U54822 ( .A1(n75071), .A2(n75056), .B(n75078), .Y(
        n75060) );
  AOI22xp33_ASAP7_75t_SL U54823 ( .A1(n76903), .A2(n77856), .B1(n76894), .B2(
        n75650), .Y(n75670) );
  OAI21xp33_ASAP7_75t_SL U54824 ( .A1(n59671), .A2(n76895), .B(n75665), .Y(
        n75668) );
  NAND3xp33_ASAP7_75t_SRAM U54825 ( .A(n76973), .B(n76972), .C(n76971), .Y(
        n76981) );
  NAND2xp33_ASAP7_75t_SL U54826 ( .A(n74791), .B(n74797), .Y(n74792) );
  AOI21xp33_ASAP7_75t_SL U54827 ( .A1(n77182), .A2(n76870), .B(n76869), .Y(
        n76871) );
  AOI22xp33_ASAP7_75t_SL U54828 ( .A1(n59673), .A2(n77873), .B1(n75558), .B2(
        n75650), .Y(n69266) );
  OA21x2_ASAP7_75t_SRAM U54829 ( .A1(n74435), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_22_), 
        .B(n74434), .Y(n74436) );
  AOI21xp33_ASAP7_75t_SL U54830 ( .A1(n76895), .A2(n57079), .B(n75665), .Y(
        n75666) );
  AOI21xp33_ASAP7_75t_SL U54831 ( .A1(n77182), .A2(n77006), .B(n77005), .Y(
        n77007) );
  INVxp67_ASAP7_75t_SL U54832 ( .A(n67113), .Y(n66510) );
  AOI21xp33_ASAP7_75t_SL U54833 ( .A1(n69265), .A2(n57079), .B(n69264), .Y(
        n69267) );
  NAND2xp33_ASAP7_75t_SL U54834 ( .A(n74794), .B(n74797), .Y(n74795) );
  INVxp33_ASAP7_75t_SL U54835 ( .A(n69265), .Y(n69261) );
  INVx2_ASAP7_75t_SL U54836 ( .A(n65308), .Y(n65331) );
  NAND2xp5_ASAP7_75t_SL U54837 ( .A(n69328), .B(n75130), .Y(n75117) );
  INVxp67_ASAP7_75t_SL U54838 ( .A(n66820), .Y(n58064) );
  INVxp67_ASAP7_75t_SL U54839 ( .A(n67187), .Y(n67192) );
  OAI21xp33_ASAP7_75t_SL U54840 ( .A1(n1600), .A2(n65322), .B(n65308), .Y(
        n65282) );
  AOI21xp33_ASAP7_75t_SL U54841 ( .A1(n77182), .A2(n76626), .B(n62299), .Y(
        n62300) );
  OAI21xp33_ASAP7_75t_SL U54842 ( .A1(n78116), .A2(n56829), .B(n78115), .Y(
        n9366) );
  OAI21xp33_ASAP7_75t_SL U54843 ( .A1(n78112), .A2(n56829), .B(n78111), .Y(
        n9365) );
  OAI21xp33_ASAP7_75t_SL U54844 ( .A1(n78108), .A2(n56829), .B(n78107), .Y(
        n9364) );
  OAI21xp33_ASAP7_75t_SL U54845 ( .A1(n78104), .A2(n56829), .B(n78103), .Y(
        n9363) );
  INVx1_ASAP7_75t_SL U54846 ( .A(n63106), .Y(n58183) );
  AOI21xp33_ASAP7_75t_SL U54847 ( .A1(n77182), .A2(n76514), .B(n76513), .Y(
        n76515) );
  OAI21xp33_ASAP7_75t_SL U54848 ( .A1(n78099), .A2(n56829), .B(n78098), .Y(
        n9362) );
  OAI21xp33_ASAP7_75t_SL U54849 ( .A1(n78087), .A2(n56829), .B(n78086), .Y(
        n9361) );
  OAI21xp33_ASAP7_75t_SL U54850 ( .A1(n78083), .A2(n56829), .B(n78082), .Y(
        n9360) );
  OAI21xp33_ASAP7_75t_SL U54851 ( .A1(n78079), .A2(n56829), .B(n78078), .Y(
        n9359) );
  INVx3_ASAP7_75t_SL U54852 ( .A(n62000), .Y(n77567) );
  NAND2xp33_ASAP7_75t_SL U54853 ( .A(n78438), .B(n74797), .Y(n62051) );
  OAI21xp33_ASAP7_75t_SL U54854 ( .A1(n78075), .A2(n56829), .B(n78074), .Y(
        n9358) );
  NAND2xp33_ASAP7_75t_SL U54855 ( .A(n78437), .B(n74797), .Y(n62050) );
  OAI21xp33_ASAP7_75t_SL U54856 ( .A1(n78071), .A2(n56829), .B(n78070), .Y(
        n9357) );
  OAI21xp5_ASAP7_75t_SL U54857 ( .A1(n73330), .A2(n73360), .B(n73329), .Y(
        n73357) );
  AOI21xp33_ASAP7_75t_SL U54858 ( .A1(n77182), .A2(n76652), .B(n62391), .Y(
        n62392) );
  AOI21xp33_ASAP7_75t_SL U54859 ( .A1(n77182), .A2(n76220), .B(n61668), .Y(
        n61669) );
  NAND2xp5_ASAP7_75t_SL U54860 ( .A(n70822), .B(n70821), .Y(n70833) );
  OAI22xp33_ASAP7_75t_SL U54861 ( .A1(n3419), .A2(n56829), .B1(n1295), .B2(
        n58399), .Y(n9377) );
  OAI22xp33_ASAP7_75t_SL U54862 ( .A1(n2843), .A2(n56829), .B1(n1290), .B2(
        n58399), .Y(n9376) );
  INVx1_ASAP7_75t_SL U54863 ( .A(n58253), .Y(n57255) );
  OAI21xp33_ASAP7_75t_SL U54864 ( .A1(n78159), .A2(n56829), .B(n78158), .Y(
        n9375) );
  OAI21xp33_ASAP7_75t_SL U54865 ( .A1(n78153), .A2(n56829), .B(n78152), .Y(
        n9374) );
  OAI21xp33_ASAP7_75t_SL U54866 ( .A1(n78147), .A2(n56829), .B(n78146), .Y(
        n9373) );
  OAI21xp33_ASAP7_75t_SL U54867 ( .A1(n78143), .A2(n56829), .B(n78142), .Y(
        n9372) );
  OAI21xp33_ASAP7_75t_SL U54868 ( .A1(n78137), .A2(n56829), .B(n78136), .Y(
        n9371) );
  OAI21xp5_ASAP7_75t_SL U54869 ( .A1(n73953), .A2(n76307), .B(n61740), .Y(
        n77904) );
  NAND2xp5_ASAP7_75t_SL U54870 ( .A(n63050), .B(n63051), .Y(n58185) );
  OAI21xp33_ASAP7_75t_SL U54871 ( .A1(n78132), .A2(n56829), .B(n78131), .Y(
        n9370) );
  INVx2_ASAP7_75t_SL U54872 ( .A(n77182), .Y(n59679) );
  OAI21xp33_ASAP7_75t_SL U54873 ( .A1(n78128), .A2(n56829), .B(n78127), .Y(
        n9369) );
  OAI21xp33_ASAP7_75t_SL U54874 ( .A1(n78124), .A2(n56829), .B(n78123), .Y(
        n9368) );
  OAI21xp33_ASAP7_75t_SL U54875 ( .A1(n65309), .A2(n65354), .B(n65308), .Y(
        n65316) );
  OAI21xp33_ASAP7_75t_SL U54876 ( .A1(n78120), .A2(n56829), .B(n78119), .Y(
        n9367) );
  INVxp67_ASAP7_75t_SL U54877 ( .A(n63368), .Y(n62950) );
  AOI21xp33_ASAP7_75t_SL U54878 ( .A1(n77182), .A2(n76689), .B(n61264), .Y(
        n61265) );
  INVx1_ASAP7_75t_SL U54879 ( .A(n67764), .Y(n58846) );
  AOI21x1_ASAP7_75t_SL U54880 ( .A1(n76835), .A2(n76834), .B(n61163), .Y(
        n76590) );
  OAI21xp33_ASAP7_75t_SL U54881 ( .A1(n1727), .A2(n59689), .B(n69342), .Y(
        n1728) );
  AND2x2_ASAP7_75t_SL U54882 ( .A(n73361), .B(n73360), .Y(n73362) );
  OAI21xp33_ASAP7_75t_SL U54883 ( .A1(n77763), .A2(n61997), .B(n61309), .Y(
        n9344) );
  OAI21xp33_ASAP7_75t_SL U54884 ( .A1(n71306), .A2(n71299), .B(n71298), .Y(
        n71300) );
  AOI21xp5_ASAP7_75t_SL U54885 ( .A1(n76264), .A2(n77031), .B(n62546), .Y(
        n77891) );
  INVxp67_ASAP7_75t_SL U54886 ( .A(n73841), .Y(n53191) );
  XNOR2xp5_ASAP7_75t_SL U54887 ( .A(n63873), .B(n58824), .Y(n63792) );
  OAI21xp33_ASAP7_75t_SL U54888 ( .A1(n1882), .A2(n59689), .B(n77409), .Y(
        n1883) );
  AOI21xp33_ASAP7_75t_SL U54889 ( .A1(n61308), .A2(n59696), .B(n61307), .Y(
        n61309) );
  OAI21xp33_ASAP7_75t_SL U54890 ( .A1(n1888), .A2(n59689), .B(n77409), .Y(
        n1889) );
  OAI21xp33_ASAP7_75t_SL U54891 ( .A1(n1879), .A2(n57073), .B(n77409), .Y(
        n1880) );
  OAI21xp33_ASAP7_75t_SL U54892 ( .A1(n1900), .A2(n59689), .B(n77409), .Y(
        n1901) );
  OAI21xp33_ASAP7_75t_SL U54893 ( .A1(n1891), .A2(n59688), .B(n77409), .Y(
        n1892) );
  AND2x2_ASAP7_75t_SL U54894 ( .A(n78440), .B(n77459), .Y(n77456) );
  OAI21xp33_ASAP7_75t_SL U54895 ( .A1(n1906), .A2(n59689), .B(n77409), .Y(
        n1907) );
  OAI21xp33_ASAP7_75t_SL U54896 ( .A1(n1894), .A2(n57074), .B(n77409), .Y(
        n1895) );
  OAI21xp33_ASAP7_75t_SL U54897 ( .A1(n1909), .A2(n57073), .B(n77409), .Y(
        n1910) );
  OAI21xp33_ASAP7_75t_SL U54898 ( .A1(n59688), .A2(n2521), .B(n77569), .Y(
        n2522) );
  OAI21xp33_ASAP7_75t_SL U54899 ( .A1(n1915), .A2(n57073), .B(n77409), .Y(
        n1916) );
  OAI21xp33_ASAP7_75t_SL U54900 ( .A1(n1903), .A2(n57073), .B(n77409), .Y(
        n1904) );
  OAI21xp33_ASAP7_75t_SL U54901 ( .A1(n1876), .A2(n57073), .B(n77409), .Y(
        n1877) );
  OAI21xp33_ASAP7_75t_SL U54902 ( .A1(n1885), .A2(n59688), .B(n77409), .Y(
        n1886) );
  OAI21xp33_ASAP7_75t_SL U54903 ( .A1(n1897), .A2(n59688), .B(n77409), .Y(
        n1898) );
  OAI21xp33_ASAP7_75t_SL U54904 ( .A1(n59688), .A2(n2047), .B(n77563), .Y(
        n2048) );
  OAI21xp33_ASAP7_75t_SL U54905 ( .A1(n1912), .A2(n57074), .B(n77409), .Y(
        n1913) );
  OAI21xp33_ASAP7_75t_SL U54906 ( .A1(n59689), .A2(n2028), .B(n77560), .Y(
        n2029) );
  OAI21xp33_ASAP7_75t_SL U54907 ( .A1(n59689), .A2(n2632), .B(n77515), .Y(
        n2633) );
  OAI21xp33_ASAP7_75t_SL U54908 ( .A1(n69283), .A2(n69260), .B(n69259), .Y(
        n69265) );
  OAI21xp33_ASAP7_75t_SL U54909 ( .A1(n59689), .A2(n2618), .B(n77519), .Y(
        n2619) );
  OAI22xp33_ASAP7_75t_SL U54910 ( .A1(n2037), .A2(n60489), .B1(n57073), .B2(
        n2026), .Y(n9197) );
  OAI21xp33_ASAP7_75t_SL U54911 ( .A1(n76906), .A2(n69263), .B(n69262), .Y(
        n69264) );
  OAI21xp33_ASAP7_75t_SL U54912 ( .A1(n57074), .A2(n2639), .B(n77513), .Y(
        n2640) );
  OAI21xp33_ASAP7_75t_SL U54913 ( .A1(n59689), .A2(n2611), .B(n77521), .Y(
        n2612) );
  OAI22xp33_ASAP7_75t_SL U54914 ( .A1(n2172), .A2(n77025), .B1(n59567), .B2(
        n57073), .Y(n77005) );
  OAI22xp33_ASAP7_75t_SL U54915 ( .A1(n2098), .A2(n77025), .B1(n57500), .B2(
        n57074), .Y(n61803) );
  OAI21xp33_ASAP7_75t_SL U54916 ( .A1(n59688), .A2(wb_insn[26]), .B(n77523), 
        .Y(n2601) );
  AOI21xp33_ASAP7_75t_SL U54917 ( .A1(n74426), .A2(n74425), .B(n74435), .Y(
        n74438) );
  NAND2xp5_ASAP7_75t_SL U54918 ( .A(n75553), .B(n75554), .Y(n75552) );
  OAI21xp33_ASAP7_75t_SL U54919 ( .A1(n74385), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_35_), .B(
        n74392), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n26) );
  OAI21xp33_ASAP7_75t_SL U54920 ( .A1(n59688), .A2(n2591), .B(n77525), .Y(
        n2592) );
  INVxp33_ASAP7_75t_SL U54921 ( .A(n77449), .Y(n77450) );
  INVxp67_ASAP7_75t_SL U54922 ( .A(n69219), .Y(n69215) );
  NOR2x1_ASAP7_75t_SL U54923 ( .A(n74391), .B(n74392), .Y(n74402) );
  INVxp67_ASAP7_75t_SL U54924 ( .A(n67189), .Y(n67169) );
  AOI21xp5_ASAP7_75t_SL U54925 ( .A1(n69219), .A2(n57079), .B(n69218), .Y(
        n69222) );
  INVxp67_ASAP7_75t_SL U54926 ( .A(n64813), .Y(n64809) );
  OAI22xp33_ASAP7_75t_SL U54927 ( .A1(n2464), .A2(n77025), .B1(n59558), .B2(
        n57073), .Y(n76869) );
  OAI22xp33_ASAP7_75t_SL U54928 ( .A1(n2148), .A2(n77025), .B1(n59556), .B2(
        n59688), .Y(n62299) );
  NAND2xp5_ASAP7_75t_SL U54929 ( .A(n73443), .B(n73442), .Y(n73444) );
  INVxp33_ASAP7_75t_SL U54930 ( .A(n77459), .Y(n77552) );
  INVxp67_ASAP7_75t_SL U54931 ( .A(n60489), .Y(n60486) );
  OAI21xp33_ASAP7_75t_SL U54932 ( .A1(n59688), .A2(n2625), .B(n77517), .Y(
        n2626) );
  OAI21xp33_ASAP7_75t_SL U54933 ( .A1(n73437), .A2(n58278), .B(n73442), .Y(
        n51956) );
  OAI22xp33_ASAP7_75t_SL U54934 ( .A1(n2110), .A2(n77025), .B1(n59543), .B2(
        n57074), .Y(n76513) );
  OAI22xp33_ASAP7_75t_SL U54935 ( .A1(n61127), .A2(n61126), .B1(n59539), .B2(
        n57074), .Y(n61128) );
  NAND2xp5_ASAP7_75t_SL U54936 ( .A(dbg_stall_i), .B(n77449), .Y(n60266) );
  INVx1_ASAP7_75t_SL U54937 ( .A(n77900), .Y(n77232) );
  OAI22xp33_ASAP7_75t_SL U54938 ( .A1(n2122), .A2(n77025), .B1(n59554), .B2(
        n57074), .Y(n62391) );
  NOR2x1_ASAP7_75t_SL U54939 ( .A(n62975), .B(n62976), .Y(n62994) );
  OAI22xp33_ASAP7_75t_SL U54940 ( .A1(n2160), .A2(n77025), .B1(n59544), .B2(
        n59689), .Y(n61668) );
  OAI22xp33_ASAP7_75t_SL U54941 ( .A1(n77026), .A2(n77025), .B1(n59552), .B2(
        n57073), .Y(n77027) );
  OAI21xp33_ASAP7_75t_SL U54942 ( .A1(n59688), .A2(n2539), .B(n77527), .Y(
        n2540) );
  OAI22xp33_ASAP7_75t_SL U54943 ( .A1(n2499), .A2(n77025), .B1(n59708), .B2(
        n57074), .Y(n61264) );
  OAI21xp33_ASAP7_75t_SL U54944 ( .A1(n1921), .A2(n57073), .B(n77409), .Y(
        n1922) );
  OA21x2_ASAP7_75t_SL U54945 ( .A1(n59689), .A2(n76220), .B(n76221), .Y(n61667) );
  OAI22xp33_ASAP7_75t_SL U54946 ( .A1(n65345), .A2(n65287), .B1(n65322), .B2(
        n65284), .Y(n65285) );
  OAI21xp33_ASAP7_75t_SL U54947 ( .A1(n1918), .A2(n57073), .B(n77409), .Y(
        n1919) );
  OAI21xp5_ASAP7_75t_SL U54948 ( .A1(n70455), .A2(n70305), .B(n70290), .Y(
        n2402) );
  OAI21xp33_ASAP7_75t_SL U54949 ( .A1(n59689), .A2(n2181), .B(n77533), .Y(
        n2182) );
  OAI21xp33_ASAP7_75t_SL U54950 ( .A1(n70182), .A2(n70181), .B(n70187), .Y(
        n3258) );
  OAI21xp33_ASAP7_75t_SL U54951 ( .A1(n2169), .A2(n57073), .B(n77534), .Y(
        n2170) );
  OAI21xp5_ASAP7_75t_SL U54952 ( .A1(n70455), .A2(n70378), .B(n70367), .Y(
        n2408) );
  OAI22xp33_ASAP7_75t_SL U54953 ( .A1(n1573), .A2(n77463), .B1(n59528), .B2(
        n57073), .Y(n73903) );
  OAI21xp33_ASAP7_75t_SL U54954 ( .A1(n59689), .A2(n2162), .B(n77536), .Y(
        n2163) );
  INVxp67_ASAP7_75t_SL U54955 ( .A(n65267), .Y(n65279) );
  OAI21xp33_ASAP7_75t_SL U54956 ( .A1(n59689), .A2(n2150), .B(n77539), .Y(
        n2151) );
  OAI21xp5_ASAP7_75t_SL U54957 ( .A1(n70455), .A2(n70480), .B(n70454), .Y(
        n2414) );
  OAI21xp5_ASAP7_75t_SL U54958 ( .A1(n70481), .A2(n70305), .B(n70304), .Y(
        n2421) );
  OAI21xp33_ASAP7_75t_SL U54959 ( .A1(n59689), .A2(n2136), .B(n77542), .Y(
        n2137) );
  OAI21xp5_ASAP7_75t_SL U54960 ( .A1(n70481), .A2(n70378), .B(n70377), .Y(
        n2431) );
  NOR2x1_ASAP7_75t_SL U54961 ( .A(n67989), .B(n67988), .Y(n57660) );
  OAI21xp5_ASAP7_75t_SL U54962 ( .A1(n70481), .A2(n70480), .B(n70479), .Y(
        n2435) );
  OAI22xp33_ASAP7_75t_SL U54963 ( .A1(n1590), .A2(n77463), .B1(n59529), .B2(
        n57074), .Y(n74108) );
  OAI21xp33_ASAP7_75t_SL U54964 ( .A1(n59689), .A2(n2124), .B(n77545), .Y(
        n2125) );
  INVx1_ASAP7_75t_SL U54965 ( .A(n68033), .Y(n57140) );
  OAI21xp33_ASAP7_75t_SL U54966 ( .A1(n76069), .A2(n76068), .B(n76067), .Y(
        n76070) );
  OAI21xp5_ASAP7_75t_SL U54967 ( .A1(n76081), .A2(n76080), .B(n76079), .Y(
        n76082) );
  INVxp67_ASAP7_75t_SL U54968 ( .A(n77025), .Y(n76810) );
  NAND2xp33_ASAP7_75t_SL U54969 ( .A(n76090), .B(n76096), .Y(n76102) );
  OAI21xp33_ASAP7_75t_SL U54970 ( .A1(n59689), .A2(n2112), .B(n77548), .Y(
        n2113) );
  NAND2xp5_ASAP7_75t_SL U54971 ( .A(n74460), .B(n74726), .Y(n74220) );
  INVxp67_ASAP7_75t_SL U54972 ( .A(n70840), .Y(n70839) );
  NOR2x1_ASAP7_75t_SL U54973 ( .A(n61990), .B(n77025), .Y(n77184) );
  XNOR2xp5_ASAP7_75t_SL U54974 ( .A(n64942), .B(n57608), .Y(n65000) );
  INVxp33_ASAP7_75t_SL U54975 ( .A(n68636), .Y(n66565) );
  OAI21xp33_ASAP7_75t_SL U54976 ( .A1(n57073), .A2(n2188), .B(n77849), .Y(
        n2189) );
  OAI21xp5_ASAP7_75t_SL U54977 ( .A1(n70409), .A2(n70305), .B(n70263), .Y(
        n2336) );
  INVxp67_ASAP7_75t_SL U54978 ( .A(n66513), .Y(n66517) );
  AOI21xp33_ASAP7_75t_SL U54979 ( .A1(n73463), .A2(n73462), .B(n73461), .Y(
        n73841) );
  OAI21xp5_ASAP7_75t_SL U54980 ( .A1(n70409), .A2(n70378), .B(n70335), .Y(
        n2346) );
  OAI21xp5_ASAP7_75t_SL U54981 ( .A1(n70409), .A2(n70480), .B(n70408), .Y(
        n2356) );
  OAI21xp5_ASAP7_75t_SL U54982 ( .A1(n70394), .A2(n70378), .B(n70324), .Y(
        n2358) );
  OAI21xp5_ASAP7_75t_SL U54983 ( .A1(n70394), .A2(n70305), .B(n70256), .Y(
        n2360) );
  OAI21xp5_ASAP7_75t_SL U54984 ( .A1(n70394), .A2(n70480), .B(n70393), .Y(
        n2366) );
  OAI21xp33_ASAP7_75t_SL U54985 ( .A1(n74430), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_21_), .B(
        n74443), .Y(n2373) );
  OAI21xp5_ASAP7_75t_SL U54986 ( .A1(n70419), .A2(n70305), .B(n70271), .Y(
        n2376) );
  OAI21xp5_ASAP7_75t_SL U54987 ( .A1(n70438), .A2(n70305), .B(n70282), .Y(
        n2386) );
  INVxp67_ASAP7_75t_SL U54988 ( .A(n62033), .Y(n9671) );
  AOI21xp5_ASAP7_75t_SL U54989 ( .A1(n76276), .A2(n77031), .B(n60888), .Y(
        n77897) );
  OAI21xp5_ASAP7_75t_SL U54990 ( .A1(n70438), .A2(n70378), .B(n70353), .Y(
        n2392) );
  OAI21xp5_ASAP7_75t_SL U54991 ( .A1(n70438), .A2(n70480), .B(n70437), .Y(
        n2398) );
  OAI21xp33_ASAP7_75t_SL U54992 ( .A1(n59689), .A2(n2090), .B(n77555), .Y(
        n2091) );
  OAI21xp33_ASAP7_75t_SL U54993 ( .A1(n59688), .A2(n2064), .B(n77558), .Y(
        n2065) );
  NAND2xp33_ASAP7_75t_SL U54994 ( .A(n77208), .B(n63712), .Y(n63714) );
  OAI22xp33_ASAP7_75t_SL U54995 ( .A1(n2071), .A2(n60489), .B1(n57073), .B2(
        n2062), .Y(n9199) );
  OAI21xp33_ASAP7_75t_SL U54996 ( .A1(n2095), .A2(n59688), .B(n77553), .Y(
        n2096) );
  OAI22xp33_ASAP7_75t_SL U54997 ( .A1(n62469), .A2(n60489), .B1(n57073), .B2(
        n2079), .Y(n9200) );
  XNOR2xp5_ASAP7_75t_SL U54998 ( .A(n64544), .B(n64543), .Y(n64592) );
  OAI21xp33_ASAP7_75t_SL U54999 ( .A1(n59688), .A2(n2466), .B(n77531), .Y(
        n2467) );
  NAND2xp5_ASAP7_75t_SL U55000 ( .A(n63722), .B(n77248), .Y(n63725) );
  OAI21xp33_ASAP7_75t_SL U55001 ( .A1(n59689), .A2(wb_insn[22]), .B(n77565), 
        .Y(n2080) );
  INVx1_ASAP7_75t_SL U55002 ( .A(n76932), .Y(n76973) );
  NAND2xp5_ASAP7_75t_SL U55003 ( .A(n71022), .B(n70979), .Y(n70980) );
  OAI22xp33_ASAP7_75t_SL U55004 ( .A1(n1692), .A2(n77463), .B1(n59486), .B2(
        n57074), .Y(n76240) );
  OAI21xp33_ASAP7_75t_SL U55005 ( .A1(n59688), .A2(n2503), .B(n77529), .Y(
        n2504) );
  OAI22xp33_ASAP7_75t_SL U55006 ( .A1(n1628), .A2(n77463), .B1(n57377), .B2(
        n57074), .Y(n74552) );
  NOR2xp33_ASAP7_75t_SL U55007 ( .A(n74976), .B(n74975), .Y(n75391) );
  INVxp33_ASAP7_75t_SL U55008 ( .A(n63343), .Y(n62951) );
  OAI21xp33_ASAP7_75t_SL U55009 ( .A1(n59689), .A2(n2100), .B(n77551), .Y(
        n2101) );
  INVxp67_ASAP7_75t_SL U55010 ( .A(n63367), .Y(n62949) );
  AND2x2_ASAP7_75t_SL U55011 ( .A(n60336), .B(n77459), .Y(n77566) );
  NAND2xp5_ASAP7_75t_SL U55012 ( .A(n59694), .B(n77459), .Y(n77537) );
  OAI22xp33_ASAP7_75t_SL U55013 ( .A1(n1658), .A2(n77463), .B1(n59533), .B2(
        n57074), .Y(n74989) );
  AOI21xp33_ASAP7_75t_SL U55014 ( .A1(n69129), .A2(n57079), .B(n69128), .Y(
        n69136) );
  NAND2xp33_ASAP7_75t_SL U55015 ( .A(n77532), .B(n59690), .Y(n77533) );
  O2A1O1Ixp33_ASAP7_75t_SL U55016 ( .A1(n76167), .A2(n76166), .B(n76165), .C(
        n76164), .Y(n76168) );
  OAI21xp33_ASAP7_75t_SL U55017 ( .A1(n76145), .A2(n76144), .B(n76143), .Y(
        n76148) );
  NAND2xp33_ASAP7_75t_SL U55018 ( .A(n74790), .B(n59692), .Y(n77534) );
  AND2x2_ASAP7_75t_SL U55019 ( .A(n61013), .B(n59692), .Y(n77182) );
  INVxp67_ASAP7_75t_SL U55020 ( .A(n76628), .Y(n77912) );
  XNOR2xp5_ASAP7_75t_SL U55021 ( .A(n68504), .B(n68503), .Y(n68528) );
  NAND2xp33_ASAP7_75t_SL U55022 ( .A(n77550), .B(n57073), .Y(n77551) );
  INVxp67_ASAP7_75t_SL U55023 ( .A(n70947), .Y(n70943) );
  NAND2xp33_ASAP7_75t_SL U55024 ( .A(n60995), .B(n59691), .Y(n77849) );
  NAND2xp33_ASAP7_75t_SL U55025 ( .A(n58331), .B(n70947), .Y(n70949) );
  NAND2xp5_ASAP7_75t_SL U55026 ( .A(n57684), .B(n57685), .Y(n57683) );
  INVxp67_ASAP7_75t_SL U55027 ( .A(n68434), .Y(n59203) );
  NAND2xp5_ASAP7_75t_SL U55028 ( .A(n71052), .B(n71021), .Y(n71037) );
  XOR2xp5_ASAP7_75t_SL U55029 ( .A(n64630), .B(n64631), .Y(n64632) );
  NAND2xp33_ASAP7_75t_SL U55030 ( .A(n77554), .B(n59690), .Y(n77555) );
  NAND2xp33_ASAP7_75t_SL U55031 ( .A(n66898), .B(n66897), .Y(n66899) );
  NAND2xp33_ASAP7_75t_SL U55032 ( .A(n77530), .B(n59690), .Y(n77531) );
  NAND2x1p5_ASAP7_75t_SL U55033 ( .A(n61058), .B(n59691), .Y(n77467) );
  NAND2xp5_ASAP7_75t_SL U55034 ( .A(n58616), .B(n57074), .Y(n73961) );
  NAND2xp33_ASAP7_75t_SL U55035 ( .A(n77544), .B(n59690), .Y(n77545) );
  NAND2xp33_ASAP7_75t_SL U55036 ( .A(n77541), .B(n59690), .Y(n77542) );
  NAND2xp5_ASAP7_75t_SL U55037 ( .A(n66583), .B(n66582), .Y(n68637) );
  XOR2xp5_ASAP7_75t_SL U55038 ( .A(n63652), .B(n63240), .Y(n63644) );
  INVxp67_ASAP7_75t_SL U55039 ( .A(n68304), .Y(n68260) );
  INVxp67_ASAP7_75t_SL U55040 ( .A(n68305), .Y(n68261) );
  NAND2x1_ASAP7_75t_SL U55041 ( .A(n61125), .B(n59692), .Y(n77025) );
  XOR2xp5_ASAP7_75t_SL U55042 ( .A(n58503), .B(n68534), .Y(n59320) );
  INVxp33_ASAP7_75t_SL U55043 ( .A(n66445), .Y(n66448) );
  NAND2xp33_ASAP7_75t_SL U55044 ( .A(n77535), .B(n59690), .Y(n77536) );
  NAND2xp5_ASAP7_75t_SL U55045 ( .A(n3132), .B(n59692), .Y(n61009) );
  NAND2xp33_ASAP7_75t_SL U55046 ( .A(n64806), .B(n59693), .Y(n64802) );
  INVxp33_ASAP7_75t_SL U55047 ( .A(n65318), .Y(n74463) );
  NAND2xp33_ASAP7_75t_SL U55048 ( .A(n77547), .B(n59690), .Y(n77548) );
  NAND2x1_ASAP7_75t_SL U55049 ( .A(n61316), .B(n59692), .Y(n77409) );
  NAND2xp33_ASAP7_75t_SL U55050 ( .A(n77913), .B(n59692), .Y(n76221) );
  NAND2xp33_ASAP7_75t_SL U55051 ( .A(n77538), .B(n59690), .Y(n77539) );
  INVx2_ASAP7_75t_SL U55052 ( .A(n76909), .Y(n75650) );
  NAND2xp33_ASAP7_75t_SL U55053 ( .A(n77528), .B(n59690), .Y(n77529) );
  NAND2xp33_ASAP7_75t_SL U55054 ( .A(n77512), .B(n59691), .Y(n77513) );
  INVxp67_ASAP7_75t_SL U55055 ( .A(n62861), .Y(n62812) );
  NAND2xp33_ASAP7_75t_SL U55056 ( .A(n76745), .B(n59690), .Y(n76805) );
  AOI21xp33_ASAP7_75t_SL U55057 ( .A1(n59621), .A2(n58579), .B(n69822), .Y(
        n2293) );
  NAND2xp33_ASAP7_75t_SL U55058 ( .A(n77514), .B(n59691), .Y(n77515) );
  NAND2xp33_ASAP7_75t_SL U55059 ( .A(n77562), .B(n57073), .Y(n77563) );
  NAND2xp33_ASAP7_75t_SL U55060 ( .A(n62866), .B(n62867), .Y(n62852) );
  NAND2xp33_ASAP7_75t_SL U55061 ( .A(n77568), .B(n59690), .Y(n77569) );
  NOR2xp33_ASAP7_75t_SL U55062 ( .A(n71274), .B(n71273), .Y(n71294) );
  AOI21xp33_ASAP7_75t_SL U55063 ( .A1(n59621), .A2(n69842), .B(n69841), .Y(
        n2291) );
  NAND2xp33_ASAP7_75t_SL U55064 ( .A(n77516), .B(n59691), .Y(n77517) );
  XNOR2xp5_ASAP7_75t_SL U55065 ( .A(n64448), .B(n57770), .Y(n64703) );
  AOI21xp5_ASAP7_75t_SL U55066 ( .A1(n71749), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_1_), .B(
        n71748), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n115) );
  NAND2xp33_ASAP7_75t_SL U55067 ( .A(n69986), .B(n69987), .Y(n69992) );
  NAND2xp5_ASAP7_75t_SL U55068 ( .A(n61302), .B(n77472), .Y(n61997) );
  AOI21xp33_ASAP7_75t_SL U55069 ( .A1(n69857), .A2(n59621), .B(n69856), .Y(
        n2289) );
  AND3x1_ASAP7_75t_SL U55070 ( .A(n59694), .B(n77579), .C(n77578), .Y(finish)
         );
  INVxp33_ASAP7_75t_SL U55071 ( .A(n77472), .Y(n61308) );
  NAND2xp33_ASAP7_75t_SL U55072 ( .A(n77518), .B(n59691), .Y(n77519) );
  NAND2xp5_ASAP7_75t_SL U55073 ( .A(n76675), .B(n59690), .Y(n77685) );
  NAND2xp33_ASAP7_75t_SL U55074 ( .A(n77526), .B(n59690), .Y(n77527) );
  NAND2xp33_ASAP7_75t_SL U55075 ( .A(n77559), .B(n59690), .Y(n77560) );
  NAND2xp33_ASAP7_75t_SL U55076 ( .A(n77202), .B(n77201), .Y(n77205) );
  AOI21xp33_ASAP7_75t_SL U55077 ( .A1(n74943), .A2(n69353), .B(n69352), .Y(
        n69354) );
  INVxp33_ASAP7_75t_SL U55078 ( .A(n64193), .Y(n64195) );
  NAND2xp5_ASAP7_75t_SL U55079 ( .A(n61122), .B(n61121), .Y(n77900) );
  NAND2xp33_ASAP7_75t_SL U55080 ( .A(n59621), .B(n70010), .Y(n69967) );
  INVxp67_ASAP7_75t_SL U55081 ( .A(n67672), .Y(n67673) );
  NAND2xp33_ASAP7_75t_SL U55082 ( .A(n77520), .B(n59691), .Y(n77521) );
  AO21x1_ASAP7_75t_SL U55083 ( .A1(n74348), .A2(n74347), .B(n74385), .Y(n74349) );
  NAND2xp33_ASAP7_75t_SL U55084 ( .A(n77522), .B(n59690), .Y(n77523) );
  NAND2xp33_ASAP7_75t_SL U55085 ( .A(n64330), .B(n59693), .Y(n64327) );
  INVx1_ASAP7_75t_SL U55086 ( .A(n67574), .Y(n67527) );
  NAND2x1_ASAP7_75t_SL U55087 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_35_), .B(
        n74385), .Y(n74392) );
  NAND2xp5_ASAP7_75t_SL U55088 ( .A(n60341), .B(n59690), .Y(n60489) );
  INVxp67_ASAP7_75t_SL U55089 ( .A(n62914), .Y(n62917) );
  NAND2xp33_ASAP7_75t_SL U55090 ( .A(n77524), .B(n59690), .Y(n77525) );
  NAND2xp5_ASAP7_75t_SL U55091 ( .A(n60340), .B(n59691), .Y(n62071) );
  OAI21xp33_ASAP7_75t_SL U55092 ( .A1(n76906), .A2(n69217), .B(n69216), .Y(
        n69218) );
  NAND2xp33_ASAP7_75t_SL U55093 ( .A(n65363), .B(n65362), .Y(n1991) );
  INVxp67_ASAP7_75t_SL U55094 ( .A(n64995), .Y(n64947) );
  NAND2xp5_ASAP7_75t_SL U55095 ( .A(n65258), .B(n65318), .Y(n65267) );
  INVxp67_ASAP7_75t_SL U55096 ( .A(n64997), .Y(n64945) );
  INVxp33_ASAP7_75t_SL U55097 ( .A(n62549), .Y(n62552) );
  INVxp33_ASAP7_75t_SL U55098 ( .A(n69352), .Y(n63703) );
  NAND2xp33_ASAP7_75t_SL U55099 ( .A(n77564), .B(n57073), .Y(n77565) );
  INVxp67_ASAP7_75t_SL U55100 ( .A(n66897), .Y(n66836) );
  INVx1_ASAP7_75t_SL U55101 ( .A(n66992), .Y(n66896) );
  NAND2xp33_ASAP7_75t_SL U55102 ( .A(n74633), .B(n57074), .Y(n74632) );
  AOI22xp5_ASAP7_75t_SL U55103 ( .A1(n71744), .A2(n71729), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_2_), .B2(
        n71749), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n116) );
  NAND2xp33_ASAP7_75t_SL U55104 ( .A(n77557), .B(n57073), .Y(n77558) );
  INVxp67_ASAP7_75t_SL U55105 ( .A(n71734), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n117) );
  INVxp67_ASAP7_75t_SL U55106 ( .A(n66366), .Y(n66367) );
  NAND2xp33_ASAP7_75t_SL U55107 ( .A(n61035), .B(n59692), .Y(n61126) );
  INVxp33_ASAP7_75t_SL U55108 ( .A(n71050), .Y(n71021) );
  AOI21xp33_ASAP7_75t_SL U55109 ( .A1(n77413), .A2(n77750), .B(n77412), .Y(
        dwb_biu_N62) );
  NAND2xp33_ASAP7_75t_SL U55110 ( .A(n70231), .B(n58553), .Y(n70230) );
  AOI21xp33_ASAP7_75t_SL U55111 ( .A1(n77486), .A2(n77485), .B(n77487), .Y(
        n77490) );
  OAI21xp5_ASAP7_75t_SL U55112 ( .A1(n58151), .A2(n68403), .B(n57053), .Y(
        n58149) );
  XOR2xp5_ASAP7_75t_SL U55113 ( .A(icqmem_adr_qmem[30]), .B(n757), .Y(n60268)
         );
  INVxp67_ASAP7_75t_SL U55114 ( .A(n62731), .Y(n62732) );
  NAND2xp5_ASAP7_75t_SL U55115 ( .A(n64859), .B(n73945), .Y(n64860) );
  NOR2xp33_ASAP7_75t_SL U55116 ( .A(n69285), .B(n69214), .Y(n74117) );
  NAND2xp5_ASAP7_75t_SL U55117 ( .A(n70975), .B(n70939), .Y(n70947) );
  INVx1_ASAP7_75t_SL U55118 ( .A(n61267), .Y(n77919) );
  AOI21xp5_ASAP7_75t_SL U55119 ( .A1(n73429), .A2(n73450), .B(n73422), .Y(
        n73432) );
  NAND2xp33_ASAP7_75t_SL U55120 ( .A(n57079), .B(n69074), .Y(n69080) );
  AOI21xp33_ASAP7_75t_SL U55121 ( .A1(n64800), .A2(n77082), .B(n64799), .Y(
        n64801) );
  INVxp67_ASAP7_75t_SL U55122 ( .A(n66722), .Y(n59347) );
  INVxp67_ASAP7_75t_SL U55123 ( .A(n71132), .Y(n71135) );
  INVxp33_ASAP7_75t_SL U55124 ( .A(n76163), .Y(n76164) );
  INVxp67_ASAP7_75t_SL U55125 ( .A(n68950), .Y(n68971) );
  INVx1_ASAP7_75t_SL U55126 ( .A(n64557), .Y(n57685) );
  INVx1_ASAP7_75t_SL U55127 ( .A(n64431), .Y(n64435) );
  NAND2xp5_ASAP7_75t_SL U55128 ( .A(n71126), .B(n71120), .Y(n71124) );
  INVxp67_ASAP7_75t_SL U55129 ( .A(n62905), .Y(n62903) );
  OAI21xp33_ASAP7_75t_SL U55130 ( .A1(n76906), .A2(n68950), .B(n68947), .Y(
        n68948) );
  INVxp67_ASAP7_75t_SL U55131 ( .A(n76654), .Y(n77909) );
  AOI21xp33_ASAP7_75t_SL U55132 ( .A1(n71030), .A2(n71029), .B(n71028), .Y(
        n71031) );
  INVx2_ASAP7_75t_SL U55133 ( .A(n58553), .Y(n59621) );
  INVxp67_ASAP7_75t_SL U55134 ( .A(n62899), .Y(n62901) );
  INVx1_ASAP7_75t_SL U55135 ( .A(n74924), .Y(n74942) );
  AOI21xp33_ASAP7_75t_SL U55136 ( .A1(n69329), .A2(n57079), .B(n69314), .Y(
        n69315) );
  INVx1_ASAP7_75t_SL U55137 ( .A(n77173), .Y(n69341) );
  OAI21xp33_ASAP7_75t_SL U55138 ( .A1(n59671), .A2(n69329), .B(n69314), .Y(
        n69317) );
  INVxp67_ASAP7_75t_SL U55139 ( .A(n68600), .Y(n57844) );
  OAI21xp33_ASAP7_75t_SL U55140 ( .A1(n57081), .A2(n69821), .B(n69820), .Y(
        n69822) );
  NOR2xp33_ASAP7_75t_SL U55141 ( .A(n58617), .B(n69329), .Y(n75123) );
  NAND2xp5_ASAP7_75t_SL U55142 ( .A(n70733), .B(n70715), .Y(n70720) );
  NAND2xp33_ASAP7_75t_SL U55143 ( .A(n69867), .B(n58553), .Y(n69868) );
  INVx1_ASAP7_75t_SL U55144 ( .A(n64059), .Y(n63854) );
  OAI22xp33_ASAP7_75t_SL U55145 ( .A1(n71733), .A2(n71788), .B1(n71745), .B2(
        n71732), .Y(n71734) );
  OAI21xp33_ASAP7_75t_SL U55146 ( .A1(n57081), .A2(n69919), .B(n69918), .Y(
        n69920) );
  INVxp67_ASAP7_75t_SL U55147 ( .A(n64058), .Y(n63856) );
  INVx1_ASAP7_75t_SL U55148 ( .A(n76873), .Y(n77917) );
  INVxp67_ASAP7_75t_SL U55149 ( .A(n73566), .Y(n73561) );
  XNOR2xp5_ASAP7_75t_SL U55150 ( .A(n65012), .B(n68224), .Y(n68280) );
  INVxp33_ASAP7_75t_SL U55151 ( .A(n73585), .Y(n73565) );
  INVx1_ASAP7_75t_SL U55152 ( .A(n75472), .Y(n58840) );
  OAI21xp33_ASAP7_75t_SL U55153 ( .A1(n74338), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_33_), .B(
        n74348), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n22) );
  INVx1_ASAP7_75t_SL U55154 ( .A(n66518), .Y(n66436) );
  INVx1_ASAP7_75t_SL U55155 ( .A(n66514), .Y(n66515) );
  INVx1_ASAP7_75t_SL U55156 ( .A(n68271), .Y(n68275) );
  OAI21xp33_ASAP7_75t_SL U55157 ( .A1(n74413), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_19_), .B(
        n74423), .Y(n2399) );
  NAND2xp33_ASAP7_75t_SL U55158 ( .A(n59628), .B(n72985), .Y(n1547) );
  INVx1_ASAP7_75t_SL U55159 ( .A(n59270), .Y(n58693) );
  NAND2xp5_ASAP7_75t_SL U55160 ( .A(n59499), .B(n76304), .Y(n61121) );
  XNOR2xp5_ASAP7_75t_SL U55161 ( .A(n63226), .B(n63225), .Y(n63625) );
  INVxp33_ASAP7_75t_SL U55162 ( .A(n66276), .Y(n66274) );
  XNOR2xp5_ASAP7_75t_SL U55163 ( .A(n63619), .B(n63618), .Y(n63623) );
  XNOR2xp5_ASAP7_75t_SL U55164 ( .A(n57438), .B(n57928), .Y(n68208) );
  OAI21xp33_ASAP7_75t_SL U55165 ( .A1(n58679), .A2(n58710), .B(n58678), .Y(
        n58682) );
  XNOR2xp5_ASAP7_75t_SL U55166 ( .A(n62937), .B(n62839), .Y(n62915) );
  INVxp67_ASAP7_75t_SL U55167 ( .A(n63232), .Y(n63119) );
  INVxp33_ASAP7_75t_SL U55168 ( .A(n4099), .Y(n75173) );
  XNOR2xp5_ASAP7_75t_SL U55169 ( .A(n66507), .B(n66435), .Y(n66518) );
  NAND2xp5_ASAP7_75t_SL U55170 ( .A(n78208), .B(n4099), .Y(icqmem_adr_qmem[29]) );
  INVxp33_ASAP7_75t_SL U55171 ( .A(n64269), .Y(n64274) );
  NAND2xp33_ASAP7_75t_SL U55172 ( .A(n70313), .B(n70372), .Y(n70312) );
  INVx1_ASAP7_75t_SL U55173 ( .A(n64665), .Y(n57141) );
  AOI211xp5_ASAP7_75t_SRAM U55174 ( .A1(n65402), .A2(n65353), .B(n65401), .C(
        n65361), .Y(n65359) );
  AOI21xp33_ASAP7_75t_SL U55175 ( .A1(n77128), .A2(n77618), .B(n61739), .Y(
        n61740) );
  AOI22xp33_ASAP7_75t_SL U55176 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[21]), .A2(n70502), .B1(
        n70521), .B2(n70372), .Y(n70012) );
  NAND2xp33_ASAP7_75t_SL U55177 ( .A(n70520), .B(n70372), .Y(n69989) );
  NAND2xp33_ASAP7_75t_SL U55178 ( .A(n73571), .B(n73573), .Y(n73563) );
  OA21x2_ASAP7_75t_SL U55179 ( .A1(n74403), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_18_), 
        .B(n74312), .Y(n74310) );
  AOI22xp33_ASAP7_75t_SL U55180 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[19]), .A2(n70502), .B1(
        n70519), .B2(n70372), .Y(n69966) );
  INVxp67_ASAP7_75t_SL U55181 ( .A(n76807), .Y(n76745) );
  NAND2xp5_ASAP7_75t_SL U55182 ( .A(n69960), .B(n69934), .Y(n69969) );
  OAI21xp33_ASAP7_75t_SL U55183 ( .A1(n76744), .A2(n77612), .B(n61375), .Y(
        n61376) );
  OAI21xp33_ASAP7_75t_SL U55184 ( .A1(n76744), .A2(n77614), .B(n61797), .Y(
        n61802) );
  INVxp67_ASAP7_75t_SL U55185 ( .A(n62998), .Y(n62713) );
  NAND2xp33_ASAP7_75t_SL U55186 ( .A(n70518), .B(n70372), .Y(n69936) );
  AO22x1_ASAP7_75t_SL U55187 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[23]), .A2(n70502), .B1(
        n70524), .B2(n70372), .Y(n70069) );
  NAND2xp33_ASAP7_75t_SL U55188 ( .A(n70497), .B(n70372), .Y(n69918) );
  NAND2xp5_ASAP7_75t_SL U55189 ( .A(n67134), .B(n67135), .Y(n58681) );
  NOR4xp25_ASAP7_75t_SL U55190 ( .A(n60170), .B(n60169), .C(n60168), .D(n60167), .Y(n60184) );
  INVx1_ASAP7_75t_SL U55191 ( .A(n68611), .Y(n68610) );
  AOI22xp33_ASAP7_75t_SL U55192 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[15]), .A2(n70502), .B1(
        n70517), .B2(n70372), .Y(n69888) );
  INVx1_ASAP7_75t_SL U55193 ( .A(n70372), .Y(n70422) );
  INVx1_ASAP7_75t_SL U55194 ( .A(n77284), .Y(n77680) );
  INVxp33_ASAP7_75t_SL U55195 ( .A(n60716), .Y(n60717) );
  INVx1_ASAP7_75t_SL U55196 ( .A(n67695), .Y(n67696) );
  NAND2xp33_ASAP7_75t_SL U55197 ( .A(n70494), .B(n70372), .Y(n69854) );
  OAI22xp33_ASAP7_75t_SL U55198 ( .A1(n59700), .A2(n77820), .B1(n57084), .B2(
        n896), .Y(n897) );
  AOI21xp33_ASAP7_75t_SL U55199 ( .A1(n77593), .A2(n77128), .B(n61564), .Y(
        n76873) );
  AOI21xp5_ASAP7_75t_SL U55200 ( .A1(n69313), .A2(n69312), .B(n69311), .Y(
        n69329) );
  NAND2xp33_ASAP7_75t_SL U55201 ( .A(n70493), .B(n70372), .Y(n69839) );
  NAND2xp5_ASAP7_75t_SL U55202 ( .A(n75772), .B(n76693), .Y(n77161) );
  NAND2xp33_ASAP7_75t_SL U55203 ( .A(n70492), .B(n70372), .Y(n69820) );
  INVx1_ASAP7_75t_SL U55204 ( .A(n77009), .Y(n77915) );
  INVxp33_ASAP7_75t_SL U55205 ( .A(n70752), .Y(n70749) );
  AOI22xp33_ASAP7_75t_SL U55206 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[10]), .A2(n70502), .B1(
        n70516), .B2(n70372), .Y(n69806) );
  OAI21xp33_ASAP7_75t_SL U55207 ( .A1(n77847), .A2(n77875), .B(n77655), .Y(
        n1505) );
  INVxp33_ASAP7_75t_SL U55208 ( .A(n64663), .Y(n64668) );
  OAI21xp33_ASAP7_75t_SL U55209 ( .A1(n77847), .A2(n77873), .B(n77661), .Y(
        n1487) );
  AO21x1_ASAP7_75t_SL U55210 ( .A1(n74326), .A2(n74325), .B(n74338), .Y(n74327) );
  INVxp33_ASAP7_75t_SL U55211 ( .A(n65353), .Y(n65334) );
  NAND2xp5_ASAP7_75t_SL U55212 ( .A(n71457), .B(n71493), .Y(n71509) );
  INVxp67_ASAP7_75t_SL U55213 ( .A(n71133), .Y(n71120) );
  INVxp67_ASAP7_75t_SL U55214 ( .A(n70875), .Y(n70879) );
  NAND2xp5_ASAP7_75t_SL U55215 ( .A(n62492), .B(n62491), .Y(n62496) );
  NAND2xp5_ASAP7_75t_SL U55216 ( .A(n71302), .B(n71253), .Y(n71260) );
  INVxp67_ASAP7_75t_SL U55217 ( .A(n62864), .Y(n62789) );
  INVx1_ASAP7_75t_SL U55218 ( .A(n67797), .Y(n57801) );
  INVxp67_ASAP7_75t_SL U55219 ( .A(n62865), .Y(n62853) );
  INVx1_ASAP7_75t_SL U55220 ( .A(n77631), .Y(n1705) );
  NAND2xp33_ASAP7_75t_SL U55221 ( .A(n71127), .B(n71126), .Y(n71128) );
  OAI21xp33_ASAP7_75t_SL U55222 ( .A1(n71952), .A2(n71445), .B(n71444), .Y(
        n71458) );
  INVxp67_ASAP7_75t_SL U55223 ( .A(n71802), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n112) );
  AOI22xp5_ASAP7_75t_SL U55224 ( .A1(n77672), .A2(n77859), .B1(n77671), .B2(
        n77668), .Y(n52475) );
  AOI22xp33_ASAP7_75t_SL U55225 ( .A1(n77672), .A2(n77856), .B1(n77671), .B2(
        n77670), .Y(n1697) );
  INVxp67_ASAP7_75t_SL U55226 ( .A(n67011), .Y(n67015) );
  INVxp67_ASAP7_75t_SL U55227 ( .A(n62931), .Y(n62798) );
  AOI21xp5_ASAP7_75t_SL U55228 ( .A1(n77618), .A2(n77675), .B(n77617), .Y(
        n1113) );
  INVxp67_ASAP7_75t_SL U55229 ( .A(n71214), .Y(n58294) );
  AOI21xp33_ASAP7_75t_SL U55230 ( .A1(n69077), .A2(n59672), .B(n69076), .Y(
        n69079) );
  INVxp33_ASAP7_75t_SL U55231 ( .A(n69077), .Y(n69074) );
  NAND2xp5_ASAP7_75t_SL U55232 ( .A(n69165), .B(n69113), .Y(n69130) );
  INVx1_ASAP7_75t_SL U55233 ( .A(n74217), .Y(n74219) );
  NAND2xp33_ASAP7_75t_SL U55234 ( .A(n71170), .B(n71169), .Y(n71267) );
  INVxp33_ASAP7_75t_SL U55235 ( .A(n71169), .Y(n71167) );
  OR4x1_ASAP7_75t_SL U55236 ( .A(n78199), .B(n78198), .C(n76976), .D(n74213), 
        .Y(n74214) );
  OAI21xp33_ASAP7_75t_SL U55237 ( .A1(n76906), .A2(n68911), .B(n68894), .Y(
        n68895) );
  NAND2xp33_ASAP7_75t_SL U55238 ( .A(n61285), .B(n61286), .Y(n61288) );
  INVxp33_ASAP7_75t_SL U55239 ( .A(n74633), .Y(n74635) );
  OAI22xp33_ASAP7_75t_SL U55240 ( .A1(n62871), .A2(n62851), .B1(n62850), .B2(
        n62869), .Y(n57990) );
  NOR2xp33_ASAP7_75t_SL U55241 ( .A(n58029), .B(n58028), .Y(n58027) );
  INVx1_ASAP7_75t_SL U55242 ( .A(n71400), .Y(n71389) );
  NAND2xp5_ASAP7_75t_SL U55243 ( .A(n71794), .B(n71796), .Y(n71788) );
  INVx1_ASAP7_75t_SL U55244 ( .A(n71129), .Y(n71110) );
  NAND2xp5_ASAP7_75t_SL U55245 ( .A(n69198), .B(n69197), .Y(n74568) );
  INVx1_ASAP7_75t_SL U55246 ( .A(n67046), .Y(n67047) );
  INVxp67_ASAP7_75t_SL U55247 ( .A(n66833), .Y(n66834) );
  NOR2x1_ASAP7_75t_SL U55248 ( .A(n59114), .B(n67378), .Y(n67767) );
  INVxp67_ASAP7_75t_SL U55249 ( .A(n73419), .Y(n73421) );
  NAND2xp5_ASAP7_75t_SL U55250 ( .A(n71022), .B(n70960), .Y(n70962) );
  AOI22xp33_ASAP7_75t_SL U55251 ( .A1(n77672), .A2(n77880), .B1(n77675), .B2(
        n77653), .Y(n1622) );
  NAND2xp5_ASAP7_75t_SL U55252 ( .A(n64595), .B(n64596), .Y(n64602) );
  NAND2xp5_ASAP7_75t_SL U55253 ( .A(n64529), .B(n64531), .Y(n64534) );
  INVxp33_ASAP7_75t_SL U55254 ( .A(n70970), .Y(n70966) );
  NOR2xp67_ASAP7_75t_SL U55255 ( .A(n67004), .B(n57547), .Y(n57546) );
  OAI21xp33_ASAP7_75t_SL U55256 ( .A1(or1200_dc_top_dirty), .A2(n61993), .B(
        n61306), .Y(n61307) );
  AOI21xp33_ASAP7_75t_SL U55257 ( .A1(n64857), .A2(n64856), .B(n64855), .Y(
        n64859) );
  INVxp67_ASAP7_75t_SL U55258 ( .A(n70857), .Y(n70842) );
  NAND2xp33_ASAP7_75t_SL U55259 ( .A(n61299), .B(n61298), .Y(n61300) );
  INVxp33_ASAP7_75t_SL U55260 ( .A(n71327), .Y(n58310) );
  NAND2xp5_ASAP7_75t_SL U55261 ( .A(n66222), .B(n66221), .Y(n74217) );
  AOI21xp5_ASAP7_75t_SL U55262 ( .A1(n75295), .A2(n69196), .B(n69199), .Y(
        n69197) );
  NAND2xp5_ASAP7_75t_SL U55263 ( .A(n66557), .B(n66319), .Y(n66320) );
  INVx1_ASAP7_75t_SL U55264 ( .A(n66813), .Y(n66762) );
  INVxp67_ASAP7_75t_SL U55265 ( .A(n73409), .Y(n73411) );
  INVx1_ASAP7_75t_SL U55266 ( .A(n63236), .Y(n63152) );
  INVxp67_ASAP7_75t_SL U55267 ( .A(n70973), .Y(n70940) );
  AOI21xp33_ASAP7_75t_SL U55268 ( .A1(n77921), .A2(n61058), .B(n61057), .Y(
        n69338) );
  AOI22xp33_ASAP7_75t_SL U55269 ( .A1(n77112), .A2(n75374), .B1(n77128), .B2(
        n77650), .Y(n75383) );
  INVxp67_ASAP7_75t_SL U55270 ( .A(n63056), .Y(n63057) );
  NAND2xp5_ASAP7_75t_SL U55271 ( .A(n69093), .B(n69092), .Y(n69113) );
  INVxp33_ASAP7_75t_SL U55272 ( .A(n71491), .Y(n71445) );
  OAI21xp33_ASAP7_75t_SL U55273 ( .A1(n63075), .A2(n63074), .B(n63073), .Y(
        n63076) );
  AOI21xp5_ASAP7_75t_SL U55274 ( .A1(n71491), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), 
        .B(n71456), .Y(n71493) );
  AOI22xp33_ASAP7_75t_SL U55275 ( .A1(n77672), .A2(n77871), .B1(n77675), .B2(
        n77662), .Y(n1603) );
  OAI21xp33_ASAP7_75t_SL U55276 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_30_), .A2(n71119), 
        .B(n59523), .Y(n71133) );
  NAND2xp5_ASAP7_75t_SL U55277 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_30_), .B(n71119), 
        .Y(n71126) );
  AOI22xp33_ASAP7_75t_SL U55278 ( .A1(n77672), .A2(n77888), .B1(n77675), .B2(
        n77650), .Y(n1668) );
  INVxp33_ASAP7_75t_SL U55279 ( .A(n70836), .Y(n70838) );
  AOI21xp33_ASAP7_75t_SL U55280 ( .A1(n64250), .A2(n77664), .B(n64249), .Y(
        n64253) );
  INVxp33_ASAP7_75t_SL U55281 ( .A(n76162), .Y(n76167) );
  AOI22xp5_ASAP7_75t_SL U55282 ( .A1(n77672), .A2(n77883), .B1(n77675), .B2(
        n77652), .Y(n1637) );
  INVxp33_ASAP7_75t_SL U55283 ( .A(n62866), .Y(n62854) );
  OAI21xp33_ASAP7_75t_SL U55284 ( .A1(n76744), .A2(n77609), .B(n62389), .Y(
        n62390) );
  INVxp67_ASAP7_75t_SL U55285 ( .A(n71303), .Y(n71256) );
  OAI21xp5_ASAP7_75t_SL U55286 ( .A1(n77672), .A2(n77648), .B(n77647), .Y(
        n1702) );
  NAND2xp33_ASAP7_75t_SL U55287 ( .A(n77128), .B(n77652), .Y(n74633) );
  AOI22xp5_ASAP7_75t_SL U55288 ( .A1(n77672), .A2(n77877), .B1(n77675), .B2(
        n58557), .Y(n1701) );
  INVxp67_ASAP7_75t_SL U55289 ( .A(n66970), .Y(n57812) );
  OAI22xp33_ASAP7_75t_SL U55290 ( .A1(n59706), .A2(n77792), .B1(n57083), .B2(
        n1187), .Y(n1188) );
  INVxp33_ASAP7_75t_SL U55291 ( .A(n71297), .Y(n71253) );
  NAND2xp33_ASAP7_75t_SL U55292 ( .A(n71236), .B(n71235), .Y(n71237) );
  INVxp67_ASAP7_75t_SL U55293 ( .A(n71236), .Y(n71218) );
  INVxp67_ASAP7_75t_SL U55294 ( .A(n77669), .Y(n77670) );
  NAND2xp5_ASAP7_75t_SL U55295 ( .A(n70873), .B(n70872), .Y(n70874) );
  INVx1_ASAP7_75t_SL U55296 ( .A(n58331), .Y(n70974) );
  INVxp33_ASAP7_75t_SL U55297 ( .A(n53458), .Y(n62799) );
  INVxp33_ASAP7_75t_SL U55298 ( .A(n75883), .Y(n75213) );
  INVxp67_ASAP7_75t_SL U55299 ( .A(n68452), .Y(n68451) );
  INVxp67_ASAP7_75t_SL U55300 ( .A(n66410), .Y(n66361) );
  NAND2xp33_ASAP7_75t_SL U55301 ( .A(n68597), .B(n68596), .Y(n68599) );
  AOI21xp33_ASAP7_75t_SL U55302 ( .A1(n77128), .A2(n77596), .B(n61461), .Y(
        n77009) );
  OAI21xp33_ASAP7_75t_SL U55303 ( .A1(n74320), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_31_), .B(
        n74326), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n18) );
  AOI21xp33_ASAP7_75t_SL U55304 ( .A1(n74405), .A2(n74404), .B(n74403), .Y(
        n74410) );
  AOI21xp33_ASAP7_75t_SL U55305 ( .A1(n69852), .A2(n69859), .B(n69851), .Y(
        n69857) );
  NAND2xp33_ASAP7_75t_SL U55306 ( .A(n76544), .B(n76543), .Y(n77284) );
  INVxp33_ASAP7_75t_SL U55307 ( .A(n77921), .Y(n61017) );
  OAI21xp33_ASAP7_75t_SL U55308 ( .A1(n60728), .A2(n61021), .B(n60715), .Y(
        n60716) );
  NAND2xp5_ASAP7_75t_SL U55309 ( .A(n71721), .B(n71798), .Y(n71745) );
  NAND2x1p5_ASAP7_75t_SL U55310 ( .A(n57936), .B(n67870), .Y(n68131) );
  XNOR2xp5_ASAP7_75t_SL U55311 ( .A(n805), .B(icqmem_adr_qmem[18]), .Y(n60169)
         );
  NAND2xp5_ASAP7_75t_SL U55312 ( .A(n73454), .B(n73453), .Y(n73466) );
  INVxp33_ASAP7_75t_SL U55313 ( .A(n4101), .Y(n75170) );
  INVxp67_ASAP7_75t_SL U55314 ( .A(n68360), .Y(n68364) );
  AO21x1_ASAP7_75t_SL U55315 ( .A1(n59700), .A2(n77805), .B(n77804), .Y(n77806) );
  AOI21xp33_ASAP7_75t_SL U55316 ( .A1(n77128), .A2(n77648), .B(n77127), .Y(
        n77131) );
  INVxp67_ASAP7_75t_SL U55317 ( .A(n68220), .Y(n65007) );
  XNOR2xp5_ASAP7_75t_SL U55318 ( .A(n58362), .B(n68219), .Y(n68273) );
  OAI21xp33_ASAP7_75t_SL U55319 ( .A1(n68222), .A2(n68221), .B(n68220), .Y(
        n68223) );
  INVxp33_ASAP7_75t_SL U55320 ( .A(n74925), .Y(n63702) );
  INVx1_ASAP7_75t_SL U55321 ( .A(n61021), .Y(n77923) );
  MAJx2_ASAP7_75t_SL U55322 ( .A(n68184), .B(n68182), .C(n68180), .Y(n59313)
         );
  INVxp67_ASAP7_75t_SL U55323 ( .A(n68612), .Y(n75067) );
  OAI21xp33_ASAP7_75t_SL U55324 ( .A1(n69910), .A2(n69886), .B(n69892), .Y(
        n69889) );
  INVxp67_ASAP7_75t_SL U55325 ( .A(n77190), .Y(n77192) );
  INVxp67_ASAP7_75t_SL U55326 ( .A(n57973), .Y(n57972) );
  AOI22xp5_ASAP7_75t_SL U55327 ( .A1(n77672), .A2(n77866), .B1(n77675), .B2(
        n77665), .Y(n1567) );
  XNOR2xp5_ASAP7_75t_SL U55328 ( .A(n769), .B(icqmem_adr_qmem[27]), .Y(n60188)
         );
  XOR2xp5_ASAP7_75t_SL U55329 ( .A(icqmem_adr_qmem[25]), .B(n777), .Y(n60183)
         );
  INVx1_ASAP7_75t_SL U55330 ( .A(n75269), .Y(n77668) );
  NAND2xp33_ASAP7_75t_SL U55331 ( .A(n71344), .B(n71386), .Y(n71348) );
  OAI21xp33_ASAP7_75t_SL U55332 ( .A1(n74409), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_17_), .B(
        n74408), .Y(n2323) );
  AOI21xp33_ASAP7_75t_SL U55333 ( .A1(n77599), .A2(n77128), .B(n61666), .Y(
        n77913) );
  NAND2xp5_ASAP7_75t_SL U55334 ( .A(n77847), .B(n77654), .Y(n77655) );
  NAND2xp5_ASAP7_75t_SL U55335 ( .A(n77999), .B(n77484), .Y(n77766) );
  NAND2xp5_ASAP7_75t_SL U55336 ( .A(n61696), .B(n61695), .Y(n77618) );
  INVxp67_ASAP7_75t_SL U55337 ( .A(n62870), .Y(n62851) );
  OAI22xp33_ASAP7_75t_SL U55338 ( .A1(n59706), .A2(n77791), .B1(n57083), .B2(
        n1192), .Y(n1193) );
  INVxp67_ASAP7_75t_SL U55339 ( .A(n66889), .Y(n66887) );
  OAI21xp33_ASAP7_75t_SL U55340 ( .A1(n76508), .A2(n76890), .B(n62402), .Y(
        n9266) );
  NAND2xp5_ASAP7_75t_SL U55341 ( .A(n69910), .B(n69886), .Y(n69892) );
  OAI21xp5_ASAP7_75t_SL U55342 ( .A1(n73479), .A2(n73478), .B(n73477), .Y(
        n12827) );
  AOI21xp33_ASAP7_75t_SL U55343 ( .A1(n73269), .A2(n73462), .B(n73214), .Y(
        n73419) );
  INVx1_ASAP7_75t_SL U55344 ( .A(n68214), .Y(n57145) );
  NOR2x1_ASAP7_75t_SL U55345 ( .A(n64940), .B(n59049), .Y(n65013) );
  INVxp67_ASAP7_75t_SL U55346 ( .A(n64348), .Y(n64074) );
  NOR3xp33_ASAP7_75t_SRAM U55347 ( .A(n65364), .B(n65337), .C(n65354), .Y(
        n65291) );
  INVxp33_ASAP7_75t_SL U55348 ( .A(n65337), .Y(n65368) );
  INVxp67_ASAP7_75t_SL U55349 ( .A(n63211), .Y(n63638) );
  INVx1_ASAP7_75t_SL U55350 ( .A(n68438), .Y(n57146) );
  OAI22xp33_ASAP7_75t_SL U55351 ( .A1(n59706), .A2(n77788), .B1(n57083), .B2(
        n1252), .Y(n1253) );
  INVxp67_ASAP7_75t_SL U55352 ( .A(n66390), .Y(n66319) );
  OAI21xp33_ASAP7_75t_SL U55353 ( .A1(n59627), .A2(n72750), .B(n72748), .Y(
        n1762) );
  AOI21xp33_ASAP7_75t_SL U55354 ( .A1(n73422), .A2(n73418), .B(n73188), .Y(
        n73409) );
  INVxp33_ASAP7_75t_SL U55355 ( .A(n4103), .Y(n75160) );
  NAND2xp5_ASAP7_75t_SL U55356 ( .A(n64106), .B(n64105), .Y(n77653) );
  INVxp67_ASAP7_75t_SL U55357 ( .A(n68407), .Y(n66936) );
  OAI22xp33_ASAP7_75t_SL U55358 ( .A1(n59706), .A2(n77790), .B1(n57083), .B2(
        n1222), .Y(n1223) );
  INVxp67_ASAP7_75t_SL U55359 ( .A(n66823), .Y(n66825) );
  INVxp33_ASAP7_75t_SL U55360 ( .A(n64464), .Y(n64430) );
  INVx2_ASAP7_75t_SL U55361 ( .A(n67731), .Y(n57147) );
  XNOR2xp5_ASAP7_75t_SL U55362 ( .A(n63016), .B(n63015), .Y(n63017) );
  OAI21xp33_ASAP7_75t_SL U55363 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_5_), .A2(n59629), .B(
        n72828), .Y(n1837) );
  INVx1_ASAP7_75t_SL U55364 ( .A(n69865), .Y(n69851) );
  INVxp67_ASAP7_75t_SL U55365 ( .A(n66950), .Y(n58125) );
  INVx2_ASAP7_75t_SL U55366 ( .A(n63818), .Y(n57148) );
  XNOR2xp5_ASAP7_75t_SL U55367 ( .A(n67053), .B(n67054), .Y(n58795) );
  OAI21xp5_ASAP7_75t_SL U55368 ( .A1(n67869), .A2(n57494), .B(n59039), .Y(
        n68132) );
  INVxp67_ASAP7_75t_SL U55369 ( .A(n66969), .Y(n66642) );
  OAI21xp33_ASAP7_75t_SL U55370 ( .A1(n75796), .A2(n76890), .B(n75028), .Y(
        n9276) );
  INVxp67_ASAP7_75t_SL U55371 ( .A(n62886), .Y(n62885) );
  OAI22xp33_ASAP7_75t_SL U55372 ( .A1(n75648), .A2(n75647), .B1(n75646), .B2(
        n75645), .Y(n76892) );
  OAI21xp33_ASAP7_75t_SL U55373 ( .A1(n77966), .A2(n61618), .B(n61074), .Y(
        n77641) );
  INVxp67_ASAP7_75t_SL U55374 ( .A(n68112), .Y(n58712) );
  INVx1_ASAP7_75t_SL U55375 ( .A(n66496), .Y(n66405) );
  NAND2xp5_ASAP7_75t_SL U55376 ( .A(n72980), .B(n72979), .Y(n72981) );
  NAND2xp5_ASAP7_75t_SL U55377 ( .A(n66382), .B(n66381), .Y(n66430) );
  INVxp67_ASAP7_75t_SL U55378 ( .A(n62823), .Y(n62828) );
  INVxp33_ASAP7_75t_SL U55379 ( .A(n66574), .Y(n66577) );
  INVx1_ASAP7_75t_SL U55380 ( .A(n62871), .Y(n62849) );
  INVx1_ASAP7_75t_SL U55381 ( .A(n62868), .Y(n62850) );
  INVxp67_ASAP7_75t_SL U55382 ( .A(n66585), .Y(n66543) );
  OAI21xp33_ASAP7_75t_SL U55383 ( .A1(n75781), .A2(n76890), .B(n62405), .Y(
        n9265) );
  INVxp33_ASAP7_75t_SL U55384 ( .A(n4093), .Y(n77507) );
  NAND2xp5_ASAP7_75t_SL U55385 ( .A(n62484), .B(n62483), .Y(n62488) );
  INVxp33_ASAP7_75t_SL U55386 ( .A(n4133), .Y(n77315) );
  NAND2xp5_ASAP7_75t_SL U55387 ( .A(n64767), .B(n64766), .Y(n77662) );
  NAND2xp33_ASAP7_75t_SL U55388 ( .A(n73451), .B(n73269), .Y(n73270) );
  INVxp67_ASAP7_75t_SL U55389 ( .A(n67079), .Y(n67090) );
  AOI22xp5_ASAP7_75t_SL U55390 ( .A1(n77672), .A2(n77896), .B1(n77675), .B2(
        n77643), .Y(n1703) );
  INVxp67_ASAP7_75t_SL U55391 ( .A(n64893), .Y(n57587) );
  INVxp67_ASAP7_75t_SL U55392 ( .A(n67540), .Y(n67550) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U55393 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_0_), .A2(n65398), .B(
        n65376), .C(n65375), .Y(n1664) );
  OAI21xp5_ASAP7_75t_SL U55394 ( .A1(n67522), .A2(n67521), .B(n67520), .Y(
        n67539) );
  INVxp67_ASAP7_75t_SL U55395 ( .A(n67159), .Y(n57659) );
  INVx1_ASAP7_75t_SL U55396 ( .A(n67487), .Y(n57765) );
  INVx1_ASAP7_75t_SL U55397 ( .A(n58757), .Y(n58756) );
  NAND2xp5_ASAP7_75t_SL U55398 ( .A(n4128), .B(n78254), .Y(icqmem_adr_qmem[15]) );
  OAI21xp33_ASAP7_75t_SL U55399 ( .A1(n75632), .A2(n60014), .B(n59988), .Y(
        n60001) );
  INVxp33_ASAP7_75t_SL U55400 ( .A(n71391), .Y(n71387) );
  INVxp67_ASAP7_75t_SL U55401 ( .A(n62149), .Y(n63700) );
  INVxp67_ASAP7_75t_SL U55402 ( .A(n71385), .Y(n71401) );
  NAND2xp33_ASAP7_75t_SL U55403 ( .A(n77432), .B(n77441), .Y(n77431) );
  NAND2xp5_ASAP7_75t_SL U55404 ( .A(n73906), .B(n75884), .Y(n73948) );
  NAND2xp33_ASAP7_75t_SL U55405 ( .A(n71453), .B(n71472), .Y(n71454) );
  OAI21xp33_ASAP7_75t_SL U55406 ( .A1(n759), .A2(n77260), .B(n60009), .Y(
        n60015) );
  OAI21xp5_ASAP7_75t_SL U55407 ( .A1(n71384), .A2(n71383), .B(n71382), .Y(
        n71404) );
  INVx1_ASAP7_75t_SL U55408 ( .A(n61304), .Y(n61993) );
  NAND2xp5_ASAP7_75t_SL U55409 ( .A(n4126), .B(n78255), .Y(icqmem_adr_qmem[16]) );
  NAND2xp5_ASAP7_75t_SL U55410 ( .A(n4112), .B(n78263), .Y(icqmem_adr_qmem[23]) );
  INVx1_ASAP7_75t_SL U55411 ( .A(n71293), .Y(n71302) );
  INVxp67_ASAP7_75t_SL U55412 ( .A(n71027), .Y(n71028) );
  OAI21xp5_ASAP7_75t_SL U55413 ( .A1(n69289), .A2(n69288), .B(n69287), .Y(
        n69291) );
  NAND2xp5_ASAP7_75t_SL U55414 ( .A(n4116), .B(n78259), .Y(icqmem_adr_qmem[21]) );
  NAND2xp5_ASAP7_75t_SL U55415 ( .A(n71308), .B(n71266), .Y(n71279) );
  INVxp67_ASAP7_75t_SL U55416 ( .A(n60014), .Y(n59989) );
  NAND2xp5_ASAP7_75t_SL U55417 ( .A(n4118), .B(n78258), .Y(icqmem_adr_qmem[20]) );
  INVx1_ASAP7_75t_SL U55418 ( .A(n70861), .Y(n70858) );
  OAI21xp33_ASAP7_75t_SL U55419 ( .A1(n71362), .A2(n71146), .B(n71118), .Y(
        n71119) );
  OAI21xp33_ASAP7_75t_SL U55420 ( .A1(n71149), .A2(n71146), .B(n70989), .Y(
        n70991) );
  NAND2xp5_ASAP7_75t_SL U55421 ( .A(n71369), .B(n71383), .Y(n71360) );
  OAI21xp33_ASAP7_75t_SL U55422 ( .A1(n71984), .A2(n71487), .B(n71486), .Y(
        n71489) );
  INVxp67_ASAP7_75t_SL U55423 ( .A(n60464), .Y(n60457) );
  AOI211xp5_ASAP7_75t_SRAM U55424 ( .A1(n65402), .A2(n65337), .B(n65401), .C(
        n65342), .Y(n65341) );
  NAND2xp5_ASAP7_75t_SL U55425 ( .A(n4124), .B(n78256), .Y(icqmem_adr_qmem[17]) );
  INVxp67_ASAP7_75t_SL U55426 ( .A(n71340), .Y(n71386) );
  AOI21xp33_ASAP7_75t_SL U55427 ( .A1(n69195), .A2(n69194), .B(n69179), .Y(
        n69180) );
  INVxp67_ASAP7_75t_SL U55428 ( .A(n59890), .Y(n61319) );
  NAND2xp33_ASAP7_75t_SL U55429 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_4_), .B(n74179), 
        .Y(n74186) );
  INVxp67_ASAP7_75t_SL U55430 ( .A(n71324), .Y(n71344) );
  NAND2xp5_ASAP7_75t_SL U55431 ( .A(n61959), .B(n61958), .Y(n61960) );
  AO21x1_ASAP7_75t_SRAM U55432 ( .A1(n74315), .A2(n74314), .B(n74320), .Y(
        n74316) );
  NAND2xp5_ASAP7_75t_SL U55433 ( .A(n61291), .B(n61290), .Y(n61298) );
  NAND2xp5_ASAP7_75t_SL U55434 ( .A(n71235), .B(n71269), .Y(n71225) );
  NAND2xp5_ASAP7_75t_SL U55435 ( .A(n4120), .B(n78188), .Y(icqmem_adr_qmem[19]) );
  NAND2xp5_ASAP7_75t_SL U55436 ( .A(n70871), .B(n70870), .Y(n70967) );
  INVxp67_ASAP7_75t_SL U55437 ( .A(n71082), .Y(n71058) );
  INVxp67_ASAP7_75t_SL U55438 ( .A(n71272), .Y(n71196) );
  INVx1_ASAP7_75t_SL U55439 ( .A(n71113), .Y(n71111) );
  INVxp67_ASAP7_75t_SL U55440 ( .A(n61842), .Y(n61850) );
  NAND2xp5_ASAP7_75t_SL U55441 ( .A(n78204), .B(n4103), .Y(icqmem_adr_qmem[27]) );
  NAND2xp5_ASAP7_75t_SL U55442 ( .A(n78205), .B(n4110), .Y(icqmem_adr_qmem[24]) );
  OA21x2_ASAP7_75t_SL U55443 ( .A1(n74394), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_16_), 
        .B(n74405), .Y(n74395) );
  NAND2xp5_ASAP7_75t_SL U55444 ( .A(n78391), .B(n71234), .Y(n71303) );
  INVx1_ASAP7_75t_SL U55445 ( .A(n71136), .Y(n71098) );
  INVxp33_ASAP7_75t_SL U55446 ( .A(n71200), .Y(n71189) );
  INVxp33_ASAP7_75t_SL U55447 ( .A(n71600), .Y(n71626) );
  INVxp67_ASAP7_75t_SL U55448 ( .A(n70743), .Y(n70744) );
  AOI21xp5_ASAP7_75t_SL U55449 ( .A1(n69710), .A2(n69709), .B(n70090), .Y(
        n69716) );
  INVxp33_ASAP7_75t_SL U55450 ( .A(n71094), .Y(n71097) );
  INVxp67_ASAP7_75t_SL U55451 ( .A(n59078), .Y(n59077) );
  INVxp67_ASAP7_75t_SL U55452 ( .A(n70800), .Y(n70802) );
  OAI22xp33_ASAP7_75t_SL U55453 ( .A1(or1200_cpu_or1200_except_n604), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n419), .B2(n59676), .Y(n61341)
         );
  OAI21xp33_ASAP7_75t_SL U55454 ( .A1(or1200_cpu_or1200_except_n643), .A2(
        n59675), .B(n64281), .Y(n64286) );
  INVxp67_ASAP7_75t_SL U55455 ( .A(n66765), .Y(n66677) );
  OAI21xp5_ASAP7_75t_SL U55456 ( .A1(n71371), .A2(n71370), .B(n71369), .Y(
        n71391) );
  INVxp33_ASAP7_75t_SL U55457 ( .A(n60301), .Y(n60265) );
  NOR2x1_ASAP7_75t_SL U55458 ( .A(n57013), .B(n59103), .Y(n66872) );
  INVxp33_ASAP7_75t_SL U55459 ( .A(n71343), .Y(n71349) );
  NAND2xp33_ASAP7_75t_SL U55460 ( .A(n59629), .B(n72829), .Y(n72828) );
  AOI21xp33_ASAP7_75t_SL U55461 ( .A1(n76713), .A2(n77619), .B(n77624), .Y(
        n62461) );
  NAND2xp5_ASAP7_75t_SL U55462 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_27_), .B(n71084), 
        .Y(n71130) );
  OAI22xp33_ASAP7_75t_SL U55463 ( .A1(or1200_cpu_spr_dat_ppc[21]), .A2(n59676), 
        .B1(or1200_cpu_or1200_except_n144), .B2(n57102), .Y(n62102) );
  INVxp67_ASAP7_75t_SL U55464 ( .A(n77126), .Y(n77127) );
  OAI22xp33_ASAP7_75t_SL U55465 ( .A1(or1200_cpu_or1200_except_n595), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n410), .B2(n59676), .Y(n62248)
         );
  OAI21xp33_ASAP7_75t_SL U55466 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_9_), .A2(n59629), .B(
        n72799), .Y(n1808) );
  NAND2xp33_ASAP7_75t_SL U55467 ( .A(n59628), .B(n72870), .Y(n72869) );
  INVxp67_ASAP7_75t_SL U55468 ( .A(n66856), .Y(n57993) );
  NAND2xp33_ASAP7_75t_SL U55469 ( .A(n71353), .B(n71049), .Y(n71082) );
  AOI21xp33_ASAP7_75t_SL U55470 ( .A1(n73905), .A2(
        or1200_cpu_or1200_except_n542), .B(n76791), .Y(n73906) );
  OAI21xp33_ASAP7_75t_SL U55471 ( .A1(n71381), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_44_), .B(n71390), 
        .Y(n71399) );
  OAI22xp33_ASAP7_75t_SL U55472 ( .A1(or1200_cpu_or1200_except_n504), .A2(
        n77032), .B1(or1200_cpu_or1200_except_n416), .B2(n59676), .Y(n62329)
         );
  NAND2xp5_ASAP7_75t_SL U55473 ( .A(n71382), .B(n71390), .Y(n71374) );
  NAND2xp5_ASAP7_75t_SL U55474 ( .A(n74923), .B(n74922), .Y(n9486) );
  INVxp33_ASAP7_75t_SL U55475 ( .A(n75611), .Y(n75613) );
  INVxp33_ASAP7_75t_SL U55476 ( .A(n68479), .Y(n68482) );
  OAI21xp33_ASAP7_75t_SL U55477 ( .A1(n76906), .A2(n69085), .B(n69075), .Y(
        n69076) );
  AOI21xp5_ASAP7_75t_SL U55478 ( .A1(n70869), .A2(n59526), .B(n70868), .Y(
        n70870) );
  AOI21xp33_ASAP7_75t_SL U55479 ( .A1(n74387), .A2(n74386), .B(n74394), .Y(
        n74396) );
  INVx1_ASAP7_75t_SL U55480 ( .A(n66590), .Y(n66562) );
  INVx1_ASAP7_75t_SL U55481 ( .A(n67294), .Y(n59084) );
  INVxp67_ASAP7_75t_SL U55482 ( .A(n68439), .Y(n57622) );
  AOI21xp5_ASAP7_75t_SL U55483 ( .A1(n75605), .A2(n75604), .B(n75603), .Y(
        n75606) );
  NAND2xp5_ASAP7_75t_SL U55484 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_37_), .B(n71224), 
        .Y(n71235) );
  OAI21xp33_ASAP7_75t_SL U55485 ( .A1(n74355), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_29_), .B(
        n74315), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n14) );
  INVxp33_ASAP7_75t_SL U55486 ( .A(n60016), .Y(n60024) );
  BUFx2_ASAP7_75t_SL U55487 ( .A(n59229), .Y(n57273) );
  INVxp67_ASAP7_75t_SL U55488 ( .A(n70908), .Y(n70965) );
  NAND2xp5_ASAP7_75t_SL U55489 ( .A(n78393), .B(n71213), .Y(n71268) );
  OAI21xp33_ASAP7_75t_SL U55490 ( .A1(n62153), .A2(n60420), .B(n77368), .Y(
        n60308) );
  INVxp33_ASAP7_75t_SL U55491 ( .A(n70903), .Y(n70904) );
  OAI22xp33_ASAP7_75t_SL U55492 ( .A1(or1200_cpu_or1200_except_n482), .A2(
        n59676), .B1(or1200_cpu_or1200_except_n126), .B2(n57102), .Y(n75697)
         );
  NOR2xp33_ASAP7_75t_SL U55493 ( .A(n57278), .B(n57299), .Y(n57609) );
  OAI22xp33_ASAP7_75t_SL U55494 ( .A1(or1200_cpu_or1200_except_n661), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n476), .B2(n59676), .Y(n75830)
         );
  NAND2xp5_ASAP7_75t_SL U55495 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_44_), .B(n71381), 
        .Y(n71383) );
  INVxp67_ASAP7_75t_SL U55496 ( .A(n53464), .Y(n76013) );
  INVx1_ASAP7_75t_SL U55497 ( .A(n75066), .Y(n57149) );
  NAND2xp33_ASAP7_75t_SL U55498 ( .A(n78224), .B(n71539), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_mul_s_exp_10_o_9_) );
  INVxp67_ASAP7_75t_SL U55499 ( .A(n68362), .Y(n66920) );
  INVxp67_ASAP7_75t_SL U55500 ( .A(n75049), .Y(n75050) );
  OAI22xp33_ASAP7_75t_SL U55501 ( .A1(or1200_cpu_or1200_except_n583), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n398), .B2(n59676), .Y(n61261)
         );
  AOI21xp33_ASAP7_75t_SL U55502 ( .A1(n71117), .A2(n71394), .B(n71116), .Y(
        n71118) );
  NAND2xp33_ASAP7_75t_SL U55503 ( .A(n65402), .B(n65302), .Y(n2476) );
  INVxp67_ASAP7_75t_SL U55504 ( .A(n68601), .Y(n57845) );
  XNOR2xp5_ASAP7_75t_SL U55505 ( .A(n66869), .B(n66868), .Y(n66703) );
  OAI22xp33_ASAP7_75t_SL U55506 ( .A1(or1200_cpu_or1200_except_n496), .A2(
        n77032), .B1(or1200_cpu_or1200_except_n404), .B2(n59676), .Y(n61394)
         );
  INVxp67_ASAP7_75t_SL U55507 ( .A(n70830), .Y(n70831) );
  NAND2xp5_ASAP7_75t_SL U55508 ( .A(n70959), .B(n70958), .Y(n71022) );
  NOR2x1_ASAP7_75t_SL U55509 ( .A(n57015), .B(n67582), .Y(n67812) );
  OAI21xp33_ASAP7_75t_SL U55510 ( .A1(n67082), .A2(n67081), .B(n67080), .Y(
        n67089) );
  INVxp67_ASAP7_75t_SL U55511 ( .A(n71296), .Y(n71266) );
  NAND2xp33_ASAP7_75t_SL U55512 ( .A(n74956), .B(n60016), .Y(n60009) );
  INVxp67_ASAP7_75t_SL U55513 ( .A(n75941), .Y(n75934) );
  NAND2xp33_ASAP7_75t_SL U55514 ( .A(n73439), .B(n73283), .Y(n73284) );
  NAND2x1p5_ASAP7_75t_SL U55515 ( .A(n57528), .B(n57526), .Y(n65004) );
  OAI21xp5_ASAP7_75t_SL U55516 ( .A1(n73428), .A2(n73431), .B(n73176), .Y(
        n73422) );
  INVx1_ASAP7_75t_SL U55517 ( .A(n64556), .Y(n57150) );
  OA21x2_ASAP7_75t_SL U55518 ( .A1(n78055), .A2(n78054), .B(n78059), .Y(n78056) );
  NAND2xp5_ASAP7_75t_SL U55519 ( .A(n69885), .B(n69914), .Y(n69886) );
  AOI21xp33_ASAP7_75t_SL U55520 ( .A1(n62292), .A2(n61374), .B(n60990), .Y(
        n60991) );
  NAND2xp33_ASAP7_75t_SL U55521 ( .A(n64442), .B(n64440), .Y(n64387) );
  AOI21xp33_ASAP7_75t_SL U55522 ( .A1(n77051), .A2(n74044), .B(n64765), .Y(
        n64766) );
  OAI21xp5_ASAP7_75t_SL U55523 ( .A1(n74053), .A2(n74190), .B(n74052), .Y(
        n74061) );
  XNOR2xp5_ASAP7_75t_SL U55524 ( .A(n64402), .B(n64541), .Y(n64403) );
  INVxp67_ASAP7_75t_SL U55525 ( .A(n66764), .Y(n66613) );
  OAI21xp33_ASAP7_75t_SL U55526 ( .A1(n74167), .A2(n74190), .B(n74172), .Y(
        n74171) );
  OAI21xp33_ASAP7_75t_SL U55527 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_6_), .A2(n74190), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_7_), .Y(n74178)
         );
  AOI21xp33_ASAP7_75t_SL U55528 ( .A1(n69837), .A2(n69836), .B(n69861), .Y(
        n69842) );
  OAI21xp33_ASAP7_75t_SL U55529 ( .A1(n74174), .A2(n74190), .B(n74173), .Y(
        n74177) );
  OAI21xp33_ASAP7_75t_SL U55530 ( .A1(n74189), .A2(n74190), .B(n74188), .Y(
        n74185) );
  NAND2xp33_ASAP7_75t_SL U55531 ( .A(n77765), .B(n77764), .Y(n77768) );
  OAI22xp33_ASAP7_75t_SL U55532 ( .A1(or1200_cpu_or1200_except_n598), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n413), .B2(n59676), .Y(n76743)
         );
  OAI21xp33_ASAP7_75t_SL U55533 ( .A1(n74390), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_15_), .B(
        n74400), .Y(n2339) );
  NAND2xp5_ASAP7_75t_SL U55534 ( .A(n73479), .B(n73478), .Y(n73477) );
  INVxp67_ASAP7_75t_SL U55535 ( .A(n66735), .Y(n66614) );
  OAI21xp5_ASAP7_75t_SL U55536 ( .A1(n67480), .A2(n63841), .B(n58179), .Y(
        n64051) );
  OAI21xp33_ASAP7_75t_SL U55537 ( .A1(or1200_cpu_spr_dat_ppc[26]), .A2(n59676), 
        .B(n64817), .Y(n64823) );
  INVxp33_ASAP7_75t_SL U55538 ( .A(n73905), .Y(n64862) );
  INVxp67_ASAP7_75t_SL U55539 ( .A(n63857), .Y(n62847) );
  OAI21xp33_ASAP7_75t_SL U55540 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_17_), .A2(n59629), .B(
        n72735), .Y(n1662) );
  INVx1_ASAP7_75t_SL U55541 ( .A(n65005), .Y(n58048) );
  NOR2x1_ASAP7_75t_SL U55542 ( .A(n64754), .B(n75605), .Y(n64755) );
  NAND2xp5_ASAP7_75t_SL U55543 ( .A(n62826), .B(n62825), .Y(n62827) );
  OAI22xp33_ASAP7_75t_SL U55544 ( .A1(or1200_cpu_spr_dat_ppc[19]), .A2(n59676), 
        .B1(or1200_cpu_or1200_except_n148), .B2(n57102), .Y(n74591) );
  OAI22xp33_ASAP7_75t_SL U55545 ( .A1(or1200_cpu_or1200_except_n510), .A2(
        n77032), .B1(or1200_cpu_or1200_except_n425), .B2(n59676), .Y(n61692)
         );
  OAI22xp33_ASAP7_75t_SL U55546 ( .A1(or1200_cpu_or1200_except_n628), .A2(
        n59675), .B1(or1200_cpu_spr_dat_ppc[17]), .B2(n59676), .Y(n75373) );
  NAND2xp5_ASAP7_75t_SL U55547 ( .A(n60836), .B(n60835), .Y(n77643) );
  NAND2xp33_ASAP7_75t_SL U55548 ( .A(n59687), .B(n78084), .Y(n557) );
  INVxp33_ASAP7_75t_SL U55549 ( .A(n78084), .Y(n78083) );
  INVxp67_ASAP7_75t_SL U55550 ( .A(n64530), .Y(n64535) );
  NAND2xp33_ASAP7_75t_SL U55551 ( .A(n59687), .B(n78088), .Y(n555) );
  INVxp33_ASAP7_75t_SL U55552 ( .A(n78088), .Y(n78087) );
  OAI22xp33_ASAP7_75t_SL U55553 ( .A1(or1200_cpu_or1200_except_n625), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n440), .B2(n59676), .Y(n62513)
         );
  NAND2xp33_ASAP7_75t_SL U55554 ( .A(n71950), .B(n71599), .Y(n71600) );
  INVx1_ASAP7_75t_SL U55555 ( .A(n64451), .Y(n64452) );
  INVx1_ASAP7_75t_SL U55556 ( .A(n76592), .Y(n76521) );
  AOI21xp33_ASAP7_75t_SL U55557 ( .A1(n77051), .A2(n74126), .B(n64104), .Y(
        n64105) );
  XNOR2xp5_ASAP7_75t_SL U55558 ( .A(n62704), .B(n62703), .Y(n62705) );
  INVxp67_ASAP7_75t_SL U55559 ( .A(n64098), .Y(n64106) );
  INVxp67_ASAP7_75t_SL U55560 ( .A(n63031), .Y(n58874) );
  INVxp67_ASAP7_75t_SL U55561 ( .A(n61841), .Y(n61851) );
  OAI22xp33_ASAP7_75t_SL U55562 ( .A1(or1200_cpu_spr_dat_ppc[31]), .A2(n59676), 
        .B1(or1200_cpu_or1200_except_n124), .B2(n57102), .Y(n61842) );
  NOR2x1_ASAP7_75t_SL U55563 ( .A(n68157), .B(n68089), .Y(n59284) );
  NAND2xp5_ASAP7_75t_SL U55564 ( .A(n76001), .B(n53464), .Y(n76002) );
  INVxp67_ASAP7_75t_SL U55565 ( .A(n71785), .Y(n71797) );
  INVxp33_ASAP7_75t_SL U55566 ( .A(n66277), .Y(n66275) );
  NAND2xp5_ASAP7_75t_SL U55567 ( .A(n74775), .B(n74774), .Y(n9488) );
  NAND2xp5_ASAP7_75t_SL U55568 ( .A(n59133), .B(n68001), .Y(n57728) );
  NAND2xp5_ASAP7_75t_SL U55569 ( .A(n74786), .B(n74785), .Y(n52469) );
  NAND2xp33_ASAP7_75t_SL U55570 ( .A(n66431), .B(n66252), .Y(n66272) );
  NAND2xp5_ASAP7_75t_SL U55571 ( .A(n74769), .B(n74768), .Y(n9489) );
  INVxp33_ASAP7_75t_SL U55572 ( .A(n66646), .Y(n66626) );
  NAND2xp5_ASAP7_75t_SL U55573 ( .A(n60579), .B(n60578), .Y(n60580) );
  NAND2xp33_ASAP7_75t_SL U55574 ( .A(n78436), .B(n76480), .Y(n76506) );
  OAI22xp33_ASAP7_75t_SL U55575 ( .A1(or1200_cpu_or1200_except_n664), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n546), .B2(n77032), .Y(n75212)
         );
  OAI22xp33_ASAP7_75t_SL U55576 ( .A1(or1200_cpu_or1200_except_n658), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n542), .B2(n77032), .Y(n73914)
         );
  AOI21xp5_ASAP7_75t_SL U55577 ( .A1(n73582), .A2(n73553), .B(n73552), .Y(
        n73558) );
  INVxp67_ASAP7_75t_SL U55578 ( .A(n71342), .Y(n71352) );
  INVxp33_ASAP7_75t_SL U55579 ( .A(n71368), .Y(n71370) );
  INVxp33_ASAP7_75t_SL U55580 ( .A(n64146), .Y(n64149) );
  OAI22xp33_ASAP7_75t_SL U55581 ( .A1(or1200_cpu_or1200_except_n622), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n518), .B2(n77032), .Y(n77055)
         );
  OAI21xp33_ASAP7_75t_SL U55582 ( .A1(n73593), .A2(n73583), .B(n73582), .Y(
        n73654) );
  NAND2xp5_ASAP7_75t_SL U55583 ( .A(n71358), .B(n71359), .Y(n71369) );
  INVxp33_ASAP7_75t_SL U55584 ( .A(n62076), .Y(n62079) );
  INVxp67_ASAP7_75t_SL U55585 ( .A(n75816), .Y(n75828) );
  INVxp33_ASAP7_75t_SL U55586 ( .A(n63234), .Y(n63235) );
  NAND2xp33_ASAP7_75t_SL U55587 ( .A(n66419), .B(n67020), .Y(n66420) );
  INVx1_ASAP7_75t_SL U55588 ( .A(n63802), .Y(n57152) );
  NAND2xp33_ASAP7_75t_SL U55589 ( .A(n66412), .B(n66423), .Y(n66486) );
  INVxp67_ASAP7_75t_SL U55590 ( .A(n71322), .Y(n71320) );
  BUFx2_ASAP7_75t_SL U55591 ( .A(n67457), .Y(n57243) );
  NAND2xp5_ASAP7_75t_SL U55592 ( .A(n71379), .B(n71378), .Y(n71380) );
  NAND2xp5_ASAP7_75t_SL U55593 ( .A(n58105), .B(n58104), .Y(n58103) );
  OAI21xp33_ASAP7_75t_SL U55594 ( .A1(n62132), .A2(n75548), .B(n62131), .Y(
        n62136) );
  OAI22xp33_ASAP7_75t_SL U55595 ( .A1(or1200_cpu_or1200_except_n640), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n530), .B2(n77032), .Y(n62103)
         );
  NAND2xp5_ASAP7_75t_SL U55596 ( .A(n70128), .B(n70127), .Y(n70129) );
  INVx1_ASAP7_75t_SL U55597 ( .A(n64450), .Y(n64453) );
  OAI21xp33_ASAP7_75t_SL U55598 ( .A1(or1200_cpu_or1200_except_n140), .A2(
        n57102), .B(n75563), .Y(n75564) );
  INVxp67_ASAP7_75t_SL U55599 ( .A(n63075), .Y(n62772) );
  INVxp33_ASAP7_75t_SL U55600 ( .A(n63072), .Y(n63074) );
  INVxp67_ASAP7_75t_SL U55601 ( .A(n62719), .Y(n62704) );
  INVxp67_ASAP7_75t_SL U55602 ( .A(n62718), .Y(n62703) );
  OAI22xp33_ASAP7_75t_SL U55603 ( .A1(n71284), .A2(n71230), .B1(n71149), .B2(
        n71262), .Y(n71116) );
  INVxp67_ASAP7_75t_SL U55604 ( .A(n62997), .Y(n62712) );
  INVxp33_ASAP7_75t_SL U55605 ( .A(n77468), .Y(n77764) );
  INVxp67_ASAP7_75t_SL U55606 ( .A(n62908), .Y(n58061) );
  OAI21xp5_ASAP7_75t_SL U55607 ( .A1(n57410), .A2(n65042), .B(n59130), .Y(
        n64559) );
  INVx2_ASAP7_75t_SL U55608 ( .A(n67005), .Y(n57153) );
  INVxp67_ASAP7_75t_SL U55609 ( .A(n68415), .Y(n66791) );
  INVxp33_ASAP7_75t_SL U55610 ( .A(n66830), .Y(n66831) );
  INVxp67_ASAP7_75t_SL U55611 ( .A(n64583), .Y(n57584) );
  INVxp33_ASAP7_75t_SL U55612 ( .A(n62896), .Y(n62895) );
  INVxp33_ASAP7_75t_SL U55613 ( .A(n75568), .Y(n64317) );
  NAND2xp33_ASAP7_75t_SL U55614 ( .A(n69902), .B(n70067), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[6]) );
  NAND2xp5_ASAP7_75t_SL U55615 ( .A(n64573), .B(n64572), .Y(n64571) );
  INVxp67_ASAP7_75t_SL U55616 ( .A(n71061), .Y(n71062) );
  NAND2xp5_ASAP7_75t_SL U55617 ( .A(n71079), .B(n71078), .Y(n71084) );
  AOI21xp33_ASAP7_75t_SL U55618 ( .A1(n75568), .A2(n75567), .B(n75882), .Y(
        n75604) );
  INVxp67_ASAP7_75t_SL U55619 ( .A(n57098), .Y(n57392) );
  INVxp67_ASAP7_75t_SL U55620 ( .A(n64349), .Y(n64073) );
  INVxp67_ASAP7_75t_SL U55621 ( .A(n66748), .Y(n58799) );
  OAI21xp5_ASAP7_75t_SL U55622 ( .A1(n71365), .A2(n71223), .B(n71222), .Y(
        n71224) );
  OA21x2_ASAP7_75t_SL U55623 ( .A1(n74350), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_14_), 
        .B(n74387), .Y(n74351) );
  INVx1_ASAP7_75t_SL U55624 ( .A(n58501), .Y(n62964) );
  AOI21xp33_ASAP7_75t_SL U55625 ( .A1(n70043), .A2(n70083), .B(n70042), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[21]) );
  INVxp67_ASAP7_75t_SL U55626 ( .A(n68117), .Y(n68122) );
  NAND2xp5_ASAP7_75t_SL U55627 ( .A(n71250), .B(n71249), .Y(n71252) );
  NAND2xp5_ASAP7_75t_SL U55628 ( .A(n76738), .B(n76737), .Y(n76742) );
  NAND2xp5_ASAP7_75t_SL U55629 ( .A(n71265), .B(n71264), .Y(n71308) );
  OAI21xp33_ASAP7_75t_SL U55630 ( .A1(n59526), .A2(n70828), .B(n70791), .Y(
        n70793) );
  INVxp67_ASAP7_75t_SL U55631 ( .A(n71290), .Y(n71288) );
  INVxp67_ASAP7_75t_SL U55632 ( .A(n67083), .Y(n67080) );
  OAI22xp33_ASAP7_75t_SL U55633 ( .A1(n71142), .A2(n71362), .B1(n71335), .B2(
        n71141), .Y(n71143) );
  NAND2xp33_ASAP7_75t_SL U55634 ( .A(n76071), .B(n68602), .Y(n59111) );
  INVxp67_ASAP7_75t_SL U55635 ( .A(n62934), .Y(n62938) );
  AO21x1_ASAP7_75t_SL U55636 ( .A1(n74370), .A2(n74356), .B(n74355), .Y(n74357) );
  NAND2xp33_ASAP7_75t_SL U55637 ( .A(n69902), .B(n70043), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[5]) );
  NAND2xp5_ASAP7_75t_SL U55638 ( .A(n59059), .B(n58501), .Y(n63014) );
  INVxp33_ASAP7_75t_SL U55639 ( .A(n63007), .Y(n63010) );
  INVxp67_ASAP7_75t_SL U55640 ( .A(n71183), .Y(n71184) );
  OAI21xp33_ASAP7_75t_SL U55641 ( .A1(n59629), .A2(n72884), .B(n72883), .Y(
        n1758) );
  INVxp33_ASAP7_75t_SL U55642 ( .A(n76193), .Y(n75974) );
  OAI22xp33_ASAP7_75t_SL U55643 ( .A1(n66085), .A2(n65869), .B1(n65868), .B2(
        n65867), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n29) );
  OAI21xp33_ASAP7_75t_SL U55644 ( .A1(n70149), .A2(n69517), .B(n69516), .Y(
        n52520) );
  INVxp67_ASAP7_75t_SL U55645 ( .A(n76594), .Y(n61573) );
  NAND2xp33_ASAP7_75t_SL U55646 ( .A(n59629), .B(n72736), .Y(n72735) );
  OAI22xp33_ASAP7_75t_SL U55647 ( .A1(or1200_cpu_or1200_except_n634), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n526), .B2(n77032), .Y(n74592)
         );
  NAND2xp33_ASAP7_75t_SL U55648 ( .A(n59628), .B(n72736), .Y(n72737) );
  AOI22xp33_ASAP7_75t_SL U55649 ( .A1(n77275), .A2(n58554), .B1(n77051), .B2(
        n76210), .Y(n61616) );
  OAI22xp33_ASAP7_75t_SL U55650 ( .A1(or1200_cpu_or1200_except_n655), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n134), .B2(n57102), .Y(n64824)
         );
  INVxp67_ASAP7_75t_SL U55651 ( .A(n67751), .Y(n67753) );
  AOI22xp33_ASAP7_75t_SL U55652 ( .A1(n63972), .A2(n58554), .B1(n77051), .B2(
        n77018), .Y(n60835) );
  NAND2xp33_ASAP7_75t_SL U55653 ( .A(n66076), .B(n65938), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n20) );
  INVxp67_ASAP7_75t_SL U55654 ( .A(n67418), .Y(n58052) );
  OAI21xp33_ASAP7_75t_SL U55655 ( .A1(n70077), .A2(n69883), .B(n69882), .Y(
        n52519) );
  NAND2xp33_ASAP7_75t_SL U55656 ( .A(n77272), .B(n77271), .Y(n77273) );
  OAI21xp33_ASAP7_75t_SL U55657 ( .A1(n59627), .A2(n72811), .B(n72810), .Y(
        n1791) );
  NAND2xp5_ASAP7_75t_SL U55658 ( .A(n75026), .B(n75027), .Y(n75029) );
  AOI21xp33_ASAP7_75t_SL U55659 ( .A1(n70029), .A2(n70028), .B(n70027), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[47]) );
  AOI21xp33_ASAP7_75t_SL U55660 ( .A1(n75747), .A2(n62292), .B(n62291), .Y(
        n62293) );
  INVxp33_ASAP7_75t_SL U55661 ( .A(n4128), .Y(n63986) );
  AOI21xp33_ASAP7_75t_SL U55662 ( .A1(n69562), .A2(n70149), .B(n69513), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[42]) );
  INVxp33_ASAP7_75t_SL U55663 ( .A(n4130), .Y(n63983) );
  NAND2xp33_ASAP7_75t_SL U55664 ( .A(n73400), .B(n73388), .Y(n73397) );
  INVxp33_ASAP7_75t_SL U55665 ( .A(n72955), .Y(n72956) );
  INVxp67_ASAP7_75t_SL U55666 ( .A(n68373), .Y(n68376) );
  NOR2xp33_ASAP7_75t_SL U55667 ( .A(n763), .B(n60029), .Y(n60016) );
  OAI21xp33_ASAP7_75t_SL U55668 ( .A1(or1200_cpu_or1200_except_n180), .A2(
        n57102), .B(n61465), .Y(n61467) );
  NAND2xp5_ASAP7_75t_SL U55669 ( .A(n61338), .B(n61337), .Y(n61340) );
  NAND2xp33_ASAP7_75t_SL U55670 ( .A(n66076), .B(n65771), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n30) );
  NAND2xp5_ASAP7_75t_SL U55671 ( .A(n65413), .B(n65559), .Y(n65445) );
  NAND2xp33_ASAP7_75t_SL U55672 ( .A(n59628), .B(n73006), .Y(n3341) );
  OAI22xp33_ASAP7_75t_SL U55673 ( .A1(or1200_cpu_or1200_except_n631), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n150), .B2(n57102), .Y(n63560)
         );
  NAND2xp5_ASAP7_75t_SL U55674 ( .A(n69747), .B(n69883), .Y(n17028) );
  NAND2xp33_ASAP7_75t_SL U55675 ( .A(n66076), .B(n65963), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n16) );
  XNOR2xp5_ASAP7_75t_SL U55676 ( .A(n61833), .B(n62454), .Y(n61117) );
  NAND2xp5_ASAP7_75t_SL U55677 ( .A(n69831), .B(n69818), .Y(n69837) );
  NAND2xp33_ASAP7_75t_SL U55678 ( .A(n76133), .B(n76132), .Y(n76135) );
  OR2x2_ASAP7_75t_SL U55679 ( .A(n75926), .B(n76003), .Y(n58297) );
  NAND2xp33_ASAP7_75t_SL U55680 ( .A(n66076), .B(n66035), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n18) );
  AOI22xp33_ASAP7_75t_SL U55681 ( .A1(or1200_cpu_or1200_fpu_zero_conv), .A2(
        n74921), .B1(n74920), .B2(or1200_cpu_or1200_fpu_zero), .Y(n74922) );
  NAND2xp33_ASAP7_75t_SL U55682 ( .A(n74083), .B(n77051), .Y(n64213) );
  AOI21xp33_ASAP7_75t_SL U55683 ( .A1(n69517), .A2(n70149), .B(n69472), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[46]) );
  INVxp67_ASAP7_75t_SL U55684 ( .A(n67516), .Y(n67522) );
  NAND2xp5_ASAP7_75t_SL U55685 ( .A(n69747), .B(n70028), .Y(n17031) );
  INVx1_ASAP7_75t_SL U55686 ( .A(n73435), .Y(n73437) );
  INVxp33_ASAP7_75t_SL U55687 ( .A(n62401), .Y(n62396) );
  NAND2xp33_ASAP7_75t_SL U55688 ( .A(n69747), .B(n69571), .Y(n17027) );
  OAI21xp33_ASAP7_75t_SL U55689 ( .A1(n70149), .A2(n69515), .B(n69514), .Y(
        n52517) );
  AOI21xp5_ASAP7_75t_SL U55690 ( .A1(n75996), .A2(n75995), .B(n75994), .Y(
        n75997) );
  INVxp67_ASAP7_75t_SL U55691 ( .A(n62459), .Y(n60883) );
  INVx1_ASAP7_75t_SL U55692 ( .A(n73388), .Y(n73354) );
  OAI21xp33_ASAP7_75t_SL U55693 ( .A1(or1200_cpu_or1200_except_n138), .A2(
        n57102), .B(n64764), .Y(n64765) );
  NAND2xp33_ASAP7_75t_SL U55694 ( .A(or1200_cpu_or1200_fpu_inf), .B(n74920), 
        .Y(n74786) );
  NOR2x1_ASAP7_75t_SL U55695 ( .A(n60299), .B(n60298), .Y(n78440) );
  NAND2xp33_ASAP7_75t_SL U55696 ( .A(n59628), .B(n73022), .Y(n3340) );
  AOI21xp33_ASAP7_75t_SL U55697 ( .A1(n74920), .A2(
        or1200_cpu_or1200_fpu_underflow), .B(n74764), .Y(n74769) );
  AOI21xp33_ASAP7_75t_SL U55698 ( .A1(n69795), .A2(n70149), .B(n69504), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[43]) );
  OAI22xp33_ASAP7_75t_SL U55699 ( .A1(or1200_cpu_or1200_except_n637), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n146), .B2(n57102), .Y(n64098)
         );
  AOI21xp33_ASAP7_75t_SL U55700 ( .A1(n60029), .A2(n763), .B(n77260), .Y(
        n60023) );
  OAI21xp33_ASAP7_75t_SL U55701 ( .A1(n59627), .A2(n72842), .B(n72841), .Y(
        n1990) );
  NOR2xp33_ASAP7_75t_SRAM U55702 ( .A(n77943), .B(n61343), .Y(n61344) );
  OAI21xp33_ASAP7_75t_SL U55703 ( .A1(n70149), .A2(n69795), .B(n69794), .Y(
        n52522) );
  NAND2xp5_ASAP7_75t_SL U55704 ( .A(n69049), .B(n68831), .Y(n68843) );
  NAND2xp33_ASAP7_75t_SL U55705 ( .A(n66076), .B(n65914), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n22) );
  NAND2xp33_ASAP7_75t_SL U55706 ( .A(or1200_cpu_or1200_fpu_snan), .B(n74920), 
        .Y(n74775) );
  NAND2xp5_ASAP7_75t_SL U55707 ( .A(n61258), .B(n61257), .Y(n61260) );
  INVxp67_ASAP7_75t_SL U55708 ( .A(n62502), .Y(n62511) );
  AOI21xp33_ASAP7_75t_SL U55709 ( .A1(n74921), .A2(
        or1200_cpu_or1200_fpu_snan_conv), .B(n74773), .Y(n74774) );
  NAND2xp5_ASAP7_75t_SL U55710 ( .A(n76101), .B(n75937), .Y(n75914) );
  OAI21xp33_ASAP7_75t_SL U55711 ( .A1(n70149), .A2(n69562), .B(n69561), .Y(
        n52521) );
  INVxp67_ASAP7_75t_SL U55712 ( .A(n78080), .Y(n78079) );
  INVxp67_ASAP7_75t_SL U55713 ( .A(n66924), .Y(n66918) );
  NAND2xp33_ASAP7_75t_SL U55714 ( .A(n59687), .B(n78080), .Y(n559) );
  INVx1_ASAP7_75t_SL U55715 ( .A(n73452), .Y(n73467) );
  OAI21xp33_ASAP7_75t_SL U55716 ( .A1(n767), .A2(n77260), .B(n60025), .Y(
        n60030) );
  AOI21xp33_ASAP7_75t_SL U55717 ( .A1(n75015), .A2(n77864), .B(n68775), .Y(
        n68776) );
  INVxp33_ASAP7_75t_SL U55718 ( .A(n73440), .Y(n73283) );
  OAI21xp33_ASAP7_75t_SL U55719 ( .A1(n59629), .A2(n72726), .B(n72725), .Y(
        n1931) );
  AOI21xp33_ASAP7_75t_SL U55720 ( .A1(n74813), .A2(n74812), .B(n74811), .Y(
        n74824) );
  OAI21xp33_ASAP7_75t_SL U55721 ( .A1(n59629), .A2(n72856), .B(n72855), .Y(
        n1979) );
  AOI21xp33_ASAP7_75t_SL U55722 ( .A1(n75015), .A2(n77862), .B(n75004), .Y(
        n75005) );
  OAI21xp33_ASAP7_75t_SL U55723 ( .A1(n59627), .A2(n72726), .B(n72724), .Y(
        n1996) );
  INVxp33_ASAP7_75t_SL U55724 ( .A(n65289), .Y(n65374) );
  NAND2xp33_ASAP7_75t_SL U55725 ( .A(n59687), .B(n78121), .Y(n543) );
  NAND2xp33_ASAP7_75t_SL U55726 ( .A(n59687), .B(n78076), .Y(n561) );
  OAI21xp33_ASAP7_75t_SL U55727 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_16_), .A2(n59629), .B(
        n72712), .Y(n1678) );
  INVxp33_ASAP7_75t_SL U55728 ( .A(n78121), .Y(n78120) );
  INVxp33_ASAP7_75t_SL U55729 ( .A(n78105), .Y(n78104) );
  AOI22xp33_ASAP7_75t_SL U55730 ( .A1(n62290), .A2(n61627), .B1(n77125), .B2(
        n62130), .Y(n61665) );
  NAND2xp33_ASAP7_75t_SL U55731 ( .A(n73441), .B(n73295), .Y(n73296) );
  INVxp33_ASAP7_75t_SL U55732 ( .A(n75068), .Y(n75069) );
  INVxp33_ASAP7_75t_SL U55733 ( .A(n74808), .Y(n74919) );
  OAI21xp33_ASAP7_75t_SL U55734 ( .A1(n59629), .A2(n72691), .B(n72690), .Y(
        n1854) );
  INVxp67_ASAP7_75t_SL U55735 ( .A(n70755), .Y(n70756) );
  INVxp33_ASAP7_75t_SL U55736 ( .A(n66572), .Y(n66546) );
  INVxp67_ASAP7_75t_SL U55737 ( .A(n63156), .Y(n62655) );
  AOI22xp33_ASAP7_75t_SL U55738 ( .A1(or1200_cpu_spr_dat_rf[10]), .A2(n59686), 
        .B1(n77587), .B2(n74034), .Y(n61757) );
  INVxp33_ASAP7_75t_SL U55739 ( .A(n66364), .Y(n66365) );
  INVxp67_ASAP7_75t_SL U55740 ( .A(n66766), .Y(n66611) );
  NAND2xp33_ASAP7_75t_SL U55741 ( .A(n59526), .B(n70846), .Y(n70845) );
  NAND2xp33_ASAP7_75t_SL U55742 ( .A(or1200_cpu_spr_dat_rf[17]), .B(n59686), 
        .Y(n75370) );
  NAND2xp33_ASAP7_75t_SL U55743 ( .A(n59687), .B(n78105), .Y(n551) );
  INVxp33_ASAP7_75t_SL U55744 ( .A(n78072), .Y(n78071) );
  NAND2xp5_ASAP7_75t_SL U55745 ( .A(n73143), .B(n73142), .Y(n73415) );
  OAI21xp33_ASAP7_75t_SL U55746 ( .A1(n72967), .A2(n72953), .B(n72952), .Y(
        n72955) );
  INVxp67_ASAP7_75t_SL U55747 ( .A(n63114), .Y(n62679) );
  AOI22xp33_ASAP7_75t_SL U55748 ( .A1(n71263), .A2(n71000), .B1(n71396), .B2(
        n70851), .Y(n70827) );
  NAND2xp5_ASAP7_75t_SL U55749 ( .A(n72968), .B(n72967), .Y(n72970) );
  NAND2xp33_ASAP7_75t_SL U55750 ( .A(n59629), .B(n72713), .Y(n72712) );
  INVxp67_ASAP7_75t_SL U55751 ( .A(n64536), .Y(n64537) );
  INVxp67_ASAP7_75t_SL U55752 ( .A(n72961), .Y(n72969) );
  NAND2xp33_ASAP7_75t_SL U55753 ( .A(n59687), .B(n78072), .Y(n563) );
  AOI21xp33_ASAP7_75t_SL U55754 ( .A1(n65925), .A2(n65980), .B(n65924), .Y(
        n65926) );
  NAND2xp33_ASAP7_75t_SL U55755 ( .A(n71315), .B(n71067), .Y(n70899) );
  NAND2xp33_ASAP7_75t_SL U55756 ( .A(n77082), .B(n75549), .Y(n75550) );
  INVxp67_ASAP7_75t_SL U55757 ( .A(n76495), .Y(n76502) );
  OAI21xp33_ASAP7_75t_SL U55758 ( .A1(or1200_cpu_or1200_except_n266), .A2(
        n58547), .B(n76500), .Y(n76501) );
  OAI21xp33_ASAP7_75t_SL U55759 ( .A1(n69952), .A2(n69998), .B(n69901), .Y(
        n69906) );
  INVx1_ASAP7_75t_SL U55760 ( .A(n73417), .Y(n73426) );
  AOI22xp33_ASAP7_75t_SL U55761 ( .A1(or1200_cpu_spr_dat_rf[11]), .A2(n59686), 
        .B1(n77587), .B2(n75531), .Y(n61690) );
  OAI22xp33_ASAP7_75t_SL U55762 ( .A1(n1499), .A2(n74916), .B1(n59544), .B2(
        n74934), .Y(n74773) );
  NAND2xp5_ASAP7_75t_SL U55763 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_4_), .B(n70716), .Y(
        n70729) );
  AOI21xp33_ASAP7_75t_SL U55764 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[23]), 
        .B(n75562), .Y(n75563) );
  INVxp67_ASAP7_75t_SL U55765 ( .A(n75806), .Y(n75807) );
  OAI22xp33_ASAP7_75t_SL U55766 ( .A1(n1496), .A2(n74916), .B1(n57500), .B2(
        n74934), .Y(n74784) );
  NAND2xp33_ASAP7_75t_SL U55767 ( .A(n59317), .B(n58479), .Y(n59316) );
  NAND2xp33_ASAP7_75t_SL U55768 ( .A(n74947), .B(n57100), .Y(n63694) );
  O2A1O1Ixp33_ASAP7_75t_SL U55769 ( .A1(n68774), .A2(n76906), .B(n68773), .C(
        n68772), .Y(n68775) );
  OAI21xp33_ASAP7_75t_SL U55770 ( .A1(n74346), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_13_), .B(
        n74384), .Y(n2369) );
  OAI22xp33_ASAP7_75t_SL U55771 ( .A1(n1519), .A2(n74916), .B1(n59567), .B2(
        n74934), .Y(n74764) );
  INVxp67_ASAP7_75t_SL U55772 ( .A(n59118), .Y(n57935) );
  INVxp67_ASAP7_75t_SL U55773 ( .A(n73451), .Y(n73455) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U55774 ( .A1(n76970), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_22_), .B(n76969), 
        .C(n76968), .Y(n76972) );
  OAI21xp33_ASAP7_75t_SL U55775 ( .A1(n69929), .A2(n70062), .B(n69928), .Y(
        n69930) );
  INVxp67_ASAP7_75t_SL U55776 ( .A(n63170), .Y(n57417) );
  NAND2xp33_ASAP7_75t_SL U55777 ( .A(n63955), .B(n57100), .Y(n63943) );
  OAI22xp33_ASAP7_75t_SL U55778 ( .A1(n1112), .A2(n74916), .B1(n59580), .B2(
        n74934), .Y(n74829) );
  OAI22xp33_ASAP7_75t_SL U55779 ( .A1(n70060), .A2(n69953), .B1(n69952), .B2(
        n70063), .Y(n69954) );
  NAND2xp5_ASAP7_75t_SL U55780 ( .A(n73199), .B(n73198), .Y(n73202) );
  NAND2xp33_ASAP7_75t_SL U55781 ( .A(n58481), .B(n62813), .Y(n62816) );
  INVxp67_ASAP7_75t_SL U55782 ( .A(n66740), .Y(n59302) );
  OAI21xp33_ASAP7_75t_SL U55783 ( .A1(n70740), .A2(n70739), .B(n70754), .Y(
        n70741) );
  AOI22xp33_ASAP7_75t_SL U55784 ( .A1(or1200_cpu_spr_dat_rf[16]), .A2(n59686), 
        .B1(n77587), .B2(n76237), .Y(n62509) );
  NAND2xp33_ASAP7_75t_SL U55785 ( .A(n74956), .B(n60031), .Y(n60025) );
  INVx1_ASAP7_75t_SL U55786 ( .A(n73295), .Y(n73445) );
  AOI21xp5_ASAP7_75t_SL U55787 ( .A1(n73400), .A2(n73399), .B(n73394), .Y(
        n73395) );
  OAI21xp5_ASAP7_75t_SL U55788 ( .A1(n72882), .A2(n72808), .B(n72807), .Y(
        n72811) );
  NAND2xp5_ASAP7_75t_SL U55789 ( .A(n73131), .B(n73130), .Y(n73435) );
  INVxp67_ASAP7_75t_SL U55790 ( .A(n66472), .Y(n66465) );
  AOI21xp33_ASAP7_75t_SL U55791 ( .A1(n61983), .A2(n75890), .B(n75806), .Y(
        n61984) );
  NAND2xp33_ASAP7_75t_SL U55792 ( .A(n70149), .B(n69570), .Y(n69514) );
  NAND2xp5_ASAP7_75t_SL U55793 ( .A(n65786), .B(n65416), .Y(n65443) );
  AOI22xp33_ASAP7_75t_SL U55794 ( .A1(n71394), .A2(n53467), .B1(n71315), .B2(
        n70909), .Y(n70791) );
  AOI21xp5_ASAP7_75t_SL U55795 ( .A1(n58759), .A2(n57667), .B(n67946), .Y(
        n58760) );
  AOI22xp33_ASAP7_75t_SL U55796 ( .A1(or1200_cpu_spr_dat_rf[7]), .A2(n59686), 
        .B1(n77587), .B2(n76736), .Y(n76737) );
  AOI22xp33_ASAP7_75t_SL U55797 ( .A1(or1200_cpu_spr_dat_rf[9]), .A2(n59686), 
        .B1(n77587), .B2(n61336), .Y(n61337) );
  AOI22xp5_ASAP7_75t_SL U55798 ( .A1(n73314), .A2(n73313), .B1(n73316), .B2(
        n73315), .Y(n73448) );
  NAND2xp33_ASAP7_75t_SL U55799 ( .A(n59629), .B(n72706), .Y(n72707) );
  NOR2xp33_ASAP7_75t_SL U55800 ( .A(n1165), .B(n62397), .Y(n62401) );
  AOI22xp33_ASAP7_75t_SL U55801 ( .A1(or1200_cpu_spr_dat_rf[13]), .A2(n59686), 
        .B1(n77587), .B2(n77219), .Y(n61071) );
  NAND2xp5_ASAP7_75t_SL U55802 ( .A(n61981), .B(n61980), .Y(n75809) );
  NAND2xp33_ASAP7_75t_SL U55803 ( .A(n59687), .B(n78125), .Y(n541) );
  NAND2xp5_ASAP7_75t_SL U55804 ( .A(n72815), .B(n72798), .Y(n72800) );
  INVxp67_ASAP7_75t_SL U55805 ( .A(n73441), .Y(n73443) );
  NOR2xp33_ASAP7_75t_SL U55806 ( .A(n60264), .B(n60263), .Y(n75770) );
  INVxp67_ASAP7_75t_SL U55807 ( .A(n78125), .Y(n78124) );
  INVx1_ASAP7_75t_SL U55808 ( .A(n66334), .Y(n58634) );
  AOI22xp33_ASAP7_75t_SL U55809 ( .A1(n58416), .A2(n64758), .B1(n65218), .B2(
        n58554), .Y(n64767) );
  INVxp67_ASAP7_75t_SL U55810 ( .A(n76114), .Y(n76115) );
  NAND2xp33_ASAP7_75t_SL U55811 ( .A(n59628), .B(n72706), .Y(n72705) );
  NAND2xp33_ASAP7_75t_SL U55812 ( .A(n73417), .B(n73416), .Y(n73188) );
  INVxp67_ASAP7_75t_SL U55813 ( .A(n64461), .Y(n64383) );
  AOI21xp5_ASAP7_75t_SL U55814 ( .A1(n73021), .A2(n73005), .B(n73004), .Y(
        n73006) );
  INVxp67_ASAP7_75t_SL U55815 ( .A(n78144), .Y(n78143) );
  NAND2xp5_ASAP7_75t_SL U55816 ( .A(n64386), .B(n64385), .Y(n64442) );
  INVxp67_ASAP7_75t_SL U55817 ( .A(n75826), .Y(n64206) );
  INVxp67_ASAP7_75t_SL U55818 ( .A(n59060), .Y(n59059) );
  AOI21xp33_ASAP7_75t_SL U55819 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[24]), 
        .B(n64763), .Y(n64764) );
  NAND2xp33_ASAP7_75t_SL U55820 ( .A(n59687), .B(n78144), .Y(n533) );
  INVxp67_ASAP7_75t_SL U55821 ( .A(n73450), .Y(n73431) );
  AOI22xp33_ASAP7_75t_SL U55822 ( .A1(n70078), .A2(n69881), .B1(n69880), .B2(
        n69879), .Y(n69882) );
  NAND2xp5_ASAP7_75t_SL U55823 ( .A(n68815), .B(n68799), .Y(n76884) );
  INVxp67_ASAP7_75t_SL U55824 ( .A(n68109), .Y(n59035) );
  NAND2xp33_ASAP7_75t_SL U55825 ( .A(n3074), .B(n78067), .Y(n77468) );
  NAND2xp33_ASAP7_75t_SL U55826 ( .A(n59687), .B(n78133), .Y(n537) );
  AOI22xp33_ASAP7_75t_SL U55827 ( .A1(n66076), .A2(n66012), .B1(n66056), .B2(
        n66086), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n17) );
  INVxp67_ASAP7_75t_SL U55828 ( .A(n78129), .Y(n78128) );
  NAND2xp33_ASAP7_75t_SL U55829 ( .A(n59687), .B(n78129), .Y(n539) );
  OAI22xp33_ASAP7_75t_SL U55830 ( .A1(or1200_cpu_or1200_except_n522), .A2(
        n77032), .B1(or1200_cpu_or1200_except_n152), .B2(n57102), .Y(n75372)
         );
  NAND2xp33_ASAP7_75t_SL U55831 ( .A(n65402), .B(n65307), .Y(n1764) );
  NOR2x1_ASAP7_75t_SL U55832 ( .A(n57004), .B(n57879), .Y(n64568) );
  INVxp67_ASAP7_75t_SL U55833 ( .A(n62692), .Y(n62694) );
  NAND2xp33_ASAP7_75t_SL U55834 ( .A(n70149), .B(n69573), .Y(n69516) );
  NAND2xp33_ASAP7_75t_SL U55835 ( .A(or1200_cpu_spr_dat_rf[5]), .B(n59686), 
        .Y(n61610) );
  AOI21xp33_ASAP7_75t_SL U55836 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[20]), 
        .B(n64102), .Y(n64103) );
  NAND2xp33_ASAP7_75t_SL U55837 ( .A(n77270), .B(n57100), .Y(n77271) );
  INVx1_ASAP7_75t_SL U55838 ( .A(n73471), .Y(n73479) );
  INVxp67_ASAP7_75t_SL U55839 ( .A(n61956), .Y(n61959) );
  INVxp67_ASAP7_75t_SL U55840 ( .A(n73428), .Y(n73430) );
  NAND2xp5_ASAP7_75t_SL U55841 ( .A(n63976), .B(n63964), .Y(n63982) );
  NAND2xp5_ASAP7_75t_SL U55842 ( .A(n72734), .B(n72868), .Y(n72736) );
  AND2x2_ASAP7_75t_SL U55843 ( .A(n66624), .B(n66658), .Y(n58223) );
  INVxp33_ASAP7_75t_SL U55844 ( .A(n75549), .Y(n64203) );
  NAND2xp33_ASAP7_75t_SL U55845 ( .A(n73042), .B(n72819), .Y(n72746) );
  OAI21xp33_ASAP7_75t_SL U55846 ( .A1(n61572), .A2(n61571), .B(n57100), .Y(
        n76594) );
  INVxp67_ASAP7_75t_SL U55847 ( .A(n64572), .Y(n64575) );
  OAI21xp33_ASAP7_75t_SL U55848 ( .A1(n69804), .A2(n69803), .B(n69835), .Y(
        n69807) );
  INVxp67_ASAP7_75t_SL U55849 ( .A(n73418), .Y(n73423) );
  NAND2xp33_ASAP7_75t_SL U55850 ( .A(n73424), .B(n73416), .Y(n73275) );
  AOI21xp33_ASAP7_75t_SL U55851 ( .A1(n75015), .A2(n77869), .B(n65157), .Y(
        n65158) );
  O2A1O1Ixp33_ASAP7_75t_SL U55852 ( .A1(n59618), .A2(n58701), .B(n58700), .C(
        n62874), .Y(n62888) );
  INVxp67_ASAP7_75t_SL U55853 ( .A(n77789), .Y(n1238) );
  AND2x2_ASAP7_75t_SL U55854 ( .A(n57939), .B(n57820), .Y(n57938) );
  OAI21xp33_ASAP7_75t_SL U55855 ( .A1(n69944), .A2(n70026), .B(n69503), .Y(
        n69504) );
  NAND2xp5_ASAP7_75t_SL U55856 ( .A(n69880), .B(n69847), .Y(n69848) );
  NAND2xp33_ASAP7_75t_SL U55857 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .B(
        n72819), .Y(n72827) );
  OAI21xp33_ASAP7_75t_SL U55858 ( .A1(n69941), .A2(n69573), .B(n69471), .Y(
        n69472) );
  NAND2xp5_ASAP7_75t_SL U55859 ( .A(n61836), .B(n75360), .Y(n75568) );
  INVx1_ASAP7_75t_SL U55860 ( .A(n62654), .Y(n62643) );
  OAI21xp33_ASAP7_75t_SL U55861 ( .A1(n65479), .A2(n65478), .B(n65477), .Y(
        n65480) );
  INVxp67_ASAP7_75t_SL U55862 ( .A(n64428), .Y(n58186) );
  INVxp67_ASAP7_75t_SL U55863 ( .A(n76159), .Y(n76161) );
  OAI21xp5_ASAP7_75t_SL U55864 ( .A1(n57244), .A2(n59638), .B(n58154), .Y(
        n66851) );
  AOI22xp33_ASAP7_75t_SL U55865 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_1_), .A2(
        n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_2_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n3) );
  INVxp67_ASAP7_75t_SL U55866 ( .A(n66701), .Y(n66702) );
  OAI22xp33_ASAP7_75t_SL U55867 ( .A1(n71018), .A2(n71362), .B1(n71335), .B2(
        n70987), .Y(n70988) );
  AOI22xp33_ASAP7_75t_SL U55868 ( .A1(n71315), .A2(n71194), .B1(n71394), .B2(
        n71073), .Y(n71079) );
  NAND2xp33_ASAP7_75t_SL U55869 ( .A(n73367), .B(n73359), .Y(n73330) );
  INVxp33_ASAP7_75t_SL U55870 ( .A(n61342), .Y(n61343) );
  NAND2xp33_ASAP7_75t_SL U55871 ( .A(n59628), .B(n72793), .Y(n72794) );
  AOI22xp33_ASAP7_75t_SL U55872 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_2_), .A2(
        n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_3_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n5) );
  NOR2xp33_ASAP7_75t_SL U55873 ( .A(n58157), .B(n67355), .Y(n58156) );
  AOI21xp5_ASAP7_75t_SL U55874 ( .A1(n73367), .A2(n73369), .B(n73328), .Y(
        n73329) );
  AOI22xp33_ASAP7_75t_SL U55875 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_3_), .A2(
        n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_4_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n7) );
  AOI22xp33_ASAP7_75t_SL U55876 ( .A1(n71263), .A2(n71210), .B1(n71394), .B2(
        n71090), .Y(n71092) );
  AOI21xp33_ASAP7_75t_SL U55877 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[28]), 
        .B(n75825), .Y(n75827) );
  AOI21xp5_ASAP7_75t_SL U55878 ( .A1(n71337), .A2(n71338), .B(n71336), .Y(
        n71342) );
  AOI22xp33_ASAP7_75t_SL U55879 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_5_), .A2(
        n74493), .B1(n57103), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_4_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n9) );
  NAND2xp5_ASAP7_75t_SL U55880 ( .A(n67596), .B(n67595), .Y(n67597) );
  INVxp33_ASAP7_75t_SL U55881 ( .A(n62959), .Y(n59463) );
  OAI21xp33_ASAP7_75t_SL U55882 ( .A1(n74371), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_27_), .B(
        n74370), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n10) );
  NAND2xp5_ASAP7_75t_SL U55883 ( .A(n71396), .B(n71140), .Y(n71106) );
  AOI22xp33_ASAP7_75t_SL U55884 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_6_), .A2(
        n74493), .B1(n57103), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_5_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n11) );
  AOI21xp33_ASAP7_75t_SL U55885 ( .A1(n67327), .A2(n67267), .B(n67255), .Y(
        n67256) );
  OAI22xp5_ASAP7_75t_SL U55886 ( .A1(n72853), .A2(n73005), .B1(n72768), .B2(
        n72816), .Y(n72726) );
  AOI21xp33_ASAP7_75t_SL U55887 ( .A1(n62130), .A2(n75876), .B(n62129), .Y(
        n62131) );
  AOI22xp33_ASAP7_75t_SL U55888 ( .A1(n71396), .A2(n71000), .B1(n71394), .B2(
        n70954), .Y(n70956) );
  AOI22xp33_ASAP7_75t_SL U55889 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_6_), .A2(
        n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_7_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n13) );
  INVxp67_ASAP7_75t_SL U55890 ( .A(n73404), .Y(n73406) );
  AOI22xp33_ASAP7_75t_SL U55891 ( .A1(or1200_cpu_spr_dat_rf[8]), .A2(n59686), 
        .B1(n77587), .B2(n76648), .Y(n62327) );
  AOI22xp33_ASAP7_75t_SL U55892 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_7_), .A2(
        n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_8_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n15) );
  NAND2xp5_ASAP7_75t_SL U55893 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_45_), .B(n71366), 
        .Y(n71382) );
  AOI21xp33_ASAP7_75t_SL U55894 ( .A1(n53310), .A2(n75957), .B(n75949), .Y(
        n75950) );
  NAND2xp5_ASAP7_75t_SL U55895 ( .A(n75032), .B(n58631), .Y(n58630) );
  AOI22xp33_ASAP7_75t_SL U55896 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_8_), .A2(
        n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_9_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n17) );
  OAI22xp33_ASAP7_75t_SL U55897 ( .A1(n70987), .A2(n71362), .B1(n71335), .B2(
        n70932), .Y(n70933) );
  AOI22xp33_ASAP7_75t_SL U55898 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_9_), .A2(
        n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_10_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n19) );
  NAND2xp33_ASAP7_75t_SL U55899 ( .A(or1200_cpu_spr_dat_rf[27]), .B(n59686), 
        .Y(n73911) );
  AOI22xp33_ASAP7_75t_SL U55900 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_10_), 
        .A2(n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_11_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n21) );
  AOI22xp33_ASAP7_75t_SL U55901 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_11_), 
        .A2(n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_12_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n23) );
  NAND2xp33_ASAP7_75t_SL U55902 ( .A(n59526), .B(n71377), .Y(n71378) );
  OR2x2_ASAP7_75t_SL U55903 ( .A(n67276), .B(n59518), .Y(n67060) );
  AOI22xp33_ASAP7_75t_SL U55904 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_12_), 
        .A2(n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_13_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n25) );
  AOI22xp33_ASAP7_75t_SL U55905 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_13_), 
        .A2(n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_14_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n27) );
  BUFx3_ASAP7_75t_SL U55906 ( .A(n67868), .Y(n57494) );
  NAND2xp5_ASAP7_75t_SL U55907 ( .A(n57562), .B(n58982), .Y(n58981) );
  OAI21xp5_ASAP7_75t_SL U55908 ( .A1(n69746), .A2(n69745), .B(n69744), .Y(
        n70028) );
  NAND2xp33_ASAP7_75t_SL U55909 ( .A(n76574), .B(n58554), .Y(n61483) );
  BUFx6f_ASAP7_75t_SL U55910 ( .A(n67975), .Y(n57156) );
  NAND2xp33_ASAP7_75t_SL U55911 ( .A(n71394), .B(n71067), .Y(n71068) );
  AOI22xp33_ASAP7_75t_SL U55912 ( .A1(or1200_cpu_spr_dat_rf[6]), .A2(n59686), 
        .B1(n77587), .B2(n76622), .Y(n62246) );
  AOI22xp33_ASAP7_75t_SL U55913 ( .A1(n71263), .A2(n71393), .B1(n71396), .B2(
        n71248), .Y(n71222) );
  AOI22xp33_ASAP7_75t_SL U55914 ( .A1(n71263), .A2(n71395), .B1(n71394), .B2(
        n71248), .Y(n71249) );
  AOI22xp33_ASAP7_75t_SL U55915 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_1_), .A2(
        n74493), .B1(n57103), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_0_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n1) );
  AO21x1_ASAP7_75t_SL U55916 ( .A1(n58336), .A2(n67869), .B(n57596), .Y(n67896) );
  NAND2xp33_ASAP7_75t_SL U55917 ( .A(n59660), .B(n67564), .Y(n67565) );
  NAND2xp5_ASAP7_75t_SL U55918 ( .A(n57927), .B(n67344), .Y(n57926) );
  BUFx4f_ASAP7_75t_SL U55919 ( .A(n67713), .Y(n57277) );
  AOI22xp33_ASAP7_75t_SL U55920 ( .A1(n71263), .A2(n71356), .B1(n71396), .B2(
        n71210), .Y(n71211) );
  INVxp33_ASAP7_75t_SL U55921 ( .A(n67621), .Y(n67623) );
  INVxp33_ASAP7_75t_SL U55922 ( .A(n75214), .Y(n75216) );
  NAND2xp33_ASAP7_75t_SL U55923 ( .A(or1200_cpu_spr_dat_rf[30]), .B(n59686), 
        .Y(n75688) );
  AOI22xp33_ASAP7_75t_SL U55924 ( .A1(or1200_cpu_spr_dat_rf[2]), .A2(n59686), 
        .B1(n77587), .B2(n78253), .Y(n61258) );
  AOI22xp5_ASAP7_75t_SL U55925 ( .A1(n73117), .A2(n73116), .B1(n73390), .B2(
        n73389), .Y(n73388) );
  NAND2xp33_ASAP7_75t_SL U55926 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_33_), .B(n71166), 
        .Y(n71179) );
  NAND2xp33_ASAP7_75t_SL U55927 ( .A(n71315), .B(n71140), .Y(n71003) );
  INVxp67_ASAP7_75t_SL U55928 ( .A(n67404), .Y(n58008) );
  INVxp67_ASAP7_75t_SL U55929 ( .A(n67381), .Y(n58793) );
  AOI22xp33_ASAP7_75t_SL U55930 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_20_), 
        .A2(n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_21_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n41) );
  INVx1_ASAP7_75t_SL U55931 ( .A(n67719), .Y(n67721) );
  AOI21xp33_ASAP7_75t_SL U55932 ( .A1(n75877), .A2(n77125), .B(n62453), .Y(
        n62458) );
  INVxp67_ASAP7_75t_SL U55933 ( .A(n68381), .Y(n66731) );
  AOI22xp33_ASAP7_75t_SL U55934 ( .A1(or1200_cpu_spr_dat_rf[3]), .A2(n59686), 
        .B1(n77587), .B2(n61464), .Y(n61465) );
  AOI21xp33_ASAP7_75t_SL U55935 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[15]), 
        .B(n77047), .Y(n77050) );
  NAND2xp33_ASAP7_75t_SL U55936 ( .A(n70149), .B(n69793), .Y(n69794) );
  INVxp67_ASAP7_75t_SL U55937 ( .A(n67825), .Y(n57815) );
  AOI22xp33_ASAP7_75t_SL U55938 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_20_), 
        .A2(n74493), .B1(n57103), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_19_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n39) );
  O2A1O1Ixp33_ASAP7_75t_SL U55939 ( .A1(n61444), .A2(n61526), .B(n61443), .C(
        n75872), .Y(n61458) );
  INVxp67_ASAP7_75t_SL U55940 ( .A(n69570), .Y(n69571) );
  AOI22xp33_ASAP7_75t_SL U55941 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_22_), 
        .A2(n74493), .B1(n57103), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_21_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n43) );
  INVxp67_ASAP7_75t_SL U55942 ( .A(n66923), .Y(n57278) );
  AOI22xp33_ASAP7_75t_SL U55943 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_18_), 
        .A2(n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_19_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n37) );
  AOI22xp33_ASAP7_75t_SL U55944 ( .A1(ic_en), .A2(n77587), .B1(n59686), .B2(
        or1200_cpu_spr_dat_rf[4]), .Y(n61391) );
  AOI22xp33_ASAP7_75t_SL U55945 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_17_), 
        .A2(n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_18_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n35) );
  INVxp67_ASAP7_75t_SL U55946 ( .A(n70126), .Y(n70127) );
  INVxp33_ASAP7_75t_SL U55947 ( .A(n60031), .Y(n60036) );
  NAND2xp5_ASAP7_75t_SL U55948 ( .A(n60051), .B(n57100), .Y(n4132) );
  NOR2xp67_ASAP7_75t_SL U55949 ( .A(n57104), .B(n58162), .Y(n67631) );
  OAI22xp33_ASAP7_75t_SL U55950 ( .A1(n59190), .A2(n67458), .B1(n67460), .B2(
        n67459), .Y(n67461) );
  AOI22xp33_ASAP7_75t_SL U55951 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_16_), 
        .A2(n74493), .B1(n57103), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_15_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n31) );
  INVxp33_ASAP7_75t_SL U55952 ( .A(n2967), .Y(n76668) );
  INVxp67_ASAP7_75t_SL U55953 ( .A(n66921), .Y(n57610) );
  AOI22xp33_ASAP7_75t_SL U55954 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_15_), 
        .A2(n74493), .B1(n57103), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_14_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n29) );
  AOI22xp33_ASAP7_75t_SL U55955 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_16_), 
        .A2(n57103), .B1(n74493), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_17_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n33) );
  AOI21xp33_ASAP7_75t_SL U55956 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[21]), 
        .B(n62099), .Y(n62100) );
  NAND2xp5_ASAP7_75t_SL U55957 ( .A(n59499), .B(n76292), .Y(n61561) );
  INVxp67_ASAP7_75t_SL U55958 ( .A(n71248), .Y(n71139) );
  INVxp67_ASAP7_75t_SL U55959 ( .A(n73557), .Y(n73659) );
  INVxp67_ASAP7_75t_SL U55960 ( .A(n72866), .Y(n72798) );
  OAI21xp33_ASAP7_75t_SL U55961 ( .A1(n71413), .A2(n28213), .B(n70711), .Y(
        n70733) );
  AOI22xp33_ASAP7_75t_SL U55962 ( .A1(n66020), .A2(n66019), .B1(n66018), .B2(
        n66017), .Y(n66033) );
  INVxp67_ASAP7_75t_SL U55963 ( .A(n66955), .Y(n66956) );
  OAI21xp33_ASAP7_75t_SL U55964 ( .A1(n70149), .A2(n69947), .B(n69812), .Y(
        n52518) );
  INVxp33_ASAP7_75t_SL U55965 ( .A(n66061), .Y(n65723) );
  OAI21xp33_ASAP7_75t_SL U55966 ( .A1(n59627), .A2(n72709), .B(n72688), .Y(
        n1616) );
  OAI21xp33_ASAP7_75t_SL U55967 ( .A1(n59526), .A2(n70813), .B(n70780), .Y(
        n70781) );
  INVxp33_ASAP7_75t_SL U55968 ( .A(n66853), .Y(n66469) );
  NAND2xp5_ASAP7_75t_SL U55969 ( .A(n72734), .B(n72878), .Y(n72706) );
  AOI21xp33_ASAP7_75t_SL U55970 ( .A1(n73393), .A2(n73392), .B(n73391), .Y(
        n73394) );
  OAI21xp33_ASAP7_75t_SL U55971 ( .A1(n77616), .A2(n76796), .B(n61702), .Y(
        n61717) );
  BUFx2_ASAP7_75t_SL U55972 ( .A(n67883), .Y(n57366) );
  INVxp67_ASAP7_75t_SL U55973 ( .A(n73247), .Y(n73250) );
  NAND2xp33_ASAP7_75t_SL U55974 ( .A(n66079), .B(n66082), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n34) );
  INVxp67_ASAP7_75t_SL U55975 ( .A(n73248), .Y(n73249) );
  AOI21xp33_ASAP7_75t_SL U55976 ( .A1(n62508), .A2(n61335), .B(n61334), .Y(
        n61338) );
  NAND2xp5_ASAP7_75t_SL U55977 ( .A(n72815), .B(n72851), .Y(n72818) );
  INVxp33_ASAP7_75t_SL U55978 ( .A(n66064), .Y(n65848) );
  INVxp67_ASAP7_75t_SL U55979 ( .A(n67474), .Y(n66781) );
  OAI21xp33_ASAP7_75t_SL U55980 ( .A1(n70135), .A2(n69983), .B(n69779), .Y(
        n69876) );
  OAI21xp33_ASAP7_75t_SL U55981 ( .A1(n62463), .A2(n62462), .B(n62466), .Y(
        n61917) );
  AOI22xp33_ASAP7_75t_SL U55982 ( .A1(n66016), .A2(n66015), .B1(n66014), .B2(
        n66013), .Y(n66034) );
  OA21x2_ASAP7_75t_SL U55983 ( .A1(n74328), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_12_), 
        .B(n74340), .Y(n74329) );
  INVxp33_ASAP7_75t_SL U55984 ( .A(n62862), .Y(n62863) );
  AOI22xp33_ASAP7_75t_SL U55985 ( .A1(n66013), .A2(n66015), .B1(n66019), .B2(
        n65878), .Y(n65769) );
  OAI21xp33_ASAP7_75t_SL U55986 ( .A1(n63595), .A2(n75602), .B(n63594), .Y(
        n63596) );
  NAND2xp5_ASAP7_75t_SL U55987 ( .A(n57321), .B(n67535), .Y(n58975) );
  NOR2x1_ASAP7_75t_SL U55988 ( .A(n62514), .B(n77113), .Y(n75360) );
  AOI21xp33_ASAP7_75t_SL U55989 ( .A1(n68970), .A2(n57079), .B(n68946), .Y(
        n68947) );
  AOI21xp33_ASAP7_75t_SL U55990 ( .A1(n65947), .A2(n65980), .B(n65946), .Y(
        n65948) );
  INVxp67_ASAP7_75t_SL U55991 ( .A(n70079), .Y(n69879) );
  INVxp33_ASAP7_75t_SL U55992 ( .A(n62843), .Y(n62784) );
  INVxp67_ASAP7_75t_SL U55993 ( .A(n64479), .Y(n64359) );
  INVx1_ASAP7_75t_SL U55994 ( .A(n66374), .Y(n66326) );
  AOI21xp33_ASAP7_75t_SL U55995 ( .A1(n73037), .A2(n72974), .B(n72973), .Y(
        n72980) );
  OAI21xp33_ASAP7_75t_SL U55996 ( .A1(n77591), .A2(n76890), .B(n62223), .Y(
        n9272) );
  INVxp67_ASAP7_75t_SL U55997 ( .A(n73253), .Y(n73256) );
  AOI22xp33_ASAP7_75t_SL U55998 ( .A1(n66064), .A2(n66086), .B1(n66085), .B2(
        n65985), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n13) );
  NAND2xp33_ASAP7_75t_SL U55999 ( .A(n64114), .B(n61942), .Y(n61944) );
  INVxp67_ASAP7_75t_SL U56000 ( .A(n62956), .Y(n62957) );
  OAI21xp33_ASAP7_75t_SL U56001 ( .A1(n70880), .A2(n71149), .B(n70738), .Y(
        n70755) );
  OAI22xp33_ASAP7_75t_SL U56002 ( .A1(n72745), .A2(n72744), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .B2(n72797), .Y(n72819) );
  AOI22xp33_ASAP7_75t_SL U56003 ( .A1(n66045), .A2(n66086), .B1(n66085), .B2(
        n66044), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n51) );
  NAND2xp5_ASAP7_75t_SL U56004 ( .A(n62726), .B(n66786), .Y(n57703) );
  INVxp67_ASAP7_75t_SL U56005 ( .A(n67386), .Y(n67241) );
  INVx1_ASAP7_75t_SL U56006 ( .A(n57242), .Y(n64685) );
  AOI22xp33_ASAP7_75t_SL U56007 ( .A1(n66042), .A2(n66085), .B1(n66086), .B2(
        n66074), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n52) );
  AOI22xp33_ASAP7_75t_SL U56008 ( .A1(n66073), .A2(n66086), .B1(n66085), .B2(
        n66041), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n53) );
  AOI22xp33_ASAP7_75t_SL U56009 ( .A1(n66038), .A2(n66085), .B1(n66086), .B2(
        n66072), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n54) );
  INVx1_ASAP7_75t_SL U56010 ( .A(n58330), .Y(n70987) );
  NAND2xp33_ASAP7_75t_SL U56011 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_), .B(
        n72824), .Y(n72825) );
  O2A1O1Ixp33_ASAP7_75t_SL U56012 ( .A1(n71620), .A2(n71619), .B(n71618), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .Y(n71621) );
  INVxp33_ASAP7_75t_SL U56013 ( .A(n76787), .Y(n76788) );
  INVxp67_ASAP7_75t_SL U56014 ( .A(n66852), .Y(n66678) );
  NAND2xp5_ASAP7_75t_SL U56015 ( .A(n73457), .B(n73458), .Y(n73428) );
  AOI21xp33_ASAP7_75t_SL U56016 ( .A1(n70078), .A2(n69509), .B(n69470), .Y(
        n69471) );
  INVxp67_ASAP7_75t_SL U56017 ( .A(n71449), .Y(n71432) );
  NAND2xp5_ASAP7_75t_SL U56018 ( .A(n69576), .B(n69575), .Y(n17033) );
  INVxp67_ASAP7_75t_SL U56019 ( .A(n70016), .Y(n69847) );
  AOI22xp33_ASAP7_75t_SL U56020 ( .A1(n66071), .A2(n66086), .B1(n66085), .B2(
        n66037), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n55) );
  OAI21xp33_ASAP7_75t_SL U56021 ( .A1(n75315), .A2(n64121), .B(n64120), .Y(
        n64138) );
  NAND2xp33_ASAP7_75t_SL U56022 ( .A(n69899), .B(n69900), .Y(n69572) );
  OAI21xp33_ASAP7_75t_SL U56023 ( .A1(n72163), .A2(n71494), .B(n71423), .Y(
        n71442) );
  OAI22xp33_ASAP7_75t_SL U56024 ( .A1(n71284), .A2(n71283), .B1(n59526), .B2(
        n71333), .Y(n71287) );
  AOI22xp33_ASAP7_75t_SL U56025 ( .A1(n66087), .A2(n66086), .B1(n66085), .B2(
        n66084), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n56) );
  NOR2xp33_ASAP7_75t_SL U56026 ( .A(n71455), .B(n71619), .Y(n71622) );
  AOI22xp33_ASAP7_75t_SL U56027 ( .A1(n66061), .A2(n66086), .B1(n66085), .B2(
        n65984), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n15) );
  OAI22xp33_ASAP7_75t_SL U56028 ( .A1(n70064), .A2(n69998), .B1(n70062), .B2(
        n69997), .Y(n69999) );
  OAI21xp33_ASAP7_75t_SL U56029 ( .A1(n74043), .A2(n74042), .B(n78096), .Y(
        n78105) );
  AOI21xp33_ASAP7_75t_SL U56030 ( .A1(n73016), .A2(n73042), .B(n73021), .Y(
        n72785) );
  NAND2xp5_ASAP7_75t_SL U56031 ( .A(n74756), .B(n74934), .Y(n74916) );
  NAND2xp33_ASAP7_75t_SL U56032 ( .A(n69977), .B(n69983), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[3]) );
  NAND2xp5_ASAP7_75t_SL U56033 ( .A(n63864), .B(n63863), .Y(n58767) );
  INVxp67_ASAP7_75t_SL U56034 ( .A(n66857), .Y(n66859) );
  NAND2xp33_ASAP7_75t_SL U56035 ( .A(n72806), .B(n72878), .Y(n72807) );
  AOI22xp33_ASAP7_75t_SL U56036 ( .A1(n65959), .A2(n66019), .B1(n66015), .B2(
        n65958), .Y(n65960) );
  NAND2xp33_ASAP7_75t_SL U56037 ( .A(n66074), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n36) );
  NAND2xp33_ASAP7_75t_SL U56038 ( .A(n66073), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n37) );
  NAND2xp33_ASAP7_75t_SL U56039 ( .A(n66072), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n38) );
  OAI21xp33_ASAP7_75t_SL U56040 ( .A1(n61955), .A2(n61954), .B(n62498), .Y(
        n62081) );
  NAND2xp33_ASAP7_75t_SL U56041 ( .A(n66071), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n39) );
  INVxp67_ASAP7_75t_SL U56042 ( .A(n61359), .Y(n61360) );
  NAND2xp33_ASAP7_75t_SL U56043 ( .A(n59656), .B(n62958), .Y(n59278) );
  AOI21xp33_ASAP7_75t_SL U56044 ( .A1(n62508), .A2(n63764), .B(n61256), .Y(
        n61257) );
  NAND2xp33_ASAP7_75t_SL U56045 ( .A(n66087), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n40) );
  NAND2xp33_ASAP7_75t_SL U56046 ( .A(n66069), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n41) );
  OAI22xp33_ASAP7_75t_SL U56047 ( .A1(n71335), .A2(n71318), .B1(n71317), .B2(
        n71316), .Y(n71319) );
  NAND2xp5_ASAP7_75t_SL U56048 ( .A(n73178), .B(n73177), .Y(n73418) );
  NAND2xp33_ASAP7_75t_SL U56049 ( .A(n66068), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n42) );
  INVxp33_ASAP7_75t_SL U56050 ( .A(n69792), .Y(n69793) );
  OAI21xp33_ASAP7_75t_SL U56051 ( .A1(n59629), .A2(n72709), .B(n72708), .Y(
        n1623) );
  NAND2xp33_ASAP7_75t_SL U56052 ( .A(n69747), .B(n69792), .Y(n17034) );
  NAND2xp33_ASAP7_75t_SL U56053 ( .A(n66067), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n43) );
  NAND2xp33_ASAP7_75t_SL U56054 ( .A(n66066), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n44) );
  AOI21xp33_ASAP7_75t_SL U56055 ( .A1(n65980), .A2(n66043), .B(n65979), .Y(
        n65982) );
  OAI21xp5_ASAP7_75t_SL U56056 ( .A1(n1830), .A2(n77214), .B(n76215), .Y(
        or1200_cpu_to_sr[5]) );
  OAI21xp33_ASAP7_75t_SL U56057 ( .A1(n75602), .A2(n64853), .B(n64852), .Y(
        n64854) );
  INVxp67_ASAP7_75t_SL U56058 ( .A(n62942), .Y(n62815) );
  INVxp67_ASAP7_75t_SL U56059 ( .A(n67916), .Y(n57454) );
  OAI21xp33_ASAP7_75t_SL U56060 ( .A1(n73040), .A2(n73039), .B(n73038), .Y(
        n73044) );
  NAND2xp33_ASAP7_75t_SL U56061 ( .A(n66062), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n46) );
  NAND2xp5_ASAP7_75t_SL U56062 ( .A(n73246), .B(n73245), .Y(n73472) );
  AOI22xp33_ASAP7_75t_SL U56063 ( .A1(n59706), .A2(dwb_adr_o[21]), .B1(n57083), 
        .B2(sbbiu_adr_sb[21]), .Y(n77789) );
  AOI21xp5_ASAP7_75t_SL U56064 ( .A1(n75019), .A2(n75018), .B(n75017), .Y(
        n75023) );
  NAND2xp33_ASAP7_75t_SL U56065 ( .A(n63980), .B(n63981), .Y(n63964) );
  INVxp67_ASAP7_75t_SL U56066 ( .A(n62352), .Y(n62385) );
  NAND2xp33_ASAP7_75t_SL U56067 ( .A(n66061), .B(n66085), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n47) );
  OAI21xp33_ASAP7_75t_SL U56068 ( .A1(n73458), .A2(n73457), .B(n73459), .Y(
        n73214) );
  INVxp67_ASAP7_75t_SL U56069 ( .A(n75948), .Y(n75953) );
  OAI22xp33_ASAP7_75t_SL U56070 ( .A1(n59706), .A2(n77784), .B1(n57083), .B2(
        n1302), .Y(n1303) );
  AOI22xp33_ASAP7_75t_SL U56071 ( .A1(n72806), .A2(n73039), .B1(n72815), .B2(
        n73041), .Y(n72793) );
  AND2x2_ASAP7_75t_SL U56072 ( .A(n77965), .B(n77250), .Y(n77051) );
  INVxp33_ASAP7_75t_SL U56073 ( .A(n66037), .Y(n65925) );
  NAND2xp33_ASAP7_75t_SL U56074 ( .A(n69984), .B(n69900), .Y(n69901) );
  NAND2xp5_ASAP7_75t_SL U56075 ( .A(n71365), .B(n71364), .Y(n71337) );
  INVxp67_ASAP7_75t_SL U56076 ( .A(n64812), .Y(n64810) );
  XNOR2xp5_ASAP7_75t_SL U56077 ( .A(n73164), .B(n73165), .Y(n73450) );
  AOI22xp33_ASAP7_75t_SL U56078 ( .A1(n70033), .A2(n70085), .B1(n69977), .B2(
        n70082), .Y(n69978) );
  INVxp33_ASAP7_75t_SL U56079 ( .A(n75548), .Y(n75551) );
  AOI22xp33_ASAP7_75t_SL U56080 ( .A1(n70033), .A2(n70032), .B1(n70031), .B2(
        n70030), .Y(n70040) );
  AOI22xp5_ASAP7_75t_SL U56081 ( .A1(n70812), .A2(n70931), .B1(n71314), .B2(
        n58330), .Y(n70846) );
  OAI21xp33_ASAP7_75t_SL U56082 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[15]), .A2(
        n74502), .B(n73145), .Y(n73279) );
  OAI22xp33_ASAP7_75t_SL U56083 ( .A1(n71318), .A2(n71149), .B1(n71284), .B2(
        n71262), .Y(n71150) );
  NAND2xp5_ASAP7_75t_SL U56084 ( .A(n73040), .B(n72760), .Y(n72840) );
  AOI21xp33_ASAP7_75t_SL U56085 ( .A1(n68774), .A2(n59674), .B(n68771), .Y(
        n68772) );
  INVxp33_ASAP7_75t_SL U56086 ( .A(n62768), .Y(n62769) );
  NAND2xp33_ASAP7_75t_SL U56087 ( .A(n60421), .B(n60422), .Y(n60310) );
  OAI21xp33_ASAP7_75t_SL U56088 ( .A1(n62128), .A2(n75316), .B(n62127), .Y(
        n62129) );
  INVxp33_ASAP7_75t_SL U56089 ( .A(n59298), .Y(n64967) );
  INVxp67_ASAP7_75t_SL U56090 ( .A(n65882), .Y(n65883) );
  NAND2xp5_ASAP7_75t_SL U56091 ( .A(n67911), .B(n59600), .Y(n66610) );
  NAND2xp33_ASAP7_75t_SL U56092 ( .A(n73286), .B(n73285), .Y(n73154) );
  OAI21xp33_ASAP7_75t_SL U56093 ( .A1(n1717), .A2(n60570), .B(n60569), .Y(
        n60571) );
  OAI21xp33_ASAP7_75t_SL U56094 ( .A1(n75313), .A2(n62541), .B(n62540), .Y(
        n62542) );
  NAND2xp5_ASAP7_75t_SL U56095 ( .A(n68886), .B(n68848), .Y(n68863) );
  NAND2xp5_ASAP7_75t_SL U56096 ( .A(n73268), .B(n73267), .Y(n73451) );
  AOI22xp33_ASAP7_75t_SL U56097 ( .A1(n71315), .A2(n71176), .B1(n71394), .B2(
        n71175), .Y(n71177) );
  AOI22xp33_ASAP7_75t_SL U56098 ( .A1(n66017), .A2(n66015), .B1(n66019), .B2(
        n66013), .Y(n65913) );
  OAI21xp5_ASAP7_75t_SL U56099 ( .A1(n72718), .A2(n72813), .B(n72717), .Y(
        n73020) );
  INVxp67_ASAP7_75t_SL U56100 ( .A(n64196), .Y(n61975) );
  AOI22xp33_ASAP7_75t_SL U56101 ( .A1(n65994), .A2(n66085), .B1(n66086), .B2(
        n66068), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n10) );
  INVx3_ASAP7_75t_SL U56102 ( .A(n67901), .Y(n57158) );
  NAND2xp33_ASAP7_75t_SL U56103 ( .A(n71263), .B(n71090), .Y(n70901) );
  INVxp33_ASAP7_75t_SL U56104 ( .A(n70738), .Y(n70739) );
  NAND2xp33_ASAP7_75t_SL U56105 ( .A(n70118), .B(n69575), .Y(n69823) );
  INVxp67_ASAP7_75t_SL U56106 ( .A(n64498), .Y(n64072) );
  AOI22xp33_ASAP7_75t_SL U56107 ( .A1(n66069), .A2(n66086), .B1(n66085), .B2(
        n65992), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n9) );
  INVxp33_ASAP7_75t_SL U56108 ( .A(n70030), .Y(n69929) );
  NAND2xp5_ASAP7_75t_SL U56109 ( .A(n69902), .B(n69956), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[2]) );
  OAI21xp5_ASAP7_75t_SL U56110 ( .A1(n60684), .A2(n61224), .B(n60683), .Y(
        n60695) );
  INVxp67_ASAP7_75t_SL U56111 ( .A(n69972), .Y(n69980) );
  INVx5_ASAP7_75t_SL U56112 ( .A(n59516), .Y(n75895) );
  INVxp67_ASAP7_75t_SL U56113 ( .A(n71019), .Y(n71067) );
  INVxp67_ASAP7_75t_SL U56114 ( .A(n73203), .Y(n73206) );
  INVxp67_ASAP7_75t_SL U56115 ( .A(n65053), .Y(n64956) );
  NAND2xp33_ASAP7_75t_SL U56116 ( .A(n69977), .B(n69900), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[0]) );
  INVxp67_ASAP7_75t_SL U56117 ( .A(n66963), .Y(n66730) );
  INVxp67_ASAP7_75t_SL U56118 ( .A(n67453), .Y(n59097) );
  INVxp67_ASAP7_75t_SL U56119 ( .A(n75217), .Y(n61663) );
  AOI21xp33_ASAP7_75t_SL U56120 ( .A1(n66059), .A2(n66028), .B(n65957), .Y(
        n65961) );
  AO21x1_ASAP7_75t_SL U56121 ( .A1(n74343), .A2(n74342), .B(n74371), .Y(n74344) );
  AOI22xp33_ASAP7_75t_SL U56122 ( .A1(n69927), .A2(n70032), .B1(n69984), .B2(
        n69926), .Y(n69928) );
  NAND2xp5_ASAP7_75t_SL U56123 ( .A(n61622), .B(n61621), .Y(n62290) );
  OAI21xp33_ASAP7_75t_SL U56124 ( .A1(n71335), .A2(n71334), .B(n71367), .Y(
        n71336) );
  NAND2xp5_ASAP7_75t_SL U56125 ( .A(n69331), .B(n60422), .Y(n60312) );
  BUFx4f_ASAP7_75t_SL U56126 ( .A(n59668), .Y(n57398) );
  INVxp67_ASAP7_75t_SL U56127 ( .A(n67359), .Y(n58054) );
  OAI21xp33_ASAP7_75t_SL U56128 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n72986), .B(n72805), .Y(n72882) );
  AOI22xp33_ASAP7_75t_SL U56129 ( .A1(n65955), .A2(n66074), .B1(n65934), .B2(
        n66014), .Y(n65935) );
  AOI21xp33_ASAP7_75t_SL U56130 ( .A1(n72876), .A2(n73003), .B(n72875), .Y(
        n72881) );
  OAI21xp33_ASAP7_75t_SL U56131 ( .A1(n72879), .A2(n72878), .B(n73031), .Y(
        n72880) );
  INVxp67_ASAP7_75t_SL U56132 ( .A(n66755), .Y(n66757) );
  AOI21xp33_ASAP7_75t_SL U56133 ( .A1(n65980), .A2(n65989), .B(n65891), .Y(
        n65893) );
  INVxp67_ASAP7_75t_SL U56134 ( .A(n67249), .Y(n58216) );
  NAND2xp5_ASAP7_75t_SL U56135 ( .A(n66232), .B(n66233), .Y(n66238) );
  INVxp67_ASAP7_75t_SL U56136 ( .A(n69815), .Y(n69953) );
  OAI21xp33_ASAP7_75t_SL U56137 ( .A1(n75620), .A2(n76890), .B(n66228), .Y(
        n9252) );
  INVxp33_ASAP7_75t_SL U56138 ( .A(n77048), .Y(n76664) );
  INVxp67_ASAP7_75t_SL U56139 ( .A(n66802), .Y(n66801) );
  INVxp67_ASAP7_75t_SL U56140 ( .A(n73164), .Y(n73166) );
  OAI21xp5_ASAP7_75t_SL U56141 ( .A1(n71076), .A2(n71103), .B(n70826), .Y(
        n71000) );
  NAND2xp5_ASAP7_75t_SL U56142 ( .A(n74738), .B(n74734), .Y(n74072) );
  OAI21xp33_ASAP7_75t_SL U56143 ( .A1(n59529), .A2(n61973), .B(n64194), .Y(
        n61974) );
  INVxp33_ASAP7_75t_SL U56144 ( .A(n59048), .Y(n59046) );
  AOI21xp33_ASAP7_75t_SL U56145 ( .A1(n66042), .A2(n66028), .B(n65933), .Y(
        n65936) );
  INVxp67_ASAP7_75t_SL U56146 ( .A(n62664), .Y(n62833) );
  NAND2xp33_ASAP7_75t_SL U56147 ( .A(n66020), .B(n66018), .Y(n65910) );
  BUFx2_ASAP7_75t_SL U56148 ( .A(n68102), .Y(n57159) );
  NAND2xp5_ASAP7_75t_SL U56149 ( .A(n64183), .B(n64182), .Y(n9255) );
  INVxp67_ASAP7_75t_SL U56150 ( .A(n68022), .Y(n67966) );
  OAI22xp5_ASAP7_75t_SL U56151 ( .A1(n59467), .A2(n58934), .B1(n67963), .B2(
        n67408), .Y(n66783) );
  NAND2xp5_ASAP7_75t_SL U56152 ( .A(n69019), .B(n69018), .Y(n69021) );
  OAI21xp33_ASAP7_75t_SL U56153 ( .A1(n71467), .A2(n71494), .B(n71466), .Y(
        n71482) );
  INVxp67_ASAP7_75t_SL U56154 ( .A(n66431), .Y(n66432) );
  AOI22xp33_ASAP7_75t_SL U56155 ( .A1(n65986), .A2(n66085), .B1(n66086), .B2(
        n66062), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n14) );
  INVxp33_ASAP7_75t_SL U56156 ( .A(n71494), .Y(n71500) );
  NAND2xp5_ASAP7_75t_SL U56157 ( .A(n63783), .B(n63903), .Y(n63784) );
  OAI21xp33_ASAP7_75t_SL U56158 ( .A1(n75602), .A2(n64796), .B(n64795), .Y(
        n64797) );
  INVx4_ASAP7_75t_SL U56159 ( .A(n57104), .Y(n59650) );
  AOI22xp33_ASAP7_75t_SL U56160 ( .A1(n66066), .A2(n66086), .B1(n66085), .B2(
        n65988), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n12) );
  NOR2x1_ASAP7_75t_SL U56161 ( .A(n74339), .B(n74340), .Y(n74350) );
  AOI22xp33_ASAP7_75t_SL U56162 ( .A1(n71263), .A2(n71174), .B1(n71396), .B2(
        n71090), .Y(n71069) );
  AOI22xp33_ASAP7_75t_SL U56163 ( .A1(n70029), .A2(n69792), .B1(n70078), .B2(
        n70016), .Y(n69503) );
  NAND2xp5_ASAP7_75t_SL U56164 ( .A(n72734), .B(n73039), .Y(n72713) );
  OA21x2_ASAP7_75t_SL U56165 ( .A1(n57221), .A2(n67062), .B(n59601), .Y(n58005) );
  AOI22xp33_ASAP7_75t_SL U56166 ( .A1(n65955), .A2(n66072), .B1(n65909), .B2(
        n66014), .Y(n65911) );
  INVxp67_ASAP7_75t_SL U56167 ( .A(n65059), .Y(n64921) );
  NAND2xp33_ASAP7_75t_SL U56168 ( .A(n71315), .B(n71175), .Y(n71070) );
  INVxp33_ASAP7_75t_SL U56169 ( .A(n78148), .Y(n78147) );
  NAND2xp33_ASAP7_75t_SL U56170 ( .A(n66028), .B(n65986), .Y(n65767) );
  OAI21xp33_ASAP7_75t_SL U56171 ( .A1(n75701), .A2(n77078), .B(n61769), .Y(
        n61770) );
  NAND2xp33_ASAP7_75t_SL U56172 ( .A(n71245), .B(n71101), .Y(n71102) );
  INVxp67_ASAP7_75t_SL U56173 ( .A(n71592), .Y(n71593) );
  NAND2xp5_ASAP7_75t_SL U56174 ( .A(n64192), .B(n64191), .Y(n64194) );
  NAND2xp33_ASAP7_75t_SL U56175 ( .A(n71394), .B(n71104), .Y(n71105) );
  AOI21xp5_ASAP7_75t_SL U56176 ( .A1(n61791), .A2(n77088), .B(n61790), .Y(
        n61792) );
  AOI22xp33_ASAP7_75t_SL U56177 ( .A1(n71396), .A2(n71104), .B1(n71263), .B2(
        n71193), .Y(n71078) );
  INVxp67_ASAP7_75t_SL U56178 ( .A(n66083), .Y(n66084) );
  OAI21xp5_ASAP7_75t_SL U56179 ( .A1(n78351), .A2(n69564), .B(n69502), .Y(
        n70016) );
  NAND2xp5_ASAP7_75t_SL U56180 ( .A(n65542), .B(n65410), .Y(n65473) );
  OAI21xp33_ASAP7_75t_SL U56181 ( .A1(n70060), .A2(n69996), .B(n69995), .Y(
        n70000) );
  AOI22xp33_ASAP7_75t_SL U56182 ( .A1(n71354), .A2(n71087), .B1(n71245), .B2(
        n71086), .Y(n71088) );
  NAND2xp33_ASAP7_75t_SL U56183 ( .A(n59628), .B(n72761), .Y(n72763) );
  INVxp67_ASAP7_75t_SL U56184 ( .A(n68018), .Y(n57432) );
  NAND2xp33_ASAP7_75t_SL U56185 ( .A(n71174), .B(n71315), .Y(n71091) );
  AOI22xp33_ASAP7_75t_SL U56186 ( .A1(n71396), .A2(n70898), .B1(n71394), .B2(
        n70897), .Y(n70900) );
  INVxp33_ASAP7_75t_SL U56187 ( .A(n78134), .Y(n78137) );
  NAND2xp5_ASAP7_75t_SL U56188 ( .A(n62292), .B(n77124), .Y(n76787) );
  AOI22xp33_ASAP7_75t_SL U56189 ( .A1(n71394), .A2(n70779), .B1(n70897), .B2(
        n71315), .Y(n70780) );
  OAI21xp5_ASAP7_75t_SL U56190 ( .A1(n59631), .A2(n73304), .B(n73302), .Y(
        n73318) );
  OAI21xp5_ASAP7_75t_SL U56191 ( .A1(n70122), .A2(n70123), .B(n70121), .Y(
        n70138) );
  OAI21xp33_ASAP7_75t_SL U56192 ( .A1(n78348), .A2(n70054), .B(n69827), .Y(
        n70085) );
  AOI21xp33_ASAP7_75t_SL U56193 ( .A1(n69767), .A2(n69766), .B(n69765), .Y(
        n69768) );
  INVxp67_ASAP7_75t_SL U56194 ( .A(n66043), .Y(n66044) );
  INVxp67_ASAP7_75t_SL U56195 ( .A(n64408), .Y(n64039) );
  AOI21xp33_ASAP7_75t_SL U56196 ( .A1(n66050), .A2(n66049), .B(n66048), .Y(
        n66054) );
  INVxp67_ASAP7_75t_SL U56197 ( .A(n64634), .Y(n57276) );
  NAND2xp5_ASAP7_75t_SL U56198 ( .A(n72876), .B(n72747), .Y(n72824) );
  NAND2xp33_ASAP7_75t_SL U56199 ( .A(n59499), .B(n76291), .Y(n60984) );
  NAND2xp5_ASAP7_75t_SL U56200 ( .A(n71263), .B(n71104), .Y(n70916) );
  INVxp33_ASAP7_75t_SL U56201 ( .A(n76048), .Y(n76050) );
  OAI21xp33_ASAP7_75t_SL U56202 ( .A1(n65970), .A2(n65864), .B(n65863), .Y(
        n65868) );
  INVxp67_ASAP7_75t_SL U56203 ( .A(n76097), .Y(n76101) );
  INVxp67_ASAP7_75t_SL U56204 ( .A(n76047), .Y(n76053) );
  OAI21xp33_ASAP7_75t_SL U56205 ( .A1(n75316), .A2(n64136), .B(n64135), .Y(
        n64137) );
  OAI21xp33_ASAP7_75t_SL U56206 ( .A1(n72886), .A2(n73008), .B(n72739), .Y(
        n72745) );
  INVxp33_ASAP7_75t_SL U56207 ( .A(n64853), .Y(n61796) );
  INVx1_ASAP7_75t_SL U56208 ( .A(n58917), .Y(n58915) );
  NAND2xp33_ASAP7_75t_SL U56209 ( .A(n59687), .B(n78148), .Y(n531) );
  NOR2x1_ASAP7_75t_SL U56210 ( .A(n60230), .B(n76658), .Y(n73963) );
  AND2x2_ASAP7_75t_SL U56211 ( .A(n70118), .B(n69511), .Y(n69459) );
  OAI21xp33_ASAP7_75t_SL U56212 ( .A1(n59671), .A2(n68912), .B(n68893), .Y(
        n68896) );
  NAND2xp33_ASAP7_75t_SL U56213 ( .A(n70118), .B(n69881), .Y(n69825) );
  AOI21xp5_ASAP7_75t_SL U56214 ( .A1(n69509), .A2(n69880), .B(n69508), .Y(
        n69510) );
  INVxp67_ASAP7_75t_SL U56215 ( .A(n53468), .Y(n76104) );
  AOI22xp33_ASAP7_75t_SL U56216 ( .A1(n70078), .A2(n69811), .B1(n69810), .B2(
        n69809), .Y(n69947) );
  NAND2xp33_ASAP7_75t_SL U56217 ( .A(n70996), .B(n71101), .Y(n70826) );
  OAI21xp33_ASAP7_75t_SL U56218 ( .A1(n1489), .A2(n61755), .B(n61333), .Y(
        n61334) );
  AOI21xp33_ASAP7_75t_SL U56219 ( .A1(n70931), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .B(n70930), .Y(
        n70986) );
  NAND2xp33_ASAP7_75t_SL U56220 ( .A(n71315), .B(n71104), .Y(n70955) );
  NAND2xp33_ASAP7_75t_SL U56221 ( .A(n60172), .B(n60171), .Y(n60182) );
  AOI21xp33_ASAP7_75t_SL U56222 ( .A1(n61624), .A2(n61623), .B(n75882), .Y(
        n61627) );
  NAND2xp33_ASAP7_75t_SL U56223 ( .A(n71263), .B(n71160), .Y(n71004) );
  OAI21xp5_ASAP7_75t_SL U56224 ( .A1(n59631), .A2(n73312), .B(n73311), .Y(
        n73315) );
  NAND2xp5_ASAP7_75t_SL U56225 ( .A(n76001), .B(n76008), .Y(n75926) );
  AOI22xp33_ASAP7_75t_SL U56226 ( .A1(n69942), .A2(n70118), .B1(n69434), .B2(
        n69809), .Y(n69515) );
  AOI21xp33_ASAP7_75t_SL U56227 ( .A1(n70851), .A2(n71263), .B(n70719), .Y(
        n70727) );
  AOI22xp33_ASAP7_75t_SL U56228 ( .A1(n71396), .A2(n70852), .B1(n71394), .B2(
        n70851), .Y(n70853) );
  AOI22xp33_ASAP7_75t_SL U56229 ( .A1(n71465), .A2(n71422), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .B2(n71421), .Y(n71423) );
  AND2x2_ASAP7_75t_SL U56230 ( .A(n62627), .B(n62628), .Y(n57518) );
  OAI21xp33_ASAP7_75t_SL U56231 ( .A1(n59630), .A2(n73185), .B(n73183), .Y(
        n73276) );
  INVxp67_ASAP7_75t_SL U56232 ( .A(n59301), .Y(n59299) );
  OAI21xp33_ASAP7_75t_SL U56233 ( .A1(n78343), .A2(n69564), .B(n69493), .Y(
        n70017) );
  NAND3xp33_ASAP7_75t_SL U56234 ( .A(n59607), .B(n75641), .C(n57078), .Y(
        n67862) );
  AOI21xp33_ASAP7_75t_SL U56235 ( .A1(n68912), .A2(n57079), .B(n68893), .Y(
        n68894) );
  INVxp33_ASAP7_75t_SL U56236 ( .A(n73311), .Y(n73307) );
  NAND2xp33_ASAP7_75t_SL U56237 ( .A(n70135), .B(n69971), .Y(n69779) );
  OAI21xp33_ASAP7_75t_SL U56238 ( .A1(n70054), .A2(n78329), .B(n69739), .Y(
        n69926) );
  OAI21xp5_ASAP7_75t_SL U56239 ( .A1(n59631), .A2(n73333), .B(n73331), .Y(
        n73350) );
  OAI21xp33_ASAP7_75t_SL U56240 ( .A1(n78334), .A2(n70054), .B(n69738), .Y(
        n69932) );
  OAI21xp33_ASAP7_75t_SL U56241 ( .A1(n78336), .A2(n70054), .B(n69764), .Y(
        n69815) );
  NAND2xp33_ASAP7_75t_SL U56242 ( .A(n59687), .B(n78109), .Y(n549) );
  INVx2_ASAP7_75t_SL U56243 ( .A(n59475), .Y(n68104) );
  AOI21xp33_ASAP7_75t_SL U56244 ( .A1(n74621), .A2(n75876), .B(n74620), .Y(
        n74622) );
  NOR2x1_ASAP7_75t_SL U56245 ( .A(n59656), .B(n59245), .Y(n57879) );
  OAI21xp33_ASAP7_75t_SL U56246 ( .A1(n75143), .A2(n77142), .B(n75142), .Y(
        n75148) );
  INVxp33_ASAP7_75t_SL U56247 ( .A(n78109), .Y(n78108) );
  INVxp67_ASAP7_75t_SL U56248 ( .A(n76282), .Y(n76286) );
  OAI22xp33_ASAP7_75t_SL U56249 ( .A1(n70059), .A2(n70062), .B1(n70064), .B2(
        n70061), .Y(n69955) );
  INVxp67_ASAP7_75t_SL U56250 ( .A(n64406), .Y(n64512) );
  NAND2xp33_ASAP7_75t_SL U56251 ( .A(n76283), .B(n76282), .Y(n76284) );
  INVxp67_ASAP7_75t_SL U56252 ( .A(n73234), .Y(n73230) );
  INVxp67_ASAP7_75t_SL U56253 ( .A(n66827), .Y(n66828) );
  OAI22xp33_ASAP7_75t_SL U56254 ( .A1(n59706), .A2(n77781), .B1(n57083), .B2(
        n1317), .Y(n1318) );
  INVx2_ASAP7_75t_SL U56255 ( .A(n58202), .Y(n57162) );
  INVxp67_ASAP7_75t_SL U56256 ( .A(n64914), .Y(n64409) );
  NAND2xp33_ASAP7_75t_SL U56257 ( .A(n70149), .B(n69940), .Y(n69812) );
  INVxp67_ASAP7_75t_SL U56258 ( .A(n71393), .Y(n71363) );
  OAI21xp33_ASAP7_75t_SL U56259 ( .A1(n59630), .A2(n73150), .B(n73146), .Y(
        n73285) );
  OAI22xp33_ASAP7_75t_SL U56260 ( .A1(n65956), .A2(n65998), .B1(n65962), .B2(
        n65996), .Y(n65933) );
  NAND2xp33_ASAP7_75t_SL U56261 ( .A(n62292), .B(n75877), .Y(n61460) );
  OAI22xp33_ASAP7_75t_SL U56262 ( .A1(n69904), .A2(n70060), .B1(n70064), .B2(
        n69997), .Y(n69905) );
  OAI21xp5_ASAP7_75t_SL U56263 ( .A1(n59630), .A2(n73221), .B(n73220), .Y(
        n73225) );
  NAND2xp33_ASAP7_75t_SL U56264 ( .A(n71396), .B(n71376), .Y(n71379) );
  AOI22xp33_ASAP7_75t_SL U56265 ( .A1(n71396), .A2(n71395), .B1(n71394), .B2(
        n71393), .Y(n71402) );
  OAI21xp33_ASAP7_75t_SL U56266 ( .A1(n64176), .A2(n76897), .B(n64173), .Y(
        n64174) );
  NAND2xp33_ASAP7_75t_SL U56267 ( .A(n70118), .B(n69811), .Y(n69451) );
  INVxp67_ASAP7_75t_SL U56268 ( .A(n73259), .Y(n73260) );
  OAI22xp33_ASAP7_75t_SL U56269 ( .A1(n66020), .A2(n65996), .B1(n66013), .B2(
        n66001), .Y(n65882) );
  INVx1_ASAP7_75t_SL U56270 ( .A(n61624), .Y(n61621) );
  INVxp67_ASAP7_75t_SL U56271 ( .A(n73151), .Y(n73145) );
  INVxp33_ASAP7_75t_SL U56272 ( .A(n69996), .Y(n69907) );
  OAI22xp33_ASAP7_75t_SL U56273 ( .A1(n66080), .A2(n66029), .B1(n65997), .B2(
        n65996), .Y(n66005) );
  OAI22xp33_ASAP7_75t_SL U56274 ( .A1(or1200_cpu_sr_15_), .A2(n77142), .B1(
        or1200_cpu_esr[15]), .B2(n58547), .Y(n2688) );
  NAND2xp33_ASAP7_75t_SL U56275 ( .A(n66079), .B(n66030), .Y(n66031) );
  INVxp67_ASAP7_75t_SL U56276 ( .A(n66001), .Y(n66018) );
  INVxp67_ASAP7_75t_SL U56277 ( .A(n66078), .Y(n66014) );
  INVxp67_ASAP7_75t_SL U56278 ( .A(n64936), .Y(n64615) );
  AOI22xp33_ASAP7_75t_SL U56279 ( .A1(n75015), .A2(n77859), .B1(n57079), .B2(
        n75014), .Y(n75025) );
  OAI21xp33_ASAP7_75t_SL U56280 ( .A1(n70060), .A2(n70059), .B(n70058), .Y(
        n70066) );
  AOI22xp33_ASAP7_75t_SL U56281 ( .A1(n72990), .A2(n72846), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .B2(n72814), .Y(n73016) );
  OAI22xp33_ASAP7_75t_SL U56282 ( .A1(n65909), .A2(n65998), .B1(n65878), .B2(
        n66078), .Y(n65879) );
  AND2x2_ASAP7_75t_SL U56283 ( .A(n67357), .B(n57428), .Y(n57355) );
  NAND2xp33_ASAP7_75t_SL U56284 ( .A(n73037), .B(n72835), .Y(n72836) );
  INVxp33_ASAP7_75t_SL U56285 ( .A(n66068), .Y(n65881) );
  AOI21xp33_ASAP7_75t_SL U56286 ( .A1(n75877), .A2(n75876), .B(n75875), .Y(
        n75878) );
  INVxp67_ASAP7_75t_SL U56287 ( .A(n72952), .Y(n72954) );
  AOI22xp33_ASAP7_75t_SL U56288 ( .A1(n71332), .A2(n71331), .B1(n58315), .B2(
        n71330), .Y(n71364) );
  AOI21xp33_ASAP7_75t_SL U56289 ( .A1(n62508), .A2(n76236), .B(n62507), .Y(
        n62510) );
  OAI21xp33_ASAP7_75t_SL U56290 ( .A1(n78427), .A2(n69925), .B(n69875), .Y(
        n69972) );
  INVxp33_ASAP7_75t_SL U56291 ( .A(n76484), .Y(n76426) );
  INVxp33_ASAP7_75t_SL U56292 ( .A(n66041), .Y(n65947) );
  NAND2xp5_ASAP7_75t_SL U56293 ( .A(n61853), .B(n77124), .Y(n62134) );
  NAND2xp33_ASAP7_75t_SL U56294 ( .A(n65980), .B(n66083), .Y(n65905) );
  AOI22xp33_ASAP7_75t_SL U56295 ( .A1(n59499), .A2(n76290), .B1(n77125), .B2(
        n61238), .Y(n61239) );
  NAND2xp33_ASAP7_75t_SL U56296 ( .A(n66028), .B(n66038), .Y(n65912) );
  NAND2xp5_ASAP7_75t_SL U56297 ( .A(n70227), .B(n70242), .Y(n3166) );
  NAND2xp5_ASAP7_75t_SL U56298 ( .A(n70243), .B(n70242), .Y(n3165) );
  OAI21xp33_ASAP7_75t_SL U56299 ( .A1(n70236), .A2(n70228), .B(n70242), .Y(
        n3168) );
  OAI21xp33_ASAP7_75t_SL U56300 ( .A1(n72874), .A2(n72846), .B(n73040), .Y(
        n72850) );
  INVx1_ASAP7_75t_SL U56301 ( .A(n73204), .Y(n73205) );
  INVx1_ASAP7_75t_SL U56302 ( .A(n76493), .Y(n76477) );
  OAI21xp33_ASAP7_75t_SL U56303 ( .A1(n72848), .A2(n72847), .B(n72962), .Y(
        n72849) );
  INVxp33_ASAP7_75t_SL U56304 ( .A(n66036), .Y(n65927) );
  NAND2xp5_ASAP7_75t_SL U56305 ( .A(n65919), .B(n65918), .Y(n66037) );
  INVxp33_ASAP7_75t_SL U56306 ( .A(n64796), .Y(n62388) );
  NAND2xp5_ASAP7_75t_SL U56307 ( .A(n72638), .B(n72637), .Y(n72639) );
  AOI21xp33_ASAP7_75t_SL U56308 ( .A1(n57079), .A2(n63900), .B(n63899), .Y(
        n63901) );
  OAI21xp33_ASAP7_75t_SL U56309 ( .A1(n74324), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_11_), .B(
        n74337), .Y(n2405) );
  AOI22xp33_ASAP7_75t_SL U56310 ( .A1(n72792), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .B1(n72990), .B2(n72835), .Y(n73041) );
  OAI21xp5_ASAP7_75t_SL U56311 ( .A1(n78333), .A2(n69564), .B(n69461), .Y(
        n69505) );
  OAI21xp5_ASAP7_75t_SL U56312 ( .A1(n68767), .A2(n68766), .B(n68790), .Y(
        n68774) );
  NOR2x1_ASAP7_75t_SL U56313 ( .A(n57110), .B(n58990), .Y(n63082) );
  INVx1_ASAP7_75t_SL U56314 ( .A(n64185), .Y(n75553) );
  OAI21xp33_ASAP7_75t_SL U56315 ( .A1(n72874), .A2(n72989), .B(n73040), .Y(
        n72875) );
  OAI21xp33_ASAP7_75t_SL U56316 ( .A1(n1533), .A2(n61755), .B(n61479), .Y(
        n61482) );
  INVx1_ASAP7_75t_SL U56317 ( .A(n73950), .Y(n73951) );
  INVx1_ASAP7_75t_SL U56318 ( .A(n64248), .Y(n61374) );
  INVxp33_ASAP7_75t_SL U56319 ( .A(n64192), .Y(n64199) );
  INVxp67_ASAP7_75t_SL U56320 ( .A(n64757), .Y(n64190) );
  OAI21xp33_ASAP7_75t_SL U56321 ( .A1(n72716), .A2(n72715), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), .Y(
        n72717) );
  OAI21xp33_ASAP7_75t_SL U56322 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n72792), .B(n72759), .Y(n72760) );
  OAI21xp33_ASAP7_75t_SL U56323 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[1]), .A2(
        n70236), .B(n70242), .Y(n3167) );
  OAI21xp5_ASAP7_75t_SL U56324 ( .A1(n78335), .A2(n69564), .B(n69487), .Y(
        n69743) );
  INVxp33_ASAP7_75t_SL U56325 ( .A(n73548), .Y(n73547) );
  INVxp67_ASAP7_75t_SL U56326 ( .A(n67971), .Y(n64933) );
  NAND2xp5_ASAP7_75t_SL U56327 ( .A(n62091), .B(n62090), .Y(n62093) );
  AOI21xp33_ASAP7_75t_SL U56328 ( .A1(n71470), .A2(n71427), .B(n71426), .Y(
        n71449) );
  AOI22xp33_ASAP7_75t_SL U56329 ( .A1(n71396), .A2(n71243), .B1(n71315), .B2(
        n71393), .Y(n71250) );
  INVx1_ASAP7_75t_SL U56330 ( .A(n65998), .Y(n66019) );
  INVxp67_ASAP7_75t_SL U56331 ( .A(n66684), .Y(n59175) );
  INVx1_ASAP7_75t_SL U56332 ( .A(n65996), .Y(n66015) );
  OAI21xp5_ASAP7_75t_SL U56333 ( .A1(n71716), .A2(n71680), .B(n71654), .Y(
        n71678) );
  NAND2xp5_ASAP7_75t_SL U56334 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), .B(
        n72730), .Y(n72731) );
  NAND2xp33_ASAP7_75t_SL U56335 ( .A(n71396), .B(n71194), .Y(n71163) );
  AOI22xp33_ASAP7_75t_SL U56336 ( .A1(n71263), .A2(n71339), .B1(n71315), .B2(
        n71243), .Y(n71164) );
  NAND2xp33_ASAP7_75t_SL U56337 ( .A(n71394), .B(n71160), .Y(n71165) );
  NAND2xp5_ASAP7_75t_SL U56338 ( .A(n61830), .B(n61763), .Y(n61721) );
  AOI21xp33_ASAP7_75t_SL U56339 ( .A1(n75747), .A2(n75876), .B(n75746), .Y(
        n75748) );
  INVx1_ASAP7_75t_SL U56340 ( .A(n67459), .Y(n67316) );
  AOI21xp5_ASAP7_75t_SL U56341 ( .A1(n66036), .A2(n66040), .B(n65704), .Y(
        n66061) );
  OAI21xp33_ASAP7_75t_SL U56342 ( .A1(n78350), .A2(n70054), .B(n69846), .Y(
        n70032) );
  OAI21xp5_ASAP7_75t_SL U56343 ( .A1(n71314), .A2(n71174), .B(n71173), .Y(
        n71212) );
  AOI21xp33_ASAP7_75t_SL U56344 ( .A1(n66231), .A2(n75030), .B(n1133), .Y(
        n66230) );
  OAI21xp33_ASAP7_75t_SL U56345 ( .A1(n65827), .A2(n66039), .B(n65826), .Y(
        n66064) );
  INVx1_ASAP7_75t_SL U56346 ( .A(n71339), .Y(n71334) );
  OAI21xp5_ASAP7_75t_SL U56347 ( .A1(n59631), .A2(n73338), .B(n73337), .Y(
        n73346) );
  OAI22xp33_ASAP7_75t_SL U56348 ( .A1(n69944), .A2(n69943), .B1(n69942), .B2(
        n70118), .Y(n69945) );
  OAI21xp5_ASAP7_75t_SL U56349 ( .A1(n78331), .A2(n70054), .B(n69733), .Y(
        n69983) );
  INVx1_ASAP7_75t_SL U56350 ( .A(n74317), .Y(n74323) );
  INVxp33_ASAP7_75t_SL U56351 ( .A(n73114), .Y(n73110) );
  INVxp67_ASAP7_75t_SL U56352 ( .A(n72974), .Y(n72864) );
  INVx1_ASAP7_75t_SL U56353 ( .A(n58425), .Y(n58141) );
  INVx1_ASAP7_75t_SL U56354 ( .A(n67410), .Y(n58934) );
  INVx1_ASAP7_75t_SL U56355 ( .A(n73254), .Y(n73255) );
  OAI22xp33_ASAP7_75t_SL U56356 ( .A1(n70064), .A2(n70063), .B1(n70062), .B2(
        n70061), .Y(n70065) );
  NAND2xp5_ASAP7_75t_SL U56357 ( .A(n73007), .B(n72989), .Y(n72776) );
  AOI21xp33_ASAP7_75t_SL U56358 ( .A1(n73037), .A2(n73036), .B(n73035), .Y(
        n73038) );
  INVxp67_ASAP7_75t_SL U56359 ( .A(n67334), .Y(n67333) );
  NAND2xp5_ASAP7_75t_SL U56360 ( .A(n75400), .B(n75399), .Y(n9254) );
  OAI21xp33_ASAP7_75t_SL U56361 ( .A1(n70114), .A2(n69499), .B(n69477), .Y(
        n69485) );
  INVxp33_ASAP7_75t_SL U56362 ( .A(n73339), .Y(n73344) );
  OAI21xp33_ASAP7_75t_SL U56363 ( .A1(n1117), .A2(n77142), .B(n75525), .Y(
        n75526) );
  NAND2xp33_ASAP7_75t_SL U56364 ( .A(n59468), .B(n62767), .Y(n62770) );
  AOI21xp33_ASAP7_75t_SL U56365 ( .A1(n62508), .A2(n73959), .B(n61756), .Y(
        n61758) );
  OAI21xp33_ASAP7_75t_SL U56366 ( .A1(n70118), .A2(n69943), .B(n69444), .Y(
        n69454) );
  INVxp33_ASAP7_75t_SL U56367 ( .A(n67071), .Y(n67072) );
  AOI21xp33_ASAP7_75t_SL U56368 ( .A1(n61953), .A2(n61952), .B(n61951), .Y(
        n62498) );
  INVxp67_ASAP7_75t_SL U56369 ( .A(n62921), .Y(n62922) );
  NOR2x1_ASAP7_75t_SL U56370 ( .A(n59493), .B(n60833), .Y(n77250) );
  OAI22xp33_ASAP7_75t_SL U56371 ( .A1(n66081), .A2(n66029), .B1(n65956), .B2(
        n66078), .Y(n65957) );
  OAI22xp33_ASAP7_75t_SL U56372 ( .A1(n70929), .A2(n71012), .B1(n70928), .B2(
        n71076), .Y(n70930) );
  NAND2xp33_ASAP7_75t_SL U56373 ( .A(n76129), .B(n58600), .Y(n76130) );
  AOI21xp33_ASAP7_75t_SL U56374 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[9]), .B(n69796), 
        .Y(n69797) );
  NOR2x1p5_ASAP7_75t_SL U56375 ( .A(n67851), .B(n59640), .Y(n58917) );
  INVx2_ASAP7_75t_SL U56376 ( .A(n75894), .Y(n75035) );
  NAND2xp33_ASAP7_75t_SL U56377 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[22]), .B(
        n59631), .Y(n73337) );
  INVx4_ASAP7_75t_SL U56378 ( .A(n59669), .Y(n59667) );
  NAND2xp33_ASAP7_75t_SL U56379 ( .A(n71799), .B(n71703), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n122) );
  INVxp67_ASAP7_75t_SL U56380 ( .A(n66070), .Y(n66087) );
  INVxp33_ASAP7_75t_SL U56381 ( .A(n74380), .Y(n74360) );
  NAND2xp5_ASAP7_75t_SL U56382 ( .A(n68936), .B(n68937), .Y(n68912) );
  OR2x2_ASAP7_75t_SL U56383 ( .A(n74065), .B(n74276), .Y(n74492) );
  OAI21xp5_ASAP7_75t_SL U56384 ( .A1(n70106), .A2(n70105), .B(n70120), .Y(
        n70108) );
  OAI21xp33_ASAP7_75t_SL U56385 ( .A1(n70788), .A2(n70737), .B(n70736), .Y(
        n70740) );
  OAI21xp33_ASAP7_75t_SL U56386 ( .A1(n73169), .A2(n58284), .B(n73168), .Y(
        n73177) );
  NAND2xp33_ASAP7_75t_SL U56387 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[1]), .B(
        n59631), .Y(n73226) );
  INVx1_ASAP7_75t_SL U56388 ( .A(n65991), .Y(n66069) );
  OAI21xp33_ASAP7_75t_SL U56389 ( .A1(n62422), .A2(n75317), .B(n61368), .Y(
        n61371) );
  INVxp33_ASAP7_75t_SL U56390 ( .A(n74247), .Y(n74248) );
  INVxp33_ASAP7_75t_SL U56391 ( .A(n74278), .Y(n74242) );
  OAI21xp33_ASAP7_75t_SL U56392 ( .A1(or1200_cpu_or1200_except_n536), .A2(
        n76724), .B(n64762), .Y(n64763) );
  NAND2xp33_ASAP7_75t_SL U56393 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[23]), .B(
        n59631), .Y(n73331) );
  OAI22xp33_ASAP7_75t_SL U56394 ( .A1(n73308), .A2(n59630), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[18]), .B2(
        n74502), .Y(n73309) );
  NAND2xp33_ASAP7_75t_SL U56395 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[13]), .B(
        n59630), .Y(n73183) );
  OAI21xp33_ASAP7_75t_SL U56396 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_1_), .A2(
        n71711), .B(n71799), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n121) );
  AOI21xp33_ASAP7_75t_SL U56397 ( .A1(n65152), .A2(n59672), .B(n65151), .Y(
        n65155) );
  INVxp67_ASAP7_75t_SL U56398 ( .A(n72729), .Y(n72730) );
  AOI21xp33_ASAP7_75t_SL U56399 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[3]), .A2(n70038), .B(n69732), .Y(n69733) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56400 ( .A1(n65710), .A2(n65709), .B(n65974), 
        .C(n65708), .Y(n65721) );
  OAI21xp33_ASAP7_75t_SL U56401 ( .A1(n71281), .A2(n71247), .B(n71246), .Y(
        n71395) );
  AOI21xp5_ASAP7_75t_SL U56402 ( .A1(n65149), .A2(n65161), .B(n65164), .Y(
        n65156) );
  INVx2_ASAP7_75t_SL U56403 ( .A(n67268), .Y(n57166) );
  NAND2xp33_ASAP7_75t_SL U56404 ( .A(n59687), .B(n77970), .Y(n3921) );
  NAND2x1p5_ASAP7_75t_SL U56405 ( .A(n58950), .B(n58949), .Y(n59663) );
  NOR2xp33_ASAP7_75t_SL U56406 ( .A(n61835), .B(n62348), .Y(n77114) );
  INVxp67_ASAP7_75t_SL U56407 ( .A(n70038), .Y(n69560) );
  NAND2xp33_ASAP7_75t_SL U56408 ( .A(n71799), .B(n71708), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n124) );
  NAND2xp33_ASAP7_75t_SL U56409 ( .A(n76911), .B(n57080), .Y(n76915) );
  NAND2xp33_ASAP7_75t_SL U56410 ( .A(n71229), .B(n71228), .Y(n70984) );
  NAND2xp5_ASAP7_75t_SL U56411 ( .A(n62229), .B(n62228), .Y(n62233) );
  BUFx3_ASAP7_75t_SL U56412 ( .A(n59484), .Y(n57425) );
  OAI22xp33_ASAP7_75t_SL U56413 ( .A1(n73111), .A2(n59630), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[24]), .B2(
        n74502), .Y(n73112) );
  INVxp33_ASAP7_75t_SL U56414 ( .A(n65968), .Y(n65720) );
  INVxp67_ASAP7_75t_SL U56415 ( .A(n70113), .Y(n70111) );
  NAND2xp5_ASAP7_75t_SL U56416 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[1]), .B(n70038), 
        .Y(n69739) );
  NAND2xp5_ASAP7_75t_SL U56417 ( .A(n76747), .B(n76746), .Y(n76750) );
  NAND2xp33_ASAP7_75t_SL U56418 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_14_), .B(n70023), .Y(
        n69473) );
  INVxp33_ASAP7_75t_SL U56419 ( .A(n71481), .Y(n71421) );
  OAI22xp33_ASAP7_75t_SL U56420 ( .A1(n59540), .A2(n61733), .B1(n74608), .B2(
        n61783), .Y(n61734) );
  NAND2xp5_ASAP7_75t_SL U56421 ( .A(n72743), .B(n72742), .Y(n72797) );
  NAND2xp5_ASAP7_75t_SL U56422 ( .A(n63522), .B(n63441), .Y(n63454) );
  NAND2xp5_ASAP7_75t_SL U56423 ( .A(n70999), .B(n70998), .Y(n71160) );
  NAND2xp5_ASAP7_75t_SL U56424 ( .A(n76786), .B(n76785), .Y(n76789) );
  INVx3_ASAP7_75t_SL U56425 ( .A(n57402), .Y(n75641) );
  NAND2xp5_ASAP7_75t_SL U56426 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[18]), .B(
        n59631), .Y(n73311) );
  INVxp33_ASAP7_75t_SL U56427 ( .A(n65476), .Y(n65539) );
  NAND2xp5_ASAP7_75t_SL U56428 ( .A(n75832), .B(n61982), .Y(n75811) );
  AOI31xp33_ASAP7_75t_SL U56429 ( .A1(n68937), .A2(n68936), .A3(n68935), .B(
        n68934), .Y(n69001) );
  NAND2xp33_ASAP7_75t_SL U56430 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[19]), .B(n70038), .Y(n69975) );
  INVxp33_ASAP7_75t_SL U56431 ( .A(n61733), .Y(n61701) );
  INVxp67_ASAP7_75t_SL U56432 ( .A(n71148), .Y(n71086) );
  OAI21xp33_ASAP7_75t_SL U56433 ( .A1(or1200_cpu_or1200_except_n528), .A2(
        n76724), .B(n64101), .Y(n64102) );
  AOI21xp5_ASAP7_75t_SL U56434 ( .A1(n65126), .A2(n65125), .B(n65144), .Y(
        n65127) );
  AOI21xp33_ASAP7_75t_SL U56435 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[5]), .B(n69737), 
        .Y(n69738) );
  OAI21xp33_ASAP7_75t_SL U56436 ( .A1(n71066), .A2(n71281), .B(n71065), .Y(
        n71174) );
  OAI21xp5_ASAP7_75t_SL U56437 ( .A1(n74156), .A2(n74766), .B(n74157), .Y(
        n74748) );
  OAI21xp33_ASAP7_75t_SL U56438 ( .A1(n75618), .A2(n78089), .B(n75617), .Y(
        n78109) );
  OAI22xp33_ASAP7_75t_SL U56439 ( .A1(n76897), .A2(n65136), .B1(n75620), .B2(
        n65182), .Y(n65137) );
  NAND2xp33_ASAP7_75t_SL U56440 ( .A(n59687), .B(n78113), .Y(n547) );
  OAI21xp33_ASAP7_75t_SL U56441 ( .A1(n75330), .A2(n77078), .B(n62120), .Y(
        n62126) );
  INVxp33_ASAP7_75t_SL U56442 ( .A(n78113), .Y(n78112) );
  NAND2xp33_ASAP7_75t_SL U56443 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[2]), .B(
        n59631), .Y(n73240) );
  NAND2xp33_ASAP7_75t_SL U56444 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_12_), .B(n69476), .Y(
        n69511) );
  NAND2xp5_ASAP7_75t_SL U56445 ( .A(n72689), .B(n72729), .Y(n72747) );
  INVxp33_ASAP7_75t_SL U56446 ( .A(n65542), .Y(n65555) );
  NAND2xp33_ASAP7_75t_SL U56447 ( .A(n59687), .B(n78117), .Y(n545) );
  OAI22xp33_ASAP7_75t_SL U56448 ( .A1(n61629), .A2(n62422), .B1(n61628), .B2(
        n62128), .Y(n61662) );
  NAND2xp5_ASAP7_75t_SL U56449 ( .A(n65403), .B(n65476), .Y(n65431) );
  BUFx3_ASAP7_75t_SL U56450 ( .A(n67846), .Y(n57167) );
  INVxp67_ASAP7_75t_SL U56451 ( .A(n62980), .Y(n62981) );
  OAI21xp5_ASAP7_75t_SL U56452 ( .A1(n61626), .A2(n61629), .B(n61625), .Y(
        n62130) );
  NOR2x1_ASAP7_75t_SL U56453 ( .A(n783), .B(n60079), .Y(n60171) );
  AOI21xp5_ASAP7_75t_SL U56454 ( .A1(n59672), .A2(n63407), .B(n63406), .Y(
        n63408) );
  INVxp33_ASAP7_75t_SL U56455 ( .A(n67964), .Y(n64396) );
  INVxp67_ASAP7_75t_SL U56456 ( .A(n78117), .Y(n78116) );
  NAND2xp33_ASAP7_75t_SL U56457 ( .A(n59656), .B(n59614), .Y(n62793) );
  NOR2x1_ASAP7_75t_SL U56458 ( .A(n66049), .B(n66052), .Y(n66085) );
  OAI21xp33_ASAP7_75t_SL U56459 ( .A1(n72874), .A2(n72971), .B(n73040), .Y(
        n72863) );
  OAI22xp33_ASAP7_75t_SL U56460 ( .A1(n71149), .A2(n70867), .B1(n71362), .B2(
        n70778), .Y(n70760) );
  INVx5_ASAP7_75t_SL U56461 ( .A(n58892), .Y(n59510) );
  OAI21xp5_ASAP7_75t_SL U56462 ( .A1(n74278), .A2(n74071), .B(n74738), .Y(
        n74224) );
  OAI21xp5_ASAP7_75t_SL U56463 ( .A1(n59630), .A2(n73163), .B(n73162), .Y(
        n73165) );
  NAND2xp33_ASAP7_75t_SL U56464 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[19]), .B(
        n59631), .Y(n73302) );
  NAND2xp5_ASAP7_75t_SL U56465 ( .A(n74277), .B(n74070), .Y(n74243) );
  INVxp33_ASAP7_75t_SL U56466 ( .A(n73207), .Y(n73212) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U56467 ( .A1(n66049), .A2(n66047), .B(n66051), .C(
        n66046), .Y(n66048) );
  NAND2xp33_ASAP7_75t_SL U56468 ( .A(n73484), .B(n59631), .Y(n73233) );
  NAND2xp33_ASAP7_75t_SL U56469 ( .A(n71799), .B(n71701), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n123) );
  INVxp33_ASAP7_75t_SL U56470 ( .A(n75517), .Y(n74031) );
  NAND3xp33_ASAP7_75t_SRAM U56471 ( .A(n78140), .B(n59687), .C(n78139), .Y(
        n535) );
  INVx1_ASAP7_75t_SL U56472 ( .A(n70932), .Y(n70898) );
  AOI21xp33_ASAP7_75t_SL U56473 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[6]), .B(n69763), 
        .Y(n69764) );
  OR2x2_ASAP7_75t_SL U56474 ( .A(n76844), .B(n77367), .Y(n77269) );
  INVxp67_ASAP7_75t_SL U56475 ( .A(n70885), .Y(n70909) );
  OAI21xp33_ASAP7_75t_SL U56476 ( .A1(n71281), .A2(n71148), .B(n71147), .Y(
        n71176) );
  OAI21xp33_ASAP7_75t_SL U56477 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_24_), .A2(
        n74298), .B(n74332), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n4) );
  AOI21xp33_ASAP7_75t_SL U56478 ( .A1(n76840), .A2(n76841), .B(n63760), .Y(
        n76517) );
  OAI21xp33_ASAP7_75t_SL U56479 ( .A1(n65964), .A2(n65816), .B(n65697), .Y(
        n66036) );
  INVx1_ASAP7_75t_SL U56480 ( .A(n70239), .Y(n70236) );
  BUFx3_ASAP7_75t_SL U56481 ( .A(n75044), .Y(n57260) );
  AOI21xp33_ASAP7_75t_SL U56482 ( .A1(n74956), .A2(n783), .B(n60079), .Y(
        n60077) );
  AOI31xp33_ASAP7_75t_SRAM U56483 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_21_), .A2(n69443), .A3(
        n70021), .B(n69442), .Y(n69444) );
  NOR3xp33_ASAP7_75t_SRAM U56484 ( .A(n75479), .B(n76486), .C(n75478), .Y(
        n75528) );
  NAND2xp33_ASAP7_75t_SL U56485 ( .A(n65402), .B(n65312), .Y(n1782) );
  OAI22xp33_ASAP7_75t_SL U56486 ( .A1(n66226), .A2(n58597), .B1(n75447), .B2(
        n76890), .Y(n9253) );
  NAND2xp5_ASAP7_75t_SL U56487 ( .A(n61520), .B(n61519), .Y(n61522) );
  AOI21xp33_ASAP7_75t_SL U56488 ( .A1(n58296), .A2(n77899), .B(n77211), .Y(
        n77213) );
  NAND2xp33_ASAP7_75t_SL U56489 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_20_), .B(n69476), .Y(
        n69469) );
  AND2x2_ASAP7_75t_SL U56490 ( .A(n77931), .B(n60551), .Y(n77052) );
  NAND2xp5_ASAP7_75t_SL U56491 ( .A(n65766), .B(n65765), .Y(n65986) );
  NAND2xp5_ASAP7_75t_SL U56492 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[5]), .B(
        n59630), .Y(n73220) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56493 ( .A1(
        or1200_cpu_or1200_mult_mac_div_cntr_1_), .A2(
        or1200_cpu_or1200_mult_mac_div_cntr_0_), .B(n61811), .C(n76631), .Y(
        or1200_cpu_or1200_mult_mac_n1105) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U56494 ( .A1(n65249), .A2(n65248), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .C(n65247), .Y(
        n65252) );
  AOI22xp33_ASAP7_75t_SL U56495 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_18_), .A2(n70023), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_19_), .B2(n69476), .Y(
        n69477) );
  OAI21xp33_ASAP7_75t_SL U56496 ( .A1(n62376), .A2(n64768), .B(n62375), .Y(
        n62379) );
  INVxp33_ASAP7_75t_SL U56497 ( .A(n77367), .Y(n77369) );
  INVxp33_ASAP7_75t_SL U56498 ( .A(n67711), .Y(n67717) );
  NAND2xp33_ASAP7_75t_SL U56499 ( .A(n59526), .B(n71333), .Y(n71338) );
  INVx1_ASAP7_75t_SL U56500 ( .A(n65980), .Y(n66065) );
  OAI22xp33_ASAP7_75t_SL U56501 ( .A1(n73008), .A2(n72965), .B1(n72859), .B2(
        n72738), .Y(n72715) );
  NAND2xp33_ASAP7_75t_SL U56502 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_6_), .B(n70023), .Y(
        n69481) );
  INVx1_ASAP7_75t_SL U56503 ( .A(n76731), .Y(n62508) );
  AOI22xp33_ASAP7_75t_SL U56504 ( .A1(n70104), .A2(n78330), .B1(n78331), .B2(
        n70038), .Y(n69767) );
  AOI22xp33_ASAP7_75t_SL U56505 ( .A1(n75649), .A2(n77880), .B1(n64179), .B2(
        n75396), .Y(n64183) );
  INVxp33_ASAP7_75t_SL U56506 ( .A(n75396), .Y(n63918) );
  INVxp67_ASAP7_75t_SL U56507 ( .A(n73036), .Y(n72837) );
  INVxp67_ASAP7_75t_SL U56508 ( .A(n65825), .Y(n65826) );
  AOI21xp33_ASAP7_75t_SL U56509 ( .A1(n75649), .A2(n77885), .B(n74978), .Y(
        n74979) );
  NAND2xp5_ASAP7_75t_SL U56510 ( .A(n72876), .B(n72751), .Y(n72839) );
  NAND2xp33_ASAP7_75t_SL U56511 ( .A(n77112), .B(n62348), .Y(n62349) );
  INVxp67_ASAP7_75t_SL U56512 ( .A(n62089), .Y(n62090) );
  INVxp67_ASAP7_75t_SL U56513 ( .A(n75984), .Y(n75979) );
  NAND2xp5_ASAP7_75t_SL U56514 ( .A(n66052), .B(n65980), .Y(n65981) );
  OAI21xp33_ASAP7_75t_SL U56515 ( .A1(or1200_cpu_or1200_except_n256), .A2(
        n76731), .B(n60830), .Y(n60832) );
  AOI21xp33_ASAP7_75t_SL U56516 ( .A1(n65074), .A2(n59674), .B(n65073), .Y(
        n64173) );
  OAI21xp33_ASAP7_75t_SL U56517 ( .A1(n75865), .A2(n74607), .B(n62439), .Y(
        n62442) );
  INVxp33_ASAP7_75t_SL U56518 ( .A(n72940), .Y(n72941) );
  NAND2xp33_ASAP7_75t_SL U56519 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .B(
        n72758), .Y(n72803) );
  AOI21xp33_ASAP7_75t_SL U56520 ( .A1(n70023), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_20_), .B(n70022), .Y(
        n70024) );
  INVxp33_ASAP7_75t_SL U56521 ( .A(n63543), .Y(n63544) );
  OAI21xp33_ASAP7_75t_SL U56522 ( .A1(n64108), .A2(n76801), .B(n61451), .Y(
        n61456) );
  O2A1O1Ixp33_ASAP7_75t_SL U56523 ( .A1(n61478), .A2(n61753), .B(n61556), .C(
        n61477), .Y(n61479) );
  OAI21xp33_ASAP7_75t_SL U56524 ( .A1(n65970), .A2(n65969), .B(n65968), .Y(
        n65976) );
  INVx1_ASAP7_75t_SL U56525 ( .A(n57107), .Y(n57171) );
  INVxp33_ASAP7_75t_SL U56526 ( .A(n75679), .Y(n75682) );
  OAI21xp33_ASAP7_75t_SL U56527 ( .A1(n65972), .A2(n65920), .B(n65888), .Y(
        n65889) );
  OAI21xp33_ASAP7_75t_SL U56528 ( .A1(n77079), .A2(n77078), .B(n77077), .Y(
        n77086) );
  INVxp67_ASAP7_75t_SL U56529 ( .A(n61182), .Y(n61235) );
  INVxp67_ASAP7_75t_SL U56530 ( .A(n66052), .Y(n65983) );
  NAND2xp5_ASAP7_75t_SL U56531 ( .A(n66022), .B(n65968), .Y(n66001) );
  OAI21xp33_ASAP7_75t_SL U56532 ( .A1(or1200_cpu_or1200_except_n260), .A2(
        n76731), .B(n62414), .Y(n62415) );
  INVxp67_ASAP7_75t_SL U56533 ( .A(n61950), .Y(n61951) );
  OAI21xp5_ASAP7_75t_SL U56534 ( .A1(n66050), .A2(n65970), .B(n65880), .Y(
        n66068) );
  INVxp67_ASAP7_75t_SL U56535 ( .A(n61955), .Y(n60784) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56536 ( .A1(
        or1200_cpu_or1200_mult_mac_div_cntr_4_), .A2(n61812), .B(n75759), .C(
        n76631), .Y(or1200_cpu_or1200_mult_mac_n1107) );
  NAND2xp5_ASAP7_75t_SL U56537 ( .A(n68793), .B(n53437), .Y(n68766) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56538 ( .A1(n65654), .A2(n65742), .B(n65653), 
        .C(n65652), .Y(n65656) );
  INVx1_ASAP7_75t_SL U56539 ( .A(n69500), .Y(n69746) );
  AND2x4_ASAP7_75t_SL U56540 ( .A(n57883), .B(n59043), .Y(n58753) );
  NAND2xp33_ASAP7_75t_SL U56541 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[15]), .B(
        n59631), .Y(n73146) );
  OAI22xp33_ASAP7_75t_SL U56542 ( .A1(n61629), .A2(n75316), .B1(n62422), .B2(
        n62128), .Y(n61112) );
  OAI21xp33_ASAP7_75t_SL U56543 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), 
        .A2(n72758), .B(n72757), .Y(n72759) );
  OAI21xp5_ASAP7_75t_SL U56544 ( .A1(n70112), .A2(n69580), .B(n69579), .Y(
        n69940) );
  NAND2xp5_ASAP7_75t_SL U56545 ( .A(n65978), .B(n65968), .Y(n65998) );
  NAND2xp5_ASAP7_75t_SL U56546 ( .A(n66024), .B(n65968), .Y(n65996) );
  NAND2xp5_ASAP7_75t_SL U56547 ( .A(n65931), .B(n65930), .Y(n66042) );
  AND4x1_ASAP7_75t_SL U56548 ( .A(n61409), .B(n60682), .C(n60681), .D(n60680), 
        .Y(n60683) );
  AOI21xp33_ASAP7_75t_SL U56549 ( .A1(n59680), .A2(n77899), .B(n77203), .Y(
        n77204) );
  OAI22xp33_ASAP7_75t_SL U56550 ( .A1(n73013), .A2(n73012), .B1(n73031), .B2(
        n73011), .Y(n73014) );
  OAI21xp33_ASAP7_75t_SL U56551 ( .A1(n66027), .A2(n65896), .B(n65968), .Y(
        n65809) );
  OAI21xp33_ASAP7_75t_SL U56552 ( .A1(n65972), .A2(n66002), .B(n65968), .Y(
        n65943) );
  NAND2xp33_ASAP7_75t_SL U56553 ( .A(n78425), .B(n70038), .Y(n69895) );
  AOI21xp33_ASAP7_75t_SL U56554 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[13]), .B(n69845), .Y(n69846) );
  OAI21xp33_ASAP7_75t_SL U56555 ( .A1(n75729), .A2(n77107), .B(n63589), .Y(
        n63590) );
  INVxp33_ASAP7_75t_SL U56556 ( .A(n65985), .Y(n65847) );
  NAND2xp5_ASAP7_75t_SL U56557 ( .A(n73551), .B(n73550), .Y(n73553) );
  AOI21xp33_ASAP7_75t_SL U56558 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[11]), .B(n69826), .Y(n69827) );
  OAI22xp33_ASAP7_75t_SL U56559 ( .A1(n63896), .A2(n63895), .B1(n74639), .B2(
        n65182), .Y(n63905) );
  NAND2xp5_ASAP7_75t_SL U56560 ( .A(n72775), .B(n72774), .Y(n72989) );
  INVxp67_ASAP7_75t_SL U56561 ( .A(n62075), .Y(n62083) );
  NAND2xp5_ASAP7_75t_SL U56562 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[24]), .B(
        n59631), .Y(n73114) );
  OAI21xp33_ASAP7_75t_SL U56563 ( .A1(n59569), .A2(n62340), .B(n62339), .Y(
        n62343) );
  AOI21xp33_ASAP7_75t_SL U56564 ( .A1(n72635), .A2(n72634), .B(n72640), .Y(
        n52526) );
  INVxp67_ASAP7_75t_SL U56565 ( .A(n65987), .Y(n66066) );
  INVxp67_ASAP7_75t_SL U56566 ( .A(n72636), .Y(n72637) );
  NAND2xp33_ASAP7_75t_SL U56567 ( .A(n78424), .B(n70038), .Y(n69923) );
  INVxp67_ASAP7_75t_SL U56568 ( .A(n62073), .Y(n62087) );
  OAI21xp33_ASAP7_75t_SL U56569 ( .A1(n77749), .A2(n61629), .B(n61081), .Y(
        n61082) );
  OAI21xp33_ASAP7_75t_SL U56570 ( .A1(n61626), .A2(n62128), .B(n61077), .Y(
        n61083) );
  OAI21xp33_ASAP7_75t_SL U56571 ( .A1(n59671), .A2(n75011), .B(n75010), .Y(
        n75001) );
  NAND2xp5_ASAP7_75t_SL U56572 ( .A(n65993), .B(n58576), .Y(n65994) );
  OAI21xp33_ASAP7_75t_SL U56573 ( .A1(or1200_cpu_or1200_mult_mac_n231), .A2(
        n77633), .B(n77632), .Y(n77634) );
  OAI21xp33_ASAP7_75t_SL U56574 ( .A1(n1496), .A2(n61755), .B(n61754), .Y(
        n61756) );
  NAND2xp33_ASAP7_75t_SL U56575 ( .A(n65955), .B(n66062), .Y(n65770) );
  NAND2xp5_ASAP7_75t_SL U56576 ( .A(n75238), .B(n75237), .Y(n75254) );
  NOR2xp33_ASAP7_75t_SRAM U56577 ( .A(or1200_cpu_or1200_except_n268), .B(
        n76731), .Y(n62325) );
  AOI21xp33_ASAP7_75t_SL U56578 ( .A1(n63557), .A2(n74986), .B(n63556), .Y(
        n63558) );
  OAI21xp33_ASAP7_75t_SL U56579 ( .A1(n78432), .A2(n70021), .B(n69422), .Y(
        n69423) );
  AOI21xp33_ASAP7_75t_SL U56580 ( .A1(n62345), .A2(n61781), .B(n61780), .Y(
        n61789) );
  INVxp33_ASAP7_75t_SL U56581 ( .A(n65971), .Y(n65915) );
  INVxp67_ASAP7_75t_SL U56582 ( .A(n76474), .Y(n76475) );
  NAND2xp33_ASAP7_75t_SL U56583 ( .A(n72990), .B(n72812), .Y(n72718) );
  NAND2xp33_ASAP7_75t_SL U56584 ( .A(n59672), .B(n64167), .Y(n63896) );
  NAND2xp5_ASAP7_75t_SL U56585 ( .A(n70244), .B(n70597), .Y(n3154) );
  AOI22xp33_ASAP7_75t_SL U56586 ( .A1(n73379), .A2(n73129), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[16]), .B2(
        n73382), .Y(n73294) );
  OAI21xp33_ASAP7_75t_SL U56587 ( .A1(n65972), .A2(n65973), .B(n65718), .Y(
        n65719) );
  OAI22xp33_ASAP7_75t_SL U56588 ( .A1(n65970), .A2(n66000), .B1(n65999), .B2(
        n65972), .Y(n65874) );
  NAND2xp33_ASAP7_75t_SL U56589 ( .A(n70571), .B(n70597), .Y(n3160) );
  OAI21xp33_ASAP7_75t_SL U56590 ( .A1(n77749), .A2(n62341), .B(n60585), .Y(
        n60588) );
  INVxp67_ASAP7_75t_SL U56591 ( .A(n70997), .Y(n70789) );
  OAI21xp33_ASAP7_75t_SL U56592 ( .A1(n61626), .A2(n62377), .B(n60586), .Y(
        n60587) );
  OAI21xp33_ASAP7_75t_SL U56593 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[7]), .A2(
        n70235), .B(n70597), .Y(n70245) );
  AOI21xp33_ASAP7_75t_SL U56594 ( .A1(n68770), .A2(n59672), .B(n68769), .Y(
        n68773) );
  INVxp67_ASAP7_75t_SL U56595 ( .A(n69464), .Y(n69465) );
  NAND2xp33_ASAP7_75t_SL U56596 ( .A(n66016), .B(n66051), .Y(n65907) );
  OAI21xp33_ASAP7_75t_SL U56597 ( .A1(n71731), .A2(n71730), .B(n71737), .Y(
        n71732) );
  NAND2xp33_ASAP7_75t_SL U56598 ( .A(n63677), .B(n59503), .Y(n63676) );
  BUFx3_ASAP7_75t_SL U56599 ( .A(n68096), .Y(n59435) );
  INVxp33_ASAP7_75t_SL U56600 ( .A(n62218), .Y(n62222) );
  AOI21xp33_ASAP7_75t_SL U56601 ( .A1(n60928), .A2(n76627), .B(n60927), .Y(
        n61182) );
  AOI22xp33_ASAP7_75t_SL U56602 ( .A1(n64119), .A2(n64839), .B1(n64293), .B2(
        n62260), .Y(n62282) );
  NAND2xp5_ASAP7_75t_SL U56603 ( .A(n60875), .B(n77087), .Y(n60880) );
  INVxp67_ASAP7_75t_SL U56604 ( .A(n75232), .Y(n75238) );
  AOI21xp5_ASAP7_75t_SL U56605 ( .A1(n75011), .A2(n57079), .B(n75010), .Y(
        n75003) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56606 ( .A1(n70104), .A2(n78427), .B(n69922), 
        .C(n70124), .Y(n69924) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U56607 ( .A1(n59540), .A2(n59580), .B(n75852), .C(
        n62445), .Y(n61733) );
  INVxp33_ASAP7_75t_SL U56608 ( .A(n65966), .Y(n65917) );
  INVxp67_ASAP7_75t_SL U56609 ( .A(n77096), .Y(n62340) );
  INVxp67_ASAP7_75t_SL U56610 ( .A(n72770), .Y(n72775) );
  BUFx3_ASAP7_75t_SL U56611 ( .A(n67610), .Y(n57274) );
  INVxp67_ASAP7_75t_SL U56612 ( .A(n72995), .Y(n72768) );
  INVx1_ASAP7_75t_SL U56613 ( .A(n59209), .Y(n57783) );
  OAI22xp33_ASAP7_75t_SL U56614 ( .A1(n63288), .A2(n76897), .B1(n77591), .B2(
        n65182), .Y(n63289) );
  NAND2xp5_ASAP7_75t_SL U56615 ( .A(n77752), .B(n77116), .Y(n60879) );
  INVxp33_ASAP7_75t_SL U56616 ( .A(n66076), .Y(n66077) );
  AOI22xp33_ASAP7_75t_SL U56617 ( .A1(n64119), .A2(n62257), .B1(n64293), .B2(
        n61785), .Y(n61786) );
  OAI21xp33_ASAP7_75t_SL U56618 ( .A1(n75317), .A2(n61626), .B(n60910), .Y(
        n60911) );
  OAI22xp33_ASAP7_75t_SL U56619 ( .A1(n73010), .A2(n72899), .B1(n73009), .B2(
        n72966), .Y(n72716) );
  BUFx4f_ASAP7_75t_SL U56620 ( .A(n67586), .Y(n57172) );
  INVxp67_ASAP7_75t_SL U56621 ( .A(n75476), .Y(n61904) );
  NAND2xp33_ASAP7_75t_SL U56622 ( .A(n71715), .B(n71799), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n125) );
  OAI21xp33_ASAP7_75t_SL U56623 ( .A1(n77749), .A2(n75314), .B(n60909), .Y(
        n60912) );
  AOI21xp33_ASAP7_75t_SL U56624 ( .A1(n75030), .A2(n62218), .B(n1175), .Y(
        n62217) );
  NAND2xp33_ASAP7_75t_SL U56625 ( .A(n59522), .B(n71039), .Y(n70718) );
  AOI22xp33_ASAP7_75t_SL U56626 ( .A1(n75705), .A2(n61782), .B1(n62274), .B2(
        n62260), .Y(n61788) );
  OAI21xp33_ASAP7_75t_SL U56627 ( .A1(n1177), .A2(n62215), .B(n62214), .Y(
        n9274) );
  OA21x2_ASAP7_75t_SL U56628 ( .A1(n78335), .A2(n70021), .B(n69460), .Y(n69461) );
  OAI22xp33_ASAP7_75t_SL U56629 ( .A1(n63463), .A2(n76897), .B1(n77295), .B2(
        n65182), .Y(n63464) );
  INVxp67_ASAP7_75t_SL U56630 ( .A(n75357), .Y(n60987) );
  OAI22xp33_ASAP7_75t_SL U56631 ( .A1(n65971), .A2(n65970), .B1(n65972), .B2(
        n65966), .Y(n65689) );
  INVxp33_ASAP7_75t_SL U56632 ( .A(n64191), .Y(n64200) );
  OAI21xp33_ASAP7_75t_SL U56633 ( .A1(n65244), .A2(n65240), .B(n65239), .Y(
        n65312) );
  OAI22xp33_ASAP7_75t_SL U56634 ( .A1(n65916), .A2(n66027), .B1(n65974), .B2(
        n65967), .Y(n65704) );
  NOR2xp33_ASAP7_75t_SL U56635 ( .A(n72635), .B(n72634), .Y(n72640) );
  NAND2xp33_ASAP7_75t_SL U56636 ( .A(n65816), .B(n66075), .Y(n65697) );
  OAI21xp33_ASAP7_75t_SL U56637 ( .A1(n1432), .A2(n57114), .B(n75402), .Y(
        n9280) );
  AOI21xp33_ASAP7_75t_SL U56638 ( .A1(n75011), .A2(n75010), .B(n75009), .Y(
        n75012) );
  OAI22xp33_ASAP7_75t_SL U56639 ( .A1(n76897), .A2(n65183), .B1(n69371), .B2(
        n65182), .Y(n65184) );
  OAI21xp33_ASAP7_75t_SL U56640 ( .A1(n63564), .A2(n61626), .B(n61179), .Y(
        n61180) );
  OAI21xp33_ASAP7_75t_SL U56641 ( .A1(n77749), .A2(n63565), .B(n61178), .Y(
        n61181) );
  INVx2_ASAP7_75t_SL U56642 ( .A(n75903), .Y(n57173) );
  NAND2xp5_ASAP7_75t_SL U56643 ( .A(n72431), .B(n72430), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n72) );
  AOI21xp33_ASAP7_75t_SL U56644 ( .A1(n59571), .A2(n76280), .B(n76288), .Y(
        n60771) );
  OAI21xp33_ASAP7_75t_SL U56645 ( .A1(n1434), .A2(n57114), .B(n66223), .Y(
        n9281) );
  OAI22xp33_ASAP7_75t_SL U56646 ( .A1(n65974), .A2(n65973), .B1(n65972), .B2(
        n65971), .Y(n65975) );
  NAND2xp33_ASAP7_75t_SL U56647 ( .A(n66017), .B(n66051), .Y(n65993) );
  NOR2x1_ASAP7_75t_SL U56648 ( .A(or1200_cpu_or1200_except_n524), .B(n75311), 
        .Y(n74593) );
  INVxp33_ASAP7_75t_SL U56649 ( .A(n76423), .Y(n76420) );
  OAI21xp33_ASAP7_75t_SL U56650 ( .A1(n1436), .A2(n57114), .B(n74078), .Y(
        n9282) );
  NAND2xp33_ASAP7_75t_SL U56651 ( .A(n77117), .B(n77116), .Y(n77118) );
  INVxp33_ASAP7_75t_SL U56652 ( .A(n63546), .Y(n63548) );
  INVx2_ASAP7_75t_SL U56653 ( .A(n63120), .Y(n57174) );
  OAI21xp33_ASAP7_75t_SL U56654 ( .A1(n78434), .A2(n70109), .B(n69447), .Y(
        n69580) );
  NAND2xp33_ASAP7_75t_SL U56655 ( .A(n73134), .B(n73382), .Y(n73135) );
  OAI22xp33_ASAP7_75t_SL U56656 ( .A1(n73009), .A2(n72787), .B1(n73010), .B2(
        n72935), .Y(n72780) );
  NAND2xp5_ASAP7_75t_SL U56657 ( .A(n66060), .B(n66076), .Y(n65980) );
  OAI21xp33_ASAP7_75t_SL U56658 ( .A1(n78429), .A2(n70109), .B(n69478), .Y(
        n69500) );
  OAI21xp33_ASAP7_75t_SL U56659 ( .A1(n1440), .A2(n57114), .B(n75404), .Y(
        n9284) );
  AOI22xp33_ASAP7_75t_SL U56660 ( .A1(n73379), .A2(n73333), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[23]), .B2(
        n73382), .Y(n73352) );
  NOR3xp33_ASAP7_75t_SRAM U56661 ( .A(n72966), .B(n72965), .C(n72964), .Y(
        n72968) );
  INVxp33_ASAP7_75t_SL U56662 ( .A(n62307), .Y(n62315) );
  NAND2xp5_ASAP7_75t_SL U56663 ( .A(n59537), .B(n61939), .Y(n62075) );
  OAI21xp33_ASAP7_75t_SL U56664 ( .A1(n1442), .A2(n57114), .B(n75401), .Y(
        n9285) );
  AOI22xp33_ASAP7_75t_SL U56665 ( .A1(n61631), .A2(n62260), .B1(n61785), .B2(
        n64219), .Y(n61110) );
  NAND2xp33_ASAP7_75t_SL U56666 ( .A(n59541), .B(n61798), .Y(n61676) );
  AOI22xp33_ASAP7_75t_SL U56667 ( .A1(n73030), .A2(n72889), .B1(n73024), .B2(
        n72908), .Y(n72804) );
  OAI22xp33_ASAP7_75t_SL U56668 ( .A1(n72859), .A2(n72788), .B1(n73008), .B2(
        n72890), .Y(n72783) );
  OAI21xp33_ASAP7_75t_SL U56669 ( .A1(n78367), .A2(n70021), .B(n70020), .Y(
        n70022) );
  OAI21xp33_ASAP7_75t_SL U56670 ( .A1(n73570), .A2(n73569), .B(n73568), .Y(
        n73580) );
  OAI21xp33_ASAP7_75t_SL U56671 ( .A1(n1444), .A2(n57114), .B(n62159), .Y(
        n9286) );
  INVxp33_ASAP7_75t_SL U56672 ( .A(n76258), .Y(n61952) );
  OAI21xp33_ASAP7_75t_SL U56673 ( .A1(n1446), .A2(n57114), .B(n64184), .Y(
        n9287) );
  OAI21xp33_ASAP7_75t_SL U56674 ( .A1(n1448), .A2(n57114), .B(n63919), .Y(
        n9288) );
  OAI21xp33_ASAP7_75t_SL U56675 ( .A1(n66027), .A2(n66026), .B(n66025), .Y(
        n66046) );
  OAI21xp33_ASAP7_75t_SL U56676 ( .A1(n74208), .A2(n66138), .B(n66164), .Y(
        n65609) );
  NAND2xp33_ASAP7_75t_SL U56677 ( .A(n66008), .B(n66051), .Y(n66009) );
  OAI21xp33_ASAP7_75t_SL U56678 ( .A1(n61626), .A2(n61703), .B(n61553), .Y(
        n74621) );
  AOI21xp5_ASAP7_75t_SL U56679 ( .A1(n61511), .A2(n62373), .B(n60676), .Y(
        n60681) );
  OAI21xp33_ASAP7_75t_SL U56680 ( .A1(n1454), .A2(n57114), .B(n75403), .Y(
        n9291) );
  NAND2xp5_ASAP7_75t_SL U56681 ( .A(n69578), .B(n69577), .Y(n69579) );
  AOI22xp33_ASAP7_75t_SL U56682 ( .A1(n75524), .A2(n75523), .B1(n77971), .B2(
        n77212), .Y(n75525) );
  INVxp67_ASAP7_75t_SL U56683 ( .A(n75310), .Y(n63547) );
  NAND2xp33_ASAP7_75t_SL U56684 ( .A(n72658), .B(n72657), .Y(n72659) );
  NAND2xp5_ASAP7_75t_SL U56685 ( .A(n61486), .B(n62288), .Y(n61446) );
  OAI21xp33_ASAP7_75t_SL U56686 ( .A1(n61639), .A2(n61417), .B(n60968), .Y(
        n60970) );
  OAI21xp33_ASAP7_75t_SL U56687 ( .A1(n78339), .A2(n70021), .B(n69448), .Y(
        n69449) );
  AOI22xp33_ASAP7_75t_SL U56688 ( .A1(n62382), .A2(n61450), .B1(n61449), .B2(
        n61448), .Y(n61451) );
  OAI21xp33_ASAP7_75t_SL U56689 ( .A1(n74353), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_9_), .B(
        n74319), .Y(n2428) );
  INVxp33_ASAP7_75t_SL U56690 ( .A(n65909), .Y(n65749) );
  INVxp33_ASAP7_75t_SL U56691 ( .A(n66039), .Y(n65949) );
  NAND2xp33_ASAP7_75t_SL U56692 ( .A(n65942), .B(n66051), .Y(n65870) );
  AOI22xp33_ASAP7_75t_SL U56693 ( .A1(n65978), .A2(n66008), .B1(n66024), .B2(
        n66006), .Y(n65941) );
  INVxp67_ASAP7_75t_SL U56694 ( .A(n63595), .Y(n61238) );
  INVxp67_ASAP7_75t_SL U56695 ( .A(n69762), .Y(n69596) );
  NAND2xp33_ASAP7_75t_SL U56696 ( .A(n65995), .B(n66051), .Y(n65940) );
  OAI22xp33_ASAP7_75t_SL U56697 ( .A1(n78430), .A2(n69564), .B1(n78355), .B2(
        n70021), .Y(n69440) );
  NAND2xp5_ASAP7_75t_SL U56698 ( .A(n72934), .B(n72933), .Y(n72945) );
  AOI22xp33_ASAP7_75t_SL U56699 ( .A1(n62382), .A2(n77589), .B1(n61449), .B2(
        n61227), .Y(n61232) );
  AOI21xp33_ASAP7_75t_SL U56700 ( .A1(n62374), .A2(n62373), .B(n62372), .Y(
        n62375) );
  AOI21xp33_ASAP7_75t_SL U56701 ( .A1(n73382), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[17]), .B(
        n73132), .Y(n73299) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56702 ( .A1(n70104), .A2(n78428), .B(n69894), 
        .C(n70124), .Y(n69896) );
  OAI22xp33_ASAP7_75t_SL U56703 ( .A1(n65974), .A2(n66011), .B1(n66027), .B2(
        n65939), .Y(n65825) );
  XNOR2xp5_ASAP7_75t_SRAM U56704 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[7]), .B(
        n74277), .Y(n74280) );
  INVx1_ASAP7_75t_SL U56705 ( .A(n76279), .Y(n62296) );
  AOI22xp33_ASAP7_75t_SL U56706 ( .A1(n66023), .A2(n65978), .B1(n66051), .B2(
        n66021), .Y(n65880) );
  OAI22xp33_ASAP7_75t_SL U56707 ( .A1(n66027), .A2(n66000), .B1(n65999), .B2(
        n65970), .Y(n65944) );
  INVxp67_ASAP7_75t_SL U56708 ( .A(n62088), .Y(n62091) );
  INVxp67_ASAP7_75t_SL U56709 ( .A(n71799), .Y(n71721) );
  OA21x2_ASAP7_75t_SL U56710 ( .A1(n78337), .A2(n70021), .B(n69486), .Y(n69487) );
  OAI21xp33_ASAP7_75t_SL U56711 ( .A1(n70232), .A2(n70224), .B(n70235), .Y(
        n70239) );
  INVx1_ASAP7_75t_SL U56712 ( .A(n76906), .Y(n59674) );
  OAI21xp33_ASAP7_75t_SL U56713 ( .A1(n61626), .A2(n64136), .B(n61401), .Y(
        n61404) );
  NOR4xp25_ASAP7_75t_SRAM U56714 ( .A(n75760), .B(n75516), .C(n75522), .D(
        n75515), .Y(n75521) );
  BUFx3_ASAP7_75t_SL U56715 ( .A(n57551), .Y(n57356) );
  AOI21xp33_ASAP7_75t_SL U56716 ( .A1(n61538), .A2(n57639), .B(n61221), .Y(
        n61222) );
  NOR2xp33_ASAP7_75t_SRAM U56717 ( .A(n78055), .B(n76844), .Y(n76845) );
  OAI22xp33_ASAP7_75t_SL U56718 ( .A1(n73008), .A2(n72909), .B1(n73009), .B2(
        n72890), .Y(n72755) );
  AOI22xp33_ASAP7_75t_SL U56719 ( .A1(n65958), .A2(n66051), .B1(n65978), .B2(
        n65954), .Y(n65931) );
  INVx1_ASAP7_75t_SL U56720 ( .A(n69564), .Y(n70023) );
  INVxp67_ASAP7_75t_SL U56721 ( .A(n72930), .Y(n72931) );
  INVxp33_ASAP7_75t_SL U56722 ( .A(n61768), .Y(n61200) );
  AOI21xp33_ASAP7_75t_SL U56723 ( .A1(n73026), .A2(n72898), .B(n72756), .Y(
        n72757) );
  OAI21xp33_ASAP7_75t_SL U56724 ( .A1(or1200_cpu_or1200_except_n520), .A2(
        n76724), .B(n62506), .Y(n62507) );
  INVxp67_ASAP7_75t_SL U56725 ( .A(n72898), .Y(n72738) );
  AOI22xp33_ASAP7_75t_SL U56726 ( .A1(n66017), .A2(n65978), .B1(n66051), .B2(
        n66020), .Y(n65765) );
  INVxp67_ASAP7_75t_SL U56727 ( .A(n60295), .Y(n60296) );
  AOI22xp33_ASAP7_75t_SL U56728 ( .A1(n59525), .A2(n73141), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[14]), .B2(
        n73382), .Y(n73282) );
  OAI22xp33_ASAP7_75t_SL U56729 ( .A1(n73010), .A2(n73023), .B1(n73009), .B2(
        n73029), .Y(n73012) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56730 ( .A1(n65803), .A2(n65802), .B(n65974), 
        .C(n65801), .Y(n65810) );
  NAND2xp5_ASAP7_75t_SL U56731 ( .A(n72451), .B(n72450), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n71) );
  OAI22xp33_ASAP7_75t_SL U56732 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_), .A2(n69564), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_3_), .B2(n70021), .Y(
        n69479) );
  INVxp67_ASAP7_75t_SL U56733 ( .A(n59657), .Y(n59125) );
  OAI21xp33_ASAP7_75t_SL U56734 ( .A1(n76906), .A2(n65074), .B(n65073), .Y(
        n64175) );
  INVxp33_ASAP7_75t_SL U56735 ( .A(n71064), .Y(n71066) );
  OAI22xp33_ASAP7_75t_SL U56736 ( .A1(n66106), .A2(n66153), .B1(n66109), .B2(
        n66122), .Y(n65521) );
  NAND2xp33_ASAP7_75t_SL U56737 ( .A(n70593), .B(n70597), .Y(n3156) );
  OAI21xp33_ASAP7_75t_SL U56738 ( .A1(n64313), .A2(n77749), .B(n60838), .Y(
        n60839) );
  INVxp33_ASAP7_75t_SL U56739 ( .A(n76288), .Y(n76283) );
  INVxp67_ASAP7_75t_SL U56740 ( .A(n66137), .Y(n65577) );
  INVxp67_ASAP7_75t_SL U56741 ( .A(n76280), .Y(n76281) );
  INVxp33_ASAP7_75t_SL U56742 ( .A(n74298), .Y(n74299) );
  INVxp33_ASAP7_75t_SL U56743 ( .A(n71424), .Y(n71425) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56744 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[16]), .A2(
        n70104), .B(n69974), .C(n70124), .Y(n69976) );
  OAI21xp33_ASAP7_75t_SL U56745 ( .A1(n66119), .A2(n66132), .B(n66118), .Y(
        n66131) );
  OAI21xp33_ASAP7_75t_SL U56746 ( .A1(n61626), .A2(n62253), .B(n60837), .Y(
        n60840) );
  NAND2xp5_ASAP7_75t_SL U56747 ( .A(n72670), .B(n72669), .Y(n72677) );
  INVxp33_ASAP7_75t_SL U56748 ( .A(n73029), .Y(n72991) );
  AOI22xp33_ASAP7_75t_SL U56749 ( .A1(n59525), .A2(n73304), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[19]), .B2(
        n73382), .Y(n73320) );
  NAND2xp33_ASAP7_75t_SL U56750 ( .A(n71209), .B(n71039), .Y(n71043) );
  NAND2xp5_ASAP7_75t_SL U56751 ( .A(n72672), .B(n72671), .Y(n72674) );
  NAND2xp5_ASAP7_75t_SL U56752 ( .A(n72269), .B(n72486), .Y(n72368) );
  NAND2xp33_ASAP7_75t_SL U56753 ( .A(n71087), .B(n71282), .Y(n71042) );
  NAND2xp33_ASAP7_75t_SL U56754 ( .A(n70587), .B(n70597), .Y(n3157) );
  INVxp33_ASAP7_75t_SL U56755 ( .A(n78138), .Y(n78140) );
  AOI31xp33_ASAP7_75t_SL U56756 ( .A1(n69762), .A2(n69761), .A3(n69760), .B(
        n69759), .Y(n69790) );
  AOI22xp33_ASAP7_75t_SL U56757 ( .A1(n71087), .A2(n71064), .B1(n71115), .B2(
        n59522), .Y(n70932) );
  NAND2xp33_ASAP7_75t_SL U56758 ( .A(n59687), .B(n77985), .Y(n3910) );
  INVxp67_ASAP7_75t_SL U56759 ( .A(n66132), .Y(n66134) );
  OAI21xp33_ASAP7_75t_SL U56760 ( .A1(n77749), .A2(n61703), .B(n61549), .Y(
        n61550) );
  NAND2xp33_ASAP7_75t_SL U56761 ( .A(n72734), .B(n72995), .Y(n72693) );
  AOI22xp33_ASAP7_75t_SL U56762 ( .A1(n59525), .A2(n73180), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[12]), .B2(
        n73382), .Y(n73274) );
  OAI21xp33_ASAP7_75t_SL U56763 ( .A1(or1200_cpu_or1200_except_n532), .A2(
        n76724), .B(n64278), .Y(n64280) );
  NAND2xp33_ASAP7_75t_SL U56764 ( .A(n70573), .B(n70597), .Y(n3159) );
  OAI21xp33_ASAP7_75t_SL U56765 ( .A1(n61626), .A2(n74619), .B(n61545), .Y(
        n61551) );
  INVxp67_ASAP7_75t_SL U56766 ( .A(n59513), .Y(n58928) );
  NAND2xp5_ASAP7_75t_SL U56767 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[7]), .B(
        n74277), .Y(n74071) );
  AOI22xp33_ASAP7_75t_SL U56768 ( .A1(n59525), .A2(n73123), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[20]), .B2(
        n73382), .Y(n73324) );
  INVxp33_ASAP7_75t_SL U56769 ( .A(n74069), .Y(n74070) );
  OAI21xp33_ASAP7_75t_SL U56770 ( .A1(n70112), .A2(n69577), .B(n70149), .Y(
        n69561) );
  INVx1_ASAP7_75t_SL U56771 ( .A(n58299), .Y(n58296) );
  AOI22xp33_ASAP7_75t_SL U56772 ( .A1(n71087), .A2(n71115), .B1(n59522), .B2(
        n71172), .Y(n71018) );
  INVxp67_ASAP7_75t_SL U56773 ( .A(n71040), .Y(n71103) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U56774 ( .A1(n70104), .A2(n78425), .B(n69949), .C(
        n69948), .Y(n69950) );
  NAND2xp5_ASAP7_75t_SL U56775 ( .A(n72240), .B(n72239), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n80) );
  OAI21xp33_ASAP7_75t_SL U56776 ( .A1(n74751), .A2(n74205), .B(n74175), .Y(
        n74176) );
  OAI21xp33_ASAP7_75t_SL U56777 ( .A1(or1200_dc_top_from_dcram_5_), .A2(n61546), .B(n61080), .Y(n61629) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56778 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_1_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_2_), .B(
        n71702), .C(n71710), .Y(n71703) );
  AOI22xp33_ASAP7_75t_SL U56779 ( .A1(n77088), .A2(n61705), .B1(n61704), .B2(
        n77117), .Y(n61715) );
  AOI21xp33_ASAP7_75t_SL U56780 ( .A1(n75342), .A2(n65159), .B(n64831), .Y(
        n64832) );
  INVxp33_ASAP7_75t_SL U56781 ( .A(n71331), .Y(n71077) );
  INVxp67_ASAP7_75t_SL U56782 ( .A(n74883), .Y(n77193) );
  OAI22xp33_ASAP7_75t_SL U56783 ( .A1(n78345), .A2(n69563), .B1(n78349), .B2(
        n69488), .Y(n69458) );
  OAI21xp33_ASAP7_75t_SL U56784 ( .A1(or1200_dc_top_from_dcram_13_), .A2(
        n61546), .B(n61076), .Y(n62128) );
  NAND2xp33_ASAP7_75t_SL U56785 ( .A(n73384), .B(n73382), .Y(n73385) );
  OAI22xp33_ASAP7_75t_SL U56786 ( .A1(n63405), .A2(n76906), .B1(n76828), .B2(
        n68787), .Y(n63406) );
  INVxp33_ASAP7_75t_SL U56787 ( .A(or1200_cpu_or1200_rf_n44), .Y(n77932) );
  OA21x2_ASAP7_75t_SL U56788 ( .A1(n78352), .A2(n70021), .B(n69501), .Y(n69502) );
  INVxp33_ASAP7_75t_SL U56789 ( .A(n64108), .Y(n64139) );
  AOI22xp33_ASAP7_75t_SL U56790 ( .A1(n76888), .A2(n77971), .B1(n63438), .B2(
        n57079), .Y(n63443) );
  AOI22xp33_ASAP7_75t_SL U56791 ( .A1(n72512), .A2(n72375), .B1(n72412), .B2(
        n72376), .Y(n72379) );
  AOI22xp33_ASAP7_75t_SL U56792 ( .A1(n71209), .A2(n70997), .B1(n70996), .B2(
        n71331), .Y(n70998) );
  NAND2xp5_ASAP7_75t_SL U56793 ( .A(n72822), .B(n72821), .Y(n72971) );
  OAI21xp33_ASAP7_75t_SL U56794 ( .A1(n74169), .A2(n74205), .B(n74175), .Y(
        n74170) );
  NAND2xp5_ASAP7_75t_SL U56795 ( .A(n63440), .B(n63439), .Y(n63441) );
  OAI22xp33_ASAP7_75t_SL U56796 ( .A1(n73027), .A2(n73010), .B1(n72859), .B2(
        n73029), .Y(n72862) );
  NAND2xp5_ASAP7_75t_SL U56797 ( .A(n72796), .B(n72795), .Y(n72975) );
  INVxp33_ASAP7_75t_SL U56798 ( .A(n71710), .Y(n71711) );
  INVxp33_ASAP7_75t_SL U56799 ( .A(n71208), .Y(n70928) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U56800 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_5_), .A2(
        n74719), .B(n74718), .C(n74717), .Y(n74720) );
  NAND2xp33_ASAP7_75t_SL U56801 ( .A(n76960), .B(n76959), .Y(n76961) );
  AOI21xp5_ASAP7_75t_SL U56802 ( .A1(n65150), .A2(n65176), .B(n65171), .Y(
        n65152) );
  NAND2xp33_ASAP7_75t_SL U56803 ( .A(n59687), .B(n78160), .Y(n527) );
  NAND2xp33_ASAP7_75t_SL U56804 ( .A(n59687), .B(n77964), .Y(n3923) );
  AND2x4_ASAP7_75t_SL U56805 ( .A(n62673), .B(n62672), .Y(n59099) );
  AOI22xp33_ASAP7_75t_SL U56806 ( .A1(n73379), .A2(n73169), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[11]), .B2(
        n73382), .Y(n73168) );
  AOI22xp33_ASAP7_75t_SL U56807 ( .A1(n73026), .A2(n72902), .B1(n73024), .B2(
        n72741), .Y(n72743) );
  INVxp33_ASAP7_75t_SL U56808 ( .A(n69913), .Y(n69657) );
  NAND2xp5_ASAP7_75t_SL U56809 ( .A(or1200_cpu_or1200_mult_mac_n64), .B(n59657), .Y(n75984) );
  INVxp67_ASAP7_75t_SL U56810 ( .A(n70110), .Y(n70120) );
  OAI21xp33_ASAP7_75t_SL U56811 ( .A1(n62254), .A2(n62253), .B(n62252), .Y(
        n64315) );
  AOI21xp33_ASAP7_75t_SL U56812 ( .A1(n74372), .A2(n74359), .B(n74358), .Y(
        n74380) );
  NOR2x1_ASAP7_75t_SL U56813 ( .A(n66269), .B(n66259), .Y(n66270) );
  AOI22xp33_ASAP7_75t_SL U56814 ( .A1(n65409), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[33]), .B1(n65553), 
        .B2(n65661), .Y(n65542) );
  BUFx2_ASAP7_75t_SL U56815 ( .A(n58844), .Y(n57402) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56816 ( .A1(n65469), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[18]), .B(n65468), 
        .C(n65467), .Y(n65470) );
  AOI22xp33_ASAP7_75t_SL U56817 ( .A1(n76763), .A2(n76762), .B1(n76761), .B2(
        n76760), .Y(n76786) );
  OAI21xp33_ASAP7_75t_SL U56818 ( .A1(n72544), .A2(n72389), .B(n72388), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n77) );
  AOI21xp33_ASAP7_75t_SL U56819 ( .A1(n73382), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[25]), .B(
        n73380), .Y(n73393) );
  NAND2x1p5_ASAP7_75t_SL U56820 ( .A(n66254), .B(n66263), .Y(n75033) );
  AOI21xp5_ASAP7_75t_SL U56821 ( .A1(n78358), .A2(n72667), .B(n72666), .Y(
        n72680) );
  INVxp33_ASAP7_75t_SL U56822 ( .A(n65995), .Y(n65997) );
  AOI22xp33_ASAP7_75t_SL U56823 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_5_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_4_), .B2(n70018), .Y(
        n69482) );
  AOI22xp33_ASAP7_75t_SL U56824 ( .A1(n75570), .A2(
        or1200_dc_top_from_dcram_17_), .B1(dwb_dat_i[17]), .B2(n75569), .Y(
        n75357) );
  AOI21xp33_ASAP7_75t_SL U56825 ( .A1(n61829), .A2(n61833), .B(n60813), .Y(
        n60814) );
  INVx1_ASAP7_75t_SL U56826 ( .A(n63809), .Y(n63807) );
  AOI22xp33_ASAP7_75t_SL U56827 ( .A1(n66022), .A2(n66047), .B1(n66016), .B2(
        n65978), .Y(n65877) );
  INVx1_ASAP7_75t_SL U56828 ( .A(n75015), .Y(n65182) );
  AOI22xp33_ASAP7_75t_SL U56829 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_11_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_10_), .B2(n70018), .Y(
        n69501) );
  NAND2xp5_ASAP7_75t_SL U56830 ( .A(n75719), .B(n75718), .Y(n75732) );
  OAI22xp33_ASAP7_75t_SL U56831 ( .A1(n75317), .A2(n61628), .B1(n62284), .B2(
        n75314), .Y(n60986) );
  AOI22xp33_ASAP7_75t_SL U56832 ( .A1(n75649), .A2(n77877), .B1(n75398), .B2(
        n75397), .Y(n75399) );
  OAI21xp33_ASAP7_75t_SL U56833 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[16]), .A2(n66160), 
        .B(n65598), .Y(n65606) );
  INVxp33_ASAP7_75t_SL U56834 ( .A(n64773), .Y(n62361) );
  OAI22xp33_ASAP7_75t_SL U56835 ( .A1(n64834), .A2(n75574), .B1(n63583), .B2(
        n77101), .Y(n63591) );
  AOI21xp33_ASAP7_75t_SL U56836 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .A2(
        n72422), .B(n72172), .Y(n72150) );
  INVxp67_ASAP7_75t_SL U56837 ( .A(n66079), .Y(n66050) );
  AOI21xp5_ASAP7_75t_SL U56838 ( .A1(n78377), .A2(n72667), .B(n72615), .Y(
        n72631) );
  OAI22xp33_ASAP7_75t_SL U56839 ( .A1(n63583), .A2(n75574), .B1(n75729), .B2(
        n77105), .Y(n60866) );
  INVxp67_ASAP7_75t_SL U56840 ( .A(n65939), .Y(n66006) );
  NAND2xp33_ASAP7_75t_SL U56841 ( .A(n62493), .B(n75030), .Y(n62495) );
  OAI22xp33_ASAP7_75t_SL U56842 ( .A1(n65974), .A2(n65953), .B1(n66027), .B2(
        n66081), .Y(n66074) );
  AOI22xp33_ASAP7_75t_SL U56843 ( .A1(or1200_dc_top_from_dcram_20_), .A2(
        n58285), .B1(n75570), .B2(or1200_dc_top_from_dcram_28_), .Y(n61401) );
  AOI22xp33_ASAP7_75t_SL U56844 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_19_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_18_), .B2(n70018), .Y(
        n70020) );
  NAND2xp33_ASAP7_75t_SL U56845 ( .A(n66235), .B(n75030), .Y(n66237) );
  OAI21xp33_ASAP7_75t_SL U56846 ( .A1(n75244), .A2(n61783), .B(n61632), .Y(
        n61642) );
  OAI22xp33_ASAP7_75t_SL U56847 ( .A1(n75317), .A2(n75316), .B1(n75315), .B2(
        n75314), .Y(n75354) );
  INVx3_ASAP7_75t_SL U56848 ( .A(n57442), .Y(n64367) );
  NAND2xp5_ASAP7_75t_SL U56849 ( .A(n73569), .B(n73570), .Y(n73568) );
  NAND2xp5_ASAP7_75t_SL U56850 ( .A(n76421), .B(n74015), .Y(n76423) );
  NAND2xp33_ASAP7_75t_SL U56851 ( .A(n78337), .B(n70018), .Y(n69455) );
  INVxp67_ASAP7_75t_SL U56852 ( .A(n60977), .Y(n77586) );
  OAI21xp33_ASAP7_75t_SL U56853 ( .A1(n75324), .A2(n77093), .B(n61103), .Y(
        n61108) );
  INVxp67_ASAP7_75t_SL U56854 ( .A(n65942), .Y(n66002) );
  OAI22xp33_ASAP7_75t_SL U56855 ( .A1(n73009), .A2(n72888), .B1(n73008), .B2(
        n72885), .Y(n72687) );
  AOI21xp33_ASAP7_75t_SL U56856 ( .A1(n75387), .A2(n75386), .B(n75390), .Y(
        n75389) );
  OAI22xp33_ASAP7_75t_SL U56857 ( .A1(n75588), .A2(n75587), .B1(n75586), .B2(
        n77103), .Y(n75598) );
  OAI21xp5_ASAP7_75t_SL U56858 ( .A1(n72694), .A2(n72888), .B(n72692), .Y(
        n72995) );
  OAI22xp33_ASAP7_75t_SL U56859 ( .A1(n65953), .A2(n65970), .B1(n65974), .B2(
        n65929), .Y(n65796) );
  INVxp67_ASAP7_75t_SL U56860 ( .A(n70232), .Y(n70593) );
  OAI22xp33_ASAP7_75t_SL U56861 ( .A1(n75348), .A2(n75347), .B1(n75346), .B2(
        n75574), .Y(n75352) );
  OAI22xp5_ASAP7_75t_SL U56862 ( .A1(n57115), .A2(n70722), .B1(n70717), .B2(
        n70993), .Y(n71039) );
  OAI22xp33_ASAP7_75t_SL U56863 ( .A1(n75350), .A2(n77103), .B1(n75349), .B2(
        n75587), .Y(n75351) );
  NOR2xp33_ASAP7_75t_SRAM U56864 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]), .B(n70104), .Y(n69922) );
  AOI21xp33_ASAP7_75t_SL U56865 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .A2(
        n72298), .B(n72172), .Y(n72138) );
  OAI22xp33_ASAP7_75t_SL U56866 ( .A1(n65969), .A2(n65972), .B1(n65974), .B2(
        n65921), .Y(n65922) );
  OAI21xp5_ASAP7_75t_SL U56867 ( .A1(n65668), .A2(n65667), .B(n76976), .Y(
        n66076) );
  INVxp67_ASAP7_75t_SL U56868 ( .A(n70175), .Y(n70178) );
  OAI21xp5_ASAP7_75t_SL U56869 ( .A1(n60877), .A2(n61078), .B(n60876), .Y(
        n77116) );
  NAND2xp33_ASAP7_75t_SL U56870 ( .A(n62382), .B(n77608), .Y(n62383) );
  AOI22xp5_ASAP7_75t_SL U56871 ( .A1(or1200_dc_top_from_dcram_31_), .A2(n75570), .B1(n61544), .B2(or1200_dc_top_from_dcram_23_), .Y(n60878) );
  INVx8_ASAP7_75t_SL U56872 ( .A(n67343), .Y(n59504) );
  AOI22xp33_ASAP7_75t_SL U56873 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_3_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_), .B2(n70018), .Y(
        n69486) );
  NOR2x1p5_ASAP7_75t_SL U56874 ( .A(n59010), .B(n59115), .Y(n64034) );
  INVxp33_ASAP7_75t_SL U56875 ( .A(n61971), .Y(n61973) );
  AOI22xp33_ASAP7_75t_SL U56876 ( .A1(n66024), .A2(n66021), .B1(n66047), .B2(
        n65978), .Y(n65908) );
  AOI22xp33_ASAP7_75t_SL U56877 ( .A1(n73024), .A2(n72889), .B1(n73030), .B2(
        n72902), .Y(n72812) );
  NAND2xp5_ASAP7_75t_SL U56878 ( .A(n73893), .B(n73892), .Y(n74277) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56879 ( .A1(n59575), .A2(n75250), .B(n75249), 
        .C(n75248), .Y(n75252) );
  INVxp67_ASAP7_75t_SL U56880 ( .A(n60973), .Y(n60928) );
  INVxp33_ASAP7_75t_SL U56881 ( .A(n72915), .Y(n72936) );
  INVxp33_ASAP7_75t_SL U56882 ( .A(n72935), .Y(n72939) );
  AOI22xp33_ASAP7_75t_SL U56883 ( .A1(dwb_dat_i[17]), .A2(n61548), .B1(n75569), 
        .B2(dwb_dat_i[25]), .Y(n60910) );
  OAI22xp33_ASAP7_75t_SL U56884 ( .A1(n63577), .A2(n77107), .B1(n64843), .B2(
        n77103), .Y(n62258) );
  INVxp33_ASAP7_75t_SL U56885 ( .A(n69862), .Y(n69660) );
  AOI22xp33_ASAP7_75t_SL U56886 ( .A1(or1200_dc_top_from_dcram_25_), .A2(
        n75570), .B1(n58285), .B2(or1200_dc_top_from_dcram_17_), .Y(n60909) );
  NOR2x1_ASAP7_75t_SL U56887 ( .A(n74359), .B(n74372), .Y(n74358) );
  NAND2xp33_ASAP7_75t_SL U56888 ( .A(n78260), .B(n77040), .Y(n60992) );
  INVxp33_ASAP7_75t_SL U56889 ( .A(n72886), .Y(n72899) );
  OAI22xp33_ASAP7_75t_SL U56890 ( .A1(n62256), .A2(n75574), .B1(n62255), .B2(
        n75587), .Y(n62259) );
  INVxp33_ASAP7_75t_SL U56891 ( .A(n75587), .Y(n61367) );
  NAND2xp33_ASAP7_75t_SL U56892 ( .A(n72907), .B(n72890), .Y(n72932) );
  OAI21xp33_ASAP7_75t_SL U56893 ( .A1(n62319), .A2(n60902), .B(n60901), .Y(
        n60903) );
  INVx1_ASAP7_75t_SL U56894 ( .A(n72888), .Y(n72965) );
  AOI31xp33_ASAP7_75t_SRAM U56895 ( .A1(n61162), .A2(
        or1200_ic_top_from_icram[22]), .A3(n22057), .B(n60403), .Y(n60404) );
  INVxp67_ASAP7_75t_SL U56896 ( .A(n60902), .Y(n60904) );
  NAND2xp5_ASAP7_75t_SL U56897 ( .A(n59557), .B(n60759), .Y(n61399) );
  INVxp67_ASAP7_75t_SL U56898 ( .A(n72947), .Y(n72948) );
  INVx1_ASAP7_75t_SL U56899 ( .A(n71800), .Y(n71720) );
  NAND2xp33_ASAP7_75t_SL U56900 ( .A(n77065), .B(n62275), .Y(n62372) );
  INVxp67_ASAP7_75t_SL U56901 ( .A(n65959), .Y(n65937) );
  OAI21xp33_ASAP7_75t_SL U56902 ( .A1(n73008), .A2(n73027), .B(n73007), .Y(
        n73013) );
  NAND2xp33_ASAP7_75t_SL U56903 ( .A(n62382), .B(n77582), .Y(n60692) );
  AOI22xp33_ASAP7_75t_SL U56904 ( .A1(n66024), .A2(n66023), .B1(n66022), .B2(
        n66021), .Y(n66025) );
  AOI22xp33_ASAP7_75t_SL U56905 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_13_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_12_), .B2(n70018), .Y(
        n69474) );
  OAI21xp5_ASAP7_75t_SL U56906 ( .A1(n68780), .A2(n68768), .B(n68777), .Y(
        n68770) );
  OAI22xp33_ASAP7_75t_SL U56907 ( .A1(n64113), .A2(n77101), .B1(n62536), .B2(
        n77103), .Y(n62537) );
  NAND2xp5_ASAP7_75t_SL U56908 ( .A(n61481), .B(n77852), .Y(n60816) );
  NAND2xp5_ASAP7_75t_SL U56909 ( .A(n74294), .B(n74296), .Y(n74729) );
  OAI22xp33_ASAP7_75t_SL U56910 ( .A1(n73010), .A2(n72913), .B1(n73009), .B2(
        n72907), .Y(n72782) );
  NAND2xp5_ASAP7_75t_SL U56911 ( .A(n69690), .B(n69689), .Y(n69698) );
  AOI22xp33_ASAP7_75t_SL U56912 ( .A1(n66022), .A2(n66008), .B1(n65995), .B2(
        n65978), .Y(n65871) );
  AOI22xp33_ASAP7_75t_SL U56913 ( .A1(or1200_dc_top_from_dcram_21_), .A2(
        n58285), .B1(n75570), .B2(or1200_dc_top_from_dcram_29_), .Y(n61077) );
  AOI22xp33_ASAP7_75t_SL U56914 ( .A1(or1200_dc_top_from_dcram_30_), .A2(
        n75570), .B1(n58285), .B2(or1200_dc_top_from_dcram_22_), .Y(n60837) );
  OAI21xp33_ASAP7_75t_SL U56915 ( .A1(n74297), .A2(n74296), .B(n74295), .Y(
        n74300) );
  OAI22xp33_ASAP7_75t_SL U56916 ( .A1(n62284), .A2(n64313), .B1(n77601), .B2(
        n76796), .Y(n62285) );
  OAI21xp33_ASAP7_75t_SL U56917 ( .A1(n60203), .A2(n60202), .B(n60201), .Y(
        n60204) );
  NAND2xp5_ASAP7_75t_SL U56918 ( .A(n77847), .B(n77852), .Y(
        or1200_cpu_or1200_rf_n44) );
  INVx1_ASAP7_75t_SL U56919 ( .A(n60741), .Y(n61798) );
  OAI22xp33_ASAP7_75t_SL U56920 ( .A1(n66081), .A2(n65970), .B1(n65974), .B2(
        n65928), .Y(n65894) );
  OAI22xp33_ASAP7_75t_SL U56921 ( .A1(n77639), .A2(n77638), .B1(n77847), .B2(
        n77637), .Y(n77640) );
  INVxp67_ASAP7_75t_SL U56922 ( .A(n77619), .Y(n77620) );
  AOI22xp33_ASAP7_75t_SL U56923 ( .A1(n77672), .A2(n77901), .B1(n77644), .B2(
        n77627), .Y(n77628) );
  INVxp33_ASAP7_75t_SL U56924 ( .A(n65934), .Y(n65897) );
  OAI21xp33_ASAP7_75t_SL U56925 ( .A1(n73916), .A2(n75840), .B(n73915), .Y(
        n75251) );
  INVx1_ASAP7_75t_SL U56926 ( .A(n72161), .Y(n72326) );
  INVxp67_ASAP7_75t_SL U56927 ( .A(n60772), .Y(n60736) );
  INVxp67_ASAP7_75t_SL U56928 ( .A(n77105), .Y(n62260) );
  OAI22xp33_ASAP7_75t_SL U56929 ( .A1(n73008), .A2(n72911), .B1(n72859), .B2(
        n72915), .Y(n72781) );
  INVxp67_ASAP7_75t_SL U56930 ( .A(n70176), .Y(n70177) );
  AOI22xp33_ASAP7_75t_SL U56931 ( .A1(dwb_dat_i[21]), .A2(n61548), .B1(n75569), 
        .B2(dwb_dat_i[29]), .Y(n61081) );
  OAI21xp33_ASAP7_75t_SL U56932 ( .A1(n76765), .A2(n75586), .B(n61879), .Y(
        n61889) );
  AOI21xp33_ASAP7_75t_SL U56933 ( .A1(n72161), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .B(
        n71904), .Y(n71905) );
  INVx1_ASAP7_75t_SL U56934 ( .A(n65887), .Y(n65973) );
  NAND2xp5_ASAP7_75t_SL U56935 ( .A(n75000), .B(n74999), .Y(n75011) );
  NAND2xp33_ASAP7_75t_SL U56936 ( .A(n66021), .B(n65978), .Y(n65737) );
  AOI22xp33_ASAP7_75t_SL U56937 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_), .B2(n70018), .Y(
        n69460) );
  INVx1_ASAP7_75t_SL U56938 ( .A(n75575), .Y(n76761) );
  OAI21xp33_ASAP7_75t_SL U56939 ( .A1(n70598), .A2(n70211), .B(n70212), .Y(
        n70244) );
  NAND2xp33_ASAP7_75t_SL U56940 ( .A(n77875), .B(n57114), .Y(n75401) );
  INVxp33_ASAP7_75t_SL U56941 ( .A(n73027), .Y(n72921) );
  NAND2xp5_ASAP7_75t_SL U56942 ( .A(n63525), .B(n63430), .Y(n63439) );
  AOI22xp33_ASAP7_75t_SL U56943 ( .A1(n62279), .A2(n75844), .B1(n61439), .B2(
        n76760), .Y(n61440) );
  AOI21xp33_ASAP7_75t_SL U56944 ( .A1(n76975), .A2(n76974), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_nan), .Y(n76980) );
  OAI22xp33_ASAP7_75t_SL U56945 ( .A1(n66107), .A2(n66144), .B1(n66104), .B2(
        n66105), .Y(n65522) );
  NOR2xp33_ASAP7_75t_SRAM U56946 ( .A(or1200_cpu_or1200_except_n512), .B(
        n76724), .Y(n62413) );
  AOI22xp33_ASAP7_75t_SL U56947 ( .A1(n66022), .A2(n66023), .B1(n66024), .B2(
        n66079), .Y(n65738) );
  OAI22xp33_ASAP7_75t_SL U56948 ( .A1(n75574), .A2(n77102), .B1(n77100), .B2(
        n77101), .Y(n61709) );
  INVxp33_ASAP7_75t_SL U56949 ( .A(n65244), .Y(n65243) );
  NAND2xp5_ASAP7_75t_SL U56950 ( .A(n65729), .B(n65728), .Y(n66026) );
  INVxp67_ASAP7_75t_SL U56951 ( .A(n64931), .Y(n59290) );
  AOI22xp33_ASAP7_75t_SL U56952 ( .A1(n75570), .A2(
        or1200_dc_top_from_dcram_22_), .B1(dwb_dat_i[22]), .B2(n75569), .Y(
        n62252) );
  AOI22xp33_ASAP7_75t_SL U56953 ( .A1(n62273), .A2(n62278), .B1(n62262), .B2(
        n64294), .Y(n61766) );
  OAI22xp33_ASAP7_75t_SL U56954 ( .A1(n75729), .A2(n77101), .B1(
        or1200_cpu_or1200_mult_mac_n193), .B2(n74606), .Y(n64849) );
  NAND2xp5_ASAP7_75t_SL U56955 ( .A(n66089), .B(n65654), .Y(n65651) );
  INVxp67_ASAP7_75t_SL U56956 ( .A(n72907), .Y(n72741) );
  AOI21xp5_ASAP7_75t_SL U56957 ( .A1(n74246), .A2(n72593), .B(n72592), .Y(
        n74727) );
  OA21x2_ASAP7_75t_SL U56958 ( .A1(n77094), .A2(n77093), .B(n77092), .Y(n77095) );
  NAND2xp33_ASAP7_75t_SL U56959 ( .A(n69489), .B(n69488), .Y(n69491) );
  OAI22xp33_ASAP7_75t_SL U56960 ( .A1(n63418), .A2(n76897), .B1(n76508), .B2(
        n68787), .Y(n63419) );
  INVxp67_ASAP7_75t_SL U56961 ( .A(n61684), .Y(n61686) );
  OAI21xp33_ASAP7_75t_SL U56962 ( .A1(or1200_cpu_or1200_mult_mac_n247), .A2(
        n74587), .B(n62098), .Y(n62099) );
  AOI21xp5_ASAP7_75t_SL U56963 ( .A1(n64294), .A2(n64293), .B(n64292), .Y(
        n64299) );
  AOI21xp33_ASAP7_75t_SL U56964 ( .A1(n72393), .A2(n72233), .B(n72232), .Y(
        n72240) );
  AOI22xp33_ASAP7_75t_SL U56965 ( .A1(n73028), .A2(n72912), .B1(n73030), .B2(
        n72893), .Y(n72795) );
  AOI22xp33_ASAP7_75t_SL U56966 ( .A1(n61425), .A2(n75322), .B1(n76749), .B2(
        n60632), .Y(n60633) );
  AOI22xp33_ASAP7_75t_SL U56967 ( .A1(n66024), .A2(n66008), .B1(n66022), .B2(
        n65995), .Y(n65846) );
  NAND2xp33_ASAP7_75t_SL U56968 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_), .B(n70109), .Y(
        n69478) );
  AOI22xp33_ASAP7_75t_SL U56969 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_18_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_17_), .B2(n70018), .Y(
        n69468) );
  OAI21xp33_ASAP7_75t_SL U56970 ( .A1(n69961), .A2(n69960), .B(n69959), .Y(
        n69962) );
  AOI22xp33_ASAP7_75t_SL U56971 ( .A1(dwb_dat_i[16]), .A2(n61548), .B1(n75569), 
        .B2(dwb_dat_i[24]), .Y(n60586) );
  AOI22xp33_ASAP7_75t_SL U56972 ( .A1(n66024), .A2(n66047), .B1(n66022), .B2(
        n66016), .Y(n65766) );
  OAI22xp33_ASAP7_75t_SL U56973 ( .A1(n75729), .A2(n75574), .B1(n77101), .B2(
        n64834), .Y(n64310) );
  OAI22xp33_ASAP7_75t_SL U56974 ( .A1(n62531), .A2(n61417), .B1(n64113), .B2(
        n61416), .Y(n61432) );
  INVxp67_ASAP7_75t_SL U56975 ( .A(n72183), .Y(n72185) );
  INVxp67_ASAP7_75t_SL U56976 ( .A(n62275), .Y(n61635) );
  OAI22xp33_ASAP7_75t_SL U56977 ( .A1(n77104), .A2(n77103), .B1(n77102), .B2(
        n77101), .Y(n77110) );
  OAI21xp5_ASAP7_75t_SL U56978 ( .A1(n68825), .A2(n74999), .B(n68824), .Y(
        n68891) );
  AOI22xp33_ASAP7_75t_SL U56979 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_4_), .A2(n70019), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_3_), .B2(n70018), .Y(
        n69448) );
  OAI22xp33_ASAP7_75t_SL U56980 ( .A1(n62525), .A2(n77093), .B1(n77099), .B2(
        n62426), .Y(n62438) );
  NAND2xp33_ASAP7_75t_SL U56981 ( .A(n61075), .B(n61078), .Y(n61076) );
  NAND2xp33_ASAP7_75t_SL U56982 ( .A(n59687), .B(n77979), .Y(n3914) );
  INVxp33_ASAP7_75t_SL U56983 ( .A(n75880), .Y(n64250) );
  INVx1_ASAP7_75t_SL U56984 ( .A(n72658), .Y(n72661) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U56985 ( .A1(n65553), .A2(n65552), .B(n65551), 
        .C(n65550), .Y(n65554) );
  AOI21xp33_ASAP7_75t_SL U56986 ( .A1(n72459), .A2(n72412), .B(n72377), .Y(
        n72184) );
  NAND2xp33_ASAP7_75t_SL U56987 ( .A(n59687), .B(n77982), .Y(n3912) );
  AOI22xp33_ASAP7_75t_SL U56988 ( .A1(n75570), .A2(
        or1200_dc_top_from_dcram_23_), .B1(dwb_dat_i[23]), .B2(n75569), .Y(
        n75572) );
  INVxp33_ASAP7_75t_SL U56989 ( .A(n61703), .Y(n61705) );
  NAND2xp33_ASAP7_75t_SL U56990 ( .A(n61079), .B(n61078), .Y(n61080) );
  OAI22xp33_ASAP7_75t_SL U56991 ( .A1(n64113), .A2(n75574), .B1(n62531), .B2(
        n77101), .Y(n62441) );
  INVx1_ASAP7_75t_SL U56992 ( .A(n69182), .Y(n76903) );
  OAI22xp33_ASAP7_75t_SL U56993 ( .A1(n76897), .A2(n63471), .B1(n77637), .B2(
        n68787), .Y(n63472) );
  NAND2xp33_ASAP7_75t_SL U56994 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_), .B(n70109), .Y(
        n69447) );
  AOI21xp33_ASAP7_75t_SL U56995 ( .A1(n72192), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .B(
        n72377), .Y(n72193) );
  OAI22xp33_ASAP7_75t_SL U56996 ( .A1(n66102), .A2(n66156), .B1(n66108), .B2(
        n66147), .Y(n65520) );
  OAI22xp33_ASAP7_75t_SL U56997 ( .A1(n64131), .A2(n77107), .B1(n64132), .B2(
        n77105), .Y(n62440) );
  AOI22xp33_ASAP7_75t_SL U56998 ( .A1(or1200_dc_top_from_dcram_19_), .A2(
        n58285), .B1(n75570), .B2(or1200_dc_top_from_dcram_27_), .Y(n61545) );
  AOI21xp33_ASAP7_75t_SL U56999 ( .A1(n74168), .A2(n74209), .B(n74752), .Y(
        n74175) );
  NAND2xp33_ASAP7_75t_SL U57000 ( .A(n77883), .B(n57114), .Y(n63919) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57001 ( .A1(n65691), .A2(n65586), .B(n65585), .C(
        n65639), .Y(n65608) );
  OAI21xp33_ASAP7_75t_SL U57002 ( .A1(n59577), .A2(n75338), .B(n62117), .Y(
        n62118) );
  INVx1_ASAP7_75t_SL U57003 ( .A(n66113), .Y(n66153) );
  AOI21xp33_ASAP7_75t_SL U57004 ( .A1(n72242), .A2(n72376), .B(n72020), .Y(
        n72032) );
  AOI22xp33_ASAP7_75t_SL U57005 ( .A1(or1200_dc_top_from_dcram_18_), .A2(
        n58285), .B1(n75570), .B2(or1200_dc_top_from_dcram_26_), .Y(n61178) );
  INVxp33_ASAP7_75t_SL U57006 ( .A(n74619), .Y(n61704) );
  INVx1_ASAP7_75t_SL U57007 ( .A(n66111), .Y(n66164) );
  OAI22xp33_ASAP7_75t_SL U57008 ( .A1(n75233), .A2(n75574), .B1(n75346), .B2(
        n77101), .Y(n62125) );
  INVxp67_ASAP7_75t_SL U57009 ( .A(n62341), .Y(n60592) );
  NAND2xp33_ASAP7_75t_SL U57010 ( .A(n77877), .B(n57114), .Y(n62159) );
  OAI21xp33_ASAP7_75t_SL U57011 ( .A1(n69832), .A2(n69831), .B(n69830), .Y(
        n69833) );
  INVxp33_ASAP7_75t_SL U57012 ( .A(n65659), .Y(n65465) );
  NAND2xp5_ASAP7_75t_SL U57013 ( .A(n77777), .B(n77776), .Y(n9342) );
  OAI22xp33_ASAP7_75t_SL U57014 ( .A1(n62123), .A2(n75587), .B1(n75240), .B2(
        n77103), .Y(n62124) );
  OAI21xp33_ASAP7_75t_SL U57015 ( .A1(n65816), .A2(n66007), .B(n65815), .Y(
        n66039) );
  NAND2xp33_ASAP7_75t_SL U57016 ( .A(n77293), .B(n77292), .Y(n78160) );
  INVxp33_ASAP7_75t_SL U57017 ( .A(n61945), .Y(n61927) );
  NAND2xp5_ASAP7_75t_SL U57018 ( .A(n61535), .B(n61534), .Y(n61536) );
  INVxp67_ASAP7_75t_SL U57019 ( .A(n72630), .Y(n72616) );
  AOI22xp33_ASAP7_75t_SL U57020 ( .A1(dwb_dat_i[18]), .A2(n61548), .B1(n75569), 
        .B2(dwb_dat_i[26]), .Y(n61179) );
  NAND2xp33_ASAP7_75t_SL U57021 ( .A(n73028), .B(n72911), .Y(n72789) );
  AOI22xp33_ASAP7_75t_SL U57022 ( .A1(n78002), .A2(n59654), .B1(n62660), .B2(
        n62659), .Y(n62662) );
  AOI31xp33_ASAP7_75t_SRAM U57023 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_6_), .A2(
        n71714), .A3(n71713), .B(n71712), .Y(n71715) );
  AOI21xp33_ASAP7_75t_SL U57024 ( .A1(n72498), .A2(n72131), .B(n72013), .Y(
        n72014) );
  AOI21xp33_ASAP7_75t_SL U57025 ( .A1(n72335), .A2(n72131), .B(n71996), .Y(
        n71997) );
  OAI22xp33_ASAP7_75t_SL U57026 ( .A1(n65518), .A2(n66160), .B1(n66103), .B2(
        n66158), .Y(n65519) );
  AOI22xp33_ASAP7_75t_SL U57027 ( .A1(n75570), .A2(
        or1200_dc_top_from_dcram_18_), .B1(dwb_dat_i[18]), .B2(n75569), .Y(
        n63595) );
  AOI21xp33_ASAP7_75t_SL U57028 ( .A1(n72513), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .B(
        n72377), .Y(n72378) );
  INVxp67_ASAP7_75t_SL U57029 ( .A(n76727), .Y(n76730) );
  INVx1_ASAP7_75t_SL U57030 ( .A(n77078), .Y(n75584) );
  NAND2xp5_ASAP7_75t_SL U57031 ( .A(n71731), .B(n71730), .Y(n71737) );
  OAI21xp33_ASAP7_75t_SL U57032 ( .A1(n73537), .A2(n73536), .B(n73544), .Y(
        n73539) );
  AOI21xp33_ASAP7_75t_SL U57033 ( .A1(n70119), .A2(n70118), .B(n70139), .Y(
        n70121) );
  OAI21xp5_ASAP7_75t_SL U57034 ( .A1(n73942), .A2(n73941), .B(n73940), .Y(
        n73943) );
  NAND2xp33_ASAP7_75t_SL U57035 ( .A(n65942), .B(n65978), .Y(n65845) );
  NAND2xp33_ASAP7_75t_SL U57036 ( .A(n66114), .B(n66113), .Y(n66132) );
  AOI21xp33_ASAP7_75t_SL U57037 ( .A1(n74956), .A2(n791), .B(n60147), .Y(
        n60066) );
  INVxp33_ASAP7_75t_SL U57038 ( .A(n69973), .Y(n69979) );
  OAI22xp33_ASAP7_75t_SL U57039 ( .A1(n74608), .A2(n74607), .B1(n77106), .B2(
        n77107), .Y(n74612) );
  OAI21xp33_ASAP7_75t_SL U57040 ( .A1(n77104), .A2(n77093), .B(n74610), .Y(
        n74611) );
  OAI22xp33_ASAP7_75t_SL U57041 ( .A1(n75590), .A2(n77103), .B1(n77102), .B2(
        n75587), .Y(n74616) );
  OAI21xp33_ASAP7_75t_SL U57042 ( .A1(n66158), .A2(n66128), .B(n66127), .Y(
        n66129) );
  OAI22xp33_ASAP7_75t_SL U57043 ( .A1(n77108), .A2(n75574), .B1(n75588), .B2(
        n77101), .Y(n74615) );
  OAI22xp33_ASAP7_75t_SL U57044 ( .A1(n66121), .A2(n66160), .B1(n66120), .B2(
        n66147), .Y(n66130) );
  BUFx6f_ASAP7_75t_SL U57045 ( .A(n59610), .Y(n57181) );
  NOR2x1_ASAP7_75t_SL U57046 ( .A(n61229), .B(n61228), .Y(n62288) );
  OAI21xp33_ASAP7_75t_SL U57047 ( .A1(n72645), .A2(n1859), .B(n72617), .Y(
        n72634) );
  NAND2xp33_ASAP7_75t_SL U57048 ( .A(n65886), .B(n65978), .Y(n65718) );
  INVxp67_ASAP7_75t_SL U57049 ( .A(n76724), .Y(n63557) );
  AOI22xp33_ASAP7_75t_SL U57050 ( .A1(n62213), .A2(n75387), .B1(n77920), .B2(
        n75649), .Y(n62214) );
  INVxp33_ASAP7_75t_SL U57051 ( .A(n75397), .Y(n62215) );
  OAI22xp33_ASAP7_75t_SL U57052 ( .A1(n75346), .A2(n61645), .B1(n61644), .B2(
        n62332), .Y(n61657) );
  NAND2xp33_ASAP7_75t_SL U57053 ( .A(n74850), .B(n74855), .Y(n74877) );
  AOI21xp33_ASAP7_75t_SL U57054 ( .A1(n72412), .A2(n72287), .B(n72410), .Y(
        n72288) );
  OAI22xp33_ASAP7_75t_SL U57055 ( .A1(n73008), .A2(n72916), .B1(n72859), .B2(
        n72937), .Y(n72770) );
  AOI21xp33_ASAP7_75t_SL U57056 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .A2(
        n72440), .B(n72172), .Y(n72159) );
  AOI21xp33_ASAP7_75t_SL U57057 ( .A1(n72412), .A2(n72390), .B(n72410), .Y(
        n72395) );
  AOI22xp33_ASAP7_75t_SL U57058 ( .A1(n73024), .A2(n72917), .B1(n73026), .B2(
        n72935), .Y(n72822) );
  OAI22xp33_ASAP7_75t_SL U57059 ( .A1(n61639), .A2(n75574), .B1(n62123), .B2(
        n77105), .Y(n61640) );
  OAI22xp33_ASAP7_75t_SL U57060 ( .A1(n66027), .A2(n65928), .B1(n65972), .B2(
        n66081), .Y(n65797) );
  AOI21xp33_ASAP7_75t_SL U57061 ( .A1(n78223), .A2(n72667), .B(n72652), .Y(
        n72671) );
  NAND2xp33_ASAP7_75t_SL U57062 ( .A(n62230), .B(n75030), .Y(n62232) );
  INVx1_ASAP7_75t_SL U57063 ( .A(n61450), .Y(n77595) );
  OAI22xp33_ASAP7_75t_SL U57064 ( .A1(n63565), .A2(n75315), .B1(n75316), .B2(
        n63564), .Y(n63593) );
  OAI22xp33_ASAP7_75t_SL U57065 ( .A1(n77106), .A2(n75574), .B1(n75573), .B2(
        n77101), .Y(n75583) );
  INVxp67_ASAP7_75t_SL U57066 ( .A(n61385), .Y(n61387) );
  NAND2xp33_ASAP7_75t_SL U57067 ( .A(n74884), .B(n74855), .Y(n74883) );
  OAI21xp33_ASAP7_75t_SL U57068 ( .A1(n63576), .A2(n63575), .B(n75332), .Y(
        n63581) );
  INVxp33_ASAP7_75t_SL U57069 ( .A(n75574), .Y(n62345) );
  OAI21xp33_ASAP7_75t_SL U57070 ( .A1(or1200_cpu_or1200_except_n544), .A2(
        n76724), .B(n75824), .Y(n75825) );
  NAND2xp33_ASAP7_75t_SL U57071 ( .A(n62485), .B(n75030), .Y(n62487) );
  AOI21xp33_ASAP7_75t_SL U57072 ( .A1(n63579), .A2(n63892), .B(n63578), .Y(
        n63580) );
  AOI21xp33_ASAP7_75t_SL U57073 ( .A1(n72412), .A2(n72273), .B(n72272), .Y(
        n72277) );
  OAI22xp33_ASAP7_75t_SL U57074 ( .A1(n65974), .A2(n65920), .B1(n66027), .B2(
        n65969), .Y(n65688) );
  NAND2xp33_ASAP7_75t_SL U57075 ( .A(n77885), .B(n57114), .Y(n74980) );
  OAI22xp33_ASAP7_75t_SL U57076 ( .A1(n64113), .A2(n75587), .B1(n75871), .B2(
        n77103), .Y(n64118) );
  INVx1_ASAP7_75t_SL U57077 ( .A(n75268), .Y(n75271) );
  NAND2xp33_ASAP7_75t_SL U57078 ( .A(n77880), .B(n75015), .Y(n64178) );
  AOI22xp33_ASAP7_75t_SL U57079 ( .A1(or1200_dc_top_from_dcram_16_), .A2(
        n58285), .B1(n75570), .B2(or1200_dc_top_from_dcram_24_), .Y(n60585) );
  INVxp33_ASAP7_75t_SL U57080 ( .A(n64097), .Y(n61824) );
  INVxp33_ASAP7_75t_SL U57081 ( .A(n63565), .Y(n61791) );
  INVxp33_ASAP7_75t_SL U57082 ( .A(n63563), .Y(n61823) );
  OAI21xp33_ASAP7_75t_SL U57083 ( .A1(n70006), .A2(n70005), .B(n70004), .Y(
        n70007) );
  NAND2xp5_ASAP7_75t_SL U57084 ( .A(n70232), .B(n70224), .Y(n70235) );
  OAI21xp33_ASAP7_75t_SL U57085 ( .A1(or1200_cpu_or1200_mult_mac_n331), .A2(
        n75738), .B(n64306), .Y(n64307) );
  OAI22xp33_ASAP7_75t_SL U57086 ( .A1(n64132), .A2(n75574), .B1(n64131), .B2(
        n77101), .Y(n64133) );
  AOI22xp33_ASAP7_75t_SL U57087 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[19]), .A2(n71013), 
        .B1(n58291), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[20]), .Y(n71012) );
  NAND2xp33_ASAP7_75t_SL U57088 ( .A(n77888), .B(n57114), .Y(n75296) );
  OAI22xp33_ASAP7_75t_SL U57089 ( .A1(n77108), .A2(n77105), .B1(n76759), .B2(
        n75587), .Y(n61708) );
  OAI22xp33_ASAP7_75t_SL U57090 ( .A1(n62422), .A2(n61703), .B1(n77592), .B2(
        n76796), .Y(n61557) );
  NOR2xp33_ASAP7_75t_SRAM U57091 ( .A(n70006), .B(n70004), .Y(n70014) );
  AOI22xp33_ASAP7_75t_SL U57092 ( .A1(n73026), .A2(n72891), .B1(n73024), .B2(
        n72916), .Y(n72796) );
  INVxp67_ASAP7_75t_SL U57093 ( .A(n65965), .Y(n65916) );
  NAND2xp33_ASAP7_75t_SL U57094 ( .A(n70112), .B(n70109), .Y(n69496) );
  AOI21xp33_ASAP7_75t_SL U57095 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .A2(
        n72322), .B(n72172), .Y(n72173) );
  OAI22xp33_ASAP7_75t_SL U57096 ( .A1(n77108), .A2(n77107), .B1(n77106), .B2(
        n77105), .Y(n77109) );
  NAND2xp33_ASAP7_75t_SL U57097 ( .A(n77871), .B(n57114), .Y(n74040) );
  AOI21xp33_ASAP7_75t_SL U57098 ( .A1(n78374), .A2(n72667), .B(n72623), .Y(
        n72624) );
  INVxp33_ASAP7_75t_SL U57099 ( .A(n77103), .Y(n61782) );
  OAI22xp33_ASAP7_75t_SL U57100 ( .A1(n78336), .A2(n70035), .B1(n78338), .B2(
        n70034), .Y(n69559) );
  AOI22xp33_ASAP7_75t_SL U57101 ( .A1(n76766), .A2(n75862), .B1(n75861), .B2(
        n75860), .Y(n75864) );
  OAI22xp33_ASAP7_75t_SL U57102 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), 
        .A2(n72904), .B1(n72993), .B2(n72901), .Y(n72727) );
  INVxp67_ASAP7_75t_SL U57103 ( .A(n61409), .Y(n61415) );
  INVx1_ASAP7_75t_SL U57104 ( .A(n72938), .Y(n72917) );
  INVx1_ASAP7_75t_SL U57105 ( .A(n62096), .Y(n75361) );
  AOI22xp33_ASAP7_75t_SL U57106 ( .A1(n73026), .A2(n72937), .B1(n73024), .B2(
        n72923), .Y(n72845) );
  INVxp67_ASAP7_75t_SL U57107 ( .A(n61106), .Y(n73941) );
  NAND2xp5_ASAP7_75t_SL U57108 ( .A(n63773), .B(n63772), .Y(n63771) );
  OAI22xp33_ASAP7_75t_SL U57109 ( .A1(n78338), .A2(n70035), .B1(n78340), .B2(
        n70034), .Y(n69796) );
  INVx1_ASAP7_75t_SL U57110 ( .A(n66022), .Y(n65970) );
  AOI21xp33_ASAP7_75t_SL U57111 ( .A1(n77039), .A2(n74584), .B(n74583), .Y(
        n74585) );
  NAND2xp33_ASAP7_75t_SL U57112 ( .A(n70073), .B(n70072), .Y(n70074) );
  OAI21xp5_ASAP7_75t_SL U57113 ( .A1(n77260), .A2(n60164), .B(n60163), .Y(
        n60165) );
  AND2x2_ASAP7_75t_SL U57114 ( .A(n72474), .B(n72511), .Y(n72375) );
  AOI21xp33_ASAP7_75t_SL U57115 ( .A1(n75847), .A2(n77701), .B(n75228), .Y(
        n75229) );
  NAND2xp5_ASAP7_75t_SL U57116 ( .A(n70453), .B(n70452), .Y(n2380) );
  OAI22xp33_ASAP7_75t_SL U57117 ( .A1(n1755), .A2(n61226), .B1(n1757), .B2(
        n76717), .Y(n77589) );
  O2A1O1Ixp33_ASAP7_75t_SL U57118 ( .A1(n61408), .A2(n61523), .B(n62761), .C(
        n61407), .Y(n61444) );
  INVxp67_ASAP7_75t_SL U57119 ( .A(n60566), .Y(n60568) );
  OAI21xp33_ASAP7_75t_SL U57120 ( .A1(n72383), .A2(n72382), .B(n72381), .Y(
        n72386) );
  INVxp67_ASAP7_75t_SL U57121 ( .A(n72381), .Y(n72377) );
  AOI21xp33_ASAP7_75t_SL U57122 ( .A1(n70002), .A2(n70048), .B(n69706), .Y(
        n69709) );
  AOI21xp33_ASAP7_75t_SL U57123 ( .A1(n76767), .A2(n77062), .B(n73924), .Y(
        n73926) );
  OAI22xp33_ASAP7_75t_SL U57124 ( .A1(n72495), .A2(n72473), .B1(n72546), .B2(
        n72471), .Y(n72217) );
  AOI21xp33_ASAP7_75t_SL U57125 ( .A1(n77070), .A2(n77705), .B(n77069), .Y(
        n77071) );
  OAI21xp33_ASAP7_75t_SL U57126 ( .A1(n74379), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_7_), .B(
        n74378), .Y(n2349) );
  AOI22xp33_ASAP7_75t_SL U57127 ( .A1(n75247), .A2(n77061), .B1(n75246), .B2(
        n75245), .Y(n75248) );
  AOI21xp5_ASAP7_75t_SL U57128 ( .A1(n64168), .A2(n65077), .B(n65075), .Y(
        n64176) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57129 ( .A1(n59575), .A2(n59549), .B(n75852), .C(
        n75589), .Y(n75249) );
  INVx1_ASAP7_75t_SL U57130 ( .A(n68787), .Y(n76888) );
  INVxp33_ASAP7_75t_SL U57131 ( .A(n61622), .Y(n61623) );
  NAND2xp5_ASAP7_75t_SL U57132 ( .A(n77429), .B(n77428), .Y(n77438) );
  AOI31xp33_ASAP7_75t_SRAM U57133 ( .A1(n65543), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .A3(n65758), 
        .B(n65437), .Y(n65438) );
  NAND2xp5_ASAP7_75t_SL U57134 ( .A(n63413), .B(n63412), .Y(n63414) );
  NOR2xp33_ASAP7_75t_SL U57135 ( .A(n60761), .B(n60760), .Y(n60762) );
  AOI21xp33_ASAP7_75t_SL U57136 ( .A1(n70302), .A2(n70387), .B(n70254), .Y(
        n2316) );
  INVxp33_ASAP7_75t_SL U57137 ( .A(n77089), .Y(n77094) );
  NAND2xp33_ASAP7_75t_SL U57138 ( .A(n74956), .B(n60124), .Y(n60132) );
  INVxp33_ASAP7_75t_SL U57139 ( .A(n66090), .Y(n65649) );
  OAI21xp33_ASAP7_75t_SL U57140 ( .A1(n74093), .A2(n74205), .B(n74092), .Y(
        n74094) );
  OAI21xp33_ASAP7_75t_SL U57141 ( .A1(n75729), .A2(n77099), .B(n75728), .Y(
        n75730) );
  NAND2xp5_ASAP7_75t_SL U57142 ( .A(n65552), .B(n65543), .Y(n65466) );
  INVxp33_ASAP7_75t_SL U57143 ( .A(n61511), .Y(n61424) );
  OAI22xp33_ASAP7_75t_SL U57144 ( .A1(dwb_dat_i[0]), .A2(n61547), .B1(
        or1200_dc_top_from_dcram_0_), .B2(n61546), .Y(n62341) );
  OAI21xp33_ASAP7_75t_SL U57145 ( .A1(n74138), .A2(n74205), .B(n74162), .Y(
        n66214) );
  INVxp33_ASAP7_75t_SL U57146 ( .A(n61494), .Y(n61416) );
  INVx1_ASAP7_75t_SL U57147 ( .A(n72992), .Y(n73023) );
  NAND2xp5_ASAP7_75t_SL U57148 ( .A(n60856), .B(n76772), .Y(n61346) );
  OAI21xp33_ASAP7_75t_SL U57149 ( .A1(n72544), .A2(n72335), .B(n72381), .Y(
        n72232) );
  AOI22xp33_ASAP7_75t_SL U57150 ( .A1(n72474), .A2(n72336), .B1(n72412), .B2(
        n72238), .Y(n72239) );
  INVxp67_ASAP7_75t_SL U57151 ( .A(n69757), .Y(n69749) );
  NAND2xp5_ASAP7_75t_SL U57152 ( .A(n61814), .B(n61813), .Y(n75815) );
  OAI21xp33_ASAP7_75t_SL U57153 ( .A1(n72064), .A2(n72106), .B(n71781), .Y(
        n71782) );
  INVxp33_ASAP7_75t_SL U57154 ( .A(n71675), .Y(n71638) );
  OAI21xp33_ASAP7_75t_SL U57155 ( .A1(n63428), .A2(n63404), .B(n63412), .Y(
        n63405) );
  OAI22xp33_ASAP7_75t_SL U57156 ( .A1(n78334), .A2(n70035), .B1(n78336), .B2(
        n70034), .Y(n69778) );
  OAI21xp33_ASAP7_75t_SL U57157 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[24]), .A2(
        n58284), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[24]), .Y(
        n73117) );
  OAI21xp5_ASAP7_75t_SL U57158 ( .A1(n72399), .A2(n72202), .B(n72082), .Y(
        n72396) );
  AOI22xp33_ASAP7_75t_SL U57159 ( .A1(n62360), .A2(n64127), .B1(n62359), .B2(
        n62518), .Y(n64773) );
  INVxp33_ASAP7_75t_SL U57160 ( .A(n70005), .Y(n69986) );
  NAND2xp5_ASAP7_75t_SL U57161 ( .A(n61818), .B(n61817), .Y(n64754) );
  NAND2xp5_ASAP7_75t_SL U57162 ( .A(n61820), .B(n61819), .Y(n75567) );
  OAI21xp33_ASAP7_75t_SL U57163 ( .A1(n72354), .A2(n72106), .B(n72052), .Y(
        n72053) );
  NAND2xp33_ASAP7_75t_SL U57164 ( .A(n65695), .B(n65694), .Y(n65696) );
  INVxp33_ASAP7_75t_SL U57165 ( .A(n73944), .Y(n73936) );
  OAI21xp5_ASAP7_75t_SL U57166 ( .A1(or1200_cpu_or1200_mult_mac_n88), .A2(
        n61826), .B(n61821), .Y(n64097) );
  INVx1_ASAP7_75t_SL U57167 ( .A(n62110), .Y(n75244) );
  INVx1_ASAP7_75t_SL U57168 ( .A(n70073), .Y(n70090) );
  INVx1_ASAP7_75t_SL U57169 ( .A(n61556), .Y(n77592) );
  INVx1_ASAP7_75t_SL U57170 ( .A(n65570), .Y(n66144) );
  OAI22xp33_ASAP7_75t_SL U57171 ( .A1(n1719), .A2(n61226), .B1(n1721), .B2(
        n76717), .Y(n77582) );
  OAI21xp33_ASAP7_75t_SL U57172 ( .A1(n62270), .A2(n62332), .B(n62269), .Y(
        n62271) );
  AOI21xp33_ASAP7_75t_SL U57173 ( .A1(n75852), .A2(n63584), .B(n77070), .Y(
        n63586) );
  INVxp67_ASAP7_75t_SL U57174 ( .A(n65945), .Y(n65864) );
  NAND2xp33_ASAP7_75t_SL U57175 ( .A(n61486), .B(n61445), .Y(n60808) );
  NAND2xp33_ASAP7_75t_SL U57176 ( .A(n73024), .B(n72893), .Y(n72766) );
  OAI22xp33_ASAP7_75t_SL U57177 ( .A1(dwb_dat_i[1]), .A2(n61547), .B1(
        or1200_dc_top_from_dcram_1_), .B2(n61546), .Y(n75314) );
  NAND2xp33_ASAP7_75t_SL U57178 ( .A(n77883), .B(n75649), .Y(n63916) );
  NAND2xp33_ASAP7_75t_SL U57179 ( .A(n61658), .B(n61494), .Y(n60941) );
  AOI22xp33_ASAP7_75t_SL U57180 ( .A1(dwb_dat_i[4]), .A2(n61546), .B1(
        or1200_dc_top_from_dcram_4_), .B2(n61547), .Y(n64121) );
  OAI22xp33_ASAP7_75t_SL U57181 ( .A1(n78344), .A2(n70035), .B1(n78348), .B2(
        n70034), .Y(n69844) );
  AOI22xp33_ASAP7_75t_SL U57182 ( .A1(dwb_dat_i[9]), .A2(n61546), .B1(
        or1200_dc_top_from_dcram_9_), .B2(n61547), .Y(n75317) );
  AOI21xp33_ASAP7_75t_SL U57183 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_), .A2(n59627), .B(
        n72612), .Y(n78358) );
  INVx1_ASAP7_75t_SL U57184 ( .A(n61990), .Y(n61316) );
  OAI21xp5_ASAP7_75t_SL U57185 ( .A1(n65818), .A2(n65703), .B(n65702), .Y(
        n65967) );
  NAND2xp33_ASAP7_75t_SL U57186 ( .A(n76779), .B(n61353), .Y(n60938) );
  AOI22xp33_ASAP7_75t_SL U57187 ( .A1(n77075), .A2(n61511), .B1(n76763), .B2(
        n76771), .Y(n61512) );
  O2A1O1Ixp33_ASAP7_75t_SL U57188 ( .A1(n71673), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_8_), .B(
        n71675), .C(n71672), .Y(n71674) );
  NOR2xp33_ASAP7_75t_SRAM U57189 ( .A(n74927), .B(n77356), .Y(n74928) );
  OAI22xp33_ASAP7_75t_SL U57190 ( .A1(n78348), .A2(n70035), .B1(n78346), .B2(
        n70034), .Y(n69845) );
  NAND2xp33_ASAP7_75t_SL U57191 ( .A(n77871), .B(n75649), .Y(n66229) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57192 ( .A1(n75245), .A2(n62133), .B(n57126), .C(
        n61864), .Y(n61867) );
  OAI22xp33_ASAP7_75t_SL U57193 ( .A1(n77639), .A2(n77604), .B1(n77847), .B2(
        n77603), .Y(n77607) );
  INVxp67_ASAP7_75t_SL U57194 ( .A(n72416), .Y(n72431) );
  NAND2xp33_ASAP7_75t_SL U57195 ( .A(n77866), .B(n75649), .Y(n66236) );
  NOR2xp67_ASAP7_75t_SL U57196 ( .A(n68810), .B(n64275), .Y(n75015) );
  INVxp67_ASAP7_75t_SL U57197 ( .A(n72446), .Y(n72447) );
  OAI22xp33_ASAP7_75t_SL U57198 ( .A1(n78346), .A2(n70035), .B1(n78350), .B2(
        n70034), .Y(n69871) );
  INVxp33_ASAP7_75t_SL U57199 ( .A(n69885), .Y(n69656) );
  NAND2xp5_ASAP7_75t_SL U57200 ( .A(n69864), .B(n69644), .Y(n69862) );
  AOI21xp5_ASAP7_75t_SL U57201 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[13]), .A2(
        n59627), .B(n72740), .Y(n72907) );
  OAI22xp33_ASAP7_75t_SL U57202 ( .A1(n77639), .A2(n77616), .B1(n77847), .B2(
        n77615), .Y(n77617) );
  INVxp67_ASAP7_75t_SL U57203 ( .A(n77656), .Y(n77657) );
  NAND3xp33_ASAP7_75t_SRAM U57204 ( .A(n75576), .B(n64776), .C(n77242), .Y(
        n62530) );
  INVxp33_ASAP7_75t_SL U57205 ( .A(n62374), .Y(n61417) );
  OAI21xp33_ASAP7_75t_SL U57206 ( .A1(or1200_cpu_or1200_mult_mac_n315), .A2(
        n77073), .B(n60812), .Y(n60813) );
  INVxp33_ASAP7_75t_SL U57207 ( .A(n62332), .Y(n62338) );
  NAND2xp33_ASAP7_75t_SL U57208 ( .A(n65678), .B(n65677), .Y(n65679) );
  OAI21xp33_ASAP7_75t_SL U57209 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[18]), .A2(
        n58284), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[18]), .Y(
        n73314) );
  INVxp33_ASAP7_75t_SL U57210 ( .A(n70034), .Y(n69874) );
  INVxp33_ASAP7_75t_SL U57211 ( .A(n72426), .Y(n72427) );
  INVxp67_ASAP7_75t_SL U57212 ( .A(n69957), .Y(n69690) );
  INVxp67_ASAP7_75t_SL U57213 ( .A(n73551), .Y(n73543) );
  OAI22xp33_ASAP7_75t_SL U57214 ( .A1(n78340), .A2(n70035), .B1(n78342), .B2(
        n70034), .Y(n69814) );
  OAI22xp33_ASAP7_75t_SL U57215 ( .A1(n78329), .A2(n70035), .B1(n78330), .B2(
        n70034), .Y(n69732) );
  NAND2xp33_ASAP7_75t_SL U57216 ( .A(n77971), .B(n75649), .Y(n62406) );
  NOR2x1_ASAP7_75t_SL U57217 ( .A(n77759), .B(n61546), .Y(n75570) );
  NAND2xp5_ASAP7_75t_SL U57218 ( .A(dwb_dat_i[15]), .B(n61546), .Y(n60876) );
  NAND2xp5_ASAP7_75t_SL U57219 ( .A(dwb_dat_i[7]), .B(n61546), .Y(n60873) );
  INVxp33_ASAP7_75t_SL U57220 ( .A(n65385), .Y(n65309) );
  NOR2x1_ASAP7_75t_SL U57221 ( .A(n77759), .B(n61547), .Y(n75569) );
  INVxp67_ASAP7_75t_SL U57222 ( .A(n69933), .Y(n69675) );
  OAI21xp33_ASAP7_75t_SL U57223 ( .A1(n65808), .A2(n65807), .B(n65706), .Y(
        n65921) );
  NAND2xp33_ASAP7_75t_SL U57224 ( .A(n77922), .B(n75649), .Y(n62211) );
  BUFx2_ASAP7_75t_SL U57225 ( .A(n57118), .Y(n57271) );
  OAI22xp33_ASAP7_75t_SL U57226 ( .A1(n78342), .A2(n70035), .B1(n78344), .B2(
        n70034), .Y(n69826) );
  NAND2xp5_ASAP7_75t_SL U57227 ( .A(n65693), .B(n65692), .Y(n65964) );
  AOI21xp33_ASAP7_75t_SL U57228 ( .A1(n77041), .A2(n69188), .B(n63551), .Y(
        n63554) );
  NAND2xp33_ASAP7_75t_SL U57229 ( .A(n77918), .B(n75649), .Y(n62216) );
  INVx1_ASAP7_75t_SL U57230 ( .A(n75648), .Y(n75030) );
  NAND2xp33_ASAP7_75t_SL U57231 ( .A(n61622), .B(n62287), .Y(n60809) );
  OAI22xp33_ASAP7_75t_SL U57232 ( .A1(n59709), .A2(n77056), .B1(n59708), .B2(
        n77062), .Y(n75575) );
  NAND2xp33_ASAP7_75t_SL U57233 ( .A(n77974), .B(n75649), .Y(n62225) );
  AOI22xp33_ASAP7_75t_SL U57234 ( .A1(n72393), .A2(n72392), .B1(n72474), .B2(
        n72391), .Y(n72394) );
  NAND2xp33_ASAP7_75t_SL U57235 ( .A(n77977), .B(n75649), .Y(n62231) );
  OAI21xp5_ASAP7_75t_SL U57236 ( .A1(n68783), .A2(n68782), .B(n68781), .Y(
        n74999) );
  INVx1_ASAP7_75t_SL U57237 ( .A(n66116), .Y(n66156) );
  NAND2xp33_ASAP7_75t_SL U57238 ( .A(n77983), .B(n75649), .Y(n62306) );
  NAND2xp5_ASAP7_75t_SL U57239 ( .A(n72266), .B(n72426), .Y(n72476) );
  NAND2xp33_ASAP7_75t_SL U57240 ( .A(n77986), .B(n75649), .Y(n62395) );
  INVxp33_ASAP7_75t_SL U57241 ( .A(n73540), .Y(n73542) );
  AOI21xp33_ASAP7_75t_SL U57242 ( .A1(n72514), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .B(
        n71881), .Y(n72161) );
  AOI21xp33_ASAP7_75t_SL U57243 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[8]), .A2(n59627), .B(n72773), .Y(n72935) );
  NAND2xp33_ASAP7_75t_SL U57244 ( .A(n77901), .B(n75649), .Y(n62480) );
  NAND2xp33_ASAP7_75t_SL U57245 ( .A(n77899), .B(n75649), .Y(n62486) );
  INVx1_ASAP7_75t_SL U57246 ( .A(n63555), .Y(n75368) );
  NOR2x1_ASAP7_75t_SL U57247 ( .A(n57340), .B(n57339), .Y(n59292) );
  OAI21xp33_ASAP7_75t_SL U57248 ( .A1(n72286), .A2(n72382), .B(n72381), .Y(
        n72410) );
  INVxp33_ASAP7_75t_SL U57249 ( .A(n74606), .Y(n63579) );
  NAND2xp33_ASAP7_75t_SL U57250 ( .A(n77893), .B(n75649), .Y(n62494) );
  OAI22xp33_ASAP7_75t_SL U57251 ( .A1(n63577), .A2(n77099), .B1(
        or1200_cpu_or1200_mult_mac_n323), .B2(n75738), .Y(n63578) );
  AOI22xp5_ASAP7_75t_SL U57252 ( .A1(n77672), .A2(n77992), .B1(n77644), .B2(
        n77610), .Y(n77611) );
  NAND2xp33_ASAP7_75t_SL U57253 ( .A(n77890), .B(n75649), .Y(n62550) );
  INVxp67_ASAP7_75t_SL U57254 ( .A(n77626), .Y(n77627) );
  NAND2xp33_ASAP7_75t_SL U57255 ( .A(n77888), .B(n75649), .Y(n75388) );
  AOI22xp33_ASAP7_75t_SL U57256 ( .A1(dwb_dat_i[12]), .A2(n61546), .B1(
        or1200_dc_top_from_dcram_12_), .B2(n61547), .Y(n64136) );
  OAI22xp33_ASAP7_75t_SL U57257 ( .A1(n72107), .A2(n72269), .B1(n72411), .B2(
        n72106), .Y(n72130) );
  INVxp67_ASAP7_75t_SL U57258 ( .A(n72469), .Y(n72458) );
  INVxp33_ASAP7_75t_SL U57259 ( .A(n60935), .Y(n60632) );
  INVx1_ASAP7_75t_SL U57260 ( .A(n65901), .Y(n65962) );
  AOI22xp33_ASAP7_75t_SL U57261 ( .A1(n66117), .A2(n66116), .B1(n66115), .B2(
        n66162), .Y(n66118) );
  INVxp67_ASAP7_75t_SL U57262 ( .A(n70035), .Y(n70057) );
  AOI22xp33_ASAP7_75t_SL U57263 ( .A1(n72474), .A2(n72468), .B1(n72412), .B2(
        n72191), .Y(n72194) );
  INVxp33_ASAP7_75t_SL U57264 ( .A(n64217), .Y(n75347) );
  AOI22xp33_ASAP7_75t_SL U57265 ( .A1(dwb_dat_i[2]), .A2(n61546), .B1(
        or1200_dc_top_from_dcram_2_), .B2(n61547), .Y(n63565) );
  NOR2x1_ASAP7_75t_SL U57266 ( .A(n74354), .B(n74378), .Y(n74353) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57267 ( .A1(n66145), .A2(n65582), .B(n66114), .C(
        n65581), .Y(n65586) );
  AOI22xp33_ASAP7_75t_SL U57268 ( .A1(n64221), .A2(n64774), .B1(n64220), .B2(
        n64219), .Y(n64228) );
  NAND2xp5_ASAP7_75t_SL U57269 ( .A(n57126), .B(n62371), .Y(n77078) );
  INVxp67_ASAP7_75t_SL U57270 ( .A(n61643), .Y(n61644) );
  NAND2xp5_ASAP7_75t_SL U57271 ( .A(n71628), .B(n71587), .Y(n71569) );
  INVxp67_ASAP7_75t_SL U57272 ( .A(n62273), .Y(n61645) );
  NAND2xp5_ASAP7_75t_SL U57273 ( .A(n70211), .B(n70598), .Y(n70212) );
  INVxp67_ASAP7_75t_SL U57274 ( .A(n77060), .Y(n62447) );
  NAND2xp33_ASAP7_75t_SL U57275 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .B(
        n72938), .Y(n72873) );
  AOI22xp33_ASAP7_75t_SL U57276 ( .A1(n77061), .A2(n64223), .B1(n64222), .B2(
        n75591), .Y(n64227) );
  OAI21xp33_ASAP7_75t_SL U57277 ( .A1(n73009), .A2(n72901), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), .Y(
        n72756) );
  AOI21xp33_ASAP7_75t_SL U57278 ( .A1(n77039), .A2(n65090), .B(n62097), .Y(
        n62098) );
  AOI21xp33_ASAP7_75t_SL U57279 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_), .A2(n59627), .B(n72613), 
        .Y(n72630) );
  INVxp67_ASAP7_75t_SL U57280 ( .A(n62287), .Y(n76748) );
  NAND2xp33_ASAP7_75t_SL U57281 ( .A(n72993), .B(n72891), .Y(n72753) );
  NAND2xp5_ASAP7_75t_SL U57282 ( .A(n59387), .B(n60779), .Y(n60783) );
  OAI22xp33_ASAP7_75t_SL U57283 ( .A1(n76770), .A2(n64843), .B1(n75713), .B2(
        n76765), .Y(n64845) );
  INVxp33_ASAP7_75t_SL U57284 ( .A(n71681), .Y(n71736) );
  INVxp67_ASAP7_75t_SL U57285 ( .A(n63900), .Y(n63895) );
  NAND2xp33_ASAP7_75t_SL U57286 ( .A(n57083), .B(sbbiu_adr_sb[3]), .Y(n77776)
         );
  INVx1_ASAP7_75t_SL U57287 ( .A(n77099), .Y(n64294) );
  OAI22xp33_ASAP7_75t_SL U57288 ( .A1(dwb_dat_i[11]), .A2(n61547), .B1(
        or1200_dc_top_from_dcram_11_), .B2(n61546), .Y(n74619) );
  AOI22xp33_ASAP7_75t_SL U57289 ( .A1(n62366), .A2(n77076), .B1(n74776), .B2(
        n61410), .Y(n60682) );
  NAND2xp5_ASAP7_75t_SL U57290 ( .A(n68812), .B(n68811), .Y(n69182) );
  AOI21xp33_ASAP7_75t_SL U57291 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[14]), .A2(
        n59627), .B(n72722), .Y(n72890) );
  AOI21xp33_ASAP7_75t_SL U57292 ( .A1(n61630), .A2(n61533), .B(n61532), .Y(
        n61534) );
  INVxp67_ASAP7_75t_SL U57293 ( .A(n65932), .Y(n65956) );
  NAND2xp33_ASAP7_75t_SL U57294 ( .A(n59687), .B(n77973), .Y(n3918) );
  OAI22xp33_ASAP7_75t_SL U57295 ( .A1(dwb_dat_i[3]), .A2(n61547), .B1(
        or1200_dc_top_from_dcram_3_), .B2(n61546), .Y(n61703) );
  AOI21xp33_ASAP7_75t_SL U57296 ( .A1(n70302), .A2(n70269), .B(n70268), .Y(
        n2332) );
  OAI22xp33_ASAP7_75t_SL U57297 ( .A1(n72278), .A2(n72462), .B1(n72415), .B2(
        n72182), .Y(n72183) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U57298 ( .A1(n66117), .A2(n65597), .B(n65596), 
        .C(n65691), .Y(n65598) );
  AOI21xp5_ASAP7_75t_SL U57299 ( .A1(n74191), .A2(n74192), .B(n74151), .Y(
        n74168) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57300 ( .A1(n72393), .A2(n72137), .B(n71830), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .Y(
        n71831) );
  OAI21xp33_ASAP7_75t_SL U57301 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), .A2(n58571), 
        .B(n65685), .Y(n65920) );
  INVx1_ASAP7_75t_SL U57302 ( .A(n75736), .Y(n64830) );
  INVxp67_ASAP7_75t_SL U57303 ( .A(n71652), .Y(n71653) );
  AOI22xp33_ASAP7_75t_SL U57304 ( .A1(n72303), .A2(n72474), .B1(n72393), .B2(
        n72137), .Y(n72139) );
  INVxp67_ASAP7_75t_SL U57305 ( .A(n62608), .Y(n58236) );
  OAI22xp33_ASAP7_75t_SL U57306 ( .A1(n78331), .A2(n70035), .B1(n78332), .B2(
        n70034), .Y(n69737) );
  INVx1_ASAP7_75t_SL U57307 ( .A(n76956), .Y(n74855) );
  AOI22xp33_ASAP7_75t_SL U57308 ( .A1(n66126), .A2(n66125), .B1(n66124), .B2(
        n66133), .Y(n66127) );
  INVxp33_ASAP7_75t_SL U57309 ( .A(n68812), .Y(n74587) );
  AOI21xp33_ASAP7_75t_SL U57310 ( .A1(n72158), .A2(n72393), .B(n72157), .Y(
        n72160) );
  OAI21xp33_ASAP7_75t_SL U57311 ( .A1(n78329), .A2(n70034), .B(n69899), .Y(
        n69765) );
  NAND2xp5_ASAP7_75t_SL U57312 ( .A(n69864), .B(n69850), .Y(n69859) );
  INVx1_ASAP7_75t_SL U57313 ( .A(n62381), .Y(n77608) );
  AOI21xp33_ASAP7_75t_SL U57314 ( .A1(n70302), .A2(n70401), .B(n70259), .Y(
        n2318) );
  INVx1_ASAP7_75t_SL U57315 ( .A(n61084), .Y(n77638) );
  OAI22xp33_ASAP7_75t_SL U57316 ( .A1(n78424), .A2(n70035), .B1(n78354), .B2(
        n70034), .Y(n69994) );
  AOI21xp33_ASAP7_75t_SL U57317 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_), .A2(n59627), .B(n72627), 
        .Y(n72658) );
  INVx1_ASAP7_75t_SL U57318 ( .A(n61445), .Y(n61447) );
  INVx1_ASAP7_75t_SL U57319 ( .A(n61831), .Y(n61358) );
  INVxp33_ASAP7_75t_SL U57320 ( .A(n66261), .Y(n66262) );
  NAND2xp5_ASAP7_75t_SL U57321 ( .A(n69885), .B(n69858), .Y(n69863) );
  OAI21xp33_ASAP7_75t_SL U57322 ( .A1(n69758), .A2(n69757), .B(n69756), .Y(
        n69759) );
  AOI22xp33_ASAP7_75t_SL U57323 ( .A1(dwb_dat_i[14]), .A2(n61546), .B1(
        or1200_dc_top_from_dcram_14_), .B2(n61547), .Y(n62253) );
  OAI21xp33_ASAP7_75t_SL U57324 ( .A1(n77108), .A2(n76770), .B(n76769), .Y(
        n76783) );
  OAI21xp33_ASAP7_75t_SL U57325 ( .A1(n61408), .A2(n61426), .B(n61202), .Y(
        n61203) );
  NAND2xp5_ASAP7_75t_SL U57326 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_4_), .B(
        n71651), .Y(n71723) );
  INVxp67_ASAP7_75t_SL U57327 ( .A(n74205), .Y(n74193) );
  INVxp33_ASAP7_75t_SL U57328 ( .A(n70019), .Y(n69488) );
  NAND2xp33_ASAP7_75t_SL U57329 ( .A(n65402), .B(n65388), .Y(n2479) );
  INVxp33_ASAP7_75t_SL U57330 ( .A(n77056), .Y(n77079) );
  OAI21xp5_ASAP7_75t_SL U57331 ( .A1(n57120), .A2(n77696), .B(n60738), .Y(
        n60775) );
  INVxp67_ASAP7_75t_SL U57332 ( .A(n75589), .Y(n64230) );
  AOI22xp33_ASAP7_75t_SL U57333 ( .A1(n76763), .A2(n62366), .B1(n62425), .B2(
        n77076), .Y(n61441) );
  AOI22xp33_ASAP7_75t_SL U57334 ( .A1(n62344), .A2(n61494), .B1(n62374), .B2(
        n62425), .Y(n60680) );
  AOI22xp33_ASAP7_75t_SL U57335 ( .A1(n72393), .A2(n72149), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B2(
        n72416), .Y(n72151) );
  INVxp33_ASAP7_75t_SL U57336 ( .A(n76772), .Y(n62276) );
  OAI21xp5_ASAP7_75t_SL U57337 ( .A1(n65785), .A2(n58419), .B(n65733), .Y(
        n66079) );
  OAI22xp33_ASAP7_75t_SL U57338 ( .A1(n78332), .A2(n70035), .B1(n78334), .B2(
        n70034), .Y(n69763) );
  OAI22xp33_ASAP7_75t_SL U57339 ( .A1(n58599), .A2(n72513), .B1(n72030), .B2(
        n72029), .Y(n72031) );
  OA21x2_ASAP7_75t_SL U57340 ( .A1(n72415), .A2(n72208), .B(n72207), .Y(n72209) );
  AOI22xp33_ASAP7_75t_SL U57341 ( .A1(dwb_dat_i[10]), .A2(n61546), .B1(
        or1200_dc_top_from_dcram_10_), .B2(n61547), .Y(n63564) );
  OAI21xp33_ASAP7_75t_SL U57342 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[29]), .A2(n58419), 
        .B(n65762), .Y(n65763) );
  NAND2xp5_ASAP7_75t_SL U57343 ( .A(n60144), .B(n60143), .Y(n60145) );
  INVxp33_ASAP7_75t_SL U57344 ( .A(n75845), .Y(n61637) );
  OAI22xp33_ASAP7_75t_SL U57345 ( .A1(dwb_dat_i[8]), .A2(n61547), .B1(
        or1200_dc_top_from_dcram_8_), .B2(n61546), .Y(n62377) );
  OAI21xp33_ASAP7_75t_SL U57346 ( .A1(n2794), .A2(n76717), .B(n61382), .Y(
        n61450) );
  INVxp67_ASAP7_75t_SL U57347 ( .A(n74701), .Y(n74707) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U57348 ( .A1(n66145), .A2(n66089), .B(n66125), 
        .C(n65642), .Y(n65589) );
  NOR2xp33_ASAP7_75t_SRAM U57349 ( .A(n69832), .B(n69830), .Y(n69836) );
  AOI22xp33_ASAP7_75t_SL U57350 ( .A1(n65658), .A2(n65453), .B1(n65452), .B2(
        n65451), .Y(n65659) );
  AOI22xp33_ASAP7_75t_SL U57351 ( .A1(dwb_dat_i[6]), .A2(n61546), .B1(
        or1200_dc_top_from_dcram_6_), .B2(n61547), .Y(n64313) );
  OAI21xp33_ASAP7_75t_SL U57352 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[11]), .A2(
        n58284), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[11]), .Y(
        n73172) );
  NOR2xp33_ASAP7_75t_SRAM U57353 ( .A(or1200_cpu_or1200_mult_mac_n147), .B(
        n63555), .Y(n61472) );
  AOI21xp33_ASAP7_75t_SL U57354 ( .A1(n77097), .A2(n75628), .B(n75736), .Y(
        n75594) );
  OA21x2_ASAP7_75t_SL U57355 ( .A1(n70530), .A2(n27502), .B(n70498), .Y(n70499) );
  INVxp67_ASAP7_75t_SL U57356 ( .A(n77041), .Y(n77633) );
  INVx1_ASAP7_75t_SL U57357 ( .A(n70048), .Y(n70071) );
  AOI21xp33_ASAP7_75t_SL U57358 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[22]), .B(n70524), .Y(
        n2254) );
  AOI22xp33_ASAP7_75t_SL U57359 ( .A1(n63451), .A2(n57121), .B1(n53430), .B2(
        n60803), .Y(n62456) );
  AOI22xp33_ASAP7_75t_SL U57360 ( .A1(n63409), .A2(n57121), .B1(n61827), .B2(
        n61348), .Y(n61831) );
  OAI21xp33_ASAP7_75t_SL U57361 ( .A1(n63328), .A2(n63327), .B(n63335), .Y(
        n63329) );
  INVxp67_ASAP7_75t_SL U57362 ( .A(n63327), .Y(n63330) );
  NOR2xp33_ASAP7_75t_SRAM U57363 ( .A(n61297), .B(n77767), .Y(n61299) );
  AOI21xp33_ASAP7_75t_SL U57364 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[13]), .B(n70495), .Y(
        n2236) );
  INVxp67_ASAP7_75t_SL U57365 ( .A(n70147), .Y(n70148) );
  INVx1_ASAP7_75t_SL U57366 ( .A(n69877), .Y(n69873) );
  OA21x2_ASAP7_75t_SL U57367 ( .A1(n70530), .A2(n27504), .B(n70522), .Y(n70523) );
  INVxp33_ASAP7_75t_SL U57368 ( .A(n60401), .Y(n59963) );
  AOI21xp33_ASAP7_75t_SL U57369 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[20]), .B(n70521), .Y(
        n2250) );
  AOI21xp33_ASAP7_75t_SL U57370 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[19]), .B(n70520), .Y(
        n2248) );
  AOI21xp33_ASAP7_75t_SL U57371 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[18]), .B(n70519), .Y(
        n2246) );
  AOI21xp33_ASAP7_75t_SL U57372 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[17]), .B(n70518), .Y(
        n2244) );
  AOI21xp33_ASAP7_75t_SL U57373 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[16]), .B(n70497), .Y(
        n2242) );
  AOI21xp33_ASAP7_75t_SL U57374 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[15]), .B(n70496), .Y(
        n2240) );
  AOI21xp33_ASAP7_75t_SL U57375 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[14]), .B(n70517), .Y(
        n2238) );
  NAND2xp33_ASAP7_75t_SL U57376 ( .A(n63282), .B(n57121), .Y(n60804) );
  AOI21xp33_ASAP7_75t_SL U57377 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[12]), .B(n70494), .Y(
        n2234) );
  AOI21xp33_ASAP7_75t_SL U57378 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[11]), .B(n70493), .Y(
        n2232) );
  AOI21xp33_ASAP7_75t_SL U57379 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[10]), .B(n70492), .Y(
        n2230) );
  AOI21xp33_ASAP7_75t_SL U57380 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[9]), .B(n70516), .Y(
        n2228) );
  NAND2xp5_ASAP7_75t_SL U57381 ( .A(n62208), .B(n62209), .Y(n75648) );
  OA21x2_ASAP7_75t_SL U57382 ( .A1(n70530), .A2(n27518), .B(n70513), .Y(n70514) );
  INVx1_ASAP7_75t_SL U57383 ( .A(n69944), .Y(n69880) );
  OA21x2_ASAP7_75t_SL U57384 ( .A1(n70530), .A2(n27519), .B(n70511), .Y(n70512) );
  INVxp33_ASAP7_75t_SL U57385 ( .A(n77080), .Y(n77084) );
  INVx1_ASAP7_75t_SL U57386 ( .A(n75882), .Y(n77112) );
  OAI21xp33_ASAP7_75t_SL U57387 ( .A1(n71629), .A2(n71613), .B(n71554), .Y(
        n71555) );
  NAND2xp33_ASAP7_75t_SL U57388 ( .A(n61678), .B(n61677), .Y(n61679) );
  OAI21xp33_ASAP7_75t_SL U57389 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[32]), .A2(n65436), 
        .B(n65435), .Y(n65437) );
  AOI21xp33_ASAP7_75t_SL U57390 ( .A1(n74209), .A2(n74091), .B(n74752), .Y(
        n74092) );
  INVxp33_ASAP7_75t_SL U57391 ( .A(n70829), .Y(n70832) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U57392 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .A2(
        n72228), .B(n72227), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .Y(
        n72229) );
  NOR2x1_ASAP7_75t_SL U57393 ( .A(n799), .B(n60140), .Y(n60149) );
  INVx1_ASAP7_75t_SL U57394 ( .A(n74752), .Y(n74162) );
  INVxp67_ASAP7_75t_SL U57395 ( .A(n72081), .Y(n72082) );
  INVx1_ASAP7_75t_SL U57396 ( .A(n70091), .Y(n70098) );
  NAND2xp33_ASAP7_75t_SL U57397 ( .A(n75855), .B(n57121), .Y(n61813) );
  NAND2xp5_ASAP7_75t_SL U57398 ( .A(n63404), .B(n63428), .Y(n63412) );
  NAND2xp5_ASAP7_75t_SL U57399 ( .A(n72078), .B(n72077), .Y(n72202) );
  AOI22xp5_ASAP7_75t_SL U57400 ( .A1(n65160), .A2(n57121), .B1(n53430), .B2(
        n64240), .Y(n64251) );
  OAI22xp33_ASAP7_75t_SL U57401 ( .A1(n70439), .A2(n70551), .B1(n74660), .B2(
        n70553), .Y(n70407) );
  NAND2xp5_ASAP7_75t_SL U57402 ( .A(n69708), .B(n69707), .Y(n70073) );
  NOR2xp33_ASAP7_75t_SRAM U57403 ( .A(n1169), .B(n61597), .Y(n61601) );
  INVxp33_ASAP7_75t_SL U57404 ( .A(n77100), .Y(n61493) );
  AOI21xp33_ASAP7_75t_SL U57405 ( .A1(n75727), .A2(n64124), .B(n64123), .Y(
        n64125) );
  INVxp33_ASAP7_75t_SL U57406 ( .A(n70006), .Y(n70008) );
  AOI21xp33_ASAP7_75t_SL U57407 ( .A1(n75705), .A2(n75861), .B(n75704), .Y(
        n75719) );
  INVxp33_ASAP7_75t_SL U57408 ( .A(n70003), .Y(n70009) );
  OAI21xp5_ASAP7_75t_SL U57409 ( .A1(n2982), .A2(n74953), .B(n60012), .Y(
        n60013) );
  AOI22xp33_ASAP7_75t_SL U57410 ( .A1(n65124), .A2(n57121), .B1(n53430), .B2(
        n64305), .Y(n64319) );
  INVxp33_ASAP7_75t_SL U57411 ( .A(n61595), .Y(n61596) );
  NAND2xp5_ASAP7_75t_SL U57412 ( .A(n60109), .B(n60108), .Y(n60112) );
  NAND2xp33_ASAP7_75t_SL U57413 ( .A(n70049), .B(n70072), .Y(n69706) );
  NAND2xp33_ASAP7_75t_SL U57414 ( .A(n58912), .B(n61406), .Y(n61407) );
  AOI21xp33_ASAP7_75t_SL U57415 ( .A1(n70447), .A2(n70545), .B(n70287), .Y(
        n2374) );
  INVxp67_ASAP7_75t_SL U57416 ( .A(n75717), .Y(n63567) );
  INVxp67_ASAP7_75t_SL U57417 ( .A(n75346), .Y(n64219) );
  NAND2xp33_ASAP7_75t_SL U57418 ( .A(n61324), .B(n76713), .Y(n61325) );
  INVx1_ASAP7_75t_SL U57419 ( .A(n72421), .Y(n72425) );
  OAI21xp33_ASAP7_75t_SL U57420 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_4_), .A2(
        n74331), .B(n74341), .Y(n2395) );
  INVxp33_ASAP7_75t_SL U57421 ( .A(n69849), .Y(n69644) );
  OAI21xp33_ASAP7_75t_SL U57422 ( .A1(n66151), .A2(n65639), .B(n65638), .Y(
        n65640) );
  OAI21xp33_ASAP7_75t_SL U57423 ( .A1(n64769), .A2(n75838), .B(n62520), .Y(
        n62521) );
  INVxp33_ASAP7_75t_SL U57424 ( .A(n61531), .Y(n60943) );
  NAND2xp5_ASAP7_75t_SL U57425 ( .A(n69641), .B(n69640), .Y(n69864) );
  INVxp67_ASAP7_75t_SL U57426 ( .A(n75833), .Y(n62536) );
  NAND2xp5_ASAP7_75t_SL U57427 ( .A(n71840), .B(n71839), .Y(n72446) );
  NOR2x1_ASAP7_75t_SL U57428 ( .A(n65680), .B(n65827), .Y(n66024) );
  OAI21xp5_ASAP7_75t_SL U57429 ( .A1(n63693), .A2(n77260), .B(n63692), .Y(
        n74947) );
  INVxp67_ASAP7_75t_SL U57430 ( .A(n75349), .Y(n61658) );
  INVxp33_ASAP7_75t_SL U57431 ( .A(n75729), .Y(n62278) );
  AOI21xp33_ASAP7_75t_SL U57432 ( .A1(n72534), .A2(n72398), .B(n72168), .Y(
        n72324) );
  NOR2x1_ASAP7_75t_SL U57433 ( .A(n75872), .B(n76775), .Y(n75736) );
  OAI21xp33_ASAP7_75t_SL U57434 ( .A1(n72355), .A2(n72017), .B(n71880), .Y(
        n71881) );
  INVxp33_ASAP7_75t_SL U57435 ( .A(n61514), .Y(n60924) );
  NAND2xp33_ASAP7_75t_SL U57436 ( .A(n61379), .B(n61677), .Y(n61380) );
  AOI21xp33_ASAP7_75t_SL U57437 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[5]), .B(n70510), .Y(
        n2220) );
  AOI21xp33_ASAP7_75t_SL U57438 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[4]), .B(n70509), .Y(
        n2218) );
  INVxp33_ASAP7_75t_SL U57439 ( .A(n77767), .Y(n77485) );
  AOI21xp33_ASAP7_75t_SL U57440 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[3]), .B(n70508), .Y(
        n2216) );
  OA21x2_ASAP7_75t_SL U57441 ( .A1(n70530), .A2(n27523), .B(n70506), .Y(n70507) );
  OA21x2_ASAP7_75t_SL U57442 ( .A1(n70530), .A2(n27524), .B(n70504), .Y(n70505) );
  INVxp67_ASAP7_75t_SL U57443 ( .A(n72397), .Y(n72414) );
  AOI22xp33_ASAP7_75t_SL U57444 ( .A1(n63315), .A2(n57121), .B1(n53430), .B2(
        n61633), .Y(n61622) );
  INVx1_ASAP7_75t_SL U57445 ( .A(n72412), .Y(n72382) );
  INVxp67_ASAP7_75t_SL U57446 ( .A(n69890), .Y(n69912) );
  AOI21xp33_ASAP7_75t_SL U57447 ( .A1(n76713), .A2(n62235), .B(n62234), .Y(
        n62242) );
  AOI22xp33_ASAP7_75t_SL U57448 ( .A1(n63334), .A2(n57121), .B1(n61827), .B2(
        n62268), .Y(n62287) );
  INVxp67_ASAP7_75t_SL U57449 ( .A(n70172), .Y(n70174) );
  OAI22xp33_ASAP7_75t_SL U57450 ( .A1(n65800), .A2(n65799), .B1(n58582), .B2(
        n65859), .Y(n65932) );
  AOI22xp33_ASAP7_75t_SL U57451 ( .A1(n63300), .A2(n57121), .B1(n61827), .B2(
        n60806), .Y(n61486) );
  AOI22xp33_ASAP7_75t_SL U57452 ( .A1(n61418), .A2(n57121), .B1(n61827), .B2(
        n60807), .Y(n61445) );
  NAND2xp5_ASAP7_75t_SL U57453 ( .A(n69655), .B(n69654), .Y(n69885) );
  NAND2xp5_ASAP7_75t_SL U57454 ( .A(n63942), .B(n63941), .Y(n63955) );
  OAI21xp33_ASAP7_75t_SL U57455 ( .A1(n65841), .A2(n65840), .B(n65687), .Y(
        n65969) );
  NOR2xp33_ASAP7_75t_SRAM U57456 ( .A(n76836), .B(n60401), .Y(n77428) );
  NAND2xp33_ASAP7_75t_SL U57457 ( .A(n75833), .B(n77061), .Y(n75834) );
  INVxp33_ASAP7_75t_SL U57458 ( .A(n63266), .Y(n63268) );
  NOR2xp33_ASAP7_75t_SRAM U57459 ( .A(n61303), .B(n68810), .Y(n77967) );
  AOI21xp33_ASAP7_75t_SL U57460 ( .A1(n72334), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .B(
        n72148), .Y(n72416) );
  NAND2xp5_ASAP7_75t_SL U57461 ( .A(n74294), .B(n74290), .Y(n72559) );
  INVxp67_ASAP7_75t_SL U57462 ( .A(n64221), .Y(n75329) );
  AOI22xp5_ASAP7_75t_SL U57463 ( .A1(n70171), .A2(n70170), .B1(n70169), .B2(
        n70185), .Y(n70186) );
  INVxp33_ASAP7_75t_SL U57464 ( .A(n76775), .Y(n77070) );
  OR3x4_ASAP7_75t_SL U57465 ( .A(n63266), .B(n63265), .C(n63264), .Y(n76897)
         );
  INVxp67_ASAP7_75t_SL U57466 ( .A(n72325), .Y(n72451) );
  OAI22xp33_ASAP7_75t_SL U57467 ( .A1(n65604), .A2(n66095), .B1(n65603), .B2(
        n66121), .Y(n65605) );
  NOR2x1p5_ASAP7_75t_SL U57468 ( .A(n63814), .B(n63654), .Y(n57644) );
  INVxp33_ASAP7_75t_SL U57469 ( .A(n64167), .Y(n64168) );
  NOR2xp33_ASAP7_75t_SRAM U57470 ( .A(n62355), .B(n62354), .Y(n62360) );
  INVxp33_ASAP7_75t_SL U57471 ( .A(n75555), .Y(n64284) );
  NAND2xp5_ASAP7_75t_SL U57472 ( .A(n76712), .B(n63253), .Y(n63254) );
  NAND2xp33_ASAP7_75t_SL U57473 ( .A(n74956), .B(n60042), .Y(n60050) );
  NAND2xp33_ASAP7_75t_SL U57474 ( .A(n72095), .B(n72242), .Y(n72106) );
  INVxp67_ASAP7_75t_SL U57475 ( .A(n72104), .Y(n72127) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U57476 ( .A1(n76954), .A2(n76953), .B(n76952), 
        .C(n76951), .Y(n76955) );
  OAI21xp33_ASAP7_75t_SL U57477 ( .A1(n74232), .A2(n74231), .B(n74273), .Y(
        n74238) );
  NAND2xp33_ASAP7_75t_SL U57478 ( .A(n75220), .B(n74594), .Y(n74606) );
  AOI21xp33_ASAP7_75t_SL U57479 ( .A1(n76753), .A2(n63453), .B(n61719), .Y(
        n61720) );
  BUFx3_ASAP7_75t_SL U57480 ( .A(n67030), .Y(n57184) );
  INVxp33_ASAP7_75t_SL U57481 ( .A(n69755), .Y(n69760) );
  AOI21xp33_ASAP7_75t_SL U57482 ( .A1(n62471), .A2(n76557), .B(n62470), .Y(
        n69344) );
  NAND2xp5_ASAP7_75t_SL U57483 ( .A(n74688), .B(n74687), .Y(n74701) );
  NAND2xp33_ASAP7_75t_SL U57484 ( .A(n69742), .B(n70078), .Y(n69745) );
  INVxp67_ASAP7_75t_SL U57485 ( .A(n74594), .Y(n64855) );
  INVx1_ASAP7_75t_SL U57486 ( .A(n75625), .Y(n77301) );
  NAND2xp33_ASAP7_75t_SL U57487 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .B(
        n72393), .Y(n72010) );
  NAND2xp5_ASAP7_75t_SL U57488 ( .A(n76458), .B(n76457), .Y(n76470) );
  OAI21x1_ASAP7_75t_SL U57489 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_22_), .A2(n69421), .B(
        n78244), .Y(n70109) );
  OAI22xp33_ASAP7_75t_SL U57490 ( .A1(n59709), .A2(n75327), .B1(n59708), .B2(
        n75326), .Y(n62110) );
  NAND2xp5_ASAP7_75t_SL U57491 ( .A(n70240), .B(n70576), .Y(n70234) );
  INVxp33_ASAP7_75t_SL U57492 ( .A(n70599), .Y(n70216) );
  OAI21xp33_ASAP7_75t_SL U57493 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[24]), .A2(n70249), 
        .B(n2456), .Y(n70248) );
  OAI22xp33_ASAP7_75t_SL U57494 ( .A1(n74645), .A2(n70553), .B1(n74691), .B2(
        n70551), .Y(n70259) );
  OAI22xp33_ASAP7_75t_SL U57495 ( .A1(n74645), .A2(n70551), .B1(n70552), .B2(
        n70553), .Y(n70254) );
  INVxp67_ASAP7_75t_SL U57496 ( .A(n70323), .Y(n2324) );
  INVxp67_ASAP7_75t_SL U57497 ( .A(n65595), .Y(n65642) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U57498 ( .A1(n72384), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        n72051), .C(n72104), .Y(n72052) );
  OAI21xp33_ASAP7_75t_SL U57499 ( .A1(n63889), .A2(n63770), .B(n63890), .Y(
        n63772) );
  NAND2xp5_ASAP7_75t_SL U57500 ( .A(n69720), .B(n69728), .Y(n69721) );
  INVxp67_ASAP7_75t_SL U57501 ( .A(n72273), .Y(n72016) );
  INVxp67_ASAP7_75t_SL U57502 ( .A(n72233), .Y(n72002) );
  INVx1_ASAP7_75t_SL U57503 ( .A(n73606), .Y(n73608) );
  AOI21xp33_ASAP7_75t_SL U57504 ( .A1(n69346), .A2(n76557), .B(n69345), .Y(
        n77133) );
  OAI22xp33_ASAP7_75t_SL U57505 ( .A1(n74654), .A2(n70553), .B1(n74664), .B2(
        n70551), .Y(n70332) );
  INVxp67_ASAP7_75t_SL U57506 ( .A(n62576), .Y(n62577) );
  NAND2xp33_ASAP7_75t_SL U57507 ( .A(n2071), .B(n61034), .Y(n61035) );
  INVxp33_ASAP7_75t_SL U57508 ( .A(n65663), .Y(n65515) );
  INVxp33_ASAP7_75t_SL U57509 ( .A(n71095), .Y(n71096) );
  NAND2xp33_ASAP7_75t_SL U57510 ( .A(n61246), .B(n76713), .Y(n61247) );
  AOI21xp33_ASAP7_75t_SL U57511 ( .A1(n72037), .A2(n72399), .B(n58599), .Y(
        n71920) );
  NAND2xp33_ASAP7_75t_SL U57512 ( .A(n65514), .B(n65663), .Y(n66090) );
  NAND2xp5_ASAP7_75t_SL U57513 ( .A(n72105), .B(n72104), .Y(n72269) );
  NAND2xp33_ASAP7_75t_SL U57514 ( .A(n74798), .B(n59168), .Y(n1512) );
  NAND2xp33_ASAP7_75t_SL U57515 ( .A(n77984), .B(n77988), .Y(n3909) );
  INVx1_ASAP7_75t_SL U57516 ( .A(n62344), .Y(n62531) );
  NAND2xp33_ASAP7_75t_SL U57517 ( .A(n75558), .B(n77041), .Y(n75559) );
  NAND2xp5_ASAP7_75t_SL U57518 ( .A(n71945), .B(n71944), .Y(n72206) );
  NOR2xp33_ASAP7_75t_SL U57519 ( .A(n58305), .B(n75737), .Y(n64217) );
  NAND2xp33_ASAP7_75t_SL U57520 ( .A(n77989), .B(n77988), .Y(n3907) );
  INVxp33_ASAP7_75t_SL U57521 ( .A(n75330), .Y(n64223) );
  NAND2xp33_ASAP7_75t_SL U57522 ( .A(n77963), .B(n77988), .Y(n3922) );
  NAND2xp33_ASAP7_75t_SL U57523 ( .A(n61381), .B(n76720), .Y(n61382) );
  NAND2xp33_ASAP7_75t_SL U57524 ( .A(n65816), .B(n66080), .Y(n65815) );
  INVxp67_ASAP7_75t_SL U57525 ( .A(n77104), .Y(n75585) );
  NAND2xp33_ASAP7_75t_SL U57526 ( .A(n77969), .B(n77988), .Y(n3920) );
  AOI21xp33_ASAP7_75t_SL U57527 ( .A1(n75727), .A2(n64240), .B(n64239), .Y(
        n64243) );
  INVxp67_ASAP7_75t_SL U57528 ( .A(n72330), .Y(n72203) );
  OAI21xp33_ASAP7_75t_SL U57529 ( .A1(n72112), .A2(n72017), .B(n71964), .Y(
        n72208) );
  AOI21xp33_ASAP7_75t_SL U57530 ( .A1(n76754), .A2(n76753), .B(n76752), .Y(
        n76756) );
  OAI21xp5_ASAP7_75t_SL U57531 ( .A1(n2979), .A2(n74953), .B(n60006), .Y(
        n60007) );
  INVxp33_ASAP7_75t_SL U57532 ( .A(n65450), .Y(n65451) );
  INVx1_ASAP7_75t_SL U57533 ( .A(n77039), .Y(n64275) );
  OR2x2_ASAP7_75t_SL U57534 ( .A(n76717), .B(n75766), .Y(n77233) );
  INVxp33_ASAP7_75t_SL U57535 ( .A(n64775), .Y(n60650) );
  INVxp67_ASAP7_75t_SL U57536 ( .A(n72588), .Y(n72591) );
  INVx1_ASAP7_75t_SL U57537 ( .A(n64295), .Y(n75576) );
  AOI21xp33_ASAP7_75t_SL U57538 ( .A1(n75727), .A2(n75579), .B(n75578), .Y(
        n75580) );
  INVxp67_ASAP7_75t_SL U57539 ( .A(n72242), .Y(n72207) );
  AOI22xp33_ASAP7_75t_SL U57540 ( .A1(n77140), .A2(n77043), .B1(n77042), .B2(
        n77041), .Y(n77044) );
  INVxp33_ASAP7_75t_SL U57541 ( .A(n61783), .Y(n76760) );
  AOI21xp33_ASAP7_75t_SL U57542 ( .A1(n76720), .A2(n61606), .B(n61605), .Y(
        n77598) );
  NAND2xp5_ASAP7_75t_SL U57543 ( .A(n61698), .B(n61697), .Y(n76772) );
  AOI22xp33_ASAP7_75t_SL U57544 ( .A1(n75847), .A2(n78002), .B1(n75592), .B2(
        n75591), .Y(n75593) );
  AOI22xp33_ASAP7_75t_SL U57545 ( .A1(n65401), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_6_), .B1(n65400), .B2(
        n65390), .Y(n1953) );
  AOI21xp33_ASAP7_75t_SL U57546 ( .A1(n76720), .A2(n76719), .B(n76718), .Y(
        n77604) );
  NAND2xp33_ASAP7_75t_SL U57547 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        n72475), .Y(n72218) );
  INVxp33_ASAP7_75t_SL U57548 ( .A(n76779), .Y(n64220) );
  OAI21xp5_ASAP7_75t_SL U57549 ( .A1(n71522), .A2(n71521), .B(n72614), .Y(
        n71523) );
  AOI21xp33_ASAP7_75t_SL U57550 ( .A1(n75833), .A2(n64771), .B(n64770), .Y(
        n64772) );
  INVxp33_ASAP7_75t_SL U57551 ( .A(n64218), .Y(n64774) );
  NAND2xp33_ASAP7_75t_SL U57552 ( .A(n65663), .B(n65517), .Y(n66158) );
  AOI21xp5_ASAP7_75t_SL U57553 ( .A1(n61315), .A2(n61314), .B(n61313), .Y(
        n61990) );
  INVx1_ASAP7_75t_SL U57554 ( .A(n72589), .Y(n74230) );
  NAND2xp33_ASAP7_75t_SL U57555 ( .A(n76714), .B(n76713), .Y(n76715) );
  OAI21xp5_ASAP7_75t_SL U57556 ( .A1(n2985), .A2(n74953), .B(n60021), .Y(
        n60022) );
  OAI21xp33_ASAP7_75t_SL U57557 ( .A1(n65761), .A2(n58419), .B(n65760), .Y(
        n66017) );
  INVxp67_ASAP7_75t_SL U57558 ( .A(n70918), .Y(n70921) );
  INVxp33_ASAP7_75t_SL U57559 ( .A(n75819), .Y(n64821) );
  OAI21xp33_ASAP7_75t_SL U57560 ( .A1(n75116), .A2(n64819), .B(n64818), .Y(
        n64820) );
  OAI22xp33_ASAP7_75t_SL U57561 ( .A1(n2335), .A2(n70551), .B1(n74691), .B2(
        n70553), .Y(n70268) );
  INVx1_ASAP7_75t_SL U57562 ( .A(n70114), .Y(n70112) );
  NAND2xp33_ASAP7_75t_SL U57563 ( .A(n64825), .B(n75727), .Y(n64827) );
  OAI21xp33_ASAP7_75t_SL U57564 ( .A1(n70124), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[1]), .B(
        n70117), .Y(n70116) );
  OAI21xp5_ASAP7_75t_SL U57565 ( .A1(n2988), .A2(n74953), .B(n60027), .Y(
        n60028) );
  INVxp67_ASAP7_75t_SL U57566 ( .A(n71704), .Y(n71706) );
  NAND2xp33_ASAP7_75t_SL U57567 ( .A(n77972), .B(n77988), .Y(n3917) );
  INVxp33_ASAP7_75t_SL U57568 ( .A(n75573), .Y(n61533) );
  NAND2xp5_ASAP7_75t_SL U57569 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[5]), .B(n73554), 
        .Y(n73572) );
  AOI22xp33_ASAP7_75t_SL U57570 ( .A1(n77285), .A2(n62409), .B1(n62408), .B2(
        n76720), .Y(n77626) );
  INVxp33_ASAP7_75t_SL U57571 ( .A(n70902), .Y(n70905) );
  AOI21xp33_ASAP7_75t_SL U57572 ( .A1(n70545), .A2(n70429), .B(n70279), .Y(
        n2334) );
  NAND2xp33_ASAP7_75t_SL U57573 ( .A(n77975), .B(n77988), .Y(n3915) );
  NAND2xp5_ASAP7_75t_SL U57574 ( .A(n71926), .B(n71925), .Y(n72195) );
  NAND2xp33_ASAP7_75t_SL U57575 ( .A(n77978), .B(n77988), .Y(n3913) );
  NAND2xp5_ASAP7_75t_SL U57576 ( .A(n63491), .B(n63510), .Y(n63492) );
  OAI21xp33_ASAP7_75t_SL U57577 ( .A1(n76537), .A2(n76557), .B(n61159), .Y(
        n77026) );
  NAND2xp33_ASAP7_75t_SL U57578 ( .A(n77981), .B(n77988), .Y(n3911) );
  AOI21xp33_ASAP7_75t_SL U57579 ( .A1(n76720), .A2(n61681), .B(n61680), .Y(
        n77616) );
  INVx1_ASAP7_75t_SL U57580 ( .A(n75727), .Y(n64785) );
  OAI21xp5_ASAP7_75t_SL U57581 ( .A1(n61699), .A2(n61698), .B(n61697), .Y(
        n75589) );
  OAI21xp33_ASAP7_75t_SL U57582 ( .A1(n73815), .A2(n73818), .B(n73795), .Y(
        n3298) );
  AOI21xp33_ASAP7_75t_SL U57583 ( .A1(n72483), .A2(n72492), .B(n72454), .Y(
        n72455) );
  NAND2xp5_ASAP7_75t_SL U57584 ( .A(n71704), .B(n71696), .Y(n71697) );
  INVxp33_ASAP7_75t_SL U57585 ( .A(n63577), .Y(n61781) );
  INVxp33_ASAP7_75t_SL U57586 ( .A(n71707), .Y(n71651) );
  INVxp33_ASAP7_75t_SL U57587 ( .A(n60140), .Y(n60124) );
  OAI21xp33_ASAP7_75t_SL U57588 ( .A1(n60402), .A2(n69331), .B(n69330), .Y(
        n60403) );
  AND2x2_ASAP7_75t_SL U57589 ( .A(n60584), .B(n60583), .Y(n61547) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57590 ( .A1(n66163), .A2(n66149), .B(n65676), .C(
        n65617), .Y(n65618) );
  NAND2xp5_ASAP7_75t_SL U57591 ( .A(n76833), .B(n76832), .Y(n76842) );
  INVxp33_ASAP7_75t_SL U57592 ( .A(n62257), .Y(n64843) );
  INVxp33_ASAP7_75t_SL U57593 ( .A(n70726), .Y(n70728) );
  NAND2xp5_ASAP7_75t_SL U57594 ( .A(n71738), .B(n71707), .Y(n71652) );
  INVxp33_ASAP7_75t_SL U57595 ( .A(n71650), .Y(n71689) );
  OA21x2_ASAP7_75t_SL U57596 ( .A1(n74333), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_5_), 
        .B(n74345), .Y(n74334) );
  NAND2xp33_ASAP7_75t_SL U57597 ( .A(n61125), .B(n61124), .Y(n61127) );
  INVxp67_ASAP7_75t_SL U57598 ( .A(n69758), .Y(n69761) );
  OAI21xp5_ASAP7_75t_SL U57599 ( .A1(n77261), .A2(n77260), .B(n77259), .Y(
        n77270) );
  INVx1_ASAP7_75t_SL U57600 ( .A(n60777), .Y(n60779) );
  OAI22xp33_ASAP7_75t_SL U57601 ( .A1(n75324), .A2(n76770), .B1(n75325), .B2(
        n75330), .Y(n75241) );
  INVxp67_ASAP7_75t_SL U57602 ( .A(n69770), .Y(n69771) );
  OAI21xp5_ASAP7_75t_SL U57603 ( .A1(n77260), .A2(n61585), .B(n61584), .Y(
        n61586) );
  OAI22xp33_ASAP7_75t_SL U57604 ( .A1(DP_OP_741J1_129_6992_n46), .A2(n70553), 
        .B1(n70552), .B2(n70551), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_N139) );
  NAND2xp33_ASAP7_75t_SL U57605 ( .A(n60563), .B(n77041), .Y(n60564) );
  INVxp33_ASAP7_75t_SL U57606 ( .A(n74361), .Y(n74363) );
  NAND2xp5_ASAP7_75t_SL U57607 ( .A(n71724), .B(n71714), .Y(n71654) );
  INVx1_ASAP7_75t_SL U57608 ( .A(n77488), .Y(n77489) );
  INVx1_ASAP7_75t_SL U57609 ( .A(n76716), .Y(n63253) );
  INVxp67_ASAP7_75t_SL U57610 ( .A(n74788), .Y(n59168) );
  NAND2xp33_ASAP7_75t_SL U57611 ( .A(n70278), .B(n70277), .Y(n70279) );
  AOI22xp33_ASAP7_75t_SL U57612 ( .A1(n72062), .A2(n72144), .B1(n72110), .B2(
        n71923), .Y(n71926) );
  INVxp67_ASAP7_75t_SL U57613 ( .A(n64132), .Y(n75844) );
  INVxp67_ASAP7_75t_SL U57614 ( .A(n76483), .Y(n76414) );
  INVxp67_ASAP7_75t_SL U57615 ( .A(n73545), .Y(n73554) );
  OAI22xp33_ASAP7_75t_SL U57616 ( .A1(n72226), .A2(n59623), .B1(n72434), .B2(
        n72228), .Y(n72135) );
  NAND2xp33_ASAP7_75t_SL U57617 ( .A(n66089), .B(n66088), .Y(n66091) );
  INVxp33_ASAP7_75t_SL U57618 ( .A(n62262), .Y(n62270) );
  INVxp67_ASAP7_75t_SL U57619 ( .A(n74148), .Y(n74149) );
  INVxp67_ASAP7_75t_SL U57620 ( .A(n76986), .Y(n1501) );
  NAND2xp5_ASAP7_75t_SL U57621 ( .A(n65507), .B(n65601), .Y(n66122) );
  AOI21xp33_ASAP7_75t_SL U57622 ( .A1(n63743), .A2(n77864), .B(n60026), .Y(
        n60027) );
  NOR2x1_ASAP7_75t_SL U57623 ( .A(n60843), .B(n62444), .Y(n77080) );
  AOI21xp33_ASAP7_75t_SL U57624 ( .A1(n73921), .A2(n61777), .B(n61776), .Y(
        n61778) );
  AND4x1_ASAP7_75t_SL U57625 ( .A(n75452), .B(n61131), .C(n60227), .D(n77850), 
        .Y(n60228) );
  INVxp67_ASAP7_75t_SL U57626 ( .A(n72558), .Y(n72548) );
  INVx1_ASAP7_75t_SL U57627 ( .A(n76753), .Y(n77073) );
  OAI22xp33_ASAP7_75t_SL U57628 ( .A1(n59622), .A2(n72337), .B1(n59623), .B2(
        n72220), .Y(n72181) );
  INVxp67_ASAP7_75t_SL U57629 ( .A(n71291), .Y(n71289) );
  AOI22xp33_ASAP7_75t_SL U57630 ( .A1(n59687), .A2(n77494), .B1(n77493), .B2(
        n77492), .Y(n6731) );
  NAND2xp5_ASAP7_75t_SL U57631 ( .A(n60920), .B(n61411), .Y(n60921) );
  OAI22xp33_ASAP7_75t_SL U57632 ( .A1(n65354), .A2(n65389), .B1(n65322), .B2(
        n65321), .Y(n65323) );
  INVxp33_ASAP7_75t_SL U57633 ( .A(n65691), .Y(n65514) );
  AOI21xp5_ASAP7_75t_SL U57634 ( .A1(n72558), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n131), .B(n72557), 
        .Y(n74290) );
  OAI22xp33_ASAP7_75t_SL U57635 ( .A1(n65793), .A2(n58419), .B1(n65822), .B2(
        n58571), .Y(n65794) );
  NAND2xp5_ASAP7_75t_SL U57636 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[1]), .B(
        n70124), .Y(n70117) );
  INVx1_ASAP7_75t_SL U57637 ( .A(n73602), .Y(n73504) );
  NAND2xp5_ASAP7_75t_SL U57638 ( .A(n70215), .B(n70214), .Y(n70599) );
  INVx1_ASAP7_75t_SL U57639 ( .A(n61215), .Y(n61428) );
  NAND2xp33_ASAP7_75t_SL U57640 ( .A(n73813), .B(n73796), .Y(n73800) );
  NAND2xp33_ASAP7_75t_SL U57641 ( .A(ic_en), .B(n58609), .Y(n60271) );
  INVxp33_ASAP7_75t_SL U57642 ( .A(n76717), .Y(n62409) );
  OAI22xp33_ASAP7_75t_SL U57643 ( .A1(n59622), .A2(n72452), .B1(n72434), .B2(
        n72338), .Y(n72300) );
  NAND2xp33_ASAP7_75t_SL U57644 ( .A(n2644), .B(n76557), .Y(n61159) );
  AOI21xp33_ASAP7_75t_SL U57645 ( .A1(n73822), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .B(
        n73734), .Y(n73735) );
  OAI22xp33_ASAP7_75t_SL U57646 ( .A1(n72479), .A2(n59624), .B1(n59623), .B2(
        n72453), .Y(n72301) );
  NAND2xp33_ASAP7_75t_SL U57647 ( .A(n57081), .B(n69786), .Y(n70513) );
  INVxp33_ASAP7_75t_SL U57648 ( .A(n71713), .Y(n71705) );
  AOI21xp5_ASAP7_75t_SL U57649 ( .A1(n72543), .A2(n72538), .B(n72537), .Y(
        n72539) );
  NAND2xp33_ASAP7_75t_SL U57650 ( .A(n78366), .B(n59629), .Y(n72690) );
  INVxp33_ASAP7_75t_SL U57651 ( .A(n70413), .Y(n70269) );
  INVx1_ASAP7_75t_SL U57652 ( .A(n69330), .Y(n77357) );
  INVxp33_ASAP7_75t_SL U57653 ( .A(n75823), .Y(n64819) );
  OAI22xp33_ASAP7_75t_SL U57654 ( .A1(n72370), .A2(n72434), .B1(n59623), .B2(
        n72371), .Y(n72356) );
  OAI22xp33_ASAP7_75t_SL U57655 ( .A1(n72506), .A2(n59624), .B1(n59622), .B2(
        n72472), .Y(n72357) );
  NAND2xp5_ASAP7_75t_SL U57656 ( .A(n77344), .B(n77353), .Y(n59158) );
  INVxp67_ASAP7_75t_SL U57657 ( .A(n70742), .Y(n70745) );
  NAND2xp33_ASAP7_75t_SL U57658 ( .A(n59687), .B(n77976), .Y(n3916) );
  NAND2xp5_ASAP7_75t_SL U57659 ( .A(n4318), .B(n4317), .Y(n77988) );
  NAND2xp33_ASAP7_75t_SL U57660 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_12_), .B(n69853), 
        .Y(n69850) );
  OAI21xp33_ASAP7_75t_SL U57661 ( .A1(n72370), .A2(n59622), .B(n72211), .Y(
        n72216) );
  NAND2xp33_ASAP7_75t_SL U57662 ( .A(n60071), .B(n60174), .Y(n60078) );
  INVxp33_ASAP7_75t_SL U57663 ( .A(n70699), .Y(n70697) );
  INVxp67_ASAP7_75t_SL U57664 ( .A(n60944), .Y(n60663) );
  NOR2xp33_ASAP7_75t_SRAM U57665 ( .A(n1378), .B(n61599), .Y(n61069) );
  NOR3xp33_ASAP7_75t_SRAM U57666 ( .A(n76954), .B(n76941), .C(n77196), .Y(
        n76952) );
  INVxp33_ASAP7_75t_SL U57667 ( .A(n62123), .Y(n75323) );
  NAND2xp33_ASAP7_75t_SL U57668 ( .A(n60043), .B(n60174), .Y(n60049) );
  INVx1_ASAP7_75t_SL U57669 ( .A(n70124), .Y(n69948) );
  AOI21xp33_ASAP7_75t_SL U57670 ( .A1(n63743), .A2(n77890), .B(n60117), .Y(
        n60118) );
  INVxp67_ASAP7_75t_SL U57671 ( .A(n75731), .Y(n73925) );
  INVxp33_ASAP7_75t_SL U57672 ( .A(n74514), .Y(n74519) );
  NAND2xp33_ASAP7_75t_SL U57673 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_10_), .B(n69628), 
        .Y(n69629) );
  AOI22xp33_ASAP7_75t_SL U57674 ( .A1(n72095), .A2(n71913), .B1(n72093), .B2(
        n71912), .Y(n71914) );
  INVxp33_ASAP7_75t_SL U57675 ( .A(n76782), .Y(n61498) );
  OA21x2_ASAP7_75t_SL U57676 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_sign_o), .A2(n74516), .B(n74514), .Y(n74515) );
  INVx1_ASAP7_75t_SL U57677 ( .A(n64834), .Y(n62274) );
  NAND2xp5_ASAP7_75t_SL U57678 ( .A(n69590), .B(n69723), .Y(n69728) );
  INVx1_ASAP7_75t_SL U57679 ( .A(n72452), .Y(n72483) );
  INVx1_ASAP7_75t_SL U57680 ( .A(n70031), .Y(n70060) );
  NAND2xp33_ASAP7_75t_SL U57681 ( .A(n78329), .B(n59629), .Y(n73045) );
  NAND2xp33_ASAP7_75t_SL U57682 ( .A(n59493), .B(n61844), .Y(n75819) );
  NAND2xp33_ASAP7_75t_SL U57683 ( .A(n65507), .B(n65691), .Y(n66150) );
  NAND2xp33_ASAP7_75t_SL U57684 ( .A(n78332), .B(n59629), .Y(n72855) );
  NAND2xp5_ASAP7_75t_SL U57685 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_4_), .B(
        n74331), .Y(n74341) );
  INVxp33_ASAP7_75t_SL U57686 ( .A(n63939), .Y(n60042) );
  NAND2xp33_ASAP7_75t_SL U57687 ( .A(n78348), .B(n59629), .Y(n72809) );
  NAND2xp33_ASAP7_75t_SL U57688 ( .A(n78328), .B(n74516), .Y(n74517) );
  INVxp33_ASAP7_75t_SL U57689 ( .A(n72322), .Y(n71907) );
  INVxp33_ASAP7_75t_SL U57690 ( .A(n70083), .Y(n69898) );
  NOR2xp33_ASAP7_75t_SRAM U57691 ( .A(n66159), .B(n65625), .Y(n65617) );
  NOR2xp33_ASAP7_75t_SRAM U57692 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .B(n65625), .Y(
        n66126) );
  INVxp33_ASAP7_75t_SL U57693 ( .A(n69853), .Y(n69640) );
  NAND2xp33_ASAP7_75t_SL U57694 ( .A(n75654), .B(n75823), .Y(n75205) );
  NAND2xp5_ASAP7_75t_SL U57695 ( .A(n73881), .B(n73880), .Y(n73891) );
  NAND2xp5_ASAP7_75t_SL U57696 ( .A(n62358), .B(n62357), .Y(n64127) );
  NAND2xp33_ASAP7_75t_SL U57697 ( .A(n71775), .B(n72334), .Y(n71776) );
  INVxp67_ASAP7_75t_SL U57698 ( .A(n58081), .Y(n62354) );
  NAND2xp33_ASAP7_75t_SL U57699 ( .A(n65674), .B(n66088), .Y(n65595) );
  INVxp33_ASAP7_75t_SL U57700 ( .A(n75522), .Y(n75523) );
  AOI21xp33_ASAP7_75t_SL U57701 ( .A1(n61245), .A2(n77622), .B(n61244), .Y(
        n76713) );
  OAI21xp33_ASAP7_75t_SL U57702 ( .A1(n72370), .A2(n59624), .B(n72167), .Y(
        n72168) );
  NAND2xp5_ASAP7_75t_SL U57703 ( .A(n75522), .B(n76498), .Y(n60230) );
  NAND2xp33_ASAP7_75t_SL U57704 ( .A(n57081), .B(n69730), .Y(n70506) );
  NAND2xp33_ASAP7_75t_SL U57705 ( .A(n60060), .B(n60174), .Y(n60067) );
  NAND2xp33_ASAP7_75t_SL U57706 ( .A(n60090), .B(n60174), .Y(n60097) );
  INVxp33_ASAP7_75t_SL U57707 ( .A(n64113), .Y(n62373) );
  OAI22xp33_ASAP7_75t_SL U57708 ( .A1(n59624), .A2(n72338), .B1(n72434), .B2(
        n72226), .Y(n72180) );
  NAND2xp5_ASAP7_75t_SL U57709 ( .A(n74779), .B(n74551), .Y(n75625) );
  NAND2xp33_ASAP7_75t_SL U57710 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .B(
        n72487), .Y(n71839) );
  NAND2xp33_ASAP7_75t_SL U57711 ( .A(n62682), .B(n75246), .Y(n75348) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57712 ( .A1(n74686), .A2(n74685), .B(n74684), .C(
        n74683), .Y(n74687) );
  INVxp33_ASAP7_75t_SL U57713 ( .A(n69736), .Y(n69587) );
  NAND2xp33_ASAP7_75t_SL U57714 ( .A(n2637), .B(n76557), .Y(n61124) );
  NAND2xp33_ASAP7_75t_SL U57715 ( .A(n72241), .B(n72514), .Y(n72376) );
  AOI21xp33_ASAP7_75t_SL U57716 ( .A1(n63743), .A2(n77866), .B(n60032), .Y(
        n60033) );
  NAND2xp33_ASAP7_75t_SL U57717 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_13_), .B(n69866), 
        .Y(n69858) );
  AOI22xp33_ASAP7_75t_SL U57718 ( .A1(n72126), .A2(n72103), .B1(n72105), .B2(
        n71965), .Y(n71969) );
  NAND2xp5_ASAP7_75t_SL U57719 ( .A(n73923), .B(n76782), .Y(n62353) );
  OAI21xp5_ASAP7_75t_SL U57720 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]), .A2(n65485), .B(
        n65666), .Y(n65663) );
  NAND2xp33_ASAP7_75t_SL U57721 ( .A(n69719), .B(n69720), .Y(n69595) );
  OAI22xp33_ASAP7_75t_SL U57722 ( .A1(n59622), .A2(n72418), .B1(n72245), .B2(
        n59623), .Y(n72236) );
  NAND2xp33_ASAP7_75t_SL U57723 ( .A(n71843), .B(n71842), .Y(n71852) );
  INVxp33_ASAP7_75t_SL U57724 ( .A(n76557), .Y(n61034) );
  INVxp33_ASAP7_75t_SL U57725 ( .A(n65601), .Y(n65603) );
  INVxp67_ASAP7_75t_SL U57726 ( .A(n76755), .Y(n61735) );
  NAND2xp33_ASAP7_75t_SL U57727 ( .A(n74231), .B(n74232), .Y(n74273) );
  AOI22xp33_ASAP7_75t_SL U57728 ( .A1(n72105), .A2(n72009), .B1(n72095), .B2(
        n71947), .Y(n71949) );
  INVx1_ASAP7_75t_SL U57729 ( .A(n75701), .Y(n64839) );
  OAI22xp33_ASAP7_75t_SL U57730 ( .A1(n72235), .A2(n72434), .B1(n59624), .B2(
        n72465), .Y(n72237) );
  INVxp33_ASAP7_75t_SL U57731 ( .A(n75590), .Y(n75592) );
  NAND2xp33_ASAP7_75t_SL U57732 ( .A(n71627), .B(n71574), .Y(n71613) );
  OAI21xp33_ASAP7_75t_SL U57733 ( .A1(n66217), .A2(n74834), .B(n74833), .Y(
        n66211) );
  INVx1_ASAP7_75t_SL U57734 ( .A(n62644), .Y(n58221) );
  INVx1_ASAP7_75t_SL U57735 ( .A(n69878), .Y(n69872) );
  INVxp33_ASAP7_75t_SL U57736 ( .A(n59971), .Y(n59972) );
  INVx1_ASAP7_75t_SL U57737 ( .A(n75838), .Y(n75591) );
  NAND2xp33_ASAP7_75t_SL U57738 ( .A(n78428), .B(n59629), .Y(n72749) );
  NAND2xp33_ASAP7_75t_SL U57739 ( .A(n65798), .B(n58419), .Y(n65683) );
  NOR2x1_ASAP7_75t_SL U57740 ( .A(n74368), .B(n74369), .Y(n74379) );
  INVxp67_ASAP7_75t_SL U57741 ( .A(n75705), .Y(n63570) );
  NAND2xp33_ASAP7_75t_SL U57742 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_18_), .B(n69682), 
        .Y(n69683) );
  INVxp67_ASAP7_75t_SL U57743 ( .A(n65389), .Y(n65390) );
  INVxp33_ASAP7_75t_SL U57744 ( .A(n69893), .Y(n69664) );
  OAI21xp33_ASAP7_75t_SL U57745 ( .A1(n73816), .A2(n73803), .B(n73802), .Y(
        n3296) );
  OAI22xp33_ASAP7_75t_SL U57746 ( .A1(n59624), .A2(n72418), .B1(n72245), .B2(
        n59622), .Y(n72189) );
  NAND2xp5_ASAP7_75t_SL U57747 ( .A(n69613), .B(n69775), .Y(n69783) );
  INVx1_ASAP7_75t_SL U57748 ( .A(n72491), .Y(n72436) );
  NAND2xp33_ASAP7_75t_SL U57749 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B(
        n70413), .Y(n70341) );
  INVx1_ASAP7_75t_SL U57750 ( .A(n65816), .Y(n65680) );
  INVxp33_ASAP7_75t_SL U57751 ( .A(n71367), .Y(n71371) );
  INVxp67_ASAP7_75t_SL U57752 ( .A(n69985), .Y(n69689) );
  NAND2xp33_ASAP7_75t_SL U57753 ( .A(n61598), .B(n61599), .Y(n60899) );
  INVx1_ASAP7_75t_SL U57754 ( .A(n74209), .Y(n74196) );
  INVxp33_ASAP7_75t_SL U57755 ( .A(n77062), .Y(n61503) );
  AOI21xp33_ASAP7_75t_SL U57756 ( .A1(n59580), .A2(n57122), .B(n62671), .Y(
        n62673) );
  INVx1_ASAP7_75t_SL U57757 ( .A(n76768), .Y(n77106) );
  OAI21xp5_ASAP7_75t_SL U57758 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .A2(
        n72039), .B(n71805), .Y(n72485) );
  OAI22xp33_ASAP7_75t_SL U57759 ( .A1(n70402), .A2(n70549), .B1(n74710), .B2(
        n70401), .Y(n70403) );
  INVxp67_ASAP7_75t_SL U57760 ( .A(n75245), .Y(n75840) );
  INVx1_ASAP7_75t_SL U57761 ( .A(n74331), .Y(n74286) );
  INVxp33_ASAP7_75t_SL U57762 ( .A(n69887), .Y(n69662) );
  AOI21xp5_ASAP7_75t_SL U57763 ( .A1(n63468), .A2(n63488), .B(n63486), .Y(
        n63469) );
  INVxp67_ASAP7_75t_SL U57764 ( .A(n76954), .Y(n74851) );
  INVxp67_ASAP7_75t_SL U57765 ( .A(n61746), .Y(n61677) );
  NAND2xp33_ASAP7_75t_SL U57766 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_22_), .B(n70068), 
        .Y(n70072) );
  OAI22xp33_ASAP7_75t_SL U57767 ( .A1(n59623), .A2(n72140), .B1(n59622), .B2(
        n72186), .Y(n72057) );
  INVxp33_ASAP7_75t_SL U57768 ( .A(n62362), .Y(n60800) );
  INVxp67_ASAP7_75t_SL U57769 ( .A(n70774), .Y(n70772) );
  INVxp67_ASAP7_75t_SL U57770 ( .A(n75588), .Y(n77075) );
  NAND2xp33_ASAP7_75t_SL U57771 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .B(
        n72440), .Y(n72078) );
  INVxp67_ASAP7_75t_SL U57772 ( .A(n70068), .Y(n69707) );
  OAI22xp33_ASAP7_75t_SL U57773 ( .A1(n59624), .A2(n72235), .B1(n72434), .B2(
        n72422), .Y(n72058) );
  NAND2xp5_ASAP7_75t_SL U57774 ( .A(n73705), .B(n73796), .Y(n73721) );
  OAI21xp33_ASAP7_75t_SL U57775 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[26]), .A2(n73874), .B(
        n3310), .Y(n73579) );
  NAND2xp33_ASAP7_75t_SL U57776 ( .A(n59558), .B(n62362), .Y(n61783) );
  AOI21xp33_ASAP7_75t_SL U57777 ( .A1(n74304), .A2(n74301), .B(n74333), .Y(
        n74335) );
  OAI22xp33_ASAP7_75t_SL U57778 ( .A1(n65786), .A2(n58418), .B1(n65785), .B2(
        n58571), .Y(n65790) );
  NAND2xp33_ASAP7_75t_SL U57779 ( .A(n72400), .B(n72153), .Y(n72077) );
  INVxp67_ASAP7_75t_SL U57780 ( .A(n70146), .Y(n70150) );
  OAI22xp33_ASAP7_75t_SL U57781 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_0_), .A2(n62059), .B1(n62064), 
        .B2(n62048), .Y(n2206) );
  INVxp33_ASAP7_75t_SL U57782 ( .A(n60311), .Y(n60424) );
  INVxp67_ASAP7_75t_SL U57783 ( .A(n69941), .Y(n70029) );
  NAND2xp33_ASAP7_75t_SL U57784 ( .A(n72241), .B(n72334), .Y(n72238) );
  INVxp67_ASAP7_75t_SL U57785 ( .A(n69798), .Y(n69828) );
  NAND2xp33_ASAP7_75t_SL U57786 ( .A(n78331), .B(n59629), .Y(n72883) );
  NAND2xp33_ASAP7_75t_SL U57787 ( .A(n72241), .B(n72487), .Y(n72273) );
  OAI22xp33_ASAP7_75t_SL U57788 ( .A1(n72479), .A2(n72503), .B1(n72507), .B2(
        n72453), .Y(n72454) );
  INVxp33_ASAP7_75t_SL U57789 ( .A(n69917), .Y(n69670) );
  NAND2xp5_ASAP7_75t_SL U57790 ( .A(n60861), .B(n76782), .Y(n64218) );
  INVxp67_ASAP7_75t_SL U57791 ( .A(n65827), .Y(n66040) );
  OAI22xp33_ASAP7_75t_SL U57792 ( .A1(n72200), .A2(n59622), .B1(n59624), .B2(
        n72270), .Y(n72081) );
  INVxp33_ASAP7_75t_SL U57793 ( .A(n72440), .Y(n71956) );
  NAND2xp5_ASAP7_75t_SL U57794 ( .A(n69713), .B(n70087), .Y(n70091) );
  INVxp33_ASAP7_75t_SL U57795 ( .A(n71505), .Y(n71429) );
  NAND2xp5_ASAP7_75t_SL U57796 ( .A(n73923), .B(n75731), .Y(n64295) );
  NAND2xp33_ASAP7_75t_SL U57797 ( .A(n65174), .B(n65170), .Y(n65180) );
  OAI22xp33_ASAP7_75t_SL U57798 ( .A1(n72235), .A2(n59623), .B1(n72434), .B2(
        n72186), .Y(n72190) );
  NAND2xp5_ASAP7_75t_SL U57799 ( .A(n71517), .B(n71516), .Y(n71521) );
  OAI21xp33_ASAP7_75t_SL U57800 ( .A1(n72532), .A2(n72531), .B(n72530), .Y(
        n72540) );
  NOR2x1_ASAP7_75t_SL U57801 ( .A(n65816), .B(n65827), .Y(n66022) );
  AOI21xp33_ASAP7_75t_SL U57802 ( .A1(n63320), .A2(n63319), .B(n63322), .Y(
        n63327) );
  NAND2xp5_ASAP7_75t_SL U57803 ( .A(n70168), .B(n70170), .Y(n70185) );
  INVxp67_ASAP7_75t_SL U57804 ( .A(n60934), .Y(n60598) );
  AOI21xp33_ASAP7_75t_SL U57805 ( .A1(n60647), .A2(n76753), .B(n60646), .Y(
        n60648) );
  INVxp67_ASAP7_75t_SL U57806 ( .A(n72470), .Y(n72192) );
  OAI22xp33_ASAP7_75t_SL U57807 ( .A1(n59622), .A2(n72226), .B1(n59624), .B2(
        n72220), .Y(n72036) );
  INVxp33_ASAP7_75t_SL U57808 ( .A(n65453), .Y(n65436) );
  NAND2xp5_ASAP7_75t_SL U57809 ( .A(n61133), .B(n77993), .Y(n75766) );
  NAND2xp5_ASAP7_75t_SL U57810 ( .A(n70158), .B(n70157), .Y(n70172) );
  OAI211xp5_ASAP7_75t_SRAM U57811 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[3]), .A2(n66157), .B(
        n65637), .C(n66161), .Y(n65638) );
  OAI22xp33_ASAP7_75t_SL U57812 ( .A1(or1200_cpu_or1200_mult_mac_n349), .A2(
        n61828), .B1(or1200_cpu_or1200_mult_mac_n66), .B2(n61826), .Y(n61837)
         );
  NAND2xp33_ASAP7_75t_SL U57813 ( .A(or1200_cpu_or1200_mult_mac_n255), .B(
        n75823), .Y(n64211) );
  NAND2xp33_ASAP7_75t_SL U57814 ( .A(n57081), .B(n70087), .Y(n70498) );
  INVxp67_ASAP7_75t_SL U57815 ( .A(n61598), .Y(n61478) );
  INVxp33_ASAP7_75t_SL U57816 ( .A(n69866), .Y(n69654) );
  AOI22xp33_ASAP7_75t_SL U57817 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .A2(
        n72298), .B1(n72400), .B2(n72228), .Y(n72037) );
  INVxp33_ASAP7_75t_SL U57818 ( .A(n77102), .Y(n61495) );
  OAI22xp33_ASAP7_75t_SL U57819 ( .A1(or1200_cpu_or1200_mult_mac_n347), .A2(
        n61828), .B1(or1200_cpu_or1200_mult_mac_n68), .B2(n61826), .Y(n75750)
         );
  NAND2xp33_ASAP7_75t_SL U57820 ( .A(n70286), .B(n70285), .Y(n70287) );
  OAI22xp33_ASAP7_75t_SL U57821 ( .A1(n59624), .A2(n72452), .B1(n59623), .B2(
        n72338), .Y(n72339) );
  OAI21xp33_ASAP7_75t_SL U57822 ( .A1(n57127), .A2(n72346), .B(n72345), .Y(
        n72480) );
  NAND2xp33_ASAP7_75t_SL U57823 ( .A(n74718), .B(n70413), .Y(n70414) );
  INVxp33_ASAP7_75t_SL U57824 ( .A(n70765), .Y(n70763) );
  NAND3xp33_ASAP7_75t_SRAM U57825 ( .A(n72403), .B(n72402), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .Y(
        n72406) );
  INVxp67_ASAP7_75t_SL U57826 ( .A(n71691), .Y(n71700) );
  INVxp33_ASAP7_75t_SL U57827 ( .A(n75240), .Y(n64222) );
  NAND2xp33_ASAP7_75t_SL U57828 ( .A(n60125), .B(n60174), .Y(n60131) );
  OAI22xp33_ASAP7_75t_SL U57829 ( .A1(n59624), .A2(n72337), .B1(n59622), .B2(
        n72220), .Y(n72136) );
  NAND2xp33_ASAP7_75t_SL U57830 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .B(
        n72322), .Y(n72407) );
  NAND2xp5_ASAP7_75t_SL U57831 ( .A(n65381), .B(n65423), .Y(n65450) );
  INVxp33_ASAP7_75t_SL U57832 ( .A(n62425), .Y(n62426) );
  NAND2xp5_ASAP7_75t_SL U57833 ( .A(n76339), .B(n64835), .Y(n64787) );
  AOI21xp33_ASAP7_75t_SL U57834 ( .A1(n73825), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .B(
        n73749), .Y(n73750) );
  AOI21xp5_ASAP7_75t_SL U57835 ( .A1(n65691), .A2(n76976), .B(n65690), .Y(
        n66060) );
  INVxp33_ASAP7_75t_SL U57836 ( .A(n70011), .Y(n69701) );
  NAND2xp33_ASAP7_75t_SL U57837 ( .A(n70358), .B(n70370), .Y(n70364) );
  INVx1_ASAP7_75t_SL U57838 ( .A(n63192), .Y(n58043) );
  NAND2xp5_ASAP7_75t_SL U57839 ( .A(n69693), .B(n70044), .Y(n70048) );
  OAI22xp33_ASAP7_75t_SL U57840 ( .A1(n72435), .A2(n59623), .B1(n72434), .B2(
        n72271), .Y(n72256) );
  OAI22xp33_ASAP7_75t_SL U57841 ( .A1(n72337), .A2(n72434), .B1(n59622), .B2(
        n72453), .Y(n72340) );
  NAND2xp5_ASAP7_75t_SL U57842 ( .A(n72527), .B(n72526), .Y(n72541) );
  NAND2xp33_ASAP7_75t_SL U57843 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_17_), .B(n69673), 
        .Y(n69674) );
  NAND2xp5_ASAP7_75t_SL U57844 ( .A(n63336), .B(n63335), .Y(n63350) );
  OAI22xp33_ASAP7_75t_SL U57845 ( .A1(n65792), .A2(n58582), .B1(n65791), .B2(
        n58418), .Y(n65795) );
  INVxp67_ASAP7_75t_SL U57846 ( .A(n70160), .Y(n70156) );
  OAI21xp33_ASAP7_75t_SL U57847 ( .A1(n3095), .A2(n77420), .B(n77419), .Y(
        n9388) );
  AOI22xp33_ASAP7_75t_SL U57848 ( .A1(n72126), .A2(n72044), .B1(n72105), .B2(
        n71911), .Y(n71915) );
  NAND2xp33_ASAP7_75t_SL U57849 ( .A(n72433), .B(n72213), .Y(n72167) );
  INVxp33_ASAP7_75t_SL U57850 ( .A(n72398), .Y(n72401) );
  OAI21xp5_ASAP7_75t_SL U57851 ( .A1(n76437), .A2(n75735), .B(n60981), .Y(
        n60982) );
  AND2x2_ASAP7_75t_SL U57852 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[22]), .B(n73047), .Y(n72685) );
  NAND2xp33_ASAP7_75t_SL U57853 ( .A(n72417), .B(n72374), .Y(n72323) );
  OAI21xp33_ASAP7_75t_SL U57854 ( .A1(n72147), .A2(n72084), .B(n58599), .Y(
        n71834) );
  OAI21xp33_ASAP7_75t_SL U57855 ( .A1(n3375), .A2(n77420), .B(n77419), .Y(
        n9387) );
  OAI21xp33_ASAP7_75t_SL U57856 ( .A1(n72113), .A2(n72112), .B(n72111), .Y(
        n72114) );
  NAND2xp33_ASAP7_75t_SL U57857 ( .A(n57561), .B(n75852), .Y(n75250) );
  NAND2xp33_ASAP7_75t_SL U57858 ( .A(n72093), .B(n72009), .Y(n71860) );
  INVx1_ASAP7_75t_SL U57859 ( .A(n70485), .Y(n70551) );
  INVx1_ASAP7_75t_SL U57860 ( .A(n71639), .Y(n71694) );
  NAND2xp5_ASAP7_75t_SL U57861 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[4]), .B(n73872), 
        .Y(n73545) );
  INVxp33_ASAP7_75t_SL U57862 ( .A(n75392), .Y(n75393) );
  NAND2xp33_ASAP7_75t_SL U57863 ( .A(n72093), .B(n71992), .Y(n71762) );
  NAND2xp5_ASAP7_75t_SL U57864 ( .A(n78184), .B(n77996), .Y(n4320) );
  NAND2xp33_ASAP7_75t_SL U57865 ( .A(n71642), .B(n71661), .Y(n71691) );
  NAND2xp33_ASAP7_75t_SL U57866 ( .A(n72286), .B(n72144), .Y(n72145) );
  NAND2xp5_ASAP7_75t_SL U57867 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_32_), .B(n59523), 
        .Y(n71170) );
  OAI22xp33_ASAP7_75t_SL U57868 ( .A1(n72119), .A2(n71979), .B1(n72067), .B2(
        n72050), .Y(n71829) );
  INVxp67_ASAP7_75t_SL U57869 ( .A(n61885), .Y(n60957) );
  NAND2xp5_ASAP7_75t_SL U57870 ( .A(n59861), .B(n75425), .Y(n59863) );
  NAND2xp5_ASAP7_75t_SL U57871 ( .A(n71702), .B(n71663), .Y(n71713) );
  INVx1_ASAP7_75t_SL U57872 ( .A(n77260), .Y(n60174) );
  NAND2xp5_ASAP7_75t_SL U57873 ( .A(n71743), .B(n71742), .Y(n71789) );
  OAI21xp33_ASAP7_75t_SL U57874 ( .A1(n3097), .A2(n61283), .B(n61282), .Y(
        n52472) );
  AOI22xp33_ASAP7_75t_SL U57875 ( .A1(n72390), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .B1(
        n71873), .B2(n72083), .Y(n72487) );
  INVxp33_ASAP7_75t_SL U57876 ( .A(n61310), .Y(n60505) );
  NAND2xp33_ASAP7_75t_SL U57877 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .B(
        n72354), .Y(n71805) );
  AOI22xp33_ASAP7_75t_SL U57878 ( .A1(n63742), .A2(n77257), .B1(n63741), .B2(
        n74956), .Y(n63746) );
  NAND2xp5_ASAP7_75t_SL U57879 ( .A(n59774), .B(n59782), .Y(n59781) );
  OAI22xp33_ASAP7_75t_SL U57880 ( .A1(n71588), .A2(n71462), .B1(n71461), .B2(
        n71460), .Y(n71463) );
  OAI21xp33_ASAP7_75t_SL U57881 ( .A1(n76460), .A2(n75735), .B(n61775), .Y(
        n61776) );
  OAI31xp33_ASAP7_75t_SRAM U57882 ( .A1(n2596), .A2(n69335), .A3(n60494), .B(
        n60493), .Y(n60496) );
  OAI22xp33_ASAP7_75t_SL U57883 ( .A1(n76764), .A2(n64769), .B1(n75700), .B2(
        n64768), .Y(n64770) );
  AOI21xp33_ASAP7_75t_SL U57884 ( .A1(n73825), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .B(
        n73804), .Y(n73805) );
  INVx1_ASAP7_75t_SL U57885 ( .A(n72583), .Y(n72585) );
  NAND2xp5_ASAP7_75t_SL U57886 ( .A(n71518), .B(n71520), .Y(n71516) );
  OAI21xp5_ASAP7_75t_SL U57887 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_4_), .A2(
        n72580), .B(n72596), .Y(n72581) );
  NAND2xp33_ASAP7_75t_SL U57888 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_16_), .B(n59523), 
        .Y(n70871) );
  INVx1_ASAP7_75t_SL U57889 ( .A(n61526), .Y(n61521) );
  NAND2xp33_ASAP7_75t_SL U57890 ( .A(n72534), .B(n72213), .Y(n72214) );
  INVxp67_ASAP7_75t_SL U57891 ( .A(n62356), .Y(n60660) );
  INVxp33_ASAP7_75t_SL U57892 ( .A(n71462), .Y(n71447) );
  NAND2xp33_ASAP7_75t_SL U57893 ( .A(n72433), .B(n72374), .Y(n72211) );
  NAND2xp33_ASAP7_75t_SL U57894 ( .A(n74213), .B(n66216), .Y(n74833) );
  AND2x2_ASAP7_75t_SRAM U57895 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[7]), .B(n73047), 
        .Y(n72771) );
  INVxp33_ASAP7_75t_SL U57896 ( .A(n75863), .Y(n75332) );
  OAI21xp33_ASAP7_75t_SL U57897 ( .A1(n72390), .A2(n72085), .B(n58599), .Y(
        n71957) );
  INVxp67_ASAP7_75t_SL U57898 ( .A(n64112), .Y(n60678) );
  OAI22xp33_ASAP7_75t_SL U57899 ( .A1(n72355), .A2(n72084), .B1(n72147), .B2(
        n72083), .Y(n71958) );
  INVx1_ASAP7_75t_SL U57900 ( .A(n77117), .Y(n62422) );
  NAND2xp33_ASAP7_75t_SL U57901 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_17_), .B(n71353), 
        .Y(n70889) );
  INVxp33_ASAP7_75t_SL U57902 ( .A(n74103), .Y(n74105) );
  OAI22xp33_ASAP7_75t_SL U57903 ( .A1(or1200_cpu_or1200_except_n242), .A2(
        n58547), .B1(n59548), .B2(n57124), .Y(n60026) );
  NAND2xp33_ASAP7_75t_SL U57904 ( .A(n62319), .B(n61242), .Y(n61598) );
  NAND2xp5_ASAP7_75t_SL U57905 ( .A(n71790), .B(n71682), .Y(n71786) );
  OAI22xp33_ASAP7_75t_SL U57906 ( .A1(n59624), .A2(n72140), .B1(n72422), .B2(
        n59622), .Y(n72470) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57907 ( .A1(n65327), .A2(n65326), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .C(n65325), .Y(
        n65329) );
  OAI21xp33_ASAP7_75t_SL U57908 ( .A1(n76791), .A2(n61364), .B(n61363), .Y(
        n61366) );
  OAI21xp33_ASAP7_75t_SL U57909 ( .A1(n74119), .A2(n59860), .B(n59859), .Y(
        n75426) );
  INVxp33_ASAP7_75t_SL U57910 ( .A(n69681), .Y(n69682) );
  OAI21xp33_ASAP7_75t_SL U57911 ( .A1(n76434), .A2(n75735), .B(n62427), .Y(
        n62428) );
  NAND2xp33_ASAP7_75t_SL U57912 ( .A(n62205), .B(n62204), .Y(n62206) );
  AOI22xp33_ASAP7_75t_SL U57913 ( .A1(n72105), .A2(n72091), .B1(n72126), .B2(
        n72090), .Y(n72097) );
  INVxp33_ASAP7_75t_SL U57914 ( .A(n68810), .Y(n68811) );
  INVxp67_ASAP7_75t_SL U57915 ( .A(n62420), .Y(n62421) );
  OAI22xp33_ASAP7_75t_SL U57916 ( .A1(or1200_cpu_or1200_except_n222), .A2(
        n58547), .B1(n59536), .B2(n57124), .Y(n60110) );
  AOI211xp5_ASAP7_75t_SL U57917 ( .A1(n59879), .A2(n59878), .B(n78001), .C(
        n60582), .Y(n60199) );
  NAND2xp33_ASAP7_75t_SL U57918 ( .A(n78333), .B(n73047), .Y(n72854) );
  OAI21xp33_ASAP7_75t_SL U57919 ( .A1(n72068), .A2(n72067), .B(n72066), .Y(
        n72071) );
  NAND2xp33_ASAP7_75t_SL U57920 ( .A(n72093), .B(n72047), .Y(n72048) );
  AO21x1_ASAP7_75t_SRAM U57921 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]), .A2(n65500), .B(
        n74894), .Y(n65501) );
  NAND2xp5_ASAP7_75t_SL U57922 ( .A(n69591), .B(n69592), .Y(n69723) );
  NAND2xp33_ASAP7_75t_SL U57923 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_0_), .B(n69718), .Y(
        n69719) );
  INVxp33_ASAP7_75t_SL U57924 ( .A(n69679), .Y(n69673) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57925 ( .A1(n61186), .A2(n61185), .B(n59443), .C(
        n61184), .Y(n61187) );
  AOI22xp33_ASAP7_75t_SL U57926 ( .A1(n72126), .A2(n72045), .B1(n72105), .B2(
        n72044), .Y(n72049) );
  OAI21xp33_ASAP7_75t_SL U57927 ( .A1(n76462), .A2(n75735), .B(n74600), .Y(
        n74602) );
  INVxp67_ASAP7_75t_SL U57928 ( .A(n64078), .Y(n64080) );
  NAND2xp5_ASAP7_75t_SL U57929 ( .A(n66189), .B(n66188), .Y(n74140) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U57930 ( .A1(n76382), .A2(n76381), .B(n76380), 
        .C(n76379), .Y(n76392) );
  OAI22xp33_ASAP7_75t_SL U57931 ( .A1(or1200_cpu_or1200_except_n240), .A2(
        n58547), .B1(n1571), .B2(n57124), .Y(n60032) );
  INVxp33_ASAP7_75t_SL U57932 ( .A(n69446), .Y(n69742) );
  NAND2xp33_ASAP7_75t_SL U57933 ( .A(n65674), .B(n65676), .Y(n65639) );
  NAND2xp5_ASAP7_75t_SL U57934 ( .A(n69612), .B(n69611), .Y(n69775) );
  AND2x2_ASAP7_75t_SL U57935 ( .A(n58084), .B(n75708), .Y(n58082) );
  INVxp33_ASAP7_75t_SL U57936 ( .A(n76387), .Y(n76388) );
  OAI21xp33_ASAP7_75t_SL U57937 ( .A1(n76399), .A2(n76398), .B(n76397), .Y(
        n76401) );
  INVxp33_ASAP7_75t_SL U57938 ( .A(n69612), .Y(n69600) );
  NAND2xp5_ASAP7_75t_SL U57939 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]), .B(n65485), .Y(
        n65666) );
  NAND2xp33_ASAP7_75t_SL U57940 ( .A(n72126), .B(n72118), .Y(n72028) );
  INVxp67_ASAP7_75t_SL U57941 ( .A(n62208), .Y(n62210) );
  INVxp33_ASAP7_75t_SL U57942 ( .A(n65676), .Y(n66088) );
  NAND2xp33_ASAP7_75t_SL U57943 ( .A(n72095), .B(n72025), .Y(n72026) );
  INVxp33_ASAP7_75t_SL U57944 ( .A(n69627), .Y(n69628) );
  OAI21xp33_ASAP7_75t_SL U57945 ( .A1(n3376), .A2(n61283), .B(n61282), .Y(
        n52473) );
  INVxp33_ASAP7_75t_SL U57946 ( .A(n72050), .Y(n71912) );
  NAND2xp33_ASAP7_75t_SL U57947 ( .A(n72126), .B(n72072), .Y(n71930) );
  AOI22xp33_ASAP7_75t_SL U57948 ( .A1(n72062), .A2(n72061), .B1(n72110), .B2(
        n72060), .Y(n72063) );
  AOI22xp33_ASAP7_75t_SL U57949 ( .A1(n72105), .A2(n71992), .B1(n72095), .B2(
        n71927), .Y(n71929) );
  INVxp67_ASAP7_75t_SL U57950 ( .A(n61845), .Y(n61844) );
  INVxp33_ASAP7_75t_SL U57951 ( .A(n61305), .Y(n61306) );
  NAND2xp5_ASAP7_75t_SL U57952 ( .A(n72043), .B(n72042), .Y(n72384) );
  OAI21xp33_ASAP7_75t_SL U57953 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n70462), .B(n70400), .Y(n70549) );
  INVxp67_ASAP7_75t_SL U57954 ( .A(n74055), .Y(n66212) );
  INVxp67_ASAP7_75t_SL U57955 ( .A(n71946), .Y(n71947) );
  NAND2xp33_ASAP7_75t_SL U57956 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_40_), .B(n71353), 
        .Y(n71265) );
  INVx2_ASAP7_75t_SL U57957 ( .A(n58609), .Y(n57189) );
  AND3x1_ASAP7_75t_SL U57958 ( .A(n77348), .B(ic_en), .C(n77833), .Y(n60282)
         );
  OAI21xp33_ASAP7_75t_SL U57959 ( .A1(n76464), .A2(n75735), .B(n64122), .Y(
        n64123) );
  AOI22xp33_ASAP7_75t_SL U57960 ( .A1(n72126), .A2(n72091), .B1(n72093), .B2(
        n72094), .Y(n71948) );
  INVx1_ASAP7_75t_SL U57961 ( .A(n77031), .Y(n73953) );
  NAND2xp33_ASAP7_75t_SL U57962 ( .A(n72645), .B(n72644), .Y(n72648) );
  INVxp33_ASAP7_75t_SL U57963 ( .A(n72025), .Y(n71965) );
  NAND2xp33_ASAP7_75t_SL U57964 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_42_), .B(n71353), 
        .Y(n71323) );
  OAI22xp33_ASAP7_75t_SL U57965 ( .A1(n77254), .A2(n77615), .B1(n59580), .B2(
        n57124), .Y(n74949) );
  NAND2xp33_ASAP7_75t_SL U57966 ( .A(n78335), .B(n73047), .Y(n72841) );
  INVx1_ASAP7_75t_SL U57967 ( .A(n70476), .Y(n70553) );
  AOI22xp33_ASAP7_75t_SL U57968 ( .A1(n72116), .A2(n72090), .B1(n72062), .B2(
        n71943), .Y(n71944) );
  INVxp33_ASAP7_75t_SL U57969 ( .A(n72086), .Y(n71942) );
  INVxp33_ASAP7_75t_SL U57970 ( .A(n72068), .Y(n71924) );
  INVx1_ASAP7_75t_SL U57971 ( .A(n75735), .Y(n64835) );
  NAND2xp5_ASAP7_75t_SL U57972 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_43_), .B(n59523), 
        .Y(n71367) );
  INVxp33_ASAP7_75t_SL U57973 ( .A(n72059), .Y(n71923) );
  INVxp33_ASAP7_75t_SL U57974 ( .A(n60325), .Y(n60326) );
  INVxp67_ASAP7_75t_SL U57975 ( .A(n75316), .Y(n77088) );
  NAND2xp5_ASAP7_75t_SL U57976 ( .A(n77354), .B(n77311), .Y(n77353) );
  OAI21xp33_ASAP7_75t_SL U57977 ( .A1(n72108), .A2(n72112), .B(n71889), .Y(
        n72170) );
  OAI21xp33_ASAP7_75t_SL U57978 ( .A1(n72086), .A2(n72112), .B(n71850), .Y(
        n71851) );
  NAND2xp5_ASAP7_75t_SL U57979 ( .A(n69712), .B(n69711), .Y(n70087) );
  INVxp33_ASAP7_75t_SL U57980 ( .A(n61726), .Y(n61504) );
  OAI21xp33_ASAP7_75t_SL U57981 ( .A1(n72068), .A2(n72085), .B(n71756), .Y(
        n71757) );
  NAND2xp33_ASAP7_75t_SL U57982 ( .A(n59550), .B(n57504), .Y(n66248) );
  NAND2xp5_ASAP7_75t_SL U57983 ( .A(n69703), .B(n69704), .Y(n70044) );
  INVxp33_ASAP7_75t_SL U57984 ( .A(n66157), .Y(n65626) );
  BUFx2_ASAP7_75t_SL U57985 ( .A(n63654), .Y(n57316) );
  OAI22xp33_ASAP7_75t_SL U57986 ( .A1(or1200_cpu_or1200_except_n220), .A2(
        n58547), .B1(n57312), .B2(n57124), .Y(n60117) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U57987 ( .A1(n73752), .A2(n73789), .B(n73699), .C(
        n73770), .Y(n73700) );
  OAI22xp33_ASAP7_75t_SL U57988 ( .A1(n59582), .A2(n57124), .B1(n77673), .B2(
        n77254), .Y(n59997) );
  NAND2xp33_ASAP7_75t_SL U57989 ( .A(n65841), .B(n65840), .Y(n65842) );
  AOI22xp33_ASAP7_75t_SL U57990 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_3_), .A2(
        n70485), .B1(n70476), .B2(n74674), .Y(n70460) );
  AOI22xp33_ASAP7_75t_SL U57991 ( .A1(n70539), .A2(n70462), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B2(
        n70461), .Y(n70463) );
  OAI22xp33_ASAP7_75t_SL U57992 ( .A1(n65788), .A2(n58419), .B1(n65787), .B2(
        n58582), .Y(n65789) );
  OAI21xp33_ASAP7_75t_SL U57993 ( .A1(n75817), .A2(n75691), .B(n75690), .Y(
        n75694) );
  NAND2xp5_ASAP7_75t_SL U57994 ( .A(n69581), .B(n69445), .Y(n69941) );
  AOI21xp33_ASAP7_75t_SL U57995 ( .A1(n74956), .A2(n76825), .B(
        or1200_cpu_or1200_genpc_pcreg_default[7]), .Y(n63734) );
  NAND2xp5_ASAP7_75t_SL U57996 ( .A(n76553), .B(n61772), .Y(n62444) );
  NAND2xp33_ASAP7_75t_SL U57997 ( .A(n73814), .B(n73811), .Y(n73777) );
  INVxp67_ASAP7_75t_SL U57998 ( .A(n72529), .Y(n72526) );
  AOI22xp33_ASAP7_75t_SL U57999 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .A2(
        n70485), .B1(n70476), .B2(n70354), .Y(n70351) );
  NAND2xp33_ASAP7_75t_SL U58000 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_2_), .B(
        n72529), .Y(n72530) );
  AOI22xp33_ASAP7_75t_SL U58001 ( .A1(n1131), .A2(n75689), .B1(n1436), .B2(
        n75203), .Y(n64210) );
  AOI22xp33_ASAP7_75t_SL U58002 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n70339), .B1(n70373), .B2(n74706), .Y(n70416) );
  NAND2xp33_ASAP7_75t_SL U58003 ( .A(n74512), .B(n2934), .Y(n74514) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58004 ( .A1(n70412), .A2(n70411), .B(n70539), .C(
        n70410), .Y(n70415) );
  NAND2xp5_ASAP7_75t_SL U58005 ( .A(n74706), .B(n70301), .Y(n70413) );
  AOI21xp33_ASAP7_75t_SL U58006 ( .A1(n73781), .A2(n73780), .B(n73779), .Y(
        n73782) );
  AOI22xp33_ASAP7_75t_SL U58007 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_7_), .A2(
        n70476), .B1(n70485), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_6_), .Y(
        n70417) );
  OAI21xp33_ASAP7_75t_SL U58008 ( .A1(n76432), .A2(n75735), .B(n61100), .Y(
        n61102) );
  NAND2xp33_ASAP7_75t_SL U58009 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_3_), .B(n59523), .Y(
        n70699) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58010 ( .A1(n65808), .A2(n65758), .B(n65757), .C(
        n65841), .Y(n65759) );
  AOI22xp33_ASAP7_75t_SL U58011 ( .A1(n1129), .A2(n75689), .B1(n1434), .B2(
        n75203), .Y(n64818) );
  INVxp67_ASAP7_75t_SL U58012 ( .A(n72543), .Y(n72549) );
  NAND2xp5_ASAP7_75t_SL U58013 ( .A(n63353), .B(n63355), .Y(n63354) );
  NOR2x1_ASAP7_75t_SL U58014 ( .A(n75872), .B(n75227), .Y(n77097) );
  AOI21xp33_ASAP7_75t_SL U58015 ( .A1(n70485), .A2(n2442), .B(n74718), .Y(
        n70374) );
  OAI21xp33_ASAP7_75t_SL U58016 ( .A1(n76448), .A2(n75735), .B(n62113), .Y(
        n62115) );
  INVxp67_ASAP7_75t_SL U58017 ( .A(n60620), .Y(n60621) );
  INVxp33_ASAP7_75t_SL U58018 ( .A(n65781), .Y(n65701) );
  AOI21xp33_ASAP7_75t_SL U58019 ( .A1(n73771), .A2(n73752), .B(n73723), .Y(
        n73803) );
  NAND2xp33_ASAP7_75t_SL U58020 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .B(
        n73826), .Y(n73759) );
  NAND2xp5_ASAP7_75t_SL U58021 ( .A(n63328), .B(n63318), .Y(n63317) );
  AOI22xp33_ASAP7_75t_SL U58022 ( .A1(n70539), .A2(n70431), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .B2(
        n70430), .Y(n70434) );
  NAND2xp33_ASAP7_75t_SL U58023 ( .A(n65681), .B(n65841), .Y(n65798) );
  NAND2xp33_ASAP7_75t_SL U58024 ( .A(n73814), .B(n73807), .Y(n73762) );
  AOI22xp33_ASAP7_75t_SL U58025 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_), .A2(
        n70476), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_16_), .B2(
        n70485), .Y(n70322) );
  NAND2xp5_ASAP7_75t_SL U58026 ( .A(n59763), .B(n59771), .Y(n59770) );
  NAND2xp33_ASAP7_75t_SL U58027 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_6_), .B(n71353), .Y(
        n70742) );
  NOR2x1_ASAP7_75t_SL U58028 ( .A(n77943), .B(n60557), .Y(n75452) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58029 ( .A1(n59706), .A2(n77775), .B(n1337), .C(
        n77774), .Y(n77777) );
  NAND2xp33_ASAP7_75t_SL U58030 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_8_), .B(n59523), .Y(
        n70765) );
  INVxp33_ASAP7_75t_SL U58031 ( .A(n70233), .Y(n70219) );
  INVx1_ASAP7_75t_SL U58032 ( .A(n70550), .Y(n70370) );
  INVx1_ASAP7_75t_SL U58033 ( .A(n70033), .Y(n70062) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58034 ( .A1(n65831), .A2(n65830), .B(n65829), 
        .C(n65828), .Y(n65836) );
  INVxp67_ASAP7_75t_SL U58035 ( .A(n70548), .Y(n70333) );
  NAND2xp33_ASAP7_75t_SL U58036 ( .A(n78352), .B(n73047), .Y(n72748) );
  INVxp33_ASAP7_75t_SL U58037 ( .A(n76751), .Y(n75220) );
  NAND2xp33_ASAP7_75t_SL U58038 ( .A(n74799), .B(n74798), .Y(n1504) );
  NAND2xp33_ASAP7_75t_SL U58039 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_9_), .B(n71353), .Y(
        n70774) );
  NOR2xp33_ASAP7_75t_SRAM U58040 ( .A(n59575), .B(n75714), .Y(n61872) );
  OAI22xp33_ASAP7_75t_SL U58041 ( .A1(n61878), .A2(n61877), .B1(n61876), .B2(
        n61875), .Y(n75586) );
  INVxp33_ASAP7_75t_SL U58042 ( .A(n4318), .Y(n77492) );
  NAND2xp5_ASAP7_75t_SL U58043 ( .A(n61857), .B(n77065), .Y(n62133) );
  OAI21xp33_ASAP7_75t_SL U58044 ( .A1(n76341), .A2(n75735), .B(n75721), .Y(
        n75725) );
  AOI21xp5_ASAP7_75t_SL U58045 ( .A1(n63542), .A2(n63533), .B(n63540), .Y(
        n63515) );
  OAI21xp5_ASAP7_75t_SL U58046 ( .A1(n62012), .A2(n75507), .B(n60643), .Y(
        n76753) );
  NAND2xp33_ASAP7_75t_SL U58047 ( .A(n59625), .B(n72374), .Y(n72402) );
  NAND2xp33_ASAP7_75t_SL U58048 ( .A(n70327), .B(n70476), .Y(n70278) );
  OAI21xp33_ASAP7_75t_SL U58049 ( .A1(n77594), .A2(n77254), .B(n61568), .Y(
        n61572) );
  NAND2xp33_ASAP7_75t_SL U58050 ( .A(n72417), .B(n72213), .Y(n72403) );
  NAND2xp33_ASAP7_75t_SL U58051 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .B(
        n70485), .Y(n70277) );
  OAI21xp33_ASAP7_75t_SL U58052 ( .A1(n73788), .A2(n73765), .B(n73764), .Y(
        n73766) );
  INVx1_ASAP7_75t_SL U58053 ( .A(n61918), .Y(n61963) );
  INVx1_ASAP7_75t_SL U58054 ( .A(n75836), .Y(n60857) );
  OAI21xp5_ASAP7_75t_SL U58055 ( .A1(n74894), .A2(n65674), .B(n65673), .Y(
        n65816) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58056 ( .A1(n72516), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_), 
        .B(n72344), .C(n72343), .Y(n72345) );
  NAND2xp33_ASAP7_75t_SL U58057 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[18]), .B(n73047), .Y(n72701) );
  INVxp67_ASAP7_75t_SL U58058 ( .A(n70450), .Y(n70365) );
  INVxp33_ASAP7_75t_SL U58059 ( .A(n75227), .Y(n76773) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58060 ( .A1(n65822), .A2(n65808), .B(n65698), .C(
        n65841), .Y(n65700) );
  INVxp67_ASAP7_75t_SL U58061 ( .A(n77370), .Y(n75765) );
  INVx1_ASAP7_75t_SL U58062 ( .A(n75325), .Y(n76766) );
  AOI21xp33_ASAP7_75t_SL U58063 ( .A1(n69419), .A2(n78357), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_20_), .Y(n69420) );
  INVxp67_ASAP7_75t_SL U58064 ( .A(n70383), .Y(n70470) );
  NAND2xp5_ASAP7_75t_SL U58065 ( .A(n70167), .B(n70166), .Y(n70170) );
  OAI21xp33_ASAP7_75t_SL U58066 ( .A1(n73789), .A2(n73788), .B(n73787), .Y(
        n73794) );
  AOI22xp33_ASAP7_75t_SL U58067 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_5_), .A2(
        n70476), .B1(n70485), .B2(n74674), .Y(n70443) );
  INVxp33_ASAP7_75t_SL U58068 ( .A(n71580), .Y(n71609) );
  AOI21xp5_ASAP7_75t_SL U58069 ( .A1(n65676), .A2(n76976), .B(n65675), .Y(
        n65827) );
  NAND2xp33_ASAP7_75t_SL U58070 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .B(
        n70485), .Y(n70286) );
  OAI21xp33_ASAP7_75t_SL U58071 ( .A1(n76459), .A2(n75735), .B(n62526), .Y(
        n62528) );
  OAI21xp33_ASAP7_75t_SL U58072 ( .A1(n70136), .A2(n70135), .B(n70134), .Y(
        n70145) );
  OAI21xp5_ASAP7_75t_SL U58073 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .A2(n57123), .B(n71919), .Y(n72228) );
  INVxp33_ASAP7_75t_SL U58074 ( .A(n70426), .Y(n70404) );
  NAND2xp33_ASAP7_75t_SL U58075 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .B(
        n70476), .Y(n70285) );
  OAI21xp33_ASAP7_75t_SL U58076 ( .A1(or1200_cpu_or1200_mult_mac_n191), .A2(
        n75723), .B(n64238), .Y(n64239) );
  NAND2xp33_ASAP7_75t_SL U58077 ( .A(n78349), .B(n73047), .Y(n72810) );
  NAND2xp33_ASAP7_75t_SL U58078 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B(
        n70432), .Y(n70433) );
  AND2x2_ASAP7_75t_SRAM U58079 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[20]), .B(n73047), .Y(n72683) );
  OAI22xp33_ASAP7_75t_SL U58080 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .A2(
        n72113), .B1(n72411), .B2(n71873), .Y(n72514) );
  AND2x2_ASAP7_75t_SL U58081 ( .A(n59625), .B(n72213), .Y(n72023) );
  NAND2xp33_ASAP7_75t_SL U58082 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_2_), .B(n71353), .Y(
        n70701) );
  AOI22xp33_ASAP7_75t_SL U58083 ( .A1(n61270), .A2(n77257), .B1(n61269), .B2(
        n74956), .Y(n61274) );
  NAND2xp5_ASAP7_75t_SL U58084 ( .A(n63324), .B(n63326), .Y(n63320) );
  NAND2xp5_ASAP7_75t_SL U58085 ( .A(n62067), .B(n62049), .Y(n62062) );
  NAND2xp33_ASAP7_75t_SL U58086 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[21]), .B(n73047), .Y(n72682) );
  NAND2xp33_ASAP7_75t_SL U58087 ( .A(n73814), .B(n73812), .Y(n73784) );
  INVxp67_ASAP7_75t_SL U58088 ( .A(n58000), .Y(n57999) );
  OAI21xp33_ASAP7_75t_SL U58089 ( .A1(n70359), .A2(n74706), .B(n70362), .Y(
        n70447) );
  NAND2xp33_ASAP7_75t_SL U58090 ( .A(n72105), .B(n71913), .Y(n71825) );
  INVxp33_ASAP7_75t_SL U58091 ( .A(n72146), .Y(n72060) );
  NAND2xp33_ASAP7_75t_SL U58092 ( .A(n1337), .B(n77775), .Y(n77774) );
  NAND2xp33_ASAP7_75t_SL U58093 ( .A(n71659), .B(n71641), .Y(n71642) );
  OAI22xp33_ASAP7_75t_SL U58094 ( .A1(n72112), .A2(n72084), .B1(n72085), .B2(
        n72087), .Y(n72003) );
  NAND2xp5_ASAP7_75t_SL U58095 ( .A(n61816), .B(n61827), .Y(n61818) );
  AOI21xp5_ASAP7_75t_SL U58096 ( .A1(n73518), .A2(n73517), .B(n73706), .Y(
        n73519) );
  INVxp33_ASAP7_75t_SL U58097 ( .A(n77417), .Y(n77420) );
  NAND2xp33_ASAP7_75t_SL U58098 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_11_), .B(n69632), 
        .Y(n69633) );
  INVxp33_ASAP7_75t_SL U58099 ( .A(n69574), .Y(n69576) );
  INVxp33_ASAP7_75t_SL U58100 ( .A(n75853), .Y(n77057) );
  NOR2xp33_ASAP7_75t_SRAM U58101 ( .A(n77278), .B(n63571), .Y(n60862) );
  NAND2xp5_ASAP7_75t_SL U58102 ( .A(n60334), .B(n60341), .Y(n60497) );
  NAND2xp33_ASAP7_75t_SL U58103 ( .A(n65513), .B(n66145), .Y(n65518) );
  INVxp33_ASAP7_75t_SL U58104 ( .A(n77850), .Y(n77842) );
  NAND2xp5_ASAP7_75t_SL U58105 ( .A(n59571), .B(n62615), .Y(n62616) );
  INVxp67_ASAP7_75t_SL U58106 ( .A(n66217), .Y(n66218) );
  INVxp33_ASAP7_75t_SL U58107 ( .A(n71661), .Y(n71695) );
  OAI21xp33_ASAP7_75t_SL U58108 ( .A1(n72399), .A2(n72224), .B(n72434), .Y(
        n72225) );
  INVxp67_ASAP7_75t_SL U58109 ( .A(n75687), .Y(n64207) );
  NAND2xp33_ASAP7_75t_SL U58110 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_9_), .B(n69622), .Y(
        n69623) );
  NAND2xp33_ASAP7_75t_SL U58111 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .B(
        n73835), .Y(n73674) );
  NAND2xp5_ASAP7_75t_SL U58112 ( .A(n74827), .B(n74738), .Y(n76985) );
  AOI21xp33_ASAP7_75t_SL U58113 ( .A1(n73786), .A2(n73778), .B(n73793), .Y(
        n73783) );
  NAND2xp33_ASAP7_75t_SL U58114 ( .A(n2609), .B(n60492), .Y(n60339) );
  OAI21xp5_ASAP7_75t_SL U58115 ( .A1(n78166), .A2(n77686), .B(n58421), .Y(
        n4317) );
  INVxp33_ASAP7_75t_SL U58116 ( .A(n71469), .Y(n71440) );
  OAI211xp5_ASAP7_75t_SRAM U58117 ( .A1(n65391), .A2(n65348), .B(n65347), .C(
        n65346), .Y(n65349) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58118 ( .A1(n71662), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_4_), .B(
        n71661), .C(n71660), .Y(n71663) );
  NAND2xp33_ASAP7_75t_SL U58119 ( .A(n65082), .B(n65089), .Y(n65085) );
  NOR2xp33_ASAP7_75t_SRAM U58120 ( .A(n58421), .B(n77496), .Y(n77499) );
  OAI22xp33_ASAP7_75t_SL U58121 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .A2(n57123), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_10_), 
        .B2(n57127), .Y(n72246) );
  AOI211xp5_ASAP7_75t_SRAM U58122 ( .A1(n74723), .A2(n74708), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .C(
        n74713), .Y(n74704) );
  NAND2xp33_ASAP7_75t_SL U58123 ( .A(n65210), .B(n77257), .Y(n60038) );
  INVx1_ASAP7_75t_SL U58124 ( .A(n72224), .Y(n72298) );
  NAND2xp33_ASAP7_75t_SL U58125 ( .A(n72126), .B(n72094), .Y(n71853) );
  NAND2xp33_ASAP7_75t_SL U58126 ( .A(n60554), .B(n60552), .Y(n61845) );
  NAND2xp33_ASAP7_75t_SL U58127 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .B(
        n73820), .Y(n73799) );
  AOI21xp33_ASAP7_75t_SL U58128 ( .A1(n71631), .A2(n71630), .B(n71553), .Y(
        n71554) );
  AOI22xp33_ASAP7_75t_SL U58129 ( .A1(n72116), .A2(n72041), .B1(n72110), .B2(
        n72040), .Y(n72042) );
  AOI21xp33_ASAP7_75t_SL U58130 ( .A1(n73822), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .B(
        n73801), .Y(n73802) );
  NAND2xp33_ASAP7_75t_SL U58131 ( .A(n72286), .B(n72109), .Y(n71975) );
  NAND2xp33_ASAP7_75t_SL U58132 ( .A(n77943), .B(n60556), .Y(n60558) );
  NAND3xp33_ASAP7_75t_SRAM U58133 ( .A(n72502), .B(n71937), .C(n72499), .Y(
        n71781) );
  NAND2xp5_ASAP7_75t_SL U58134 ( .A(n77338), .B(n77348), .Y(n4152) );
  NAND2xp33_ASAP7_75t_SL U58135 ( .A(n75846), .B(n53430), .Y(n61814) );
  NAND2xp5_ASAP7_75t_SL U58136 ( .A(n62203), .B(n75405), .Y(n62208) );
  INVxp33_ASAP7_75t_SL U58137 ( .A(n66115), .Y(n65604) );
  NAND2xp33_ASAP7_75t_SL U58138 ( .A(n62319), .B(n75687), .Y(n61132) );
  INVxp67_ASAP7_75t_SL U58139 ( .A(n61628), .Y(n61449) );
  NAND2xp5_ASAP7_75t_SL U58140 ( .A(n78245), .B(n62066), .Y(n62049) );
  NAND2xp33_ASAP7_75t_SL U58141 ( .A(n73786), .B(n73785), .Y(n73787) );
  NAND2xp33_ASAP7_75t_SL U58142 ( .A(n72110), .B(n72117), .Y(n72019) );
  NAND2xp5_ASAP7_75t_SL U58143 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_1_), .B(
        n71649), .Y(n71682) );
  INVx1_ASAP7_75t_SL U58144 ( .A(n65486), .Y(n65485) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58145 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .A2(n72367), .B(n72517), .C(n71951), .Y(n71864) );
  INVxp33_ASAP7_75t_SL U58146 ( .A(n72285), .Y(n72287) );
  NAND3xp33_ASAP7_75t_SRAM U58147 ( .A(n75507), .B(n75506), .C(n75505), .Y(
        n75510) );
  OAI22xp33_ASAP7_75t_SL U58148 ( .A1(n57125), .A2(n72164), .B1(n72163), .B2(
        n57123), .Y(n72165) );
  NAND2xp33_ASAP7_75t_SL U58149 ( .A(n72286), .B(n72090), .Y(n72274) );
  NAND2xp33_ASAP7_75t_SL U58150 ( .A(n72105), .B(n71966), .Y(n71901) );
  NAND2xp33_ASAP7_75t_SL U58151 ( .A(n72116), .B(n72065), .Y(n71756) );
  NAND2xp5_ASAP7_75t_SL U58152 ( .A(n71497), .B(n71631), .Y(n71580) );
  INVx1_ASAP7_75t_SL U58153 ( .A(n77066), .Y(n75852) );
  INVxp33_ASAP7_75t_SL U58154 ( .A(n72045), .Y(n71818) );
  AOI22xp33_ASAP7_75t_SL U58155 ( .A1(n77696), .A2(n77253), .B1(n63743), .B2(
        n77992), .Y(n61272) );
  INVx1_ASAP7_75t_SL U58156 ( .A(n75689), .Y(n75818) );
  NOR2x1_ASAP7_75t_SL U58157 ( .A(n77410), .B(n78166), .Y(n77996) );
  NAND2xp5_ASAP7_75t_SL U58158 ( .A(n70218), .B(n70237), .Y(n70233) );
  INVx1_ASAP7_75t_SL U58159 ( .A(n77340), .Y(n77305) );
  OAI21xp33_ASAP7_75t_SL U58160 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .A2(
        n71898), .B(n71816), .Y(n72044) );
  OAI22xp33_ASAP7_75t_SL U58161 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .A2(
        n70382), .B1(n70350), .B2(n70349), .Y(n70432) );
  AOI21xp5_ASAP7_75t_SL U58162 ( .A1(n74019), .A2(n76406), .B(n76410), .Y(
        n74020) );
  NAND2xp33_ASAP7_75t_SL U58163 ( .A(n72062), .B(n72038), .Y(n71814) );
  NAND2xp33_ASAP7_75t_SL U58164 ( .A(n73786), .B(n73763), .Y(n73764) );
  OAI22xp33_ASAP7_75t_SL U58165 ( .A1(n57125), .A2(n72318), .B1(n72317), .B2(
        n57123), .Y(n72291) );
  NAND2xp33_ASAP7_75t_SL U58166 ( .A(n72987), .B(n73011), .Y(n72719) );
  INVxp67_ASAP7_75t_SL U58167 ( .A(n72120), .Y(n72121) );
  OAI21xp33_ASAP7_75t_SL U58168 ( .A1(n70399), .A2(n70398), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .Y(
        n70400) );
  NAND2xp5_ASAP7_75t_SL U58169 ( .A(n74894), .B(n74747), .Y(n74203) );
  OAI21xp33_ASAP7_75t_SL U58170 ( .A1(n72341), .A2(n72367), .B(n57123), .Y(
        n72344) );
  INVxp67_ASAP7_75t_SL U58171 ( .A(n72103), .Y(n72107) );
  NAND2xp33_ASAP7_75t_SL U58172 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B(
        n70401), .Y(n70547) );
  AOI22xp33_ASAP7_75t_SL U58173 ( .A1(n73663), .A2(n73772), .B1(n73662), .B2(
        n73771), .Y(n73630) );
  AOI22xp33_ASAP7_75t_SL U58174 ( .A1(n73786), .A2(n73754), .B1(n73785), .B2(
        n73780), .Y(n73760) );
  OAI22xp33_ASAP7_75t_SL U58175 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .A2(
        n73789), .B1(n73752), .B2(n73751), .Y(n73807) );
  NAND2xp33_ASAP7_75t_SL U58176 ( .A(n73752), .B(n73785), .Y(n73699) );
  AOI22xp33_ASAP7_75t_SL U58177 ( .A1(n72095), .A2(n72094), .B1(n72093), .B2(
        n72092), .Y(n72096) );
  NOR2x1_ASAP7_75t_SL U58178 ( .A(n70253), .B(n70252), .Y(n70476) );
  INVxp33_ASAP7_75t_SL U58179 ( .A(n62066), .Y(n62068) );
  NAND2xp33_ASAP7_75t_SL U58180 ( .A(n76356), .B(n76355), .Y(n76361) );
  INVxp67_ASAP7_75t_SL U58181 ( .A(n75847), .Y(n75319) );
  AOI21xp33_ASAP7_75t_SL U58182 ( .A1(n73993), .A2(n76364), .B(n76378), .Y(
        n73996) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58183 ( .A1(n74680), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .C(
        n70360), .Y(n70361) );
  AOI22xp33_ASAP7_75t_SL U58184 ( .A1(n73663), .A2(n73778), .B1(n73662), .B2(
        n73781), .Y(n73678) );
  NAND2xp5_ASAP7_75t_SL U58185 ( .A(n72769), .B(n73011), .Y(n72696) );
  AO21x1_ASAP7_75t_SL U58186 ( .A1(n76669), .A2(n76674), .B(n76676), .Y(n76670) );
  NAND2xp5_ASAP7_75t_SL U58187 ( .A(n59582), .B(n75486), .Y(n61810) );
  INVxp67_ASAP7_75t_SL U58188 ( .A(n70534), .Y(n70446) );
  OAI21xp33_ASAP7_75t_SL U58189 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .A2(
        n73722), .B(n73626), .Y(n73811) );
  NOR2xp33_ASAP7_75t_SRAM U58190 ( .A(n74710), .B(n74709), .Y(n74712) );
  NAND2xp33_ASAP7_75t_SL U58191 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_4_), .B(n69606), .Y(
        n69607) );
  INVxp67_ASAP7_75t_SL U58192 ( .A(n65782), .Y(n65727) );
  OAI22xp33_ASAP7_75t_SL U58193 ( .A1(n73791), .A2(n73835), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[18]), .B2(n59704), .Y(
        n73779) );
  NAND2xp33_ASAP7_75t_SL U58194 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_5_), .B(n69603), .Y(
        n69604) );
  AOI22xp33_ASAP7_75t_SL U58195 ( .A1(n73786), .A2(n73772), .B1(n73780), .B2(
        n73771), .Y(n73776) );
  NAND2xp33_ASAP7_75t_SL U58196 ( .A(n77752), .B(n75876), .Y(n75315) );
  OAI21xp33_ASAP7_75t_SL U58197 ( .A1(n65613), .A2(n65646), .B(n65612), .Y(
        n66154) );
  NAND2xp5_ASAP7_75t_SL U58198 ( .A(n71433), .B(n71469), .Y(n71462) );
  NAND2xp33_ASAP7_75t_SL U58199 ( .A(n72110), .B(n72038), .Y(n71909) );
  NAND2xp5_ASAP7_75t_SL U58200 ( .A(n77757), .B(n75876), .Y(n75316) );
  AOI22xp33_ASAP7_75t_SL U58201 ( .A1(n72116), .A2(n72045), .B1(n72062), .B2(
        n72041), .Y(n71910) );
  INVxp67_ASAP7_75t_SL U58202 ( .A(n62012), .Y(n75509) );
  INVxp67_ASAP7_75t_SL U58203 ( .A(n75817), .Y(n75203) );
  NOR3xp33_ASAP7_75t_SRAM U58204 ( .A(n76408), .B(n76407), .C(n76406), .Y(
        n76415) );
  NAND2xp5_ASAP7_75t_SL U58205 ( .A(or1200_cpu_or1200_fpu_result_conv[3]), .B(
        n77090), .Y(n61554) );
  OAI22xp33_ASAP7_75t_SL U58206 ( .A1(n57125), .A2(n72154), .B1(n72141), .B2(
        n57123), .Y(n72133) );
  INVxp67_ASAP7_75t_SL U58207 ( .A(n75702), .Y(n60627) );
  INVxp33_ASAP7_75t_SL U58208 ( .A(n76396), .Y(n76397) );
  INVx1_ASAP7_75t_SL U58209 ( .A(n72645), .Y(n72667) );
  NAND2xp5_ASAP7_75t_SL U58210 ( .A(n74828), .B(n2935), .Y(n2934) );
  NAND2xp5_ASAP7_75t_SL U58211 ( .A(n76334), .B(n74019), .Y(n76413) );
  NAND2xp33_ASAP7_75t_SL U58212 ( .A(n72116), .B(n72092), .Y(n71850) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58213 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]), .A2(n65549), 
        .B(n65548), .C(n65547), .Y(n65550) );
  INVxp33_ASAP7_75t_SL U58214 ( .A(n76395), .Y(n76398) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58215 ( .A1(n57083), .A2(n77773), .B(dwb_adr_o[2]), .C(n77771), .Y(n77772) );
  NAND2xp5_ASAP7_75t_SL U58216 ( .A(n73778), .B(n73780), .Y(n73746) );
  INVxp33_ASAP7_75t_SL U58217 ( .A(n74511), .Y(n74512) );
  INVx1_ASAP7_75t_SL U58218 ( .A(n62418), .Y(n76712) );
  NAND2xp33_ASAP7_75t_SL U58219 ( .A(n72110), .B(n72090), .Y(n71842) );
  OR2x2_ASAP7_75t_SL U58220 ( .A(n58084), .B(n63571), .Y(n58081) );
  NOR3xp33_ASAP7_75t_SRAM U58221 ( .A(n70473), .B(n70472), .C(n70487), .Y(
        n70410) );
  NAND2xp33_ASAP7_75t_SL U58222 ( .A(n72620), .B(n72645), .Y(n72617) );
  NAND2xp33_ASAP7_75t_SL U58223 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .B(
        n73827), .Y(n73769) );
  INVxp67_ASAP7_75t_SL U58224 ( .A(n72046), .Y(n72047) );
  AOI21xp33_ASAP7_75t_SL U58225 ( .A1(n2759), .A2(n77793), .B(n60276), .Y(
        n9479) );
  OAI21xp33_ASAP7_75t_SL U58226 ( .A1(n77310), .A2(n22057), .B(ic_en), .Y(
        n77311) );
  OAI22xp33_ASAP7_75t_SL U58227 ( .A1(n72316), .A2(n57123), .B1(n72317), .B2(
        n57127), .Y(n72251) );
  NAND2xp5_ASAP7_75t_SL U58228 ( .A(n74269), .B(n74067), .Y(n74102) );
  AOI21xp33_ASAP7_75t_SL U58229 ( .A1(n61429), .A2(n62762), .B(n75456), .Y(
        n60922) );
  AOI21xp33_ASAP7_75t_SL U58230 ( .A1(n2763), .A2(n60280), .B(n60279), .Y(
        n9480) );
  AOI21xp33_ASAP7_75t_SL U58231 ( .A1(n2765), .A2(n60280), .B(n60279), .Y(
        n9481) );
  AND3x1_ASAP7_75t_SL U58232 ( .A(n60670), .B(n3123), .C(n57318), .Y(n60671)
         );
  INVxp67_ASAP7_75t_SL U58233 ( .A(n60799), .Y(n60626) );
  O2A1O1Ixp33_ASAP7_75t_SL U58234 ( .A1(n59778), .A2(n59777), .B(
        or1200_dc_top_tag_19_), .C(n59776), .Y(n59779) );
  INVxp67_ASAP7_75t_SL U58235 ( .A(n69190), .Y(n69179) );
  OAI22xp33_ASAP7_75t_SL U58236 ( .A1(n57125), .A2(n72316), .B1(n72308), .B2(
        n57123), .Y(n72243) );
  NAND2xp33_ASAP7_75t_SL U58237 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .B(
        n73820), .Y(n73719) );
  NAND2xp33_ASAP7_75t_SL U58238 ( .A(n63387), .B(n63386), .Y(n63393) );
  OAI22xp33_ASAP7_75t_SL U58239 ( .A1(n72122), .A2(n71979), .B1(n72046), .B2(
        n72067), .Y(n71980) );
  NOR2xp33_ASAP7_75t_SRAM U58240 ( .A(n77349), .B(n77348), .Y(n77351) );
  INVxp33_ASAP7_75t_SL U58241 ( .A(n74954), .Y(n74955) );
  NOR2xp33_ASAP7_75t_SRAM U58242 ( .A(n57082), .B(n63571), .Y(n60659) );
  OAI21xp33_ASAP7_75t_SL U58243 ( .A1(n65354), .A2(n65399), .B(n65333), .Y(
        n65335) );
  NAND2xp5_ASAP7_75t_SL U58244 ( .A(or1200_cpu_or1200_mult_mac_div_free), .B(
        n75486), .Y(n63248) );
  OAI22xp33_ASAP7_75t_SL U58245 ( .A1(n72162), .A2(n57123), .B1(n72164), .B2(
        n57127), .Y(n72155) );
  INVxp67_ASAP7_75t_SL U58246 ( .A(n62638), .Y(n58203) );
  NAND2xp5_ASAP7_75t_SL U58247 ( .A(n61855), .B(n60618), .Y(n61526) );
  NAND2xp33_ASAP7_75t_SL U58248 ( .A(n72093), .B(n72120), .Y(n71967) );
  NAND2xp33_ASAP7_75t_SL U58249 ( .A(or1200_cpu_or1200_fpu_result_conv[5]), 
        .B(n77090), .Y(n61652) );
  OAI21xp33_ASAP7_75t_SL U58250 ( .A1(n65629), .A2(n65745), .B(n65572), .Y(
        n66098) );
  NAND2xp5_ASAP7_75t_SL U58251 ( .A(n72584), .B(n74235), .Y(n72583) );
  INVxp33_ASAP7_75t_SL U58252 ( .A(n62013), .Y(n60643) );
  NAND2xp33_ASAP7_75t_SL U58253 ( .A(n72095), .B(n71966), .Y(n71968) );
  AOI21xp5_ASAP7_75t_SL U58254 ( .A1(n63415), .A2(n63433), .B(n63431), .Y(
        n63416) );
  NAND2xp5_ASAP7_75t_SL U58255 ( .A(n74125), .B(n59759), .Y(n59757) );
  OAI22xp33_ASAP7_75t_SL U58256 ( .A1(n72154), .A2(n57123), .B1(n72163), .B2(
        n57127), .Y(n72142) );
  AOI21xp5_ASAP7_75t_SL U58257 ( .A1(n75428), .A2(n59788), .B(n59787), .Y(
        n59790) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58258 ( .A1(n74661), .A2(n74660), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_7_), .C(
        n74659), .Y(n74676) );
  NAND2xp33_ASAP7_75t_SL U58259 ( .A(n63730), .B(n77257), .Y(n63733) );
  NAND2xp5_ASAP7_75t_SL U58260 ( .A(n73772), .B(n73780), .Y(n73731) );
  NAND2xp5_ASAP7_75t_SL U58261 ( .A(n70081), .B(n69897), .Y(n70153) );
  INVx1_ASAP7_75t_SL U58262 ( .A(n76796), .Y(n62382) );
  OAI21xp5_ASAP7_75t_SL U58263 ( .A1(n63390), .A2(n63386), .B(n63387), .Y(
        n63326) );
  OAI22xp33_ASAP7_75t_SL U58264 ( .A1(n72079), .A2(n57123), .B1(n72132), .B2(
        n57127), .Y(n72055) );
  NAND2xp5_ASAP7_75t_SL U58265 ( .A(n65858), .B(n65409), .Y(n65660) );
  AOI22xp33_ASAP7_75t_SL U58266 ( .A1(n72110), .A2(n72285), .B1(n72116), .B2(
        n72061), .Y(n71938) );
  NAND2xp5_ASAP7_75t_SL U58267 ( .A(n63571), .B(n64780), .Y(n61876) );
  NAND2xp33_ASAP7_75t_SL U58268 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .B(
        n73830), .Y(n73627) );
  NAND2xp33_ASAP7_75t_SL U58269 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .B(
        n72224), .Y(n72176) );
  AND2x2_ASAP7_75t_SRAM U58270 ( .A(n72286), .B(n72040), .Y(n71916) );
  INVxp33_ASAP7_75t_SL U58271 ( .A(n73876), .Y(n73879) );
  NOR2xp33_ASAP7_75t_SRAM U58272 ( .A(n76404), .B(n76344), .Y(n76348) );
  INVxp33_ASAP7_75t_SL U58273 ( .A(n77348), .Y(n77306) );
  NAND2xp5_ASAP7_75t_SL U58274 ( .A(n73488), .B(n73490), .Y(n73872) );
  OAI22xp33_ASAP7_75t_SL U58275 ( .A1(n57125), .A2(n71984), .B1(n71953), .B2(
        n57123), .Y(n71954) );
  NAND2xp33_ASAP7_75t_SL U58276 ( .A(n78365), .B(n2935), .Y(n1521) );
  NAND2xp33_ASAP7_75t_SL U58277 ( .A(n61145), .B(n61144), .Y(n62070) );
  AOI21xp33_ASAP7_75t_SL U58278 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_4_), .A2(n65357), .B(
        n65356), .Y(n65358) );
  NAND2xp33_ASAP7_75t_SL U58279 ( .A(n1121), .B(n75689), .Y(n75690) );
  INVxp67_ASAP7_75t_SL U58280 ( .A(n72064), .Y(n72144) );
  NOR2x1_ASAP7_75t_SL U58281 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_6_), .B(n65347), .Y(
        n65326) );
  INVxp67_ASAP7_75t_SL U58282 ( .A(n69927), .Y(n70064) );
  INVxp33_ASAP7_75t_SL U58283 ( .A(n63527), .Y(n63529) );
  OAI22xp33_ASAP7_75t_SL U58284 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_), 
        .A2(n57123), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .B2(n57127), .Y(n72187) );
  INVxp33_ASAP7_75t_SL U58285 ( .A(n72535), .Y(n72532) );
  NAND2xp5_ASAP7_75t_SL U58286 ( .A(or1200_cpu_or1200_fpu_result_conv[4]), .B(
        n77090), .Y(n61453) );
  NAND2xp5_ASAP7_75t_SL U58287 ( .A(n65088), .B(n65087), .Y(n63542) );
  NAND2xp33_ASAP7_75t_SL U58288 ( .A(n72093), .B(n72069), .Y(n71928) );
  INVxp67_ASAP7_75t_SL U58289 ( .A(n71979), .Y(n71911) );
  AOI22xp33_ASAP7_75t_SL U58290 ( .A1(n72116), .A2(n72040), .B1(n72286), .B2(
        n72041), .Y(n71806) );
  NAND2xp33_ASAP7_75t_SL U58291 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_19_), .B(n69687), 
        .Y(n69688) );
  NAND2xp33_ASAP7_75t_SL U58292 ( .A(n72110), .B(n72109), .Y(n72111) );
  INVxp33_ASAP7_75t_SL U58293 ( .A(n76439), .Y(n61419) );
  OAI21xp5_ASAP7_75t_SL U58294 ( .A1(n70310), .A2(n70349), .B(n70309), .Y(
        n70484) );
  AOI21xp5_ASAP7_75t_SL U58295 ( .A1(n63435), .A2(n63434), .B(n63456), .Y(
        n63436) );
  INVx1_ASAP7_75t_SL U58296 ( .A(n69747), .Y(n69581) );
  INVxp33_ASAP7_75t_SL U58297 ( .A(n70204), .Y(n70208) );
  NOR2x1_ASAP7_75t_SL U58298 ( .A(n60625), .B(n60624), .Y(n75227) );
  OAI22xp33_ASAP7_75t_SL U58299 ( .A1(n73646), .A2(n73715), .B1(n73645), .B2(
        n73765), .Y(n73647) );
  AOI21xp33_ASAP7_75t_SL U58300 ( .A1(n2589), .A2(n60725), .B(n60724), .Y(
        n77457) );
  INVxp33_ASAP7_75t_SL U58301 ( .A(n62200), .Y(n62207) );
  INVxp67_ASAP7_75t_SL U58302 ( .A(n72547), .Y(n72536) );
  OR2x2_ASAP7_75t_SL U58303 ( .A(n60628), .B(n78182), .Y(n61828) );
  OAI22xp33_ASAP7_75t_SL U58304 ( .A1(n72346), .A2(n57123), .B1(n72360), .B2(
        n57127), .Y(n72264) );
  OAI22xp33_ASAP7_75t_SL U58305 ( .A1(n74706), .A2(n70369), .B1(n70368), .B2(
        n70398), .Y(n70461) );
  NAND2xp5_ASAP7_75t_SL U58306 ( .A(n74461), .B(n74715), .Y(n74221) );
  INVxp33_ASAP7_75t_SL U58307 ( .A(n72663), .Y(n72651) );
  NAND2xp33_ASAP7_75t_SL U58308 ( .A(n75453), .B(n60546), .Y(n60547) );
  OAI21xp33_ASAP7_75t_SL U58309 ( .A1(n78244), .A2(n71512), .B(n71511), .Y(
        n71520) );
  INVxp33_ASAP7_75t_SL U58310 ( .A(n73594), .Y(n73534) );
  NAND2xp33_ASAP7_75t_SL U58311 ( .A(n74696), .B(n74670), .Y(n74679) );
  OAI22xp33_ASAP7_75t_SL U58312 ( .A1(n72319), .A2(n57123), .B1(n72318), .B2(
        n57127), .Y(n72320) );
  INVxp67_ASAP7_75t_SL U58313 ( .A(n60963), .Y(n60619) );
  INVxp33_ASAP7_75t_SL U58314 ( .A(n61856), .Y(n61698) );
  NAND2xp33_ASAP7_75t_SL U58315 ( .A(n72126), .B(n72120), .Y(n71900) );
  NAND2xp33_ASAP7_75t_SL U58316 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_6_), .B(n69611), .Y(
        n69599) );
  OAI21xp33_ASAP7_75t_SL U58317 ( .A1(n71566), .A2(n71565), .B(n71564), .Y(
        n71572) );
  NAND2xp33_ASAP7_75t_SL U58318 ( .A(n73488), .B(n73871), .Y(n73489) );
  INVxp67_ASAP7_75t_SL U58319 ( .A(n74134), .Y(n74145) );
  AOI21xp5_ASAP7_75t_SL U58320 ( .A1(n74757), .A2(n75455), .B(n74771), .Y(
        n74779) );
  INVxp33_ASAP7_75t_SL U58321 ( .A(n70222), .Y(n70226) );
  AOI21xp33_ASAP7_75t_SL U58322 ( .A1(n63283), .A2(n63303), .B(n63304), .Y(
        n63284) );
  OAI22xp33_ASAP7_75t_SL U58323 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .A2(
        n73740), .B1(n58619), .B2(n73755), .Y(n73741) );
  NAND2xp33_ASAP7_75t_SL U58324 ( .A(n72110), .B(n71973), .Y(n71974) );
  FAx1_ASAP7_75t_SL U58325 ( .A(or1200_dc_top_tag_18_), .B(n59750), .CI(n59749), .CON(), .SN(n59755) );
  INVxp33_ASAP7_75t_SL U58326 ( .A(n69625), .Y(n69622) );
  OAI21xp33_ASAP7_75t_SL U58327 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_), 
        .A2(n57125), .B(n72177), .Y(n72179) );
  OAI21xp33_ASAP7_75t_SL U58328 ( .A1(n58422), .A2(n72319), .B(n71750), .Y(
        n71751) );
  NAND2xp33_ASAP7_75t_SL U58329 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_ine_o), 
        .B(n74759), .Y(n1534) );
  AOI21xp33_ASAP7_75t_SL U58330 ( .A1(n73682), .A2(n73681), .B(n73752), .Y(
        n73684) );
  OAI22xp33_ASAP7_75t_SL U58331 ( .A1(n72079), .A2(n57125), .B1(n72080), .B2(
        n57127), .Y(n72034) );
  INVxp67_ASAP7_75t_SL U58332 ( .A(n77997), .Y(n77999) );
  OAI21xp5_ASAP7_75t_SL U58333 ( .A1(n76976), .A2(n65672), .B(n65671), .Y(
        n65830) );
  NAND2xp5_ASAP7_75t_SL U58334 ( .A(n76886), .B(n68881), .Y(n68889) );
  INVxp67_ASAP7_75t_SL U58335 ( .A(n59716), .Y(n59714) );
  INVxp67_ASAP7_75t_SL U58336 ( .A(n68887), .Y(n68888) );
  INVxp67_ASAP7_75t_SL U58337 ( .A(n61998), .Y(n61284) );
  INVxp67_ASAP7_75t_SL U58338 ( .A(n73136), .Y(n73132) );
  INVxp33_ASAP7_75t_SL U58339 ( .A(n69642), .Y(n69632) );
  OAI21xp33_ASAP7_75t_SL U58340 ( .A1(or1200_cpu_or1200_mult_mac_n389), .A2(
        or1200_cpu_or1200_mult_mac_n243), .B(n69208), .Y(n69285) );
  INVxp33_ASAP7_75t_SL U58341 ( .A(n63897), .Y(n63902) );
  OAI21xp33_ASAP7_75t_SL U58342 ( .A1(n64172), .A2(n64171), .B(n65098), .Y(
        n65093) );
  AOI22xp33_ASAP7_75t_SL U58343 ( .A1(n66182), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[24]), .B1(n65592), 
        .B2(n66145), .Y(n65509) );
  INVx1_ASAP7_75t_SL U58344 ( .A(n75861), .Y(n76770) );
  INVxp33_ASAP7_75t_SL U58345 ( .A(n62292), .Y(n61241) );
  INVx1_ASAP7_75t_SL U58346 ( .A(n60818), .Y(n60556) );
  OAI21xp33_ASAP7_75t_SL U58347 ( .A1(n58422), .A2(n72348), .B(n71870), .Y(
        n71871) );
  INVxp67_ASAP7_75t_SL U58348 ( .A(n60494), .Y(n60340) );
  AOI21xp33_ASAP7_75t_SL U58349 ( .A1(n62065), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_s_state), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_start_i), .Y(n62057) );
  NAND2xp33_ASAP7_75t_SL U58350 ( .A(n3078), .B(n60490), .Y(n62007) );
  INVxp33_ASAP7_75t_SL U58351 ( .A(n65602), .Y(n65513) );
  OAI21xp33_ASAP7_75t_SL U58352 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .A2(
        n71849), .B(n71817), .Y(n72045) );
  INVx2_ASAP7_75t_SL U58353 ( .A(n62629), .Y(n57195) );
  NOR2xp33_ASAP7_75t_SRAM U58354 ( .A(n77410), .B(n59886), .Y(n59887) );
  NAND2xp33_ASAP7_75t_SL U58355 ( .A(n70296), .B(n69379), .Y(n69380) );
  OAI21xp33_ASAP7_75t_SL U58356 ( .A1(n2455), .A2(n70531), .B(n2456), .Y(
        n69381) );
  NAND2xp33_ASAP7_75t_SL U58357 ( .A(n65831), .B(n65808), .Y(n65777) );
  NAND2xp33_ASAP7_75t_SL U58358 ( .A(n59567), .B(n61087), .Y(n76764) );
  NAND2xp33_ASAP7_75t_SL U58359 ( .A(n75456), .B(n76404), .Y(n1523) );
  AOI22xp33_ASAP7_75t_SL U58360 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_2_), .A2(n65357), .B1(
        n65346), .B2(n65339), .Y(n65340) );
  OAI21xp33_ASAP7_75t_SL U58361 ( .A1(n72263), .A2(n57127), .B(n72249), .Y(
        n72333) );
  INVxp33_ASAP7_75t_SL U58362 ( .A(n70708), .Y(n70724) );
  INVx1_ASAP7_75t_SL U58363 ( .A(n72508), .Y(n72492) );
  AO21x1_ASAP7_75t_SRAM U58364 ( .A1(n70296), .A2(n70531), .B(n70477), .Y(
        n9559) );
  INVxp33_ASAP7_75t_SL U58365 ( .A(n74926), .Y(n69347) );
  INVxp67_ASAP7_75t_SL U58366 ( .A(n75424), .Y(n75428) );
  AOI21xp5_ASAP7_75t_SL U58367 ( .A1(n59869), .A2(n69366), .B(n59868), .Y(
        n75193) );
  AOI22xp33_ASAP7_75t_SL U58368 ( .A1(n65357), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_3_), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_20_), .B2(n65401), .Y(
        n65333) );
  NAND2xp33_ASAP7_75t_SL U58369 ( .A(n63720), .B(n74926), .Y(n63721) );
  INVxp33_ASAP7_75t_SL U58370 ( .A(n69977), .Y(n69952) );
  INVxp33_ASAP7_75t_SL U58371 ( .A(n63388), .Y(n63391) );
  NAND2xp5_ASAP7_75t_SL U58372 ( .A(n74499), .B(n69524), .Y(n69897) );
  NOR2xp33_ASAP7_75t_SRAM U58373 ( .A(n71984), .B(n57127), .Y(n71934) );
  OAI22xp33_ASAP7_75t_SL U58374 ( .A1(n72219), .A2(n57125), .B1(n72234), .B2(
        n57127), .Y(n72199) );
  OAI21xp33_ASAP7_75t_SL U58375 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .A2(
        n71877), .B(n71771), .Y(n72146) );
  NAND2xp5_ASAP7_75t_SL U58376 ( .A(n57083), .B(n77750), .Y(n77761) );
  NAND2xp5_ASAP7_75t_SL U58377 ( .A(n60278), .B(n60275), .Y(n60276) );
  INVxp33_ASAP7_75t_SL U58378 ( .A(n65628), .Y(n65569) );
  INVxp67_ASAP7_75t_SL U58379 ( .A(n77251), .Y(n61169) );
  NAND2xp33_ASAP7_75t_SL U58380 ( .A(n59182), .B(n59583), .Y(n61725) );
  OAI21xp33_ASAP7_75t_SL U58381 ( .A1(n59853), .A2(n74123), .B(n59852), .Y(
        n59858) );
  NAND2xp33_ASAP7_75t_SL U58382 ( .A(n59567), .B(n62359), .Y(n75702) );
  NAND2xp33_ASAP7_75t_SL U58383 ( .A(n59443), .B(n61488), .Y(n61490) );
  OAI22xp33_ASAP7_75t_SL U58384 ( .A1(n72005), .A2(n57125), .B1(n72054), .B2(
        n57127), .Y(n72008) );
  INVxp33_ASAP7_75t_SL U58385 ( .A(n60306), .Y(n59964) );
  OAI21xp5_ASAP7_75t_SL U58386 ( .A1(n74549), .A2(n74548), .B(n74547), .Y(
        n74827) );
  NAND2xp5_ASAP7_75t_SL U58387 ( .A(n68943), .B(n68942), .Y(n68992) );
  INVxp67_ASAP7_75t_SL U58388 ( .A(n61209), .Y(n61225) );
  NAND2xp33_ASAP7_75t_SL U58389 ( .A(n63533), .B(n63539), .Y(n65082) );
  OAI21xp33_ASAP7_75t_SL U58390 ( .A1(n73618), .A2(n73808), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .Y(
        n73650) );
  INVxp67_ASAP7_75t_SL U58391 ( .A(n72017), .Y(n72117) );
  NOR2xp33_ASAP7_75t_SRAM U58392 ( .A(n62020), .B(n62019), .Y(n62021) );
  INVxp33_ASAP7_75t_SL U58393 ( .A(n74459), .Y(n74725) );
  AOI21xp33_ASAP7_75t_SL U58394 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[9]), .A2(
        n73156), .B(n73070), .Y(n73068) );
  NAND2xp5_ASAP7_75t_SL U58395 ( .A(n74832), .B(n74831), .Y(n1502) );
  INVxp67_ASAP7_75t_SL U58396 ( .A(n60491), .Y(n60358) );
  OAI22xp33_ASAP7_75t_SL U58397 ( .A1(n73791), .A2(n73790), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[17]), .B2(n59704), .Y(
        n73792) );
  INVxp33_ASAP7_75t_SL U58398 ( .A(n69691), .Y(n69687) );
  NAND2xp33_ASAP7_75t_SL U58399 ( .A(n63723), .B(n74926), .Y(n63724) );
  AOI21xp5_ASAP7_75t_SL U58400 ( .A1(n65526), .A2(n65525), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_nan), .Y(n65532) );
  NAND2xp5_ASAP7_75t_SL U58401 ( .A(n70223), .B(n70222), .Y(n70241) );
  INVxp67_ASAP7_75t_SL U58402 ( .A(n68951), .Y(n68946) );
  NAND2xp5_ASAP7_75t_SL U58403 ( .A(n69435), .B(n69430), .Y(n69431) );
  INVx1_ASAP7_75t_SL U58404 ( .A(n61648), .Y(n60670) );
  OAI21xp33_ASAP7_75t_SL U58405 ( .A1(n65530), .A2(n74132), .B(n76976), .Y(
        n65531) );
  NAND2xp33_ASAP7_75t_SL U58406 ( .A(n78244), .B(n70154), .Y(n70157) );
  INVxp33_ASAP7_75t_SL U58407 ( .A(n61855), .Y(n60617) );
  INVxp33_ASAP7_75t_SL U58408 ( .A(n76613), .Y(n76614) );
  NAND2xp33_ASAP7_75t_SL U58409 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[8]), .B(n65808), .Y(
        n65698) );
  NAND2xp33_ASAP7_75t_SL U58410 ( .A(n73686), .B(n73716), .Y(n73646) );
  NAND2xp33_ASAP7_75t_SL U58411 ( .A(n73244), .B(n74502), .Y(n73243) );
  O2A1O1Ixp33_ASAP7_75t_SL U58412 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .A2(
        n71952), .B(n57125), .C(n71931), .Y(n71867) );
  NAND2xp33_ASAP7_75t_SL U58413 ( .A(n2951), .B(n74831), .Y(n74780) );
  NAND2xp33_ASAP7_75t_SL U58414 ( .A(n73180), .B(n74502), .Y(n73179) );
  INVxp67_ASAP7_75t_SL U58415 ( .A(n65526), .Y(n65492) );
  AOI21xp33_ASAP7_75t_SL U58416 ( .A1(n73637), .A2(n73636), .B(n73752), .Y(
        n73638) );
  INVxp33_ASAP7_75t_SL U58417 ( .A(n77851), .Y(n60577) );
  INVxp67_ASAP7_75t_SL U58418 ( .A(n77931), .Y(n77166) );
  OAI21xp33_ASAP7_75t_SL U58419 ( .A1(n70568), .A2(n70223), .B(n70238), .Y(
        n70571) );
  NAND2xp5_ASAP7_75t_SL U58420 ( .A(n60572), .B(n60544), .Y(n77164) );
  OAI21xp33_ASAP7_75t_SL U58421 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_5_), .A2(n66166), 
        .B(n66110), .Y(n66165) );
  NOR2xp33_ASAP7_75t_SRAM U58422 ( .A(n62026), .B(n63245), .Y(n62029) );
  INVxp67_ASAP7_75t_SL U58423 ( .A(n73386), .Y(n73380) );
  NAND2xp33_ASAP7_75t_SL U58424 ( .A(n73028), .B(n72964), .Y(n72689) );
  NAND2xp5_ASAP7_75t_SL U58425 ( .A(n70326), .B(n70325), .Y(n70369) );
  OAI21xp33_ASAP7_75t_SL U58426 ( .A1(n70308), .A2(n70307), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .Y(
        n70309) );
  NAND2xp33_ASAP7_75t_SL U58427 ( .A(n73185), .B(n74502), .Y(n73184) );
  NAND2xp33_ASAP7_75t_SL U58428 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .B(n71514), .Y(
        n71511) );
  NOR4xp25_ASAP7_75t_SRAM U58429 ( .A(n65456), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[36]), .C(n65455), 
        .D(n65454), .Y(n65464) );
  NAND2xp33_ASAP7_75t_SL U58430 ( .A(n74706), .B(n70397), .Y(n70368) );
  NAND2xp5_ASAP7_75t_SL U58431 ( .A(n65495), .B(n65483), .Y(n65486) );
  OAI21xp33_ASAP7_75t_SL U58432 ( .A1(n66181), .A2(n65681), .B(n65594), .Y(
        n66120) );
  NAND2xp33_ASAP7_75t_SL U58433 ( .A(n73333), .B(n74502), .Y(n73332) );
  NAND2xp5_ASAP7_75t_SL U58434 ( .A(n73081), .B(n73094), .Y(n73097) );
  INVxp67_ASAP7_75t_SL U58435 ( .A(n70539), .Y(n70471) );
  NAND2xp33_ASAP7_75t_SL U58436 ( .A(n73123), .B(n74502), .Y(n73122) );
  INVxp67_ASAP7_75t_SL U58437 ( .A(n60102), .Y(n59954) );
  INVxp67_ASAP7_75t_SL U58438 ( .A(n72528), .Y(n72525) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58439 ( .A1(n74669), .A2(n74668), .B(n74667), 
        .C(n74666), .Y(n74670) );
  NAND2xp5_ASAP7_75t_SL U58440 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_3_), .B(
        n72582), .Y(n72595) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58441 ( .A1(n61030), .A2(n61145), .B(n2814), .C(
        n61029), .Y(n61033) );
  OAI21xp33_ASAP7_75t_SL U58442 ( .A1(n76405), .A2(n76346), .B(n76338), .Y(
        n76410) );
  INVxp67_ASAP7_75t_SL U58443 ( .A(n71815), .Y(n71816) );
  INVx1_ASAP7_75t_SL U58444 ( .A(n73869), .Y(n73888) );
  BUFx2_ASAP7_75t_SL U58445 ( .A(n59108), .Y(n57457) );
  NAND2xp5_ASAP7_75t_SL U58446 ( .A(n61995), .B(n59877), .Y(n59891) );
  NOR2xp33_ASAP7_75t_SL U58447 ( .A(n71560), .B(n71565), .Y(n71631) );
  OAI21xp33_ASAP7_75t_SL U58448 ( .A1(n2335), .A2(n70540), .B(n70283), .Y(
        n70284) );
  NAND2xp5_ASAP7_75t_SL U58449 ( .A(n73673), .B(n73672), .Y(n73835) );
  NAND2xp5_ASAP7_75t_SL U58450 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_3_), .B(
        n71662), .Y(n71661) );
  INVxp33_ASAP7_75t_SL U58451 ( .A(n77918), .Y(n76688) );
  OAI22xp33_ASAP7_75t_SL U58452 ( .A1(n65853), .A2(n65546), .B1(n65421), .B2(
        n65420), .Y(n65422) );
  INVxp67_ASAP7_75t_SL U58453 ( .A(n71787), .Y(n71742) );
  NAND2xp33_ASAP7_75t_SL U58454 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[4]), .B(n66199), .Y(
        n65540) );
  INVxp33_ASAP7_75t_SL U58455 ( .A(n76364), .Y(n76365) );
  INVxp33_ASAP7_75t_SL U58456 ( .A(n71662), .Y(n71641) );
  OAI21xp33_ASAP7_75t_SL U58457 ( .A1(n59443), .A2(n62432), .B(n62431), .Y(
        n75862) );
  INVx1_ASAP7_75t_SL U58458 ( .A(n62202), .Y(n75405) );
  INVxp33_ASAP7_75t_SL U58459 ( .A(n74846), .Y(n74847) );
  NAND2xp5_ASAP7_75t_SL U58460 ( .A(n70396), .B(n70395), .Y(n70462) );
  NAND2xp33_ASAP7_75t_SL U58461 ( .A(n73304), .B(n74502), .Y(n73303) );
  AOI21xp5_ASAP7_75t_SL U58462 ( .A1(n66210), .A2(n74835), .B(n66209), .Y(
        n66217) );
  INVxp33_ASAP7_75t_SL U58463 ( .A(n76377), .Y(n76382) );
  INVxp33_ASAP7_75t_SL U58464 ( .A(n76384), .Y(n76369) );
  INVxp67_ASAP7_75t_SL U58465 ( .A(n76368), .Y(n76370) );
  INVxp67_ASAP7_75t_SL U58466 ( .A(n70397), .Y(n70399) );
  OAI21xp33_ASAP7_75t_SL U58467 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .A2(n65483), .B(
        n74133), .Y(n65484) );
  NOR2xp33_ASAP7_75t_SRAM U58468 ( .A(n76363), .B(n76367), .Y(n73982) );
  INVxp33_ASAP7_75t_SL U58469 ( .A(n76354), .Y(n76355) );
  INVx1_ASAP7_75t_SL U58470 ( .A(n70272), .Y(n70252) );
  NAND2xp5_ASAP7_75t_SL U58471 ( .A(n77623), .B(n60554), .Y(n61243) );
  NAND2xp33_ASAP7_75t_SL U58472 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .B(
        n70359), .Y(n70360) );
  NAND2xp5_ASAP7_75t_SL U58473 ( .A(n71647), .B(n71648), .Y(n71790) );
  INVxp67_ASAP7_75t_SL U58474 ( .A(n74745), .Y(n74746) );
  NAND2xp33_ASAP7_75t_SL U58475 ( .A(n73159), .B(n74502), .Y(n73158) );
  NAND2xp33_ASAP7_75t_SL U58476 ( .A(n71515), .B(n71514), .Y(n71518) );
  AOI31xp33_ASAP7_75t_SRAM U58477 ( .A1(n2600), .A2(n2693), .A3(n2972), .B(
        n60102), .Y(n60104) );
  NAND2xp33_ASAP7_75t_SL U58478 ( .A(n75851), .B(n75850), .Y(n76345) );
  NAND2xp33_ASAP7_75t_SL U58479 ( .A(n64208), .B(n60554), .Y(n77622) );
  INVxp33_ASAP7_75t_SL U58480 ( .A(n76338), .Y(n76407) );
  INVxp33_ASAP7_75t_SL U58481 ( .A(n69614), .Y(n69603) );
  NAND2xp5_ASAP7_75t_SL U58482 ( .A(n69439), .B(n70154), .Y(n2935) );
  AOI21xp33_ASAP7_75t_SL U58483 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .A2(
        n71849), .B(n71848), .Y(n72092) );
  OAI21xp33_ASAP7_75t_SL U58484 ( .A1(n70317), .A2(n70488), .B(n70298), .Y(
        n70299) );
  INVxp67_ASAP7_75t_SL U58485 ( .A(n74713), .Y(n74722) );
  NAND2xp33_ASAP7_75t_SL U58486 ( .A(n73896), .B(n73890), .Y(n74067) );
  INVxp33_ASAP7_75t_SL U58487 ( .A(n69605), .Y(n69606) );
  NAND2xp33_ASAP7_75t_SL U58488 ( .A(n73119), .B(n74502), .Y(n73118) );
  INVxp33_ASAP7_75t_SL U58489 ( .A(n59722), .Y(n59723) );
  OAI21xp33_ASAP7_75t_SL U58490 ( .A1(n66186), .A2(n66179), .B(n74136), .Y(
        n66189) );
  NOR2xp33_ASAP7_75t_SRAM U58491 ( .A(dwb_adr_o[2]), .B(n77773), .Y(n77771) );
  NAND2xp5_ASAP7_75t_SL U58492 ( .A(n60503), .B(n60502), .Y(n60504) );
  NAND2xp33_ASAP7_75t_SL U58493 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_0_), .B(n69582), .Y(
        n17036) );
  AOI22xp33_ASAP7_75t_SL U58494 ( .A1(n66182), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]), .B1(n65587), 
        .B2(n66145), .Y(n65516) );
  INVxp33_ASAP7_75t_SL U58495 ( .A(n77937), .Y(n60543) );
  INVxp33_ASAP7_75t_SL U58496 ( .A(n61010), .Y(n61011) );
  NOR3xp33_ASAP7_75t_SRAM U58497 ( .A(n77937), .B(n59493), .C(n61064), .Y(
        n61065) );
  INVx1_ASAP7_75t_SL U58498 ( .A(n73788), .Y(n73780) );
  OAI21xp33_ASAP7_75t_SL U58499 ( .A1(n65420), .A2(n65407), .B(n65406), .Y(
        n65411) );
  OAI21xp33_ASAP7_75t_SL U58500 ( .A1(n74377), .A2(n74744), .B(n74376), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_N86) );
  INVxp33_ASAP7_75t_SL U58501 ( .A(n64282), .Y(n77659) );
  INVxp67_ASAP7_75t_SL U58502 ( .A(n77125), .Y(n76801) );
  OAI21xp33_ASAP7_75t_SL U58503 ( .A1(n75198), .A2(n59494), .B(n60017), .Y(
        n60010) );
  OAI21xp33_ASAP7_75t_SL U58504 ( .A1(n75675), .A2(n59494), .B(n60017), .Y(
        n60003) );
  OAI21xp33_ASAP7_75t_SL U58505 ( .A1(n77177), .A2(n59494), .B(n60017), .Y(
        n60018) );
  AOI21xp33_ASAP7_75t_SL U58506 ( .A1(n77646), .A2(n77645), .B(n77644), .Y(
        n77647) );
  INVx1_ASAP7_75t_SL U58507 ( .A(n75318), .Y(n76450) );
  OAI21xp33_ASAP7_75t_SL U58508 ( .A1(n74660), .A2(n70488), .B(n70423), .Y(
        n70424) );
  INVxp67_ASAP7_75t_SL U58509 ( .A(n76381), .Y(n61099) );
  INVxp67_ASAP7_75t_SL U58510 ( .A(n70487), .Y(n70541) );
  INVx1_ASAP7_75t_SL U58511 ( .A(n73981), .Y(n76436) );
  INVxp33_ASAP7_75t_SL U58512 ( .A(n77064), .Y(n77067) );
  INVx1_ASAP7_75t_SL U58513 ( .A(n73032), .Y(n73007) );
  INVxp33_ASAP7_75t_SL U58514 ( .A(n72734), .Y(n72808) );
  INVx1_ASAP7_75t_SL U58515 ( .A(n77600), .Y(n77980) );
  INVx1_ASAP7_75t_SL U58516 ( .A(n77019), .Y(n77896) );
  NAND2xp33_ASAP7_75t_SL U58517 ( .A(n61028), .B(n61311), .Y(n61029) );
  AOI22xp33_ASAP7_75t_SL U58518 ( .A1(n74686), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_), .B2(
        n70543), .Y(n70276) );
  INVxp67_ASAP7_75t_SL U58519 ( .A(n61318), .Y(n59877) );
  INVxp33_ASAP7_75t_SL U58520 ( .A(n61507), .Y(n61508) );
  NAND2xp5_ASAP7_75t_SL U58521 ( .A(n70281), .B(n70280), .Y(n70438) );
  NAND2xp33_ASAP7_75t_SL U58522 ( .A(n70327), .B(n70445), .Y(n70273) );
  NAND2xp5_ASAP7_75t_SL U58523 ( .A(n70270), .B(n70288), .Y(n70481) );
  NAND2xp33_ASAP7_75t_SL U58524 ( .A(n70327), .B(n74686), .Y(n70298) );
  INVxp33_ASAP7_75t_SL U58525 ( .A(n74025), .Y(n74021) );
  INVx1_ASAP7_75t_SL U58526 ( .A(n75700), .Y(n76767) );
  NAND2xp33_ASAP7_75t_SL U58527 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .B(
        n70348), .Y(n70350) );
  NAND2xp5_ASAP7_75t_SL U58528 ( .A(n70311), .B(n70445), .Y(n70482) );
  NAND2xp5_ASAP7_75t_SL U58529 ( .A(n70261), .B(n70280), .Y(n70409) );
  OAI22xp33_ASAP7_75t_SL U58530 ( .A1(n65761), .A2(n65646), .B1(n65758), .B2(
        n66181), .Y(n65627) );
  INVx1_ASAP7_75t_SL U58531 ( .A(n72095), .Y(n72122) );
  INVxp33_ASAP7_75t_SL U58532 ( .A(n76406), .Y(n76337) );
  INVxp67_ASAP7_75t_SL U58533 ( .A(n72093), .Y(n72119) );
  NAND2xp5_ASAP7_75t_SL U58534 ( .A(n68940), .B(n69053), .Y(n68893) );
  OAI22xp33_ASAP7_75t_SL U58535 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_), .A2(
        n59633), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_24_), .B2(
        n70488), .Y(n70307) );
  NAND2xp33_ASAP7_75t_SL U58536 ( .A(n65378), .B(n65419), .Y(n65456) );
  INVxp33_ASAP7_75t_SL U58537 ( .A(n76427), .Y(n74026) );
  INVxp67_ASAP7_75t_SL U58538 ( .A(n76366), .Y(n76435) );
  INVxp67_ASAP7_75t_SL U58539 ( .A(n76444), .Y(n76446) );
  INVx1_ASAP7_75t_SL U58540 ( .A(n74004), .Y(n74599) );
  AOI22xp33_ASAP7_75t_SL U58541 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[20]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[20]), 
        .B2(n74538), .Y(n74228) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58542 ( .A1(n2499), .A2(n69335), .B(n62018), .C(
        n62017), .Y(n62023) );
  AOI22xp33_ASAP7_75t_SL U58543 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[11]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[11]), 
        .B2(n74538), .Y(n74388) );
  INVxp67_ASAP7_75t_SL U58544 ( .A(n76671), .Y(n76669) );
  INVxp33_ASAP7_75t_SL U58545 ( .A(n74771), .Y(n74759) );
  INVxp67_ASAP7_75t_SL U58546 ( .A(n61012), .Y(n61001) );
  INVxp33_ASAP7_75t_SL U58547 ( .A(n66208), .Y(n66210) );
  NAND2xp5_ASAP7_75t_SL U58548 ( .A(n73889), .B(n74066), .Y(n74269) );
  AOI22xp33_ASAP7_75t_SL U58549 ( .A1(n70542), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_15_), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_16_), .B2(
        n74686), .Y(n70357) );
  INVxp67_ASAP7_75t_SL U58550 ( .A(n74008), .Y(n74012) );
  NAND2xp33_ASAP7_75t_SL U58551 ( .A(n2335), .B(n70543), .Y(n70319) );
  NAND2xp33_ASAP7_75t_SL U58552 ( .A(n70354), .B(n70543), .Y(n70356) );
  AOI22xp33_ASAP7_75t_SL U58553 ( .A1(n70542), .A2(n74691), .B1(n74645), .B2(
        n74686), .Y(n70320) );
  NAND3xp33_ASAP7_75t_SRAM U58554 ( .A(n74665), .B(n2345), .C(n74664), .Y(
        n74669) );
  INVxp33_ASAP7_75t_SL U58555 ( .A(n73786), .Y(n73692) );
  NAND2xp5_ASAP7_75t_SL U58556 ( .A(n77338), .B(n77345), .Y(n59950) );
  NAND2xp33_ASAP7_75t_SL U58557 ( .A(n74644), .B(n70543), .Y(n70315) );
  AOI22xp33_ASAP7_75t_SL U58558 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[17]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[17]), 
        .B2(n74538), .Y(n74428) );
  AOI22xp33_ASAP7_75t_SL U58559 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_19_), .A2(
        n70542), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .B2(
        n74686), .Y(n70316) );
  AOI22xp33_ASAP7_75t_SL U58560 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[4]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[4]), 
        .B2(n74538), .Y(n74381) );
  AOI22xp33_ASAP7_75t_SL U58561 ( .A1(n70542), .A2(n74657), .B1(n74646), .B2(
        n74686), .Y(n70392) );
  NAND2xp33_ASAP7_75t_SL U58562 ( .A(n2442), .B(n70543), .Y(n70391) );
  INVx1_ASAP7_75t_SL U58563 ( .A(n73645), .Y(n73662) );
  NOR2x1_ASAP7_75t_SL U58564 ( .A(n57083), .B(n61281), .Y(n77773) );
  AOI22xp33_ASAP7_75t_SL U58565 ( .A1(n70542), .A2(n74646), .B1(n70379), .B2(
        n74686), .Y(n70381) );
  INVxp33_ASAP7_75t_SL U58566 ( .A(n77063), .Y(n77068) );
  INVxp67_ASAP7_75t_SL U58567 ( .A(n73983), .Y(n76360) );
  INVxp67_ASAP7_75t_SL U58568 ( .A(n73977), .Y(n76358) );
  AOI22xp33_ASAP7_75t_SL U58569 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_16_), .A2(
        n70542), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_), .B2(
        n74686), .Y(n70346) );
  NAND2xp33_ASAP7_75t_SL U58570 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_15_), .B(
        n70543), .Y(n70347) );
  NAND2xp33_ASAP7_75t_SL U58571 ( .A(n65311), .B(n65400), .Y(n65241) );
  INVx1_ASAP7_75t_SL U58572 ( .A(n74639), .Y(n77883) );
  AOI22xp33_ASAP7_75t_SL U58573 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[3]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[3]), 
        .B2(n74538), .Y(n74376) );
  OAI21xp33_ASAP7_75t_SL U58574 ( .A1(n74643), .A2(n70488), .B(n70336), .Y(
        n70337) );
  NAND2xp5_ASAP7_75t_SL U58575 ( .A(n61031), .B(n60720), .Y(n60718) );
  INVxp33_ASAP7_75t_SL U58576 ( .A(n75720), .Y(n76341) );
  INVxp67_ASAP7_75t_SL U58577 ( .A(n74756), .Y(n74753) );
  INVxp67_ASAP7_75t_SL U58578 ( .A(n74900), .Y(n76948) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58579 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_1_), 
        .A2(n74820), .B(n74819), .C(n74818), .Y(n74821) );
  OAI22xp33_ASAP7_75t_SL U58580 ( .A1(n65758), .A2(n65646), .B1(n65583), .B2(
        n66181), .Y(n66123) );
  INVxp33_ASAP7_75t_SL U58581 ( .A(n74166), .Y(n74167) );
  INVxp67_ASAP7_75t_SL U58582 ( .A(n72105), .Y(n72027) );
  INVx1_ASAP7_75t_SL U58583 ( .A(n77971), .Y(n77615) );
  INVx1_ASAP7_75t_SL U58584 ( .A(n77591), .Y(n77916) );
  INVxp67_ASAP7_75t_SL U58585 ( .A(n74693), .Y(n74642) );
  INVxp67_ASAP7_75t_SL U58586 ( .A(n65419), .Y(n65461) );
  INVx1_ASAP7_75t_SL U58587 ( .A(n77597), .Y(n77977) );
  INVx1_ASAP7_75t_SL U58588 ( .A(n74984), .Y(n77885) );
  INVx1_ASAP7_75t_SL U58589 ( .A(n75781), .Y(n77968) );
  NAND4xp25_ASAP7_75t_SRAM U58590 ( .A(n65419), .B(n65544), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[35]), .D(n65745), 
        .Y(n65406) );
  INVxp67_ASAP7_75t_SL U58591 ( .A(n65670), .Y(n66145) );
  NAND2xp5_ASAP7_75t_SL U58592 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_6_), .B(n74166), 
        .Y(n74174) );
  NAND2xp33_ASAP7_75t_SL U58593 ( .A(n3309), .B(n73686), .Y(n73788) );
  INVx1_ASAP7_75t_SL U58594 ( .A(n76508), .Y(n77992) );
  AOI22xp33_ASAP7_75t_SL U58595 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[19]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[19]), 
        .B2(n74538), .Y(n74446) );
  INVxp33_ASAP7_75t_SL U58596 ( .A(n66196), .Y(n65553) );
  AOI21xp33_ASAP7_75t_SL U58597 ( .A1(n74822), .A2(n76494), .B(n74810), .Y(
        n74812) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58598 ( .A1(n74654), .A2(n74653), .B(n74652), 
        .C(n74651), .Y(n74658) );
  INVxp67_ASAP7_75t_SL U58599 ( .A(n74013), .Y(n76399) );
  NAND2xp33_ASAP7_75t_SL U58600 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_24_), .B(
        n74686), .Y(n70283) );
  INVx1_ASAP7_75t_SL U58601 ( .A(n75022), .Y(n75013) );
  INVxp67_ASAP7_75t_SL U58602 ( .A(n73994), .Y(n76394) );
  NAND2xp5_ASAP7_75t_SL U58603 ( .A(n70270), .B(n70280), .Y(n70419) );
  AOI22xp33_ASAP7_75t_SL U58604 ( .A1(n70542), .A2(n74644), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_19_), .B2(
        n74686), .Y(n70326) );
  INVxp67_ASAP7_75t_SL U58605 ( .A(n73985), .Y(n76386) );
  INVxp33_ASAP7_75t_SL U58606 ( .A(n60572), .Y(n60574) );
  NAND2xp33_ASAP7_75t_SL U58607 ( .A(n73340), .B(n59525), .Y(n73343) );
  NAND2xp5_ASAP7_75t_SL U58608 ( .A(n70289), .B(n70288), .Y(n70455) );
  NAND2xp33_ASAP7_75t_SL U58609 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[1]), .B(n59521), .Y(
        n69592) );
  OAI22xp33_ASAP7_75t_SL U58610 ( .A1(n65367), .A2(n65393), .B1(n65402), .B2(
        n65397), .Y(n65369) );
  INVxp33_ASAP7_75t_SL U58611 ( .A(n76333), .Y(n76335) );
  AOI22xp33_ASAP7_75t_SL U58612 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[29]), .A2(n65634), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[27]), .B2(n66182), .Y(n65622) );
  INVx1_ASAP7_75t_SL U58613 ( .A(n77295), .Y(n77901) );
  NAND2xp33_ASAP7_75t_SL U58614 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .B(
        n70445), .Y(n70293) );
  NAND2xp33_ASAP7_75t_SL U58615 ( .A(DP_OP_741J1_129_6992_n46), .B(n74686), 
        .Y(n70265) );
  INVxp33_ASAP7_75t_SL U58616 ( .A(n71683), .Y(n71684) );
  OAI21xp33_ASAP7_75t_SL U58617 ( .A1(n2335), .A2(n70488), .B(n74706), .Y(
        n70291) );
  INVxp33_ASAP7_75t_SL U58618 ( .A(n78055), .Y(n76848) );
  NAND2xp33_ASAP7_75t_SL U58619 ( .A(n74706), .B(n70348), .Y(n70310) );
  INVxp33_ASAP7_75t_SL U58620 ( .A(n61311), .Y(n60344) );
  AOI22xp33_ASAP7_75t_SL U58621 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[5]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[5]), 
        .B2(n74538), .Y(n74366) );
  INVxp33_ASAP7_75t_SL U58622 ( .A(n77425), .Y(n60333) );
  INVxp33_ASAP7_75t_SL U58623 ( .A(n70646), .Y(n70644) );
  AOI22xp33_ASAP7_75t_SL U58624 ( .A1(n70542), .A2(n2442), .B1(n74657), .B2(
        n74686), .Y(n70396) );
  INVxp67_ASAP7_75t_SL U58625 ( .A(n65529), .Y(n65481) );
  XNOR2xp5_ASAP7_75t_SRAM U58626 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[1]), .B(
        n74066), .Y(n74068) );
  NAND2xp5_ASAP7_75t_SL U58627 ( .A(n70289), .B(n70280), .Y(n70394) );
  AOI22xp33_ASAP7_75t_SL U58628 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[18]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[18]), 
        .B2(n74538), .Y(n74439) );
  NAND2xp33_ASAP7_75t_SL U58629 ( .A(n65383), .B(n65400), .Y(n65382) );
  NAND2xp33_ASAP7_75t_SL U58630 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[6]), .B(n59520), .Y(
        n69611) );
  OAI22xp33_ASAP7_75t_SL U58631 ( .A1(n70327), .A2(n70488), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .B2(
        n70440), .Y(n70328) );
  INVxp67_ASAP7_75t_SL U58632 ( .A(n74098), .Y(n72578) );
  NAND2xp5_ASAP7_75t_SL U58633 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .B(
        n70543), .Y(n70397) );
  INVxp67_ASAP7_75t_SL U58634 ( .A(n66119), .Y(n65582) );
  OAI21xp33_ASAP7_75t_SL U58635 ( .A1(or1200_cpu_or1200_genpc_pcreg_default[2]), .A2(or1200_cpu_or1200_genpc_pcreg_default[3]), .B(n61577), .Y(n61585) );
  NAND2xp33_ASAP7_75t_SL U58636 ( .A(n60980), .B(n60845), .Y(n76352) );
  NAND2xp33_ASAP7_75t_SL U58637 ( .A(n72611), .B(n71538), .Y(n72646) );
  OAI21xp33_ASAP7_75t_SL U58638 ( .A1(n73618), .A2(n73831), .B(n73797), .Y(
        n73703) );
  INVx1_ASAP7_75t_SL U58639 ( .A(n76828), .Y(n77986) );
  INVxp67_ASAP7_75t_SL U58640 ( .A(n68823), .Y(n68785) );
  INVx1_ASAP7_75t_SL U58641 ( .A(n77646), .Y(n77893) );
  OAI22xp33_ASAP7_75t_SL U58642 ( .A1(n65853), .A2(n65646), .B1(n65743), .B2(
        n66181), .Y(n65599) );
  NAND2xp5_ASAP7_75t_SL U58643 ( .A(n72579), .B(n74098), .Y(n72582) );
  NAND2xp5_ASAP7_75t_SL U58644 ( .A(n69189), .B(n69193), .Y(n69181) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58645 ( .A1(n59527), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .C(
        n72248), .Y(n72249) );
  NAND2xp33_ASAP7_75t_SL U58646 ( .A(n59881), .B(n60293), .Y(n60196) );
  NOR2x1_ASAP7_75t_SL U58647 ( .A(n74755), .B(n60690), .Y(n77090) );
  INVxp33_ASAP7_75t_SL U58648 ( .A(n73491), .Y(n73503) );
  INVxp67_ASAP7_75t_SL U58649 ( .A(n60198), .Y(n59886) );
  INVxp67_ASAP7_75t_SL U58650 ( .A(n66138), .Y(n66110) );
  NAND2xp33_ASAP7_75t_SL U58651 ( .A(n65392), .B(n65394), .Y(n65355) );
  NAND2xp33_ASAP7_75t_SL U58652 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[44]), .B(n66182), 
        .Y(n65503) );
  NAND2xp5_ASAP7_75t_SL U58653 ( .A(n69425), .B(n78244), .Y(n69443) );
  INVx1_ASAP7_75t_SL U58654 ( .A(n63508), .Y(n63491) );
  NAND2xp5_ASAP7_75t_SL U58655 ( .A(or1200_cpu_or1200_mult_mac_n135), .B(
        n75759), .Y(n63245) );
  INVxp67_ASAP7_75t_SL U58656 ( .A(n74770), .Y(n74831) );
  OAI22xp33_ASAP7_75t_SL U58657 ( .A1(n58400), .A2(n73739), .B1(n73755), .B2(
        n58622), .Y(n73714) );
  OAI21xp33_ASAP7_75t_SL U58658 ( .A1(n65494), .A2(n65493), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]), .Y(n76978) );
  INVxp33_ASAP7_75t_SL U58659 ( .A(n63719), .Y(n63720) );
  INVxp33_ASAP7_75t_SL U58660 ( .A(n69279), .Y(n69276) );
  INVxp33_ASAP7_75t_SL U58661 ( .A(n62430), .Y(n60661) );
  INVxp33_ASAP7_75t_SL U58662 ( .A(n74938), .Y(n74939) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58663 ( .A1(n69282), .A2(n69281), .B(n69280), .C(
        n69279), .Y(n69286) );
  NOR2x1_ASAP7_75t_SL U58664 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_4_), .B(n65394), .Y(
        n65391) );
  INVxp33_ASAP7_75t_SL U58665 ( .A(n63519), .Y(n63521) );
  INVxp33_ASAP7_75t_SL U58666 ( .A(n61577), .Y(n61569) );
  NOR2xp33_ASAP7_75t_SRAM U58667 ( .A(n57082), .B(n61539), .Y(n61525) );
  NAND2xp5_ASAP7_75t_SL U58668 ( .A(n77208), .B(n69350), .Y(n69349) );
  NAND2xp33_ASAP7_75t_SL U58669 ( .A(or1200_cpu_spr_dat_rf[1]), .B(n61056), 
        .Y(n61055) );
  INVxp67_ASAP7_75t_SL U58670 ( .A(n70385), .Y(n69379) );
  NAND2xp33_ASAP7_75t_SL U58671 ( .A(n65257), .B(n65402), .Y(n2475) );
  INVx1_ASAP7_75t_SL U58672 ( .A(n74079), .Y(n77869) );
  OAI21xp33_ASAP7_75t_SL U58673 ( .A1(n58619), .A2(n73739), .B(n73724), .Y(
        n73727) );
  NAND2xp33_ASAP7_75t_SL U58674 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_0_), .B(n65402), .Y(
        n2018) );
  AOI21xp33_ASAP7_75t_SL U58675 ( .A1(n69355), .A2(n59729), .B(n59728), .Y(
        n59731) );
  INVx1_ASAP7_75t_SL U58676 ( .A(n77890), .Y(n76235) );
  AOI22xp33_ASAP7_75t_SL U58677 ( .A1(n70583), .A2(n70582), .B1(n70581), .B2(
        n70580), .Y(n70584) );
  INVx2_ASAP7_75t_SL U58678 ( .A(n59646), .Y(n57196) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58679 ( .A1(n59527), .A2(n72350), .B(n72367), .C(
        n72349), .Y(n72353) );
  NAND4xp25_ASAP7_75t_SRAM U58680 ( .A(n59405), .B(n59575), .C(n59573), .D(
        n59563), .Y(n61405) );
  NAND2xp5_ASAP7_75t_SL U58681 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[23]), .B(n59521), .Y(
        n69711) );
  OAI21xp33_ASAP7_75t_SL U58682 ( .A1(n63776), .A2(n63775), .B(n63774), .Y(
        n64171) );
  OAI21xp5_ASAP7_75t_SL U58683 ( .A1(n73640), .A2(n73639), .B(n73752), .Y(
        n73808) );
  INVxp67_ASAP7_75t_SL U58684 ( .A(n60573), .Y(n60544) );
  INVxp33_ASAP7_75t_SL U58685 ( .A(n72411), .Y(n71973) );
  INVx1_ASAP7_75t_SL U58686 ( .A(n65346), .Y(n65354) );
  NAND2x1p5_ASAP7_75t_SL U58687 ( .A(n63176), .B(n63179), .Y(n63173) );
  INVx1_ASAP7_75t_SL U58688 ( .A(n75620), .Y(n77873) );
  INVx1_ASAP7_75t_SL U58689 ( .A(n59852), .Y(n59787) );
  AOI21xp33_ASAP7_75t_SL U58690 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_2_), .A2(n65365), .B(
        n65338), .Y(n65339) );
  INVxp33_ASAP7_75t_SL U58691 ( .A(n65616), .Y(n65566) );
  NAND2x1p5_ASAP7_75t_SL U58692 ( .A(n60595), .B(n57649), .Y(n60915) );
  INVx1_ASAP7_75t_SL U58693 ( .A(n73829), .Y(n73834) );
  AOI22xp33_ASAP7_75t_SL U58694 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[21]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[21]), 
        .B2(n74538), .Y(n74455) );
  NAND2xp33_ASAP7_75t_SL U58695 ( .A(n73373), .B(n73379), .Y(n73376) );
  INVxp33_ASAP7_75t_SL U58696 ( .A(n75774), .Y(n76245) );
  NAND2xp33_ASAP7_75t_SL U58697 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[24]), .B(n70528), .Y(
        n70501) );
  OAI21xp5_ASAP7_75t_SL U58698 ( .A1(n60260), .A2(n60259), .B(
        or1200_cpu_or1200_except_delayed_iee[2]), .Y(n60264) );
  AOI31xp33_ASAP7_75t_SRAM U58699 ( .A1(n59520), .A2(n57081), .A3(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[26]), .B(n70527), .Y(
        n2262) );
  NAND2xp5_ASAP7_75t_SL U58700 ( .A(n73487), .B(n73491), .Y(n73530) );
  INVxp67_ASAP7_75t_SL U58701 ( .A(n61913), .Y(n59017) );
  INVxp67_ASAP7_75t_SL U58702 ( .A(n68990), .Y(n69051) );
  INVxp67_ASAP7_75t_SL U58703 ( .A(n73770), .Y(n73705) );
  INVx1_ASAP7_75t_SL U58704 ( .A(n77254), .Y(n63743) );
  INVxp67_ASAP7_75t_SL U58705 ( .A(n75710), .Y(n62433) );
  NAND2xp33_ASAP7_75t_SL U58706 ( .A(n65264), .B(n65402), .Y(n1550) );
  INVxp33_ASAP7_75t_SL U58707 ( .A(n73611), .Y(n73612) );
  NAND2xp33_ASAP7_75t_SL U58708 ( .A(n65274), .B(n65402), .Y(n1556) );
  INVxp67_ASAP7_75t_SL U58709 ( .A(n77922), .Y(n77583) );
  NAND2xp33_ASAP7_75t_SL U58710 ( .A(n75416), .B(n65204), .Y(n65208) );
  NAND2xp33_ASAP7_75t_SL U58711 ( .A(n60954), .B(n62595), .Y(n60974) );
  OAI22xp33_ASAP7_75t_SL U58712 ( .A1(n65831), .A2(n65646), .B1(n65833), .B2(
        n66181), .Y(n65575) );
  INVx1_ASAP7_75t_SL U58713 ( .A(n65393), .Y(n65401) );
  INVxp33_ASAP7_75t_SL U58714 ( .A(n71931), .Y(n71933) );
  INVxp67_ASAP7_75t_SL U58715 ( .A(n74500), .Y(n69524) );
  AOI21xp33_ASAP7_75t_SL U58716 ( .A1(n63427), .A2(n63426), .B(n63425), .Y(
        n63526) );
  INVxp67_ASAP7_75t_SL U58717 ( .A(n61058), .Y(n60728) );
  AOI21xp5_ASAP7_75t_SL U58718 ( .A1(n78095), .A2(n59797), .B(n69357), .Y(
        n59801) );
  INVx1_ASAP7_75t_SL U58719 ( .A(n69107), .Y(n69111) );
  NAND2xp33_ASAP7_75t_SL U58720 ( .A(n75441), .B(n75440), .Y(n75443) );
  INVx1_ASAP7_75t_SL U58721 ( .A(n69361), .Y(n78094) );
  INVxp67_ASAP7_75t_SL U58722 ( .A(n77920), .Y(n77585) );
  NAND2xp33_ASAP7_75t_SL U58723 ( .A(n63302), .B(n63301), .Y(n63386) );
  INVxp33_ASAP7_75t_SL U58724 ( .A(n73831), .Y(n73790) );
  NAND2xp5_ASAP7_75t_SL U58725 ( .A(n74137), .B(n65495), .Y(n74134) );
  OAI21xp33_ASAP7_75t_SL U58726 ( .A1(n3327), .A2(n58619), .B(n73632), .Y(
        n73635) );
  INVx1_ASAP7_75t_SL U58727 ( .A(n77603), .Y(n77983) );
  INVxp67_ASAP7_75t_SL U58728 ( .A(n69204), .Y(n69206) );
  NAND2xp5_ASAP7_75t_SL U58729 ( .A(n70223), .B(n70568), .Y(n70238) );
  INVxp67_ASAP7_75t_SL U58730 ( .A(n73715), .Y(n73717) );
  INVxp33_ASAP7_75t_SL U58731 ( .A(n60503), .Y(n60370) );
  AOI22xp33_ASAP7_75t_SL U58732 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[14]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[14]), 
        .B2(n74538), .Y(n74411) );
  INVx2_ASAP7_75t_SL U58733 ( .A(n58547), .Y(n57198) );
  INVx1_ASAP7_75t_SL U58734 ( .A(n77594), .Y(n77974) );
  AND2x2_ASAP7_75t_SL U58735 ( .A(n59994), .B(n77210), .Y(n77253) );
  INVxp67_ASAP7_75t_SL U58736 ( .A(n68943), .Y(n68945) );
  AOI21xp33_ASAP7_75t_SL U58737 ( .A1(n61293), .A2(dc_en), .B(n77410), .Y(
        n61297) );
  INVxp33_ASAP7_75t_SL U58738 ( .A(n60720), .Y(n60721) );
  NAND2xp5_ASAP7_75t_SL U58739 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[21]), .B(n59521), .Y(
        n69704) );
  INVxp33_ASAP7_75t_SL U58740 ( .A(n65400), .Y(n65360) );
  INVxp67_ASAP7_75t_SL U58741 ( .A(n70675), .Y(n70658) );
  AND2x2_ASAP7_75t_SL U58742 ( .A(n58289), .B(n58290), .Y(n60554) );
  INVx1_ASAP7_75t_SL U58743 ( .A(n75431), .Y(n77877) );
  NAND2xp33_ASAP7_75t_SL U58744 ( .A(n65268), .B(n65402), .Y(n1580) );
  AOI21xp5_ASAP7_75t_SL U58745 ( .A1(n63286), .A2(n63308), .B(n63285), .Y(
        n63287) );
  NAND2xp5_ASAP7_75t_SL U58746 ( .A(n1938), .B(n76544), .Y(n74935) );
  AOI22xp33_ASAP7_75t_SL U58747 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[13]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[13]), 
        .B2(n74538), .Y(n74406) );
  NAND2xp33_ASAP7_75t_SL U58748 ( .A(n65301), .B(n65400), .Y(n65253) );
  NOR2x1_ASAP7_75t_SL U58749 ( .A(n59928), .B(n59927), .Y(n64208) );
  AOI22xp33_ASAP7_75t_SL U58750 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[12]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[12]), 
        .B2(n74538), .Y(n74397) );
  AOI22xp33_ASAP7_75t_SL U58751 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[16]), .A2(
        n78437), .B1(or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[16]), 
        .B2(n74538), .Y(n74420) );
  INVx1_ASAP7_75t_SL U58752 ( .A(n77637), .Y(n77899) );
  INVxp67_ASAP7_75t_SL U58753 ( .A(n72806), .Y(n72816) );
  NAND2xp5_ASAP7_75t_SL U58754 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_2_), .B(n74894), .Y(
        n65673) );
  INVxp67_ASAP7_75t_SL U58755 ( .A(n78244), .Y(n69582) );
  AOI21xp33_ASAP7_75t_SL U58756 ( .A1(n59732), .A2(n59824), .B(n74118), .Y(
        n59734) );
  INVx1_ASAP7_75t_SL U58757 ( .A(n72433), .Y(n59623) );
  NAND2xp5_ASAP7_75t_SL U58758 ( .A(n61158), .B(n61139), .Y(n60494) );
  INVx1_ASAP7_75t_SL U58759 ( .A(n72853), .Y(n72815) );
  NAND2xp33_ASAP7_75t_SL U58760 ( .A(n73133), .B(n73379), .Y(n73136) );
  NOR2xp33_ASAP7_75t_SRAM U58761 ( .A(n2814), .B(n60503), .Y(n62019) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58762 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_2_), .A2(n65524), 
        .B(n65523), .C(n66138), .Y(n65535) );
  INVxp33_ASAP7_75t_SL U58763 ( .A(n77223), .Y(n78150) );
  INVxp33_ASAP7_75t_SL U58764 ( .A(n77864), .Y(n75796) );
  INVxp33_ASAP7_75t_SL U58765 ( .A(n77880), .Y(n74127) );
  INVxp67_ASAP7_75t_SL U58766 ( .A(n77862), .Y(n77177) );
  INVx1_ASAP7_75t_SL U58767 ( .A(n77854), .Y(n77673) );
  INVxp67_ASAP7_75t_SL U58768 ( .A(n77866), .Y(n69371) );
  INVxp33_ASAP7_75t_SL U58769 ( .A(n77888), .Y(n75302) );
  AOI21xp33_ASAP7_75t_SL U58770 ( .A1(n71567), .A2(n72319), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .Y(n71545) );
  INVxp67_ASAP7_75t_SL U58771 ( .A(n75653), .Y(n75140) );
  INVxp33_ASAP7_75t_SL U58772 ( .A(n76200), .Y(n76611) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58773 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .B(n65459), 
        .C(n65458), .Y(n65460) );
  NOR2xp33_ASAP7_75t_SRAM U58774 ( .A(n65631), .B(n65653), .Y(n65632) );
  INVxp67_ASAP7_75t_SL U58775 ( .A(n71332), .Y(n71355) );
  NAND2xp5_ASAP7_75t_SL U58776 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_), .B(
        n74064), .Y(n72594) );
  NOR2xp33_ASAP7_75t_SRAM U58777 ( .A(n65630), .B(n65629), .Y(n65633) );
  NAND2xp33_ASAP7_75t_SL U58778 ( .A(n71568), .B(n71567), .Y(n71570) );
  INVxp67_ASAP7_75t_SL U58779 ( .A(n75651), .Y(n75134) );
  NAND2xp5_ASAP7_75t_SL U58780 ( .A(n73595), .B(n73605), .Y(n73611) );
  INVx1_ASAP7_75t_SL U58781 ( .A(n74213), .Y(n74158) );
  NAND2xp33_ASAP7_75t_SL U58782 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .B(n58611), .Y(n71896) );
  INVxp67_ASAP7_75t_SL U58783 ( .A(n70569), .Y(n70221) );
  INVxp67_ASAP7_75t_SL U58784 ( .A(n76904), .Y(n76905) );
  AOI21xp33_ASAP7_75t_SL U58785 ( .A1(or1200_cpu_or1200_mult_mac_n401), .A2(
        n69324), .B(n69323), .Y(n69325) );
  INVxp33_ASAP7_75t_SL U58786 ( .A(n72361), .Y(n72248) );
  NAND2xp33_ASAP7_75t_SL U58787 ( .A(n69322), .B(n69321), .Y(n69327) );
  INVxp67_ASAP7_75t_SL U58788 ( .A(n75129), .Y(n75132) );
  INVxp67_ASAP7_75t_SL U58789 ( .A(n75127), .Y(n69328) );
  INVxp67_ASAP7_75t_SL U58790 ( .A(n59850), .Y(n59825) );
  INVx1_ASAP7_75t_SL U58791 ( .A(n72147), .Y(n72116) );
  OAI22xp33_ASAP7_75t_SL U58792 ( .A1(n75653), .A2(n75652), .B1(
        or1200_cpu_or1200_mult_mac_n409), .B2(n75654), .Y(n75656) );
  INVxp67_ASAP7_75t_SL U58793 ( .A(n72126), .Y(n72067) );
  NAND2xp5_ASAP7_75t_SL U58794 ( .A(n4042), .B(n4041), .Y(n77971) );
  INVxp67_ASAP7_75t_SL U58795 ( .A(n70133), .Y(n70134) );
  INVxp33_ASAP7_75t_SL U58796 ( .A(n70578), .Y(n70577) );
  NAND2xp5_ASAP7_75t_SL U58797 ( .A(n72573), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_0_), .Y(
        n72575) );
  INVx1_ASAP7_75t_SL U58798 ( .A(n77752), .Y(n61626) );
  AOI21xp33_ASAP7_75t_SL U58799 ( .A1(n3321), .A2(n59705), .B(n73797), .Y(
        n73798) );
  NAND3xp33_ASAP7_75t_SRAM U58800 ( .A(n62142), .B(n2589), .C(n2814), .Y(
        n61142) );
  NAND2xp33_ASAP7_75t_SL U58801 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .B(n71888), .Y(n71773) );
  INVxp33_ASAP7_75t_SL U58802 ( .A(n59990), .Y(n59992) );
  INVxp67_ASAP7_75t_SL U58803 ( .A(n76201), .Y(n76859) );
  INVxp67_ASAP7_75t_SL U58804 ( .A(n69203), .Y(n69196) );
  INVxp33_ASAP7_75t_SL U58805 ( .A(n70168), .Y(n70165) );
  INVxp67_ASAP7_75t_SL U58806 ( .A(n71670), .Y(n71636) );
  INVxp67_ASAP7_75t_SL U58807 ( .A(n76627), .Y(n57229) );
  OAI22xp33_ASAP7_75t_SL U58808 ( .A1(n71671), .A2(n71670), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_8_), .B2(
        n71669), .Y(n71672) );
  NAND2xp33_ASAP7_75t_SL U58809 ( .A(n65822), .B(n65537), .Y(n65541) );
  INVxp33_ASAP7_75t_SL U58810 ( .A(n70694), .Y(n70642) );
  OAI21xp33_ASAP7_75t_SL U58811 ( .A1(or1200_cpu_or1200_mult_mac_n243), .A2(
        n69201), .B(n74569), .Y(n69202) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U58812 ( .A1(n59527), .A2(n72054), .B(n72033), .C(
        n72367), .Y(n72035) );
  INVxp67_ASAP7_75t_SL U58813 ( .A(n71772), .Y(n71775) );
  NAND2xp33_ASAP7_75t_SL U58814 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_), 
        .B(n71888), .Y(n71803) );
  NOR2x1_ASAP7_75t_SL U58815 ( .A(n61806), .B(n61807), .Y(n61911) );
  NAND2xp5_ASAP7_75t_SL U58816 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_3_), .B(n74902), 
        .Y(n74900) );
  NOR2x1p5_ASAP7_75t_SL U58817 ( .A(n59709), .B(n61921), .Y(n58168) );
  INVxp33_ASAP7_75t_SL U58818 ( .A(n61031), .Y(n61032) );
  INVxp67_ASAP7_75t_SL U58819 ( .A(n72293), .Y(n72295) );
  INVx3_ASAP7_75t_SL U58820 ( .A(n58169), .Y(n57199) );
  NAND2xp33_ASAP7_75t_SL U58821 ( .A(n72367), .B(n72196), .Y(n72177) );
  INVx1_ASAP7_75t_SL U58822 ( .A(n61140), .Y(n61158) );
  INVxp67_ASAP7_75t_SL U58823 ( .A(n72342), .Y(n72343) );
  NAND2xp5_ASAP7_75t_SL U58824 ( .A(n69248), .B(n69249), .Y(n69216) );
  INVxp33_ASAP7_75t_SL U58825 ( .A(n64324), .Y(n60691) );
  NOR2xp33_ASAP7_75t_SRAM U58826 ( .A(n74496), .B(n74495), .Y(n74498) );
  NAND2xp5_ASAP7_75t_SL U58827 ( .A(n70168), .B(n70167), .Y(n70155) );
  INVx1_ASAP7_75t_SL U58828 ( .A(n72085), .Y(n72110) );
  NAND2xp33_ASAP7_75t_SL U58829 ( .A(n2616), .B(n60343), .Y(n60351) );
  NAND2xp5_ASAP7_75t_SL U58830 ( .A(n65631), .B(n65469), .Y(n66196) );
  AOI31xp33_ASAP7_75t_SRAM U58831 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .A2(n71984), .A3(n71995), .B(n71606), .Y(n71607) );
  AOI21xp33_ASAP7_75t_SL U58832 ( .A1(n73753), .A2(n59705), .B(n73793), .Y(
        n73761) );
  NAND2xp33_ASAP7_75t_SL U58833 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_), 
        .B(n71888), .Y(n71878) );
  INVxp67_ASAP7_75t_SL U58834 ( .A(n59945), .Y(n77013) );
  NAND2xp5_ASAP7_75t_SL U58835 ( .A(n69248), .B(n69247), .Y(n69250) );
  AND2x2_ASAP7_75t_SL U58836 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .B(
        n72517), .Y(n72364) );
  INVxp33_ASAP7_75t_SL U58837 ( .A(n60860), .Y(n60861) );
  INVxp33_ASAP7_75t_SL U58838 ( .A(n74064), .Y(n72597) );
  OAI21xp5_ASAP7_75t_SL U58839 ( .A1(n63977), .A2(n63976), .B(n63975), .Y(
        n63978) );
  NAND2xp5_ASAP7_75t_SL U58840 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[16]), .B(n70676), 
        .Y(n70677) );
  NAND2xp33_ASAP7_75t_SL U58841 ( .A(n76619), .B(n62263), .Y(n76792) );
  INVxp67_ASAP7_75t_SL U58842 ( .A(n77483), .Y(n61302) );
  INVx1_ASAP7_75t_SL U58843 ( .A(n59856), .Y(n59794) );
  INVx1_ASAP7_75t_SL U58844 ( .A(n61539), .Y(n57200) );
  INVx1_ASAP7_75t_SL U58845 ( .A(n74496), .Y(n69522) );
  INVx1_ASAP7_75t_SL U58846 ( .A(n77082), .Y(n76791) );
  INVx1_ASAP7_75t_SL U58847 ( .A(n59864), .Y(n78095) );
  NAND2xp5_ASAP7_75t_SL U58848 ( .A(n59799), .B(n59798), .Y(n69361) );
  NAND2xp5_ASAP7_75t_SL U58849 ( .A(n74731), .B(n74302), .Y(n73856) );
  NAND2xp33_ASAP7_75t_SL U58850 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_3_), .B(n66136), .Y(
        n66135) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58851 ( .A1(n71495), .A2(n72080), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_), 
        .C(n72141), .Y(n71499) );
  INVxp67_ASAP7_75t_SL U58852 ( .A(n57407), .Y(n59492) );
  INVxp67_ASAP7_75t_SL U58853 ( .A(n69527), .Y(n69528) );
  INVx1_ASAP7_75t_SL U58854 ( .A(n63125), .Y(n57201) );
  NAND2xp5_ASAP7_75t_SL U58855 ( .A(n3092), .B(n61285), .Y(n61318) );
  NAND2xp5_ASAP7_75t_SL U58856 ( .A(n74529), .B(n74530), .Y(n74771) );
  NAND2xp33_ASAP7_75t_SL U58857 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .B(n58447), .Y(n72021) );
  NAND2xp33_ASAP7_75t_SL U58858 ( .A(ic_en), .B(n77354), .Y(n77501) );
  NAND2xp33_ASAP7_75t_SL U58859 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[0]), .B(
        n70581), .Y(n70585) );
  NAND2xp33_ASAP7_75t_SL U58860 ( .A(n77011), .B(n77015), .Y(n77223) );
  INVxp33_ASAP7_75t_SL U58861 ( .A(n69426), .Y(n69429) );
  INVxp67_ASAP7_75t_SL U58862 ( .A(n69437), .Y(n69427) );
  NAND2xp33_ASAP7_75t_SL U58863 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_35_), 
        .B(n58447), .Y(n72100) );
  INVxp33_ASAP7_75t_SL U58864 ( .A(n71434), .Y(n71632) );
  INVxp67_ASAP7_75t_SL U58865 ( .A(n72962), .Y(n72879) );
  INVxp33_ASAP7_75t_SL U58866 ( .A(n61285), .Y(n77486) );
  INVxp33_ASAP7_75t_SL U58867 ( .A(n73529), .Y(n73531) );
  INVxp33_ASAP7_75t_SL U58868 ( .A(n74461), .Y(n74716) );
  NAND2xp33_ASAP7_75t_SL U58869 ( .A(n69368), .B(n69369), .Y(n74938) );
  NAND2xp33_ASAP7_75t_SL U58870 ( .A(n74206), .B(n74834), .Y(n65490) );
  BUFx2_ASAP7_75t_SL U58871 ( .A(n74744), .Y(n57202) );
  INVxp33_ASAP7_75t_SL U58872 ( .A(n76547), .Y(n59721) );
  AND2x2_ASAP7_75t_SL U58873 ( .A(n57561), .B(n77722), .Y(n57560) );
  INVxp33_ASAP7_75t_SL U58874 ( .A(n59843), .Y(n59813) );
  INVxp67_ASAP7_75t_SL U58875 ( .A(n69369), .Y(n69350) );
  INVxp67_ASAP7_75t_SL U58876 ( .A(n59941), .Y(n76550) );
  INVxp67_ASAP7_75t_SL U58877 ( .A(n57327), .Y(n57326) );
  NOR2xp33_ASAP7_75t_SRAM U58878 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .B(
        n71882), .Y(n71886) );
  NAND2xp5_ASAP7_75t_SL U58879 ( .A(n71529), .B(n72650), .Y(n71534) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U58880 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_13_), 
        .A2(n72313), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_), 
        .C(n71446), .Y(n71450) );
  NAND2xp5_ASAP7_75t_SL U58881 ( .A(n71536), .B(n72649), .Y(n71531) );
  INVx1_ASAP7_75t_SL U58882 ( .A(n73813), .Y(n73816) );
  NAND2xp5_ASAP7_75t_SL U58883 ( .A(n78367), .B(n69435), .Y(n69436) );
  INVxp67_ASAP7_75t_SL U58884 ( .A(n70572), .Y(n70574) );
  NOR2xp33_ASAP7_75t_SRAM U58885 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .B(
        n71856), .Y(n71859) );
  INVxp33_ASAP7_75t_SL U58886 ( .A(n77751), .Y(n60591) );
  INVxp33_ASAP7_75t_SL U58887 ( .A(n59866), .Y(n75191) );
  NAND2xp33_ASAP7_75t_SL U58888 ( .A(n77708), .B(n77755), .Y(n77754) );
  INVxp33_ASAP7_75t_SL U58889 ( .A(n59935), .Y(n76638) );
  INVx1_ASAP7_75t_SL U58890 ( .A(n74189), .Y(n66220) );
  INVxp33_ASAP7_75t_SL U58891 ( .A(n60844), .Y(n60845) );
  INVxp67_ASAP7_75t_SL U58892 ( .A(n76453), .Y(n64289) );
  INVxp67_ASAP7_75t_SL U58893 ( .A(n71550), .Y(n71563) );
  INVx1_ASAP7_75t_SL U58894 ( .A(n62254), .Y(n77757) );
  AOI22xp33_ASAP7_75t_SL U58895 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_), 
        .A2(n59527), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .B2(n72517), .Y(n72006) );
  AND3x1_ASAP7_75t_SL U58896 ( .A(n65537), .B(n65822), .C(n65821), .Y(n65403)
         );
  INVxp67_ASAP7_75t_SL U58897 ( .A(n58276), .Y(n57389) );
  INVxp67_ASAP7_75t_SL U58898 ( .A(n59429), .Y(n57388) );
  INVxp33_ASAP7_75t_SL U58899 ( .A(n59775), .Y(n59777) );
  NOR2xp33_ASAP7_75t_SRAM U58900 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .B(
        n71874), .Y(n71876) );
  NOR2xp33_ASAP7_75t_SL U58901 ( .A(n59552), .B(n62762), .Y(n73992) );
  NAND2xp5_ASAP7_75t_SL U58902 ( .A(n73818), .B(n73817), .Y(n73829) );
  INVxp33_ASAP7_75t_SL U58903 ( .A(n61646), .Y(n60920) );
  NAND2xp5_ASAP7_75t_SL U58904 ( .A(n59526), .B(n70694), .Y(n70646) );
  NAND2xp5_ASAP7_75t_SL U58905 ( .A(n76657), .B(n77210), .Y(n76503) );
  AOI21xp33_ASAP7_75t_SL U58906 ( .A1(n59698), .A2(n71365), .B(n70676), .Y(
        n70643) );
  INVxp67_ASAP7_75t_SL U58907 ( .A(n71473), .Y(n71490) );
  INVxp67_ASAP7_75t_SL U58908 ( .A(n77756), .Y(n77729) );
  INVx1_ASAP7_75t_SL U58909 ( .A(n59934), .Y(n76639) );
  INVxp67_ASAP7_75t_SL U58910 ( .A(n71446), .Y(n71476) );
  INVxp33_ASAP7_75t_SL U58911 ( .A(n60954), .Y(n60930) );
  NAND2xp5_ASAP7_75t_SL U58912 ( .A(n69351), .B(n69369), .Y(n60218) );
  NOR2x1p5_ASAP7_75t_SL U58913 ( .A(n60919), .B(n64617), .Y(n60946) );
  INVx1_ASAP7_75t_SL U58914 ( .A(n76657), .Y(n77678) );
  NAND2xp33_ASAP7_75t_SL U58915 ( .A(n72341), .B(n71888), .Y(n71832) );
  INVx1_ASAP7_75t_SL U58916 ( .A(n77015), .Y(n77014) );
  NAND2xp5_ASAP7_75t_SL U58917 ( .A(n60246), .B(n60245), .Y(n60260) );
  INVxp33_ASAP7_75t_SL U58918 ( .A(n72502), .Y(n72482) );
  NAND2xp33_ASAP7_75t_SL U58919 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_), 
        .B(n58611), .Y(n71813) );
  INVxp67_ASAP7_75t_SL U58920 ( .A(n73865), .Y(n73889) );
  INVxp67_ASAP7_75t_SL U58921 ( .A(n73501), .Y(n73487) );
  INVx1_ASAP7_75t_SL U58922 ( .A(n77349), .Y(n77337) );
  INVxp33_ASAP7_75t_SL U58923 ( .A(n59926), .Y(n77150) );
  NAND2xp5_ASAP7_75t_SL U58924 ( .A(n61145), .B(n61030), .Y(n60500) );
  INVx1_ASAP7_75t_SL U58925 ( .A(n72546), .Y(n72443) );
  NAND2xp5_ASAP7_75t_SL U58926 ( .A(n73864), .B(n73865), .Y(n73890) );
  NOR2xp33_ASAP7_75t_SRAM U58927 ( .A(n65758), .B(n65653), .Y(n65576) );
  INVx1_ASAP7_75t_SL U58928 ( .A(n75632), .Y(n60002) );
  NAND2xp5_ASAP7_75t_SL U58929 ( .A(n73485), .B(n73499), .Y(n73533) );
  INVxp33_ASAP7_75t_SL U58930 ( .A(n73541), .Y(n73538) );
  INVxp33_ASAP7_75t_SL U58931 ( .A(n62590), .Y(n62595) );
  NAND2xp5_ASAP7_75t_SL U58932 ( .A(n59700), .B(n60277), .Y(n59953) );
  OAI21xp33_ASAP7_75t_SL U58933 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[24]), .A2(
        n73115), .B(n73103), .Y(n73101) );
  INVxp33_ASAP7_75t_SL U58934 ( .A(n73372), .Y(n73374) );
  OAI21xp33_ASAP7_75t_SL U58935 ( .A1(n73333), .A2(n73100), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[23]), .Y(
        n73102) );
  INVxp33_ASAP7_75t_SL U58936 ( .A(n73147), .Y(n73148) );
  INVx1_ASAP7_75t_SL U58937 ( .A(n73100), .Y(n73341) );
  INVxp33_ASAP7_75t_SL U58938 ( .A(n59855), .Y(n59851) );
  NAND2xp5_ASAP7_75t_SL U58939 ( .A(n78435), .B(n65398), .Y(n65322) );
  INVx1_ASAP7_75t_SL U58940 ( .A(n69048), .Y(n68844) );
  NAND2xp33_ASAP7_75t_SL U58941 ( .A(n69061), .B(n69060), .Y(n69062) );
  INVxp67_ASAP7_75t_SL U58942 ( .A(n59764), .Y(n59728) );
  NOR2x1_ASAP7_75t_SL U58943 ( .A(n78435), .B(n65398), .Y(n65400) );
  INVxp33_ASAP7_75t_SL U58944 ( .A(n59821), .Y(n59732) );
  INVxp33_ASAP7_75t_SL U58945 ( .A(n70371), .Y(n70467) );
  INVxp33_ASAP7_75t_SL U58946 ( .A(n75143), .Y(n75144) );
  NAND2xp5_ASAP7_75t_SL U58947 ( .A(n63375), .B(n63306), .Y(n63286) );
  INVx1_ASAP7_75t_SL U58948 ( .A(n73086), .Y(n73084) );
  NAND2xp33_ASAP7_75t_SL U58949 ( .A(n63274), .B(n63273), .Y(n63301) );
  INVxp33_ASAP7_75t_SL U58950 ( .A(n62056), .Y(n62055) );
  NAND2xp33_ASAP7_75t_SL U58951 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_state), 
        .B(n62056), .Y(n62061) );
  NAND2xp5_ASAP7_75t_SL U58952 ( .A(n76937), .B(n76936), .Y(n76958) );
  INVx1_ASAP7_75t_SL U58953 ( .A(n63302), .Y(n63304) );
  INVx1_ASAP7_75t_SL U58954 ( .A(n63374), .Y(n63382) );
  NAND2xp5_ASAP7_75t_SL U58955 ( .A(n63307), .B(n63306), .Y(n63383) );
  OAI21xp33_ASAP7_75t_SL U58956 ( .A1(n73078), .A2(n73134), .B(n73077), .Y(
        n73080) );
  INVxp67_ASAP7_75t_SL U58957 ( .A(n73085), .Y(n73082) );
  AOI21xp33_ASAP7_75t_SL U58958 ( .A1(or1200_cpu_or1200_mult_mac_n203), .A2(
        n75508), .B(n76883), .Y(n68817) );
  NAND2xp5_ASAP7_75t_SL U58959 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[24]), .B(n70526), .Y(
        n70500) );
  INVxp33_ASAP7_75t_SL U58960 ( .A(n63385), .Y(n63396) );
  INVxp67_ASAP7_75t_SL U58961 ( .A(n73103), .Y(n73104) );
  AOI21xp33_ASAP7_75t_SL U58962 ( .A1(n63379), .A2(n63378), .B(n63377), .Y(
        n63380) );
  INVxp33_ASAP7_75t_SL U58963 ( .A(n63424), .Y(n63413) );
  INVxp33_ASAP7_75t_SL U58964 ( .A(n69356), .Y(n69359) );
  INVxp33_ASAP7_75t_SL U58965 ( .A(n69357), .Y(n69358) );
  NAND2xp5_ASAP7_75t_SL U58966 ( .A(n63502), .B(n63505), .Y(n63470) );
  OAI21xp33_ASAP7_75t_SL U58967 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[6]), .A2(
        n73264), .B(n73049), .Y(n73056) );
  INVx1_ASAP7_75t_SL U58968 ( .A(n70542), .Y(n70488) );
  NAND2xp33_ASAP7_75t_SL U58969 ( .A(n63503), .B(n63502), .Y(n63519) );
  INVxp67_ASAP7_75t_SL U58970 ( .A(n73053), .Y(n73050) );
  OAI21xp33_ASAP7_75t_SL U58971 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .A2(
        n70540), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .Y(
        n70329) );
  INVx1_ASAP7_75t_SL U58972 ( .A(n63777), .Y(n63776) );
  NAND2xp33_ASAP7_75t_SL U58973 ( .A(n63778), .B(n63777), .Y(n63779) );
  INVxp33_ASAP7_75t_SL U58974 ( .A(n64170), .Y(n63783) );
  AOI21xp33_ASAP7_75t_SL U58975 ( .A1(n73728), .A2(n59705), .B(n73793), .Y(
        n73733) );
  INVxp67_ASAP7_75t_SL U58976 ( .A(n65092), .Y(n63894) );
  INVxp33_ASAP7_75t_SL U58977 ( .A(n75775), .Y(n75776) );
  INVxp67_ASAP7_75t_SL U58978 ( .A(n69171), .Y(n69087) );
  OAI22xp33_ASAP7_75t_SL U58979 ( .A1(n58423), .A2(n73725), .B1(n58400), .B2(
        n73755), .Y(n73726) );
  INVxp33_ASAP7_75t_SL U58980 ( .A(n76198), .Y(n76612) );
  NAND2xp5_ASAP7_75t_SL U58981 ( .A(n74706), .B(n70386), .Y(n70487) );
  AND2x2_ASAP7_75t_SL U58982 ( .A(n77481), .B(n77480), .Y(n77482) );
  OAI21xp33_ASAP7_75t_SL U58983 ( .A1(n70486), .A2(n70540), .B(n70457), .Y(
        n70458) );
  AOI21xp33_ASAP7_75t_SL U58984 ( .A1(or1200_cpu_or1200_mult_mac_n183), .A2(
        n65095), .B(n65094), .Y(n65096) );
  INVx1_ASAP7_75t_SL U58985 ( .A(n74671), .Y(n74698) );
  INVxp67_ASAP7_75t_SL U58986 ( .A(n73037), .Y(n73002) );
  AOI21xp33_ASAP7_75t_SL U58987 ( .A1(n68940), .A2(n68939), .B(n69052), .Y(
        n68987) );
  NAND2xp5_ASAP7_75t_SL U58988 ( .A(n70229), .B(n70371), .Y(n59520) );
  INVx1_ASAP7_75t_SL U58989 ( .A(n73028), .Y(n73009) );
  INVx1_ASAP7_75t_SL U58990 ( .A(n73030), .Y(n73010) );
  INVx1_ASAP7_75t_SL U58991 ( .A(n62553), .Y(n57345) );
  INVxp67_ASAP7_75t_SL U58992 ( .A(n68877), .Y(n69054) );
  INVxp67_ASAP7_75t_SL U58993 ( .A(n72987), .Y(n73017) );
  INVxp67_ASAP7_75t_SL U58994 ( .A(n57082), .Y(n59379) );
  NAND2xp5_ASAP7_75t_SL U58995 ( .A(n70255), .B(n70281), .Y(n70385) );
  INVx1_ASAP7_75t_SL U58996 ( .A(n62738), .Y(n59397) );
  INVxp33_ASAP7_75t_SL U58997 ( .A(n65332), .Y(n65338) );
  INVx1_ASAP7_75t_SL U58998 ( .A(n68941), .Y(n69053) );
  INVx1_ASAP7_75t_SL U58999 ( .A(n59865), .Y(n75188) );
  INVx1_ASAP7_75t_SL U59000 ( .A(n69366), .Y(n75792) );
  OAI21xp33_ASAP7_75t_SL U59001 ( .A1(or1200_cpu_or1200_mult_mac_n355), .A2(
        or1200_cpu_or1200_mult_mac_n209), .B(n68862), .Y(n68884) );
  OAI21xp33_ASAP7_75t_SL U59002 ( .A1(n72621), .A2(n72620), .B(n72619), .Y(
        n72622) );
  NOR2x1_ASAP7_75t_SL U59003 ( .A(n69521), .B(n69520), .Y(n78243) );
  NOR2x1_ASAP7_75t_SL U59004 ( .A(n69409), .B(n69408), .Y(n78244) );
  INVxp67_ASAP7_75t_SL U59005 ( .A(n77160), .Y(n77199) );
  INVx1_ASAP7_75t_SL U59006 ( .A(n69056), .Y(n69016) );
  INVx1_ASAP7_75t_SL U59007 ( .A(n68874), .Y(n69050) );
  AOI21xp33_ASAP7_75t_SL U59008 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_), .A2(n78371), .B(n72600), 
        .Y(n72601) );
  OAI21xp33_ASAP7_75t_SL U59009 ( .A1(or1200_cpu_or1200_mult_mac_n365), .A2(
        n76721), .B(n68986), .Y(n68990) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U59010 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_1_), .A2(n78435), .B(
        n65366), .C(n65365), .Y(n65397) );
  OAI21xp33_ASAP7_75t_SL U59011 ( .A1(n68842), .A2(n68841), .B(n69048), .Y(
        n68876) );
  INVxp67_ASAP7_75t_SL U59012 ( .A(n62142), .Y(n62145) );
  NAND2xp5_ASAP7_75t_SL U59013 ( .A(n59105), .B(n76673), .Y(n62570) );
  INVxp33_ASAP7_75t_SL U59014 ( .A(n73383), .Y(n73384) );
  NAND2xp33_ASAP7_75t_SL U59015 ( .A(n73833), .B(n59632), .Y(n73669) );
  INVxp67_ASAP7_75t_SL U59016 ( .A(n75016), .Y(n75017) );
  NAND2xp5_ASAP7_75t_SL U59017 ( .A(n75008), .B(n75007), .Y(n75022) );
  NAND2xp5_ASAP7_75t_SL U59018 ( .A(n65144), .B(n65143), .Y(n65163) );
  INVxp67_ASAP7_75t_SL U59019 ( .A(n73208), .Y(n73209) );
  INVxp67_ASAP7_75t_SL U59020 ( .A(n74892), .Y(n74765) );
  AOI21xp33_ASAP7_75t_SL U59021 ( .A1(n73743), .A2(n59705), .B(n73793), .Y(
        n73748) );
  INVxp33_ASAP7_75t_SL U59022 ( .A(n69166), .Y(n69167) );
  INVxp33_ASAP7_75t_SL U59023 ( .A(n70386), .Y(n70402) );
  INVx1_ASAP7_75t_SL U59024 ( .A(n76491), .Y(n74822) );
  OAI22xp33_ASAP7_75t_SL U59025 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_), .A2(
        n70440), .B1(n70264), .B2(n74672), .Y(n70267) );
  INVxp67_ASAP7_75t_SL U59026 ( .A(n73257), .Y(n73258) );
  INVxp67_ASAP7_75t_SL U59027 ( .A(n61312), .Y(n62144) );
  NAND2xp5_ASAP7_75t_SL U59028 ( .A(n69173), .B(n69166), .Y(n69131) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U59029 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_0_), 
        .A2(or1200_cpu_or1200_fpu_b_is_zero), .B(n74815), .C(
        or1200_cpu_or1200_fpu_a_is_zero), .Y(n74820) );
  INVxp33_ASAP7_75t_SL U59030 ( .A(n70229), .Y(n70247) );
  OAI21xp33_ASAP7_75t_SL U59031 ( .A1(or1200_cpu_or1200_mult_mac_n195), .A2(
        n68791), .B(n68790), .Y(n68792) );
  NAND2xp5_ASAP7_75t_SL U59032 ( .A(n68794), .B(n68790), .Y(n65181) );
  INVxp67_ASAP7_75t_SL U59033 ( .A(n63397), .Y(n63336) );
  OAI21xp33_ASAP7_75t_SL U59034 ( .A1(n70540), .A2(n74662), .B(n70306), .Y(
        n70349) );
  NAND2xp33_ASAP7_75t_SL U59035 ( .A(n69166), .B(n69165), .Y(n69170) );
  OAI211xp5_ASAP7_75t_SRAM U59036 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_31_), .A2(n76983), .B(
        n76982), .C(n78251), .Y(n76984) );
  INVxp33_ASAP7_75t_SL U59037 ( .A(n68794), .Y(n68767) );
  NAND2xp5_ASAP7_75t_SL U59038 ( .A(n59881), .B(n59775), .Y(n75672) );
  NAND2xp33_ASAP7_75t_SL U59039 ( .A(n75008), .B(n75010), .Y(n68825) );
  INVxp67_ASAP7_75t_SL U59040 ( .A(n68796), .Y(n68797) );
  INVxp33_ASAP7_75t_SL U59041 ( .A(n77426), .Y(n60379) );
  AOI21xp33_ASAP7_75t_SL U59042 ( .A1(or1200_cpu_or1200_mult_mac_n337), .A2(
        n65165), .B(n65164), .Y(n65166) );
  INVxp67_ASAP7_75t_SL U59043 ( .A(n69191), .Y(n69193) );
  NAND2xp33_ASAP7_75t_SL U59044 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .B(
        n70542), .Y(n70348) );
  INVxp33_ASAP7_75t_SL U59045 ( .A(n60273), .Y(n77793) );
  INVx1_ASAP7_75t_SL U59046 ( .A(n77639), .Y(n77644) );
  INVxp33_ASAP7_75t_SL U59047 ( .A(n70260), .Y(n70261) );
  NAND2xp33_ASAP7_75t_SL U59048 ( .A(n74047), .B(n74081), .Y(n61839) );
  INVxp67_ASAP7_75t_SL U59049 ( .A(n73817), .Y(n73797) );
  INVxp33_ASAP7_75t_SL U59050 ( .A(n71548), .Y(n71558) );
  INVx1_ASAP7_75t_SL U59051 ( .A(n57404), .Y(n62008) );
  NAND2xp5_ASAP7_75t_SL U59052 ( .A(n1983), .B(n60217), .Y(n69369) );
  INVx1_ASAP7_75t_SL U59053 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .Y(
        n72175) );
  AND2x2_ASAP7_75t_SL U59054 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .B(
        n72399), .Y(n72417) );
  NAND2xp33_ASAP7_75t_SL U59055 ( .A(n1832), .B(n77460), .Y(n69351) );
  NAND2xp5_ASAP7_75t_SL U59056 ( .A(or1200_cpu_or1200_mult_mac_n327), .B(
        n65079), .Y(n65091) );
  INVxp33_ASAP7_75t_SL U59057 ( .A(n65145), .Y(n65133) );
  NAND2xp5_ASAP7_75t_SL U59058 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .B(
        n72241), .Y(n72147) );
  OAI21xp33_ASAP7_75t_SL U59059 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .A2(
        n72054), .B(n71822), .Y(n71856) );
  NAND2xp5_ASAP7_75t_SL U59060 ( .A(n1918), .B(n59575), .Y(n59870) );
  NAND2xp33_ASAP7_75t_SL U59061 ( .A(or1200_cpu_or1200_mult_mac_n329), .B(
        n65090), .Y(n65141) );
  INVxp33_ASAP7_75t_SL U59062 ( .A(n71561), .Y(n71562) );
  INVxp33_ASAP7_75t_SL U59063 ( .A(n71560), .Y(n71566) );
  NOR2x1_ASAP7_75t_SL U59064 ( .A(n76826), .B(n59955), .Y(n77210) );
  INVx1_ASAP7_75t_SL U59065 ( .A(n63767), .Y(n63768) );
  NOR2xp33_ASAP7_75t_SRAM U59066 ( .A(n59527), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_), 
        .Y(n72361) );
  NAND2xp5_ASAP7_75t_SL U59067 ( .A(n1798), .B(n75763), .Y(n60216) );
  INVx6_ASAP7_75t_SL U59068 ( .A(n59441), .Y(n59442) );
  INVx1_ASAP7_75t_SL U59069 ( .A(n59705), .Y(n59704) );
  OAI21xp33_ASAP7_75t_SL U59070 ( .A1(n65079), .A2(n65078), .B(n65077), .Y(
        n65080) );
  AOI21xp33_ASAP7_75t_SL U59071 ( .A1(n78336), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[4]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[6]), .Y(n69550)
         );
  AND2x2_ASAP7_75t_SL U59072 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .B(
        n72400), .Y(n72433) );
  NAND2xp5_ASAP7_75t_SL U59073 ( .A(n72544), .B(n72534), .Y(n72507) );
  NAND2xp33_ASAP7_75t_SL U59074 ( .A(n77288), .B(n77227), .Y(n60843) );
  NAND2xp5_ASAP7_75t_SL U59075 ( .A(or1200_cpu_or1200_mult_mac_n195), .B(
        n68791), .Y(n74997) );
  NAND2xp33_ASAP7_75t_SL U59076 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[4]), .B(n65479), .Y(
        n65418) );
  INVxp67_ASAP7_75t_SL U59077 ( .A(n73866), .Y(n73867) );
  NAND2xp5_ASAP7_75t_SL U59078 ( .A(or1200_cpu_or1200_mult_mac_n343), .B(
        n75854), .Y(n75016) );
  NAND2xp33_ASAP7_75t_SL U59079 ( .A(or1200_cpu_or1200_mult_mac_n197), .B(
        n75855), .Y(n75018) );
  INVxp67_ASAP7_75t_SL U59080 ( .A(n71459), .Y(n71588) );
  INVx1_ASAP7_75t_SL U59081 ( .A(n73597), .Y(n73605) );
  INVx1_ASAP7_75t_SL U59082 ( .A(n59561), .Y(n75456) );
  INVxp67_ASAP7_75t_SL U59083 ( .A(n75006), .Y(n75007) );
  NAND2xp5_ASAP7_75t_SL U59084 ( .A(n66170), .B(n66169), .Y(n66177) );
  NAND2xp5_ASAP7_75t_SL U59085 ( .A(n66172), .B(n66171), .Y(n66176) );
  NAND2xp5_ASAP7_75t_SL U59086 ( .A(n66174), .B(n66173), .Y(n66175) );
  NOR2xp33_ASAP7_75t_SRAM U59087 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_), 
        .B(n72360), .Y(n71502) );
  INVxp67_ASAP7_75t_SL U59088 ( .A(n73024), .Y(n72859) );
  NAND2xp33_ASAP7_75t_SL U59089 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_10_), 
        .B(n72362), .Y(n71446) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U59090 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_), 
        .A2(n72162), .B(n72164), .C(n71586), .Y(n71427) );
  INVxp67_ASAP7_75t_SL U59091 ( .A(n71525), .Y(n71528) );
  NAND2xp5_ASAP7_75t_SL U59092 ( .A(or1200_cpu_or1200_mult_mac_n199), .B(
        n68789), .Y(n68796) );
  INVx1_ASAP7_75t_SL U59093 ( .A(n71433), .Y(n71591) );
  NAND2xp5_ASAP7_75t_SL U59094 ( .A(n73040), .B(n72994), .Y(n72962) );
  NAND2xp5_ASAP7_75t_SL U59095 ( .A(n71525), .B(n72641), .Y(n71524) );
  NAND2xp5_ASAP7_75t_SL U59096 ( .A(or1200_cpu_or1200_mult_mac_n345), .B(
        n75219), .Y(n68816) );
  OAI21xp33_ASAP7_75t_SL U59097 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[3]), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[4]), .B(
        n70588), .Y(n70578) );
  NAND2xp5_ASAP7_75t_SL U59098 ( .A(n68879), .B(n68821), .Y(n68815) );
  INVx1_ASAP7_75t_SL U59099 ( .A(n66184), .Y(n66178) );
  NOR3xp33_ASAP7_75t_SRAM U59100 ( .A(n69335), .B(n62052), .C(n2499), .Y(
        n62018) );
  INVxp67_ASAP7_75t_SL U59101 ( .A(n75008), .Y(n68784) );
  INVxp33_ASAP7_75t_SL U59102 ( .A(n62014), .Y(n62015) );
  NAND2xp5_ASAP7_75t_SL U59103 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39), .B(n74063), .Y(n72564) );
  INVxp33_ASAP7_75t_SL U59104 ( .A(n65496), .Y(n65491) );
  NAND2xp33_ASAP7_75t_SL U59105 ( .A(n65507), .B(n74169), .Y(n65494) );
  INVxp67_ASAP7_75t_SL U59106 ( .A(n70588), .Y(n70589) );
  NOR2xp33_ASAP7_75t_SRAM U59107 ( .A(n78248), .B(n78249), .Y(n76982) );
  NAND2xp5_ASAP7_75t_SL U59108 ( .A(DP_OP_741J1_129_6992_n46), .B(n70228), .Y(
        n70569) );
  INVx1_ASAP7_75t_SL U59109 ( .A(n71549), .Y(n71552) );
  NAND2xp5_ASAP7_75t_SL U59110 ( .A(or1200_cpu_or1200_mult_mac_n189), .B(
        n65140), .Y(n65161) );
  INVxp33_ASAP7_75t_SL U59111 ( .A(n74157), .Y(n74767) );
  AND2x2_ASAP7_75t_SL U59112 ( .A(n74468), .B(n74467), .Y(n74469) );
  NAND2xp33_ASAP7_75t_SL U59113 ( .A(or1200_cpu_or1200_mult_mac_n333), .B(
        n75557), .Y(n65143) );
  INVx1_ASAP7_75t_SL U59114 ( .A(n59547), .Y(n77722) );
  NAND2xp5_ASAP7_75t_SL U59115 ( .A(or1200_cpu_or1200_mult_mac_n187), .B(
        n65146), .Y(n65162) );
  INVxp33_ASAP7_75t_SL U59116 ( .A(n71601), .Y(n71625) );
  NAND2xp33_ASAP7_75t_SL U59117 ( .A(n72262), .B(n71950), .Y(n71602) );
  INVx1_ASAP7_75t_SL U59118 ( .A(n65175), .Y(n65151) );
  INVx1_ASAP7_75t_SL U59119 ( .A(n72643), .Y(n72649) );
  NAND2xp5_ASAP7_75t_SL U59120 ( .A(n74475), .B(n74474), .Y(n74481) );
  INVx1_ASAP7_75t_SL U59121 ( .A(n72654), .Y(n72650) );
  NAND2xp33_ASAP7_75t_SL U59122 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_), 
        .B(n72341), .Y(n71620) );
  INVxp33_ASAP7_75t_SL U59123 ( .A(n77759), .Y(n60689) );
  NOR4xp25_ASAP7_75t_SRAM U59124 ( .A(n74652), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_19_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .Y(
        n74648) );
  NAND2xp33_ASAP7_75t_SL U59125 ( .A(n65176), .B(n65175), .Y(n65177) );
  INVxp67_ASAP7_75t_SL U59126 ( .A(n74087), .Y(n74088) );
  A2O1A1Ixp33_ASAP7_75t_SRAM U59127 ( .A1(n74662), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .B(
        n74644), .C(n74643), .Y(n74653) );
  NAND2xp33_ASAP7_75t_SL U59128 ( .A(n2442), .B(n74657), .Y(n74667) );
  NAND2xp5_ASAP7_75t_SL U59129 ( .A(n65787), .B(n65479), .Y(n65404) );
  OAI21xp33_ASAP7_75t_SL U59130 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_), 
        .A2(n72310), .B(n72317), .Y(n71567) );
  INVx1_ASAP7_75t_SL U59131 ( .A(n72976), .Y(n72769) );
  AOI21xp33_ASAP7_75t_SL U59132 ( .A1(n65742), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[45]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[47]), .Y(n65435) );
  NAND2xp5_ASAP7_75t_SL U59133 ( .A(or1200_cpu_or1200_mult_mac_n193), .B(
        n65159), .Y(n68794) );
  INVx2_ASAP7_75t_SL U59134 ( .A(n59539), .Y(n77701) );
  NAND2xp33_ASAP7_75t_SL U59135 ( .A(n66089), .B(n65457), .Y(n65420) );
  NAND2xp5_ASAP7_75t_SL U59136 ( .A(or1200_cpu_or1200_mult_mac_n191), .B(
        n65160), .Y(n68793) );
  INVx1_ASAP7_75t_SL U59137 ( .A(n68779), .Y(n68769) );
  INVxp67_ASAP7_75t_SL U59138 ( .A(n74834), .Y(n74054) );
  NAND2xp33_ASAP7_75t_SL U59139 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_), 
        .B(n72212), .Y(n71420) );
  INVxp33_ASAP7_75t_SL U59140 ( .A(n71627), .Y(n71573) );
  INVx1_ASAP7_75t_SL U59141 ( .A(n71576), .Y(n71455) );
  NAND2xp5_ASAP7_75t_SL U59142 ( .A(n65449), .B(n65447), .Y(n66195) );
  NAND2xp5_ASAP7_75t_SL U59143 ( .A(n71501), .B(n71478), .Y(n71468) );
  NAND2xp33_ASAP7_75t_SL U59144 ( .A(n65784), .B(n65823), .Y(n65538) );
  INVx1_ASAP7_75t_SL U59145 ( .A(n68820), .Y(n75010) );
  NAND2xp33_ASAP7_75t_SL U59146 ( .A(n72350), .B(n71576), .Y(n71417) );
  NAND2xp5_ASAP7_75t_SL U59147 ( .A(n68778), .B(n68777), .Y(n68783) );
  INVx1_ASAP7_75t_SL U59148 ( .A(n72112), .Y(n72062) );
  NAND2xp5_ASAP7_75t_SL U59149 ( .A(or1200_cpu_or1200_mult_mac_n273), .B(
        n63263), .Y(n63264) );
  NAND2xp5_ASAP7_75t_SL U59150 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[26]), .B(
        n73377), .Y(n73106) );
  BUFx2_ASAP7_75t_SL U59151 ( .A(n78184), .Y(n59696) );
  OAI22xp33_ASAP7_75t_SL U59152 ( .A1(n72360), .A2(n58422), .B1(n71890), .B2(
        n72365), .Y(n71838) );
  NAND2xp5_ASAP7_75t_SL U59153 ( .A(n63276), .B(n63275), .Y(n63306) );
  NAND2xp33_ASAP7_75t_SL U59154 ( .A(n59558), .B(n59567), .Y(n60860) );
  NAND2xp5_ASAP7_75t_SL U59155 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_), .B(n78363), .Y(
        n72606) );
  OAI22xp33_ASAP7_75t_SL U59156 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_), .A2(n78361), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_), .B2(n78363), .Y(
        n72607) );
  NAND2xp33_ASAP7_75t_SL U59157 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_), .B(n78381), .Y(
        n72605) );
  INVxp33_ASAP7_75t_SL U59158 ( .A(n2616), .Y(n61136) );
  INVx1_ASAP7_75t_SL U59159 ( .A(n2814), .Y(n60369) );
  INVx1_ASAP7_75t_SL U59160 ( .A(n63307), .Y(n63285) );
  NAND2xp33_ASAP7_75t_SL U59161 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_), .B(n78378), .Y(n72603)
         );
  OAI22xp33_ASAP7_75t_SL U59162 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[19]), .A2(
        n73304), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[20]), .B2(
        n73123), .Y(n73079) );
  OAI21xp33_ASAP7_75t_SL U59163 ( .A1(n2517), .A2(
        or1200_cpu_or1200_except_n586), .B(n63752), .Y(n76578) );
  INVxp33_ASAP7_75t_SL U59164 ( .A(n62036), .Y(n62045) );
  INVxp67_ASAP7_75t_SL U59165 ( .A(n63752), .Y(n63753) );
  OAI21xp33_ASAP7_75t_SL U59166 ( .A1(n2499), .A2(
        or1200_cpu_or1200_except_n589), .B(n63751), .Y(n76588) );
  NAND2xp33_ASAP7_75t_SL U59167 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_30_), .B(n78382), .Y(n72611)
         );
  OAI21xp33_ASAP7_75t_SL U59168 ( .A1(n2464), .A2(
        or1200_cpu_or1200_except_n592), .B(n63750), .Y(n77267) );
  NAND2xp5_ASAP7_75t_SL U59169 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[0]), .B(
        n73231), .Y(n73484) );
  INVxp33_ASAP7_75t_SL U59170 ( .A(n62060), .Y(n62042) );
  INVxp67_ASAP7_75t_SL U59171 ( .A(n60875), .Y(n77749) );
  INVxp67_ASAP7_75t_SL U59172 ( .A(n63750), .Y(n63755) );
  INVx1_ASAP7_75t_SL U59173 ( .A(n62067), .Y(n62064) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U59174 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .A2(
        n72234), .B(n71807), .C(n71894), .Y(n71810) );
  NAND2xp5_ASAP7_75t_SL U59175 ( .A(n63908), .B(n63907), .Y(n63915) );
  INVx1_ASAP7_75t_SL U59176 ( .A(n63305), .Y(n63389) );
  INVx1_ASAP7_75t_SL U59177 ( .A(n72286), .Y(n72355) );
  NAND2xp33_ASAP7_75t_SL U59178 ( .A(n63759), .B(n76841), .Y(n63758) );
  NAND2xp5_ASAP7_75t_SL U59179 ( .A(n63309), .B(n63308), .Y(n63374) );
  INVxp33_ASAP7_75t_SL U59180 ( .A(n63909), .Y(n63913) );
  NAND2xp5_ASAP7_75t_SL U59181 ( .A(n72620), .B(n72621), .Y(n72619) );
  INVxp67_ASAP7_75t_SL U59182 ( .A(n63977), .Y(n63979) );
  OAI21xp33_ASAP7_75t_SL U59183 ( .A1(n2637), .A2(
        or1200_cpu_or1200_except_n622), .B(n64000), .Y(n63995) );
  INVxp67_ASAP7_75t_SL U59184 ( .A(n70996), .Y(n70929) );
  NAND2xp5_ASAP7_75t_SL U59185 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[24]), .B(
        n73115), .Y(n73105) );
  NAND2xp5_ASAP7_75t_SL U59186 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[22]), .B(
        n73340), .Y(n73100) );
  INVx1_ASAP7_75t_SL U59187 ( .A(n58622), .Y(n59632) );
  INVx1_ASAP7_75t_SL U59188 ( .A(n58400), .Y(n57204) );
  AOI22xp33_ASAP7_75t_SL U59189 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[19]), .A2(
        n73304), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[18]), .B2(
        n73312), .Y(n73090) );
  INVx1_ASAP7_75t_SL U59190 ( .A(n58619), .Y(n57205) );
  NAND2xp5_ASAP7_75t_SL U59191 ( .A(n60701), .B(n60700), .Y(n60706) );
  OAI21xp33_ASAP7_75t_SL U59192 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[7]), .A2(
        n70205), .B(n70206), .Y(n70202) );
  INVx1_ASAP7_75t_SL U59193 ( .A(n59574), .Y(n75890) );
  NAND2xp5_ASAP7_75t_SL U59194 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[26]), .B(
        n73373), .Y(n73372) );
  NAND2xp33_ASAP7_75t_SL U59195 ( .A(n73623), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .Y(
        n73698) );
  INVxp67_ASAP7_75t_SL U59196 ( .A(n71883), .Y(n71885) );
  NAND2xp5_ASAP7_75t_SL U59197 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[25]), .B(
        n73381), .Y(n73383) );
  INVxp67_ASAP7_75t_SL U59198 ( .A(n59258), .Y(n59255) );
  INVxp67_ASAP7_75t_SL U59199 ( .A(n65396), .Y(n65365) );
  NAND2xp5_ASAP7_75t_SL U59200 ( .A(n73619), .B(n73618), .Y(n73689) );
  AOI21xp5_ASAP7_75t_SL U59201 ( .A1(n60225), .A2(supv), .B(n59921), .Y(n59925) );
  NAND2xp33_ASAP7_75t_SL U59202 ( .A(n2596), .B(n2609), .Y(n61031) );
  INVx1_ASAP7_75t_SL U59203 ( .A(n2037), .Y(n61314) );
  NAND2xp5_ASAP7_75t_SL U59204 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .B(
        n71873), .Y(n72085) );
  INVxp67_ASAP7_75t_SL U59205 ( .A(n2609), .Y(n61154) );
  NAND2xp5_ASAP7_75t_SL U59206 ( .A(n78439), .B(n60225), .Y(n60226) );
  NAND2xp33_ASAP7_75t_SL U59207 ( .A(n2589), .B(n61028), .Y(n60338) );
  NAND2xp5_ASAP7_75t_SL U59208 ( .A(n60994), .B(n60993), .Y(n61000) );
  NAND2xp5_ASAP7_75t_SL U59209 ( .A(or1200_cpu_or1200_mult_mac_n311), .B(
        n63452), .Y(n63506) );
  NAND2xp5_ASAP7_75t_SL U59210 ( .A(or1200_cpu_or1200_mult_mac_n165), .B(
        n63451), .Y(n63520) );
  NAND2xp5_ASAP7_75t_SL U59211 ( .A(n69543), .B(n69540), .Y(n69527) );
  NAND2xp5_ASAP7_75t_SL U59212 ( .A(or1200_cpu_or1200_mult_mac_n313), .B(
        n63489), .Y(n63505) );
  NAND2xp5_ASAP7_75t_SL U59213 ( .A(or1200_cpu_or1200_mult_mac_n167), .B(
        n63490), .Y(n63502) );
  OAI21xp5_ASAP7_75t_SL U59214 ( .A1(n63490), .A2(n63489), .B(n63488), .Y(
        n63540) );
  NAND2xp5_ASAP7_75t_SL U59215 ( .A(or1200_cpu_or1200_mult_mac_n169), .B(
        n63483), .Y(n63503) );
  NAND2xp5_ASAP7_75t_SL U59216 ( .A(or1200_cpu_or1200_mult_mac_n315), .B(
        n63485), .Y(n63504) );
  NOR2xp33_ASAP7_75t_SRAM U59217 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .B(n65249), .Y(
        n65247) );
  NAND2xp5_ASAP7_75t_SL U59218 ( .A(n70622), .B(n70621), .Y(n70627) );
  NOR2xp33_ASAP7_75t_SRAM U59219 ( .A(n59562), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .Y(n65563) );
  NAND2xp5_ASAP7_75t_SL U59220 ( .A(n69390), .B(n69392), .Y(n69428) );
  NAND2xp5_ASAP7_75t_SL U59221 ( .A(n69393), .B(n69388), .Y(n69438) );
  NAND2xp5_ASAP7_75t_SL U59222 ( .A(n69386), .B(n69400), .Y(n69437) );
  NAND2xp5_ASAP7_75t_SL U59223 ( .A(n70620), .B(n70619), .Y(n70628) );
  INVx1_ASAP7_75t_SL U59224 ( .A(n73008), .Y(n73026) );
  NAND2xp5_ASAP7_75t_SL U59225 ( .A(n65238), .B(n65396), .Y(n65332) );
  NAND2xp5_ASAP7_75t_SL U59226 ( .A(or1200_cpu_or1200_mult_mac_n319), .B(
        n63536), .Y(n63775) );
  NAND2xp5_ASAP7_75t_SL U59227 ( .A(or1200_cpu_or1200_mult_mac_n173), .B(
        n63537), .Y(n63778) );
  INVxp67_ASAP7_75t_SL U59228 ( .A(n59549), .Y(n57561) );
  INVxp33_ASAP7_75t_SL U59229 ( .A(n69540), .Y(n69542) );
  INVxp33_ASAP7_75t_SL U59230 ( .A(n69545), .Y(n69546) );
  NAND2xp5_ASAP7_75t_SL U59231 ( .A(or1200_cpu_or1200_mult_mac_n321), .B(
        n75367), .Y(n63774) );
  NAND2xp5_ASAP7_75t_SL U59232 ( .A(n70637), .B(n70636), .Y(n70639) );
  INVx1_ASAP7_75t_SL U59233 ( .A(n65258), .Y(n65260) );
  NAND2xp5_ASAP7_75t_SL U59234 ( .A(or1200_cpu_or1200_mult_mac_n175), .B(
        n75341), .Y(n63777) );
  OAI21xp33_ASAP7_75t_SL U59235 ( .A1(n63537), .A2(n63536), .B(n63535), .Y(
        n63538) );
  OAI21xp5_ASAP7_75t_SL U59236 ( .A1(n70635), .A2(n70634), .B(n70633), .Y(
        n70640) );
  INVxp67_ASAP7_75t_SL U59237 ( .A(n63534), .Y(n63541) );
  INVx1_ASAP7_75t_SL U59238 ( .A(n74741), .Y(n74538) );
  AND3x1_ASAP7_75t_SL U59239 ( .A(n59993), .B(n2598), .C(n2691), .Y(n59994) );
  INVx2_ASAP7_75t_SL U59240 ( .A(n58808), .Y(n57206) );
  NAND2xp33_ASAP7_75t_SL U59241 ( .A(n59702), .B(n59995), .Y(n75143) );
  NAND2xp5_ASAP7_75t_SL U59242 ( .A(n74533), .B(n74532), .Y(n74549) );
  NAND2xp33_ASAP7_75t_SL U59243 ( .A(n2596), .B(n2616), .Y(n59958) );
  INVxp67_ASAP7_75t_SL U59244 ( .A(n63887), .Y(n63890) );
  INVx1_ASAP7_75t_SL U59245 ( .A(n2589), .Y(n62024) );
  INVxp33_ASAP7_75t_SL U59246 ( .A(n69395), .Y(n69396) );
  NAND2xp5_ASAP7_75t_SL U59247 ( .A(or1200_cpu_or1200_mult_mac_n325), .B(
        n74584), .Y(n65092) );
  INVx1_ASAP7_75t_SL U59248 ( .A(n72534), .Y(n72434) );
  NAND2xp5_ASAP7_75t_SL U59249 ( .A(or1200_cpu_or1200_mult_mac_n383), .B(
        n69163), .Y(n69189) );
  INVxp67_ASAP7_75t_SL U59250 ( .A(n64000), .Y(n64002) );
  AND3x1_ASAP7_75t_SL U59251 ( .A(ic_en), .B(n2779), .C(n2777), .Y(n77312) );
  INVx1_ASAP7_75t_SL U59252 ( .A(n63399), .Y(n63319) );
  INVx1_ASAP7_75t_SL U59253 ( .A(n64265), .Y(n75416) );
  NAND2xp5_ASAP7_75t_SL U59254 ( .A(n2814), .B(n61028), .Y(n77426) );
  OAI21xp33_ASAP7_75t_SL U59255 ( .A1(n2678), .A2(
        or1200_cpu_or1200_except_n640), .B(n65201), .Y(n75414) );
  NAND2xp33_ASAP7_75t_SL U59256 ( .A(n59702), .B(n59974), .Y(n75632) );
  NAND2xp5_ASAP7_75t_SL U59257 ( .A(or1200_cpu_or1200_mult_mac_n147), .B(
        n63300), .Y(n63324) );
  NAND2xp5_ASAP7_75t_SL U59258 ( .A(n59562), .B(n74050), .Y(n65646) );
  NAND2xp33_ASAP7_75t_SL U59259 ( .A(n75540), .B(n65201), .Y(n65202) );
  INVxp67_ASAP7_75t_SL U59260 ( .A(n75543), .Y(n65205) );
  NAND2xp5_ASAP7_75t_SL U59261 ( .A(n62221), .B(n62220), .Y(n62219) );
  INVxp33_ASAP7_75t_SL U59262 ( .A(n60854), .Y(n61699) );
  NAND2xp33_ASAP7_75t_SL U59263 ( .A(n59702), .B(n60172), .Y(n65213) );
  INVx2_ASAP7_75t_SL U59264 ( .A(n58608), .Y(n57207) );
  INVx1_ASAP7_75t_SL U59265 ( .A(n77309), .Y(n77310) );
  INVxp67_ASAP7_75t_SL U59266 ( .A(n63372), .Y(n63341) );
  OAI21xp33_ASAP7_75t_SL U59267 ( .A1(or1200_cpu_or1200_except_n661), .A2(
        or1200_cpu_or1200_except_n664), .B(n2037), .Y(n77386) );
  NAND2xp5_ASAP7_75t_SL U59268 ( .A(n63340), .B(n63339), .Y(n63379) );
  INVx1_ASAP7_75t_SL U59269 ( .A(n72495), .Y(n72510) );
  OAI22xp33_ASAP7_75t_SL U59270 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[14]), .A2(
        n73140), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[13]), .B2(
        n73071), .Y(n73072) );
  INVx1_ASAP7_75t_SL U59271 ( .A(n63426), .Y(n63404) );
  OAI21xp33_ASAP7_75t_SL U59272 ( .A1(n76754), .A2(n76722), .B(n63376), .Y(
        n63377) );
  AOI22xp33_ASAP7_75t_SL U59273 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[13]), .A2(
        n73071), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[12]), .B2(
        n73064), .Y(n73065) );
  NAND2xp5_ASAP7_75t_SL U59274 ( .A(n69547), .B(n69541), .Y(n74495) );
  INVxp33_ASAP7_75t_SL U59275 ( .A(n66180), .Y(n65524) );
  NAND2xp5_ASAP7_75t_SL U59276 ( .A(or1200_cpu_or1200_mult_mac_n161), .B(
        n63422), .Y(n63525) );
  NAND2xp5_ASAP7_75t_SL U59277 ( .A(n78364), .B(n69545), .Y(n74496) );
  NAND2xp5_ASAP7_75t_SL U59278 ( .A(n69533), .B(n69538), .Y(n69526) );
  INVxp67_ASAP7_75t_SL U59279 ( .A(n63457), .Y(n63434) );
  INVxp67_ASAP7_75t_SL U59280 ( .A(n63522), .Y(n63437) );
  NAND2xp5_ASAP7_75t_SL U59281 ( .A(or1200_cpu_or1200_except_delayed_iee[1]), 
        .B(n78253), .Y(or1200_cpu_or1200_except_n1696) );
  NAND2xp5_ASAP7_75t_SL U59282 ( .A(n2761), .B(n59947), .Y(n59948) );
  INVxp67_ASAP7_75t_SL U59283 ( .A(n69108), .Y(n69091) );
  NAND2xp5_ASAP7_75t_SL U59284 ( .A(n1915), .B(n59573), .Y(n59867) );
  NAND2xp33_ASAP7_75t_SL U59285 ( .A(n73042), .B(n72994), .Y(n72848) );
  OAI21xp33_ASAP7_75t_SL U59286 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[4]), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .B(
        n73709), .Y(n73755) );
  NAND2xp5_ASAP7_75t_SL U59287 ( .A(or1200_cpu_or1200_mult_mac_n395), .B(
        n69256), .Y(n69253) );
  NAND2xp5_ASAP7_75t_SL U59288 ( .A(n3313), .B(n73728), .Y(n73501) );
  NAND2xp5_ASAP7_75t_SL U59289 ( .A(or1200_cpu_or1200_mult_mac_n229), .B(
        n69109), .Y(n69165) );
  INVx1_ASAP7_75t_SL U59290 ( .A(n74710), .Y(n74718) );
  NAND2xp5_ASAP7_75t_SL U59291 ( .A(or1200_cpu_or1200_mult_mac_n223), .B(
        n69022), .Y(n69060) );
  NOR2xp33_ASAP7_75t_SRAM U59292 ( .A(n69278), .B(n69277), .Y(n69280) );
  NOR2x1_ASAP7_75t_SL U59293 ( .A(n2450), .B(n69583), .Y(n70229) );
  NAND2xp5_ASAP7_75t_SL U59294 ( .A(or1200_cpu_or1200_mult_mac_n375), .B(
        n69110), .Y(n69169) );
  INVxp67_ASAP7_75t_SL U59295 ( .A(n75662), .Y(n75125) );
  NAND2xp5_ASAP7_75t_SL U59296 ( .A(n1879), .B(n59574), .Y(n59866) );
  NAND2xp5_ASAP7_75t_SL U59297 ( .A(or1200_cpu_or1200_mult_mac_n387), .B(
        n69188), .Y(n74569) );
  NAND2xp5_ASAP7_75t_SL U59298 ( .A(n77247), .B(n74933), .Y(n77435) );
  INVx1_ASAP7_75t_SL U59299 ( .A(n69282), .Y(n69275) );
  NAND2xp5_ASAP7_75t_SL U59300 ( .A(n3310), .B(n73690), .Y(n73486) );
  NAND2xp5_ASAP7_75t_SL U59301 ( .A(n75120), .B(n75119), .Y(n75124) );
  INVx1_ASAP7_75t_SL U59302 ( .A(n74686), .Y(n59633) );
  NAND2xp5_ASAP7_75t_SL U59303 ( .A(n2437), .B(n70546), .Y(n70253) );
  O2A1O1Ixp5_ASAP7_75t_SRAM U59304 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_), .A2(
        n74659), .B(n70456), .C(n74682), .Y(n70459) );
  NAND2xp5_ASAP7_75t_SL U59305 ( .A(or1200_cpu_or1200_mult_mac_n207), .B(
        n68847), .Y(n69048) );
  NOR3xp33_ASAP7_75t_SRAM U59306 ( .A(n76935), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_9_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_2_), .Y(n76936)
         );
  NAND2xp5_ASAP7_75t_SL U59307 ( .A(or1200_cpu_or1200_mult_mac_n371), .B(
        n69024), .Y(n69066) );
  NAND2xp5_ASAP7_75t_SL U59308 ( .A(or1200_cpu_or1200_mult_mac_n217), .B(
        n68938), .Y(n68986) );
  NAND2xp5_ASAP7_75t_SL U59309 ( .A(or1200_cpu_or1200_mult_mac_n377), .B(
        n69126), .Y(n69168) );
  AOI21xp33_ASAP7_75t_SL U59310 ( .A1(or1200_cpu_or1200_mult_mac_n259), .A2(
        or1200_cpu_or1200_mult_mac_n405), .B(n75121), .Y(n75122) );
  NAND2xp5_ASAP7_75t_SL U59311 ( .A(or1200_cpu_or1200_mult_mac_n359), .B(
        n68892), .Y(n68940) );
  NAND2xp5_ASAP7_75t_SL U59312 ( .A(or1200_cpu_or1200_mult_mac_n411), .B(
        n76894), .Y(n76904) );
  INVx1_ASAP7_75t_SL U59313 ( .A(n69273), .Y(n69259) );
  NAND2xp33_ASAP7_75t_SL U59314 ( .A(n69243), .B(n69242), .Y(n69257) );
  OAI21xp33_ASAP7_75t_SL U59315 ( .A1(n68933), .A2(n68932), .B(n68931), .Y(
        n68934) );
  INVxp67_ASAP7_75t_SL U59316 ( .A(n76911), .Y(n76901) );
  NAND2xp33_ASAP7_75t_SL U59317 ( .A(n3310), .B(n73667), .Y(n73520) );
  AOI21xp33_ASAP7_75t_SL U59318 ( .A1(or1200_cpu_or1200_mult_mac_n367), .A2(
        or1200_cpu_or1200_mult_mac_n221), .B(n68997), .Y(n68998) );
  AOI21xp33_ASAP7_75t_SL U59319 ( .A1(n73743), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[21]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[23]), .Y(n73517) );
  NAND2xp5_ASAP7_75t_SL U59320 ( .A(or1200_cpu_or1200_mult_mac_n361), .B(
        n68932), .Y(n68939) );
  NAND2xp5_ASAP7_75t_SL U59321 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B(
        n70466), .Y(n70535) );
  INVxp67_ASAP7_75t_SL U59322 ( .A(n71645), .Y(n71655) );
  NAND2xp5_ASAP7_75t_SL U59323 ( .A(n73492), .B(n73493), .Y(n73525) );
  NAND2xp5_ASAP7_75t_SL U59324 ( .A(or1200_cpu_or1200_mult_mac_n393), .B(
        n69220), .Y(n69248) );
  INVx1_ASAP7_75t_SL U59325 ( .A(n69278), .Y(n69212) );
  NAND2xp5_ASAP7_75t_SL U59326 ( .A(or1200_cpu_or1200_mult_mac_n221), .B(
        n68985), .Y(n69059) );
  NAND2xp5_ASAP7_75t_SL U59327 ( .A(or1200_cpu_or1200_mult_mac_n373), .B(
        n69084), .Y(n69171) );
  NAND2xp5_ASAP7_75t_SL U59328 ( .A(or1200_cpu_or1200_mult_mac_n247), .B(
        n69243), .Y(n69249) );
  NOR2xp33_ASAP7_75t_SRAM U59329 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_5_), .B(
        n71692), .Y(n71693) );
  NAND2xp5_ASAP7_75t_SL U59330 ( .A(or1200_cpu_or1200_mult_mac_n205), .B(
        n68830), .Y(n69049) );
  NOR2xp33_ASAP7_75t_SRAM U59331 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .B(n65327), .Y(
        n65325) );
  NAND2xp5_ASAP7_75t_SL U59332 ( .A(or1200_cpu_or1200_mult_mac_n379), .B(
        n69124), .Y(n69173) );
  INVx1_ASAP7_75t_SL U59333 ( .A(n60192), .Y(n60193) );
  INVx1_ASAP7_75t_SL U59334 ( .A(n73814), .Y(n73818) );
  NAND2xp5_ASAP7_75t_SL U59335 ( .A(or1200_cpu_or1200_mult_mac_n391), .B(
        n74114), .Y(n69247) );
  NAND2xp33_ASAP7_75t_SL U59336 ( .A(or1200_cpu_or1200_mult_mac_n365), .B(
        n76721), .Y(n68989) );
  INVx1_ASAP7_75t_SL U59337 ( .A(n73498), .Y(n73485) );
  NAND2xp33_ASAP7_75t_SL U59338 ( .A(or1200_cpu_or1200_mult_mac_n251), .B(
        n69270), .Y(n69321) );
  NAND2xp5_ASAP7_75t_SL U59339 ( .A(n2589), .B(n2609), .Y(n61140) );
  INVxp67_ASAP7_75t_SL U59340 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .Y(
        n70483) );
  NAND2xp5_ASAP7_75t_SL U59341 ( .A(or1200_cpu_or1200_mult_mac_n409), .B(
        n75654), .Y(n75655) );
  NAND2xp5_ASAP7_75t_SL U59342 ( .A(or1200_cpu_or1200_mult_mac_n349), .B(
        n68814), .Y(n69065) );
  NAND2xp33_ASAP7_75t_SL U59343 ( .A(n73690), .B(n59705), .Y(n73691) );
  NAND2xp33_ASAP7_75t_SL U59344 ( .A(n71667), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_6_), .Y(
        n71665) );
  NAND2xp33_ASAP7_75t_SL U59345 ( .A(or1200_cpu_or1200_mult_mac_n253), .B(
        n69309), .Y(n69322) );
  NAND2xp5_ASAP7_75t_SL U59346 ( .A(dbg_adr_i[15]), .B(n77847), .Y(n77639) );
  INVx1_ASAP7_75t_SL U59347 ( .A(n77847), .Y(n77672) );
  NAND2xp33_ASAP7_75t_SL U59348 ( .A(n62477), .B(dbg_dat_i[4]), .Y(n4071) );
  NAND2xp33_ASAP7_75t_SL U59349 ( .A(n62477), .B(dbg_dat_i[7]), .Y(n4058) );
  NAND2xp33_ASAP7_75t_SL U59350 ( .A(n62477), .B(dbg_dat_i[9]), .Y(n4050) );
  NAND2xp33_ASAP7_75t_SL U59351 ( .A(n62477), .B(dbg_dat_i[6]), .Y(n4062) );
  NAND2xp33_ASAP7_75t_SL U59352 ( .A(n62477), .B(dbg_dat_i[10]), .Y(n4046) );
  INVx1_ASAP7_75t_SL U59353 ( .A(or1200_cpu_or1200_mult_mac_mul_stall_count_1_), .Y(n62025) );
  INVxp67_ASAP7_75t_SL U59354 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_45_), .Y(n69686) );
  INVxp67_ASAP7_75t_SL U59355 ( .A(or1200_cpu_or1200_fpu_b_is_inf), .Y(n74814)
         );
  INVxp67_ASAP7_75t_SL U59356 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[19]), .Y(n69685) );
  INVx1_ASAP7_75t_SL U59357 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[7]), .Y(
        n27738) );
  INVx1_ASAP7_75t_SL U59358 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_7_), .Y(n78341) );
  NAND2xp5_ASAP7_75t_SL U59359 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_in_00), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2), .Y(n65530) );
  INVx1_ASAP7_75t_SL U59360 ( .A(n1135), .Y(n66227) );
  INVx1_ASAP7_75t_SL U59361 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[19]), .Y(n78356) );
  INVx1_ASAP7_75t_SL U59362 ( .A(n1153), .Y(n62492) );
  INVxp67_ASAP7_75t_SL U59363 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[20]), .Y(n70950) );
  INVx1_ASAP7_75t_SL U59364 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[8]), .Y(
        n70211) );
  INVx1_ASAP7_75t_SL U59365 ( .A(n1821), .Y(n76514) );
  INVx1_ASAP7_75t_SL U59366 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[6]), .Y(
        n27735) );
  INVxp67_ASAP7_75t_SL U59367 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_24_), .Y(n66209) );
  INVx1_ASAP7_75t_SL U59368 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[0]), .Y(n74749) );
  INVx1_ASAP7_75t_SL U59369 ( .A(n2804), .Y(n76689) );
  INVx1_ASAP7_75t_SL U59370 ( .A(n1147), .Y(n75390) );
  INVx1_ASAP7_75t_SL U59371 ( .A(or1200_cpu_or1200_mult_mac_n375), .Y(n69109)
         );
  INVxp33_ASAP7_75t_SL U59372 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_2_), .Y(n66185) );
  INVxp67_ASAP7_75t_SL U59373 ( .A(n2703), .Y(n77404) );
  INVx1_ASAP7_75t_SL U59374 ( .A(or1200_cpu_or1200_except_n419), .Y(n76249) );
  INVx1_ASAP7_75t_SL U59375 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_8_), .Y(n78343) );
  INVxp67_ASAP7_75t_SL U59376 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[6]), .Y(
        n70609) );
  INVx1_ASAP7_75t_SL U59377 ( .A(n1131), .Y(n66232) );
  INVxp33_ASAP7_75t_SL U59378 ( .A(or1200_cpu_or1200_mult_mac_n381), .Y(n69174) );
  INVx1_ASAP7_75t_SL U59379 ( .A(or1200_cpu_or1200_rf_addra_last_0_), .Y(
        n77958) );
  INVxp33_ASAP7_75t_SL U59380 ( .A(n1155), .Y(n62485) );
  INVxp67_ASAP7_75t_SL U59381 ( .A(n2713), .Y(n60417) );
  INVxp67_ASAP7_75t_SL U59382 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_41_), .Y(n69647) );
  INVx1_ASAP7_75t_SL U59383 ( .A(or1200_cpu_or1200_except_n416), .Y(n76643) );
  NAND2xp33_ASAP7_75t_SL U59384 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[2]), .Y(n65489) );
  INVx1_ASAP7_75t_SL U59385 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[9]), .Y(
        n70213) );
  INVx1_ASAP7_75t_SL U59386 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), .Y(
        n72993) );
  INVx1_ASAP7_75t_SL U59387 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]), .Y(n74750) );
  INVx1_ASAP7_75t_SL U59388 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[6]), .Y(n74169) );
  INVx1_ASAP7_75t_SL U59389 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[16]), .Y(n70881) );
  NAND2xp5_ASAP7_75t_SL U59390 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), .Y(
        n73008) );
  INVx1_ASAP7_75t_SL U59391 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[3]), .Y(n78332)
         );
  INVx1_ASAP7_75t_SL U59392 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[21]), .Y(n70983) );
  INVxp67_ASAP7_75t_SL U59393 ( .A(or1200_cpu_or1200_except_n200), .Y(n61165)
         );
  INVxp67_ASAP7_75t_SL U59394 ( .A(n986), .Y(iwb_adr_o[27]) );
  INVx1_ASAP7_75t_SL U59395 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_0_), .Y(n74835)
         );
  INVx1_ASAP7_75t_SL U59396 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_6_), .Y(
        n74368) );
  INVxp33_ASAP7_75t_SL U59397 ( .A(or1200_cpu_or1200_except_n563), .Y(n63707)
         );
  INVxp67_ASAP7_75t_SL U59398 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[5]), .Y(n65784) );
  INVxp33_ASAP7_75t_SL U59399 ( .A(n748), .Y(n76734) );
  INVxp67_ASAP7_75t_SL U59400 ( .A(n2575), .Y(n77930) );
  INVx1_ASAP7_75t_SL U59401 ( .A(n2596), .Y(n61145) );
  INVx1_ASAP7_75t_SL U59402 ( .A(n2733), .Y(n77375) );
  INVx1_ASAP7_75t_SL U59403 ( .A(n2711), .Y(n60412) );
  INVx1_ASAP7_75t_SL U59404 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[5]), .Y(
        n27733) );
  INVx1_ASAP7_75t_SL U59405 ( .A(or1200_cpu_or1200_mult_mac_n363), .Y(n68938)
         );
  INVxp33_ASAP7_75t_SL U59406 ( .A(n1151), .Y(n62493) );
  INVxp67_ASAP7_75t_SL U59407 ( .A(n2854), .Y(n65274) );
  INVx1_ASAP7_75t_SL U59408 ( .A(or1200_cpu_or1200_except_n270), .Y(n76708) );
  INVxp67_ASAP7_75t_SL U59409 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[15]), .Y(n69646) );
  INVxp67_ASAP7_75t_SL U59410 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_), .Y(n78362) );
  INVx1_ASAP7_75t_SL U59411 ( .A(n1674), .Y(n75376) );
  INVx1_ASAP7_75t_SL U59412 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[2]), .Y(
        n70223) );
  INVx1_ASAP7_75t_SL U59413 ( .A(or1200_cpu_or1200_rf_addra_last_4_), .Y(
        n77934) );
  INVxp67_ASAP7_75t_SL U59414 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_in_00), .Y(n65488) );
  INVx1_ASAP7_75t_SL U59415 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[9]), .Y(n65822) );
  INVx1_ASAP7_75t_SL U59416 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_10_), .Y(n78349) );
  INVxp67_ASAP7_75t_SL U59417 ( .A(n2721), .Y(n60511) );
  INVx1_ASAP7_75t_SL U59418 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[4]), .Y(
        n70218) );
  INVx1_ASAP7_75t_SL U59419 ( .A(or1200_cpu_or1200_rf_addra_last_2_), .Y(
        n77944) );
  INVx1_ASAP7_75t_SL U59420 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[15]), .Y(n70863) );
  INVxp67_ASAP7_75t_SL U59421 ( .A(or1200_cpu_or1200_except_n565), .Y(n63723)
         );
  INVx1_ASAP7_75t_SL U59422 ( .A(or1200_cpu_or1200_mult_mac_n177), .Y(n63892)
         );
  INVx1_ASAP7_75t_SL U59423 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[18]), .Y(n70910) );
  AND3x1_ASAP7_75t_SL U59424 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_3_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_5_), .Y(
        n70554) );
  INVx1_ASAP7_75t_SL U59425 ( .A(n2709), .Y(n60482) );
  INVx1_ASAP7_75t_SL U59426 ( .A(n3138), .Y(n78162) );
  INVx1_ASAP7_75t_SL U59427 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[10]), .Y(n70786) );
  INVxp67_ASAP7_75t_SL U59428 ( .A(n2542), .Y(n77526) );
  INVxp67_ASAP7_75t_SL U59429 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[30]), .Y(n78191) );
  INVx1_ASAP7_75t_SL U59430 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_3_), .Y(n66179) );
  INVx1_ASAP7_75t_SL U59431 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[3]), .Y(n70709) );
  INVxp67_ASAP7_75t_SL U59432 ( .A(or1200_cpu_or1200_except_n583), .Y(n76565)
         );
  INVx1_ASAP7_75t_SL U59433 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[22]), .Y(n70994) );
  NAND2xp33_ASAP7_75t_SL U59434 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_1_), .B(n2491), .Y(
        n74157) );
  INVx1_ASAP7_75t_SL U59435 ( .A(or1200_cpu_or1200_rf_addra_last_3_), .Y(
        n77940) );
  NAND2xp5_ASAP7_75t_SL U59436 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[4]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[3]), .Y(
        n70588) );
  INVx1_ASAP7_75t_SL U59437 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_4_), .Y(n74142) );
  INVx1_ASAP7_75t_SL U59438 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_state), .Y(n59698) );
  INVx1_ASAP7_75t_SL U59439 ( .A(or1200_cpu_or1200_except_n520), .Y(n76232) );
  INVxp33_ASAP7_75t_SL U59440 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[3]), .Y(
        n70583) );
  INVx1_ASAP7_75t_SL U59441 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[0]), .Y(
        n70228) );
  INVxp67_ASAP7_75t_SL U59442 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[23]), .Y(n70995) );
  INVxp67_ASAP7_75t_SL U59443 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[18]), .Y(
        n73308) );
  INVxp67_ASAP7_75t_SL U59444 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2), .Y(n66197) );
  INVx1_ASAP7_75t_SL U59445 ( .A(n2723), .Y(n78010) );
  INVx1_ASAP7_75t_SL U59446 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_5_), .Y(n74147) );
  INVx1_ASAP7_75t_SL U59447 ( .A(or1200_cpu_or1200_rf_addra_last_1_), .Y(
        n77949) );
  INVx1_ASAP7_75t_SL U59448 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_2_), .Y(
        n70566) );
  INVx1_ASAP7_75t_SL U59449 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[11]), .Y(n70809) );
  INVx1_ASAP7_75t_SL U59450 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[7]), .Y(
        n70613) );
  INVx1_ASAP7_75t_SL U59451 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[19]), .Y(
        n73304) );
  INVxp67_ASAP7_75t_SL U59452 ( .A(or1200_cpu_or1200_mult_mac_n349), .Y(n75508) );
  INVx1_ASAP7_75t_SL U59453 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[18]), .Y(n69937) );
  INVx1_ASAP7_75t_SL U59454 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[6]), .Y(
        n70215) );
  INVx1_ASAP7_75t_SL U59455 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[9]), .Y(
        n73159) );
  INVx1_ASAP7_75t_SL U59456 ( .A(or1200_cpu_or1200_mult_mac_n229), .Y(n69110)
         );
  INVx1_ASAP7_75t_SL U59457 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[18]), .Y(
        n73312) );
  INVx1_ASAP7_75t_SL U59458 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[14]), .Y(n70850) );
  INVxp67_ASAP7_75t_SL U59459 ( .A(n995), .Y(iwb_adr_o[28]) );
  NAND2xp33_ASAP7_75t_SL U59460 ( .A(or1200_cpu_or1200_mult_mac_n235), .B(
        or1200_cpu_or1200_mult_mac_n381), .Y(n69209) );
  INVx1_ASAP7_75t_SL U59461 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[5]), .Y(n70722) );
  NAND2xp5_ASAP7_75t_SL U59462 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[1]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[2]), .Y(
        n70579) );
  INVxp67_ASAP7_75t_SL U59463 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[5]), .Y(
        n73222) );
  INVx1_ASAP7_75t_SL U59464 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[14]), .Y(
        n73141) );
  INVxp67_ASAP7_75t_SL U59465 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[15]), .Y(
        n73144) );
  INVx1_ASAP7_75t_SL U59466 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[8]), .Y(n70767) );
  INVx1_ASAP7_75t_SL U59467 ( .A(or1200_cpu_or1200_except_n401), .Y(n76858) );
  INVx1_ASAP7_75t_SL U59468 ( .A(or1200_cpu_or1200_except_n494), .Y(n76857) );
  INVx1_ASAP7_75t_SL U59469 ( .A(or1200_cpu_or1200_except_n410), .Y(n76617) );
  INVxp67_ASAP7_75t_SL U59470 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[26]), .Y(n28180)
         );
  INVxp67_ASAP7_75t_SL U59471 ( .A(n3134), .Y(n77421) );
  INVx1_ASAP7_75t_SL U59472 ( .A(or1200_cpu_or1200_mult_mac_n237), .Y(n69163)
         );
  INVx1_ASAP7_75t_SL U59473 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_), .Y(n78434) );
  INVx1_ASAP7_75t_SL U59474 ( .A(n2707), .Y(n60473) );
  INVx1_ASAP7_75t_SL U59475 ( .A(n2727), .Y(n78016) );
  INVxp67_ASAP7_75t_SL U59476 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[19]), .Y(n28173)
         );
  INVxp67_ASAP7_75t_SL U59477 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_43_), .Y(n69672) );
  INVx1_ASAP7_75t_SL U59478 ( .A(DP_OP_741J1_129_6992_n46), .Y(n70311) );
  INVxp67_ASAP7_75t_SL U59479 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_21_), .Y(n69693) );
  INVx1_ASAP7_75t_SL U59480 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]), .Y(n74751) );
  INVx1_ASAP7_75t_SL U59481 ( .A(or1200_cpu_or1200_except_n274), .Y(n76217) );
  INVxp67_ASAP7_75t_SL U59482 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[12]), .Y(n28166)
         );
  AND3x1_ASAP7_75t_SL U59483 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_24_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_0_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]), .Y(n66168) );
  INVx1_ASAP7_75t_SL U59484 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_20_), .Y(
        n74422) );
  INVxp67_ASAP7_75t_SL U59485 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[3]), .Y(n28201) );
  INVxp67_ASAP7_75t_SL U59486 ( .A(n2717), .Y(n60518) );
  NAND2xp33_ASAP7_75t_SL U59487 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_expa_ff), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_r_a), .Y(n4743) );
  INVx1_ASAP7_75t_SL U59488 ( .A(n3132), .Y(n61125) );
  INVxp67_ASAP7_75t_SL U59489 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[8]), .Y(
        n73194) );
  INVxp67_ASAP7_75t_SL U59490 ( .A(n1141), .Y(n64181) );
  INVxp67_ASAP7_75t_SL U59491 ( .A(or1200_cpu_or1200_mult_mac_n159), .Y(n63410) );
  INVxp33_ASAP7_75t_SL U59492 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_0_), .Y(n27421) );
  INVx1_ASAP7_75t_SL U59493 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[13]), .Y(n70843) );
  INVx1_ASAP7_75t_SL U59494 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_7_), .Y(n74173) );
  INVx1_ASAP7_75t_SL U59495 ( .A(n2729), .Y(n78019) );
  INVx1_ASAP7_75t_SL U59496 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_0_), .Y(n78429) );
  INVxp33_ASAP7_75t_SL U59497 ( .A(or1200_cpu_or1200_mult_mac_n223), .Y(n69023) );
  INVxp67_ASAP7_75t_SL U59498 ( .A(n2524), .Y(n77568) );
  INVx1_ASAP7_75t_SL U59499 ( .A(or1200_cpu_or1200_except_n498), .Y(n77277) );
  INVxp67_ASAP7_75t_SL U59500 ( .A(or1200_cpu_or1200_except_n252), .Y(n76236)
         );
  INVx1_ASAP7_75t_SL U59501 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .Y(
        n72999) );
  INVx1_ASAP7_75t_SL U59502 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_22_), .Y(
        n74442) );
  INVx1_ASAP7_75t_SL U59503 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[6]), .Y(n70735) );
  INVx1_ASAP7_75t_SL U59504 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[7]), .Y(n70759) );
  INVx1_ASAP7_75t_SL U59505 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[17]), .Y(n69919) );
  INVx1_ASAP7_75t_SL U59506 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[0]), .Y(n27066) );
  INVx1_ASAP7_75t_SL U59507 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .Y(
        n73042) );
  NAND2xp5_ASAP7_75t_SL U59508 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_2_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_3_), .Y(n66206) );
  INVx1_ASAP7_75t_SL U59509 ( .A(n1844), .Y(n76220) );
  INVx1_ASAP7_75t_SL U59510 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[1]), .Y(n27067) );
  INVx1_ASAP7_75t_SL U59511 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[9]), .Y(n27075) );
  INVxp67_ASAP7_75t_SL U59512 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_46_), .Y(n69694) );
  NAND2xp5_ASAP7_75t_SL U59513 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_1_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_0_), .Y(n74087) );
  INVx1_ASAP7_75t_SL U59514 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_24_), .Y(
        n74448) );
  INVx1_ASAP7_75t_SL U59515 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[2]), .Y(n27068) );
  INVx1_ASAP7_75t_SL U59516 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[3]), .Y(n27069) );
  INVx1_ASAP7_75t_SL U59517 ( .A(or1200_cpu_or1200_except_n496), .Y(n76999) );
  INVx1_ASAP7_75t_SL U59518 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[20]), .Y(n69990) );
  INVx1_ASAP7_75t_SL U59519 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[22]), .Y(
        n73340) );
  INVx1_ASAP7_75t_SL U59520 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[8]), .Y(n27074) );
  INVx1_ASAP7_75t_SL U59521 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[4]), .Y(n27070) );
  NAND2xp5_ASAP7_75t_SL U59522 ( .A(or1200_cpu_or1200_mult_mac_n241), .B(
        or1200_cpu_or1200_mult_mac_n387), .Y(n74571) );
  INVx1_ASAP7_75t_SL U59523 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[5]), .Y(n27071) );
  INVx1_ASAP7_75t_SL U59524 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_12_), .Y(n78351) );
  INVx1_ASAP7_75t_SL U59525 ( .A(or1200_cpu_or1200_except_n404), .Y(n76997) );
  INVx1_ASAP7_75t_SL U59526 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[6]), .Y(n27072) );
  INVxp67_ASAP7_75t_SL U59527 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[17]), .Y(
        n73076) );
  INVx1_ASAP7_75t_SL U59528 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_exp[7]), .Y(n27073) );
  INVxp67_ASAP7_75t_SL U59529 ( .A(DP_OP_742J1_130_9702_n59), .Y(n70570) );
  INVx1_ASAP7_75t_SL U59530 ( .A(or1200_cpu_or1200_mult_mac_n227), .Y(n69084)
         );
  INVxp33_ASAP7_75t_SL U59531 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_16_), .Y(n69671) );
  INVxp67_ASAP7_75t_SL U59532 ( .A(n1815), .Y(n61327) );
  INVxp67_ASAP7_75t_SL U59533 ( .A(n2052), .Y(n74024) );
  INVx1_ASAP7_75t_SL U59534 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_21_), .Y(n76945)
         );
  INVx1_ASAP7_75t_SL U59535 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[20]), .Y(
        n73123) );
  NAND2xp5_ASAP7_75t_SL U59536 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[6]), .Y(n65496) );
  INVxp33_ASAP7_75t_SL U59537 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_26_), 
        .Y(n74508) );
  INVx1_ASAP7_75t_SL U59538 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_22_), .Y(n78365) );
  INVxp67_ASAP7_75t_SL U59539 ( .A(or1200_cpu_or1200_except_n186), .Y(n77236)
         );
  INVx1_ASAP7_75t_SL U59540 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_8_), .Y(
        n74354) );
  INVx1_ASAP7_75t_SL U59541 ( .A(or1200_cpu_or1200_mult_mac_n239), .Y(n75363)
         );
  INVxp33_ASAP7_75t_SL U59542 ( .A(n2693), .Y(n61041) );
  INVxp67_ASAP7_75t_SL U59543 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[3]), .Y(n74138) );
  INVx1_ASAP7_75t_SL U59544 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[0]), .Y(n27027) );
  INVxp67_ASAP7_75t_SL U59545 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_44_), .Y(n69680) );
  NAND2xp5_ASAP7_75t_SL U59546 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_16_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_17_), .Y(n76947)
         );
  INVx1_ASAP7_75t_SL U59547 ( .A(or1200_cpu_or1200_except_n407), .Y(n76210) );
  INVx1_ASAP7_75t_SL U59548 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_13_), .Y(n78352) );
  INVx1_ASAP7_75t_SL U59549 ( .A(or1200_cpu_or1200_except_n502), .Y(n76704) );
  INVx1_ASAP7_75t_SL U59550 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[4]), .Y(n70717) );
  INVx1_ASAP7_75t_SL U59551 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_10_), .Y(
        n74318) );
  INVxp67_ASAP7_75t_SL U59552 ( .A(n1658), .Y(n63601) );
  INVx1_ASAP7_75t_SL U59553 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[12]), .Y(n70823) );
  INVxp33_ASAP7_75t_SL U59554 ( .A(or1200_cpu_or1200_fpu_snan_conv), .Y(n74803) );
  INVx1_ASAP7_75t_SL U59555 ( .A(n2731), .Y(n78025) );
  INVx1_ASAP7_75t_SL U59556 ( .A(or1200_cpu_or1200_except_n592), .Y(n77275) );
  INVxp67_ASAP7_75t_SL U59557 ( .A(n2705), .Y(n60328) );
  INVx1_ASAP7_75t_SL U59558 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_15_), .Y(n76941)
         );
  INVx1_ASAP7_75t_SL U59559 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_11_), .Y(n78347) );
  INVx1_ASAP7_75t_SL U59560 ( .A(n2191), .Y(n60995) );
  INVx1_ASAP7_75t_SL U59561 ( .A(or1200_cpu_or1200_except_n413), .Y(n76700) );
  INVxp67_ASAP7_75t_SL U59562 ( .A(or1200_cpu_or1200_if_insn_saved[22]), .Y(
        n60402) );
  NAND2xp5_ASAP7_75t_SL U59563 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_11_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_12_), .Y(n66205)
         );
  INVx1_ASAP7_75t_SL U59564 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_12_), .Y(
        n74336) );
  INVx1_ASAP7_75t_SL U59565 ( .A(n2725), .Y(n78013) );
  INVxp67_ASAP7_75t_SL U59566 ( .A(n2715), .Y(n60526) );
  INVx1_ASAP7_75t_SL U59567 ( .A(n1127), .Y(n75026) );
  NOR4xp25_ASAP7_75t_SRAM U59568 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_3_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_5_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_10_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_18_), .Y(n76940)
         );
  INVxp67_ASAP7_75t_SL U59569 ( .A(or1200_cpu_or1200_except_n184), .Y(n77168)
         );
  INVxp33_ASAP7_75t_SL U59570 ( .A(or1200_cpu_or1200_mult_mac_n389), .Y(n69201) );
  NAND2xp33_ASAP7_75t_SL U59571 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .Y(
        n72996) );
  INVx1_ASAP7_75t_SL U59572 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[7]), .Y(
        n73193) );
  NAND2xp5_ASAP7_75t_SL U59573 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_10_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_7_), .Y(n66204)
         );
  INVx1_ASAP7_75t_SL U59574 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_14_), .Y(
        n74383) );
  INVxp67_ASAP7_75t_SL U59575 ( .A(n2719), .Y(n60531) );
  INVx1_ASAP7_75t_SL U59576 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[9]), .Y(n70776) );
  INVx1_ASAP7_75t_SL U59577 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[24]), .Y(
        n73115) );
  INVxp67_ASAP7_75t_SL U59578 ( .A(n968), .Y(iwb_adr_o[25]) );
  INVxp67_ASAP7_75t_SL U59579 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[16]), .Y(n69666) );
  NAND2xp5_ASAP7_75t_SL U59580 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_4_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_5_), .Y(n66203)
         );
  INVx1_ASAP7_75t_SL U59581 ( .A(n1139), .Y(n75398) );
  INVx1_ASAP7_75t_SL U59582 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_16_), .Y(
        n74399) );
  INVxp67_ASAP7_75t_SL U59583 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[19]), .Y(n70911) );
  INVx1_ASAP7_75t_SL U59584 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[17]), .Y(n70893) );
  INVx1_ASAP7_75t_SL U59585 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[23]), .Y(
        n73333) );
  NAND2xp5_ASAP7_75t_SL U59586 ( .A(n1934), .B(n1774), .Y(n58632) );
  INVxp67_ASAP7_75t_SL U59587 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_42_), .Y(n69667) );
  INVxp67_ASAP7_75t_SL U59588 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[45]), .Y(n28197)
         );
  INVx1_ASAP7_75t_SL U59589 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_18_), .Y(
        n74307) );
  INVxp67_ASAP7_75t_SL U59590 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[43]), .Y(n28205)
         );
  INVx1_ASAP7_75t_SL U59591 ( .A(or1200_cpu_or1200_except_n398), .Y(n76680) );
  INVxp67_ASAP7_75t_SL U59592 ( .A(n1149), .Y(n74974) );
  INVxp33_ASAP7_75t_SL U59593 ( .A(or1200_cpu_or1200_mult_mac_n361), .Y(n68933) );
  INVxp67_ASAP7_75t_SL U59594 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[41]), .Y(n28194)
         );
  INVx1_ASAP7_75t_SL U59595 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[13]), .Y(
        n73185) );
  INVxp33_ASAP7_75t_SL U59596 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[13]), .Y(
        n73071) );
  INVxp67_ASAP7_75t_SL U59597 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[42]), .Y(n28195)
         );
  INVxp67_ASAP7_75t_SL U59598 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[44]), .Y(n28196)
         );
  INVxp67_ASAP7_75t_SL U59599 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[12]), .Y(n65792) );
  INVx1_ASAP7_75t_SL U59600 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_), .Y(
        n73040) );
  INVxp67_ASAP7_75t_SL U59601 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_37_), .Y(n78392) );
  INVxp67_ASAP7_75t_SL U59602 ( .A(n1247), .Y(dwb_adr_o[19]) );
  INVx1_ASAP7_75t_SL U59603 ( .A(or1200_cpu_or1200_except_n482), .Y(n75674) );
  INVxp67_ASAP7_75t_SL U59604 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[46]), .Y(n28206)
         );
  INVx1_ASAP7_75t_SL U59605 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_36_), .Y(n78393) );
  INVxp33_ASAP7_75t_SL U59606 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[10]), .Y(n65791) );
  INVx1_ASAP7_75t_SL U59607 ( .A(or1200_cpu_or1200_except_n467), .Y(n74083) );
  INVxp33_ASAP7_75t_SL U59608 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[11]), .Y(n65793) );
  INVx1_ASAP7_75t_SL U59609 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[10]), .Y(
        n73161) );
  INVx1_ASAP7_75t_SL U59610 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[1]), .Y(n27028) );
  INVx1_ASAP7_75t_SL U59611 ( .A(or1200_cpu_or1200_except_n550), .Y(n76928) );
  INVxp67_ASAP7_75t_SL U59612 ( .A(n2628), .Y(n77516) );
  INVx1_ASAP7_75t_SL U59613 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[2]), .Y(n27029) );
  INVx1_ASAP7_75t_SL U59614 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[3]), .Y(n27030) );
  INVxp33_ASAP7_75t_SL U59615 ( .A(n2664), .Y(n60516) );
  INVx1_ASAP7_75t_SL U59616 ( .A(or1200_cpu_or1200_except_n546), .Y(n75200) );
  INVx1_ASAP7_75t_SL U59617 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[4]), .Y(n27031) );
  INVxp67_ASAP7_75t_SL U59618 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_35_), .Y(n78394) );
  INVx1_ASAP7_75t_SL U59619 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[5]), .Y(n27032) );
  INVxp33_ASAP7_75t_SL U59620 ( .A(or1200_cpu_or1200_mult_mac_n191), .Y(n65165) );
  INVx1_ASAP7_75t_SL U59621 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[7]), .Y(n27034) );
  INVx1_ASAP7_75t_SL U59622 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[8]), .Y(n27035) );
  INVx1_ASAP7_75t_SL U59623 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_34_), .Y(n78225) );
  INVxp67_ASAP7_75t_SL U59624 ( .A(n1257), .Y(dwb_adr_o[17]) );
  INVx1_ASAP7_75t_SL U59625 ( .A(or1200_cpu_or1200_except_n540), .Y(n69373) );
  INVxp67_ASAP7_75t_SL U59626 ( .A(or1200_cpu_or1200_mult_mac_n397), .Y(n69270) );
  INVx1_ASAP7_75t_SL U59627 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[9]), .Y(n27036) );
  INVxp67_ASAP7_75t_SL U59628 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_33_), .Y(n78395) );
  INVx1_ASAP7_75t_SL U59629 ( .A(n1082), .Y(n78060) );
  INVx1_ASAP7_75t_SL U59630 ( .A(n1310), .Y(n77989) );
  INVx1_ASAP7_75t_SL U59631 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[4]), .Y(n65787) );
  INVx1_ASAP7_75t_SL U59632 ( .A(or1200_cpu_spr_dat_ppc[31]), .Y(n76922) );
  INVxp67_ASAP7_75t_SL U59633 ( .A(n1195), .Y(n78069) );
  INVx1_ASAP7_75t_SL U59634 ( .A(or1200_cpu_or1200_except_n536), .Y(n74047) );
  INVx1_ASAP7_75t_SL U59635 ( .A(or1200_cpu_or1200_except_n538), .Y(n74081) );
  INVxp33_ASAP7_75t_SL U59636 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[16]), .Y(n65783) );
  INVxp33_ASAP7_75t_SL U59637 ( .A(n799), .Y(n60125) );
  INVx1_ASAP7_75t_SL U59638 ( .A(n1305), .Y(n77963) );
  INVx1_ASAP7_75t_SL U59639 ( .A(or1200_cpu_or1200_except_delayed_tee[2]), .Y(
        n60233) );
  INVx1_ASAP7_75t_SL U59640 ( .A(n3012), .Y(n64013) );
  INVx1_ASAP7_75t_SL U59641 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[12]), .Y(
        n73180) );
  INVx1_ASAP7_75t_SL U59642 ( .A(or1200_cpu_or1200_except_n282), .Y(n62156) );
  INVx1_ASAP7_75t_SL U59643 ( .A(n1300), .Y(n77969) );
  INVx1_ASAP7_75t_SL U59644 ( .A(n1737), .Y(n78260) );
  INVx1_ASAP7_75t_SL U59645 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[13]), .Y(n78428) );
  INVxp67_ASAP7_75t_SL U59646 ( .A(n1200), .Y(n78073) );
  INVx1_ASAP7_75t_SL U59647 ( .A(n2785), .Y(n61381) );
  INVx1_ASAP7_75t_SL U59648 ( .A(or1200_cpu_or1200_except_n522), .Y(n75312) );
  INVx1_ASAP7_75t_SL U59649 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1[2]), .Y(n27433) );
  INVxp67_ASAP7_75t_SL U59650 ( .A(n3426), .Y(n76836) );
  INVxp67_ASAP7_75t_SL U59651 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_32_), .Y(n78396) );
  NAND2xp5_ASAP7_75t_SL U59652 ( .A(n2117), .B(n2105), .Y(n60854) );
  INVxp67_ASAP7_75t_SL U59653 ( .A(n2469), .Y(n77530) );
  INVx1_ASAP7_75t_SL U59654 ( .A(or1200_cpu_or1200_except_n512), .Y(n77288) );
  NAND2xp33_ASAP7_75t_SL U59655 ( .A(n2970), .B(n2691), .Y(n59959) );
  INVxp33_ASAP7_75t_SL U59656 ( .A(n2598), .Y(n76672) );
  INVxp33_ASAP7_75t_SL U59657 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[34]), .Y(n65711) );
  INVx1_ASAP7_75t_SL U59658 ( .A(or1200_cpu_or1200_except_n514), .Y(n77227) );
  INVxp33_ASAP7_75t_SL U59659 ( .A(n3045), .Y(n76831) );
  INVx1_ASAP7_75t_SL U59660 ( .A(or1200_cpu_or1200_except_n510), .Y(n76553) );
  INVx1_ASAP7_75t_SL U59661 ( .A(n3078), .Y(n61028) );
  INVxp67_ASAP7_75t_SL U59662 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_30_), .Y(n78397) );
  INVx1_ASAP7_75t_SL U59663 ( .A(or1200_cpu_or1200_except_n506), .Y(n76253) );
  INVxp67_ASAP7_75t_SL U59664 ( .A(n2621), .Y(n77518) );
  INVx1_ASAP7_75t_SL U59665 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_4_), .Y(n28213) );
  INVxp33_ASAP7_75t_SL U59666 ( .A(n1582), .Y(n65268) );
  INVxp33_ASAP7_75t_SL U59667 ( .A(or1200_cpu_or1200_mult_mac_n104), .Y(n60803) );
  INVxp67_ASAP7_75t_SL U59668 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[21]), .Y(n28175)
         );
  INVxp67_ASAP7_75t_SL U59669 ( .A(n1207), .Y(dwb_adr_o[27]) );
  INVx1_ASAP7_75t_SL U59670 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[37]), .Y(n65745) );
  INVx1_ASAP7_75t_SL U59671 ( .A(or1200_cpu_or1200_mult_mac_n307), .Y(n63422)
         );
  INVxp67_ASAP7_75t_SL U59672 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[22]), .Y(n28176)
         );
  INVx1_ASAP7_75t_SL U59673 ( .A(n1330), .Y(n77975) );
  INVxp33_ASAP7_75t_SL U59674 ( .A(or1200_cpu_or1200_mult_mac_n108), .Y(n61764) );
  INVxp67_ASAP7_75t_SL U59675 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[23]), .Y(n28177)
         );
  INVx1_ASAP7_75t_SL U59676 ( .A(or1200_cpu_or1200_mult_mac_n315), .Y(n63483)
         );
  INVxp33_ASAP7_75t_SL U59677 ( .A(or1200_cpu_or1200_mult_mac_n100), .Y(n60811) );
  INVxp67_ASAP7_75t_SL U59678 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_3_), .Y(n78423) );
  INVxp67_ASAP7_75t_SL U59679 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[24]), .Y(n28178)
         );
  INVxp67_ASAP7_75t_SL U59680 ( .A(n1212), .Y(dwb_adr_o[26]) );
  INVx1_ASAP7_75t_SL U59681 ( .A(or1200_cpu_or1200_mult_mac_n313), .Y(n63490)
         );
  INVxp67_ASAP7_75t_SL U59682 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[25]), .Y(n28179)
         );
  INVxp67_ASAP7_75t_SL U59683 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_2_), .Y(n78228) );
  INVxp67_ASAP7_75t_SL U59684 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[27]), .Y(n28181)
         );
  INVx1_ASAP7_75t_SL U59685 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_1_), .Y(n28210) );
  INVxp67_ASAP7_75t_SL U59686 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[28]), .Y(n28182)
         );
  INVxp67_ASAP7_75t_SL U59687 ( .A(n1217), .Y(dwb_adr_o[25]) );
  INVxp67_ASAP7_75t_SL U59688 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[29]), .Y(n28183)
         );
  INVx1_ASAP7_75t_SL U59689 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_0_), .Y(n78421) );
  INVxp33_ASAP7_75t_SL U59690 ( .A(n971), .Y(n78039) );
  INVxp67_ASAP7_75t_SL U59691 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[30]), .Y(n28184)
         );
  INVxp67_ASAP7_75t_SL U59692 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[46]), .Y(n65742) );
  INVxp67_ASAP7_75t_SL U59693 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[31]), .Y(n28185)
         );
  INVxp67_ASAP7_75t_SL U59694 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_45_), .Y(n78385) );
  INVx1_ASAP7_75t_SL U59695 ( .A(n1325), .Y(n77978) );
  INVxp33_ASAP7_75t_SL U59696 ( .A(or1200_cpu_or1200_mult_mac_n289), .Y(n60805) );
  INVxp67_ASAP7_75t_SL U59697 ( .A(n1227), .Y(dwb_adr_o[23]) );
  INVxp33_ASAP7_75t_SL U59698 ( .A(n3423), .Y(n60589) );
  INVx1_ASAP7_75t_SL U59699 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_16_), .Y(n78431) );
  INVxp67_ASAP7_75t_SL U59700 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_44_), .Y(n78386) );
  NAND2xp5_ASAP7_75t_SL U59701 ( .A(n2807), .B(n2581), .Y(n60685) );
  INVxp67_ASAP7_75t_SL U59702 ( .A(or1200_cpu_or1200_mult_mac_n311), .Y(n63451) );
  INVxp33_ASAP7_75t_SL U59703 ( .A(or1200_cpu_or1200_mult_mac_n126), .Y(n60965) );
  INVxp67_ASAP7_75t_SL U59704 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[32]), .Y(n28186)
         );
  INVxp33_ASAP7_75t_SL U59705 ( .A(or1200_cpu_or1200_mult_mac_n287), .Y(n60647) );
  INVxp67_ASAP7_75t_SL U59706 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[33]), .Y(n28187)
         );
  INVx1_ASAP7_75t_SL U59707 ( .A(n2567), .Y(n60686) );
  INVxp33_ASAP7_75t_SL U59708 ( .A(or1200_cpu_or1200_mult_mac_n128), .Y(n60631) );
  INVx1_ASAP7_75t_SL U59709 ( .A(n1320), .Y(n77981) );
  INVxp67_ASAP7_75t_SL U59710 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_42_), .Y(n78388) );
  NAND2xp5_ASAP7_75t_SL U59711 ( .A(n2843), .B(n3419), .Y(n77759) );
  INVxp67_ASAP7_75t_SL U59712 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[34]), .Y(n28188)
         );
  INVx1_ASAP7_75t_SL U59713 ( .A(or1200_cpu_or1200_mult_mac_n297), .Y(n63315)
         );
  INVxp67_ASAP7_75t_SL U59714 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[35]), .Y(n28189)
         );
  INVxp33_ASAP7_75t_SL U59715 ( .A(or1200_cpu_or1200_mult_mac_n118), .Y(n61633) );
  INVx1_ASAP7_75t_SL U59716 ( .A(or1200_cpu_spr_dat_ppc[29]), .Y(n75197) );
  INVxp67_ASAP7_75t_SL U59717 ( .A(or1200_cpu_or1200_mult_mac_n299), .Y(n63334) );
  INVx1_ASAP7_75t_SL U59718 ( .A(or1200_cpu_or1200_mult_mac_n231), .Y(n69126)
         );
  INVxp67_ASAP7_75t_SL U59719 ( .A(n1232), .Y(dwb_adr_o[22]) );
  INVxp67_ASAP7_75t_SL U59720 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[36]), .Y(n28190)
         );
  INVx1_ASAP7_75t_SL U59721 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[8]), .Y(n65821) );
  INVxp33_ASAP7_75t_SL U59722 ( .A(or1200_cpu_or1200_mult_mac_n116), .Y(n62268) );
  INVxp67_ASAP7_75t_SL U59723 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[37]), .Y(n28191)
         );
  INVx1_ASAP7_75t_SL U59724 ( .A(or1200_cpu_or1200_mult_mac_n179), .Y(n74584)
         );
  INVxp67_ASAP7_75t_SL U59725 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[6]), .Y(n65824) );
  INVx1_ASAP7_75t_SL U59726 ( .A(or1200_cpu_or1200_mult_mac_n293), .Y(n63300)
         );
  INVx1_ASAP7_75t_SL U59727 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[2]), .Y(n65786) );
  INVxp67_ASAP7_75t_SL U59728 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_41_), .Y(n78389) );
  INVxp33_ASAP7_75t_SL U59729 ( .A(or1200_cpu_or1200_mult_mac_n122), .Y(n60806) );
  INVxp67_ASAP7_75t_SL U59730 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[38]), .Y(n28208)
         );
  INVxp67_ASAP7_75t_SL U59731 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[1]), .Y(n65785) );
  INVx1_ASAP7_75t_SL U59732 ( .A(n1352), .Y(n74581) );
  INVx1_ASAP7_75t_SL U59733 ( .A(n1315), .Y(n77984) );
  INVxp67_ASAP7_75t_SL U59734 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_40_), .Y(n78390) );
  INVxp33_ASAP7_75t_SL U59735 ( .A(or1200_cpu_or1200_mult_mac_n295), .Y(n61418) );
  INVxp67_ASAP7_75t_SL U59736 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[40]), .Y(n28193)
         );
  INVx1_ASAP7_75t_SL U59737 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[3]), .Y(n65788) );
  INVxp67_ASAP7_75t_SL U59738 ( .A(n1242), .Y(dwb_adr_o[20]) );
  INVxp33_ASAP7_75t_SL U59739 ( .A(or1200_cpu_or1200_mult_mac_n120), .Y(n60807) );
  INVxp67_ASAP7_75t_SL U59740 ( .A(n2642), .Y(n77512) );
  INVxp33_ASAP7_75t_SL U59741 ( .A(n2455), .Y(n70296) );
  INVxp67_ASAP7_75t_SL U59742 ( .A(n811), .Y(n59982) );
  INVx1_ASAP7_75t_SL U59743 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_13_), .Y(n78413) );
  INVx1_ASAP7_75t_SL U59744 ( .A(n819), .Y(n60157) );
  INVx1_ASAP7_75t_SL U59745 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[2]), .Y(
        n73244) );
  INVx1_ASAP7_75t_SL U59746 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_14_), .Y(n78412) );
  INVxp33_ASAP7_75t_SL U59747 ( .A(or1200_cpu_or1200_mult_mac_n189), .Y(n64761) );
  INVx1_ASAP7_75t_SL U59748 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_15_), .Y(n78411) );
  INVx1_ASAP7_75t_SL U59749 ( .A(or1200_cpu_or1200_except_n526), .Y(n74578) );
  INVx1_ASAP7_75t_SL U59750 ( .A(n795), .Y(n59984) );
  INVxp67_ASAP7_75t_SL U59751 ( .A(n1265), .Y(n78135) );
  INVxp67_ASAP7_75t_SL U59752 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_16_), .Y(n78410) );
  INVxp67_ASAP7_75t_SL U59753 ( .A(n3027), .Y(n60162) );
  INVx1_ASAP7_75t_SL U59754 ( .A(n787), .Y(n60053) );
  INVx1_ASAP7_75t_SL U59755 ( .A(or1200_cpu_or1200_mult_mac_n181), .Y(n65079)
         );
  INVxp67_ASAP7_75t_SL U59756 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[3]), .Y(
        n73238) );
  INVxp67_ASAP7_75t_SL U59757 ( .A(n1260), .Y(n78130) );
  INVxp67_ASAP7_75t_SL U59758 ( .A(n1225), .Y(n78102) );
  INVx1_ASAP7_75t_SL U59759 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[8]), .Y(
        n73211) );
  INVxp67_ASAP7_75t_SL U59760 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_17_), .Y(n78409) );
  INVx1_ASAP7_75t_SL U59761 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[1]), .Y(n73601)
         );
  INVx1_ASAP7_75t_SL U59762 ( .A(n1038), .Y(n78047) );
  INVx1_ASAP7_75t_SL U59763 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_18_), .Y(n78408) );
  INVxp67_ASAP7_75t_SL U59764 ( .A(n1255), .Y(n78126) );
  INVx1_ASAP7_75t_SL U59765 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_26_), .Y(n78400) );
  NAND2xp33_ASAP7_75t_SL U59766 ( .A(n3337), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .Y(
        n73709) );
  INVxp67_ASAP7_75t_SL U59767 ( .A(n1282), .Y(dwb_adr_o[12]) );
  INVxp67_ASAP7_75t_SL U59768 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[24]), .Y(n78194) );
  INVxp67_ASAP7_75t_SL U59769 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_2_), .Y(n70255) );
  INVx1_ASAP7_75t_SL U59770 ( .A(or1200_cpu_spr_dat_ppc[20]), .Y(n74126) );
  INVxp33_ASAP7_75t_SL U59771 ( .A(or1200_cpu_or1200_except_n120), .Y(n77443)
         );
  INVxp67_ASAP7_75t_SL U59772 ( .A(n1230), .Y(n78106) );
  INVxp67_ASAP7_75t_SL U59773 ( .A(n1250), .Y(n78122) );
  NAND2xp5_ASAP7_75t_SL U59774 ( .A(or1200_cpu_or1200_mult_mac_n217), .B(
        or1200_cpu_or1200_mult_mac_n363), .Y(n69000) );
  INVx1_ASAP7_75t_SL U59775 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[4]), .Y(
        n73219) );
  INVx1_ASAP7_75t_SL U59776 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_25_), .Y(n78401) );
  INVx1_ASAP7_75t_SL U59777 ( .A(n2587), .Y(n63267) );
  INVxp67_ASAP7_75t_SL U59778 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .Y(n65857) );
  INVx1_ASAP7_75t_SL U59779 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_19_), .Y(n78407) );
  INVx1_ASAP7_75t_SL U59780 ( .A(or1200_cpu_or1200_mult_mac_n203), .Y(n68814)
         );
  INVx1_ASAP7_75t_SL U59781 ( .A(n2994), .Y(n65220) );
  INVx1_ASAP7_75t_SL U59782 ( .A(n1060), .Y(n78051) );
  INVxp67_ASAP7_75t_SL U59783 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[6]), .Y(
        n73264) );
  INVxp67_ASAP7_75t_SL U59784 ( .A(n1245), .Y(n78118) );
  INVx1_ASAP7_75t_SL U59785 ( .A(n1049), .Y(n78049) );
  INVx1_ASAP7_75t_SL U59786 ( .A(or1200_cpu_or1200_except_n276), .Y(n77002) );
  INVxp33_ASAP7_75t_SL U59787 ( .A(n2451), .Y(n69376) );
  INVx1_ASAP7_75t_SL U59788 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[16]), .Y(
        n73129) );
  INVxp67_ASAP7_75t_SL U59789 ( .A(n2581), .Y(n60841) );
  INVx1_ASAP7_75t_SL U59790 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_20_), .Y(n78406) );
  INVx1_ASAP7_75t_SL U59791 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_24_), .Y(n78402) );
  INVxp67_ASAP7_75t_SL U59792 ( .A(n1235), .Y(n78110) );
  INVxp33_ASAP7_75t_SL U59793 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_20_), .Y(n65297) );
  INVxp67_ASAP7_75t_SL U59794 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]), .Y(n65833) );
  INVx1_ASAP7_75t_SL U59795 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_21_), .Y(n78405) );
  INVxp67_ASAP7_75t_SL U59796 ( .A(or1200_cpu_or1200_except_n244), .Y(n60020)
         );
  INVxp67_ASAP7_75t_SL U59797 ( .A(n1240), .Y(n78114) );
  INVx2_ASAP7_75t_SL U59798 ( .A(n2456), .Y(n70477) );
  INVx1_ASAP7_75t_SL U59799 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_23_), .Y(n78403) );
  INVx1_ASAP7_75t_SL U59800 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_22_), .Y(n78404) );
  INVxp33_ASAP7_75t_SL U59801 ( .A(or1200_cpu_or1200_genpc_pcreg_default[6]), 
        .Y(n61171) );
  INVxp67_ASAP7_75t_SL U59802 ( .A(n3051), .Y(n61174) );
  INVx1_ASAP7_75t_SL U59803 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[6]), .Y(
        n73265) );
  INVx1_ASAP7_75t_SL U59804 ( .A(or1200_cpu_or1200_except_n508), .Y(n75783) );
  INVxp67_ASAP7_75t_SL U59805 ( .A(n3015), .Y(n60139) );
  INVxp67_ASAP7_75t_SL U59806 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[38]), .Y(n65804) );
  INVxp67_ASAP7_75t_SL U59807 ( .A(n1267), .Y(dwb_adr_o[15]) );
  INVx1_ASAP7_75t_SL U59808 ( .A(or1200_cpu_or1200_except_n504), .Y(n76851) );
  INVxp67_ASAP7_75t_SL U59809 ( .A(n2635), .Y(n77514) );
  INVxp67_ASAP7_75t_SL U59810 ( .A(n2129), .Y(n60614) );
  INVxp67_ASAP7_75t_SL U59811 ( .A(n1205), .Y(n78077) );
  INVxp67_ASAP7_75t_SL U59812 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[25]), .Y(n78193) );
  INVx1_ASAP7_75t_SL U59813 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_29_), .Y(n78398) );
  INVx1_ASAP7_75t_SL U59814 ( .A(n2141), .Y(n60855) );
  INVx1_ASAP7_75t_SL U59815 ( .A(or1200_cpu_or1200_except_n500), .Y(n76619) );
  INVxp67_ASAP7_75t_SL U59816 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[10]), .Y(
        n73163) );
  INVx1_ASAP7_75t_SL U59817 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[1]), .Y(
        n27713) );
  INVxp67_ASAP7_75t_SL U59818 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_sign), .Y(n28160) );
  INVxp67_ASAP7_75t_SL U59819 ( .A(n1285), .Y(n78156) );
  NAND2xp33_ASAP7_75t_SL U59820 ( .A(or1200_cpu_or1200_mult_mac_n253), .B(
        or1200_cpu_or1200_mult_mac_n399), .Y(n69312) );
  INVx1_ASAP7_75t_SL U59821 ( .A(or1200_cpu_or1200_except_n516), .Y(n77021) );
  INVxp67_ASAP7_75t_SL U59822 ( .A(or1200_cpu_or1200_genpc_pcreg_default[4]), 
        .Y(n61168) );
  INVxp67_ASAP7_75t_SL U59823 ( .A(n3417), .Y(n59995) );
  INVx1_ASAP7_75t_SL U59824 ( .A(or1200_cpu_or1200_except_n518), .Y(n77153) );
  INVx1_ASAP7_75t_SL U59825 ( .A(or1200_cpu_or1200_except_n532), .Y(n75449) );
  INVx1_ASAP7_75t_SL U59826 ( .A(or1200_cpu_or1200_except_n534), .Y(n75622) );
  INVxp67_ASAP7_75t_SL U59827 ( .A(n1272), .Y(dwb_adr_o[14]) );
  INVx1_ASAP7_75t_SL U59828 ( .A(or1200_cpu_or1200_except_n548), .Y(n75686) );
  INVx1_ASAP7_75t_SL U59829 ( .A(n2464), .Y(n69335) );
  INVxp67_ASAP7_75t_SL U59830 ( .A(n1608), .Y(n74074) );
  INVxp67_ASAP7_75t_SL U59831 ( .A(or1200_cpu_or1200_mult_mac_n399), .Y(n69309) );
  INVxp67_ASAP7_75t_SL U59832 ( .A(n1280), .Y(n78151) );
  INVx1_ASAP7_75t_SL U59833 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_28_), .Y(n78399) );
  INVx1_ASAP7_75t_SL U59834 ( .A(n1071), .Y(n78053) );
  INVx1_ASAP7_75t_SL U59835 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[1]), .Y(
        n73227) );
  INVx1_ASAP7_75t_SL U59836 ( .A(or1200_cpu_or1200_except_n246), .Y(n75208) );
  INVx1_ASAP7_75t_SL U59837 ( .A(n2791), .Y(n77006) );
  INVxp67_ASAP7_75t_SL U59838 ( .A(n1628), .Y(n64154) );
  INVx1_ASAP7_75t_SL U59839 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[11]), .Y(
        n73169) );
  INVx1_ASAP7_75t_SL U59840 ( .A(or1200_cpu_or1200_mult_mac_n255), .Y(n69324)
         );
  INVxp67_ASAP7_75t_SL U59841 ( .A(n1210), .Y(n78081) );
  INVxp67_ASAP7_75t_SL U59842 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[2]), .Y(
        n73241) );
  INVx1_ASAP7_75t_SL U59843 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[16]), .Y(n78425) );
  INVxp67_ASAP7_75t_SL U59844 ( .A(n1275), .Y(n78145) );
  INVxp67_ASAP7_75t_SL U59845 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_1_), .Y(n78326) );
  INVxp33_ASAP7_75t_SL U59846 ( .A(n1016), .Y(n78044) );
  INVx2_ASAP7_75t_SL U59847 ( .A(n59697), .Y(n57211) );
  AND3x1_ASAP7_75t_SL U59848 ( .A(or1200_cpu_or1200_genpc_pcreg_default[7]), 
        .B(or1200_cpu_or1200_genpc_pcreg_default[6]), .C(
        or1200_cpu_or1200_genpc_pcreg_default[4]), .Y(n59979) );
  INVx1_ASAP7_75t_SL U59849 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_7_), .Y(n78419) );
  INVxp67_ASAP7_75t_SL U59850 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_8_), .Y(n78418) );
  INVxp67_ASAP7_75t_SL U59851 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[1]), .Y(
        n73229) );
  INVx1_ASAP7_75t_SL U59852 ( .A(or1200_cpu_or1200_genpc_pcreg_default[3]), 
        .Y(n61167) );
  INVxp67_ASAP7_75t_SL U59853 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_9_), .Y(n78417) );
  INVxp67_ASAP7_75t_SL U59854 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_0_), .Y(n78247) );
  INVx1_ASAP7_75t_SL U59855 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_10_), .Y(n78416) );
  INVxp67_ASAP7_75t_SL U59856 ( .A(n1215), .Y(n78085) );
  INVx1_ASAP7_75t_SL U59857 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[9]), .Y(
        n73156) );
  INVx1_ASAP7_75t_SL U59858 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_11_), .Y(n78415) );
  INVxp33_ASAP7_75t_SL U59859 ( .A(or1200_cpu_or1200_except_n202), .Y(n63731)
         );
  INVx1_ASAP7_75t_SL U59860 ( .A(n1339), .Y(dwb_adr_o[2]) );
  INVx1_ASAP7_75t_SL U59861 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[3]), .Y(
        n73239) );
  INVxp67_ASAP7_75t_SL U59862 ( .A(n1270), .Y(n78141) );
  INVx1_ASAP7_75t_SL U59863 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_12_), .Y(n78414) );
  INVx1_ASAP7_75t_SL U59864 ( .A(or1200_cpu_or1200_except_n431), .Y(n77224) );
  INVxp67_ASAP7_75t_SL U59865 ( .A(n3048), .Y(n63730) );
  INVx1_ASAP7_75t_SL U59866 ( .A(or1200_cpu_spr_dat_ppc[24]), .Y(n74044) );
  INVxp67_ASAP7_75t_SL U59867 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[20]), .Y(n28174)
         );
  INVx1_ASAP7_75t_SL U59868 ( .A(or1200_cpu_or1200_mult_mac_n265), .Y(n76894)
         );
  INVx1_ASAP7_75t_SL U59869 ( .A(or1200_cpu_or1200_except_n440), .Y(n76230) );
  INVxp67_ASAP7_75t_SL U59870 ( .A(or1200_cpu_or1200_mult_mac_n301), .Y(n76754) );
  INVx1_ASAP7_75t_SL U59871 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .Y(n65454) );
  INVx1_ASAP7_75t_SL U59872 ( .A(or1200_cpu_or1200_mult_mac_n241), .Y(n69188)
         );
  INVxp33_ASAP7_75t_SL U59873 ( .A(n852), .Y(n78026) );
  INVx1_ASAP7_75t_SL U59874 ( .A(n1159), .Y(n62404) );
  INVx1_ASAP7_75t_SL U59875 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[25]), .Y(
        n73381) );
  INVx1_ASAP7_75t_SL U59876 ( .A(n1104), .Y(n78064) );
  INVxp33_ASAP7_75t_SL U59877 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .Y(n65630) );
  NOR3xp33_ASAP7_75t_SRAM U59878 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_17_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_), 
        .C(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_22_), 
        .Y(n71430) );
  INVx1_ASAP7_75t_SL U59879 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_qnan_d), .Y(n74889) );
  INVxp33_ASAP7_75t_SL U59880 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_inf_d), .Y(n76974) );
  INVxp33_ASAP7_75t_SL U59881 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]), .Y(n65635) );
  INVx1_ASAP7_75t_SL U59882 ( .A(or1200_cpu_or1200_except_n524), .Y(n74986) );
  INVx1_ASAP7_75t_SL U59883 ( .A(or1200_cpu_spr_dat_ppc[17]), .Y(n75301) );
  INVx1_ASAP7_75t_SL U59884 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_4_), .Y(n78335) );
  INVx1_ASAP7_75t_SL U59885 ( .A(n2741), .Y(n61024) );
  INVx1_ASAP7_75t_SL U59886 ( .A(or1200_cpu_or1200_mult_mac_n225), .Y(n69024)
         );
  INVx1_ASAP7_75t_SL U59887 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[14]), .Y(
        n73140) );
  INVx1_ASAP7_75t_SL U59888 ( .A(or1200_cpu_or1200_except_n446), .Y(n74983) );
  INVx1_ASAP7_75t_SL U59889 ( .A(n1167), .Y(n62302) );
  INVx1_ASAP7_75t_SL U59890 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_5_), .Y(n78337) );
  INVx1_ASAP7_75t_SL U59891 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[4]), .Y(
        n73217) );
  INVx1_ASAP7_75t_SL U59892 ( .A(n2743), .Y(n61591) );
  INVx1_ASAP7_75t_SL U59893 ( .A(or1200_cpu_spr_dat_ppc[19]), .Y(n74576) );
  INVxp33_ASAP7_75t_SL U59894 ( .A(n1095), .Y(n63688) );
  INVxp67_ASAP7_75t_SL U59895 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_23_), .Y(n69713) );
  INVxp33_ASAP7_75t_SL U59896 ( .A(n2678), .Y(n60524) );
  NOR2xp33_ASAP7_75t_SRAM U59897 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_12_), .Y(
        n74668) );
  AND3x1_ASAP7_75t_SL U59898 ( .A(n2107), .B(n2119), .C(n78439), .Y(n59932) );
  INVxp67_ASAP7_75t_SL U59899 ( .A(n2865), .Y(n65257) );
  INVxp33_ASAP7_75t_SL U59900 ( .A(n1084), .Y(n63689) );
  INVx1_ASAP7_75t_SL U59901 ( .A(n1175), .Y(n62221) );
  INVx1_ASAP7_75t_SL U59902 ( .A(n1173), .Y(n62220) );
  INVx1_ASAP7_75t_SL U59903 ( .A(n2997), .Y(n65210) );
  INVx1_ASAP7_75t_SL U59904 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[35]), .Y(n65743) );
  INVx1_ASAP7_75t_SL U59905 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_18_), .Y(n78355) );
  INVx1_ASAP7_75t_SL U59906 ( .A(or1200_cpu_or1200_except_n528), .Y(n74129) );
  INVx1_ASAP7_75t_SL U59907 ( .A(or1200_cpu_or1200_except_n236), .Y(n64758) );
  INVx1_ASAP7_75t_SL U59908 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[36]), .Y(n65853) );
  INVx1_ASAP7_75t_SL U59909 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[26]), .Y(
        n73377) );
  INVx1_ASAP7_75t_SL U59910 ( .A(n2745), .Y(n60893) );
  INVx1_ASAP7_75t_SL U59911 ( .A(or1200_cpu_spr_dat_ppc[21]), .Y(n75430) );
  INVx1_ASAP7_75t_SL U59912 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[33]), .Y(n65858) );
  NAND2xp5_ASAP7_75t_SL U59913 ( .A(or1200_cpu_or1200_fpu_fpu_op_valid_re_r), 
        .B(or1200_cpu_or1200_fpu_fpu_op_r_3_), .Y(n76492) );
  AOI21xp33_ASAP7_75t_SL U59914 ( .A1(n1426), .A2(n1428), .B(dbg_stall_i), .Y(
        n62198) );
  INVx1_ASAP7_75t_SL U59915 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_19_), .Y(n78357) );
  INVxp33_ASAP7_75t_SL U59916 ( .A(n823), .Y(n60043) );
  INVx1_ASAP7_75t_SL U59917 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_2_), .Y(n78436) );
  INVxp67_ASAP7_75t_SL U59918 ( .A(n2506), .Y(n77528) );
  INVx1_ASAP7_75t_SL U59919 ( .A(n3030), .Y(n63968) );
  INVx1_ASAP7_75t_SL U59920 ( .A(or1200_cpu_spr_dat_ppc[22]), .Y(n75446) );
  INVx1_ASAP7_75t_SL U59921 ( .A(n1426), .Y(n62201) );
  INVx1_ASAP7_75t_SL U59922 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_6_), .Y(n78339) );
  INVx1_ASAP7_75t_SL U59923 ( .A(n2735), .Y(n60397) );
  INVx1_ASAP7_75t_SL U59924 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[2]), .Y(n70705) );
  INVxp67_ASAP7_75t_SL U59925 ( .A(or1200_cpu_or1200_except_n262), .Y(n75474)
         );
  INVx1_ASAP7_75t_SL U59926 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[18]), .Y(n65631) );
  INVx1_ASAP7_75t_SL U59927 ( .A(n1157), .Y(n62484) );
  INVx1_ASAP7_75t_SL U59928 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[4]), .Y(
        n27731) );
  INVx1_ASAP7_75t_SL U59929 ( .A(or1200_cpu_or1200_mult_mac_n155), .Y(n76722)
         );
  INVx1_ASAP7_75t_SL U59930 ( .A(or1200_cpu_or1200_except_n422), .Y(n75780) );
  INVx1_ASAP7_75t_SL U59931 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_9_), .Y(n78345) );
  INVx1_ASAP7_75t_SL U59932 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[3]), .Y(
        n27729) );
  INVxp67_ASAP7_75t_SL U59933 ( .A(n1161), .Y(n62399) );
  INVx1_ASAP7_75t_SL U59934 ( .A(or1200_cpu_or1200_mult_mac_n219), .Y(n76721)
         );
  INVx1_ASAP7_75t_SL U59935 ( .A(n1163), .Y(n62400) );
  INVxp67_ASAP7_75t_SL U59936 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_ine_o), 
        .Y(n27728) );
  INVxp67_ASAP7_75t_SL U59937 ( .A(n2976), .Y(n59998) );
  INVx3_ASAP7_75t_SL U59938 ( .A(n59528), .Y(n57212) );
  NOR2xp33_ASAP7_75t_SRAM U59939 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[44]), .Y(n65459) );
  INVx1_ASAP7_75t_SL U59940 ( .A(or1200_cpu_or1200_except_n425), .Y(n76551) );
  INVx1_ASAP7_75t_SL U59941 ( .A(n831), .Y(n77802) );
  INVx1_ASAP7_75t_SL U59942 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_6_), .Y(n74172) );
  INVx1_ASAP7_75t_SL U59943 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[1]), .Y(n70691) );
  INVxp33_ASAP7_75t_SL U59944 ( .A(n1165), .Y(n62305) );
  INVx1_ASAP7_75t_SL U59945 ( .A(n2687), .Y(n76736) );
  INVx1_ASAP7_75t_SL U59946 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[22]), .Y(n70045) );
  INVx1_ASAP7_75t_SL U59947 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_N398), .Y(n74208) );
  INVxp33_ASAP7_75t_SL U59948 ( .A(or1200_cpu_or1200_mult_mac_n377), .Y(n69127) );
  INVxp67_ASAP7_75t_SL U59949 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[0]), .Y(n70687) );
  INVx1_ASAP7_75t_SL U59950 ( .A(or1200_cpu_or1200_except_n428), .Y(n77291) );
  INVx1_ASAP7_75t_SL U59951 ( .A(n2737), .Y(n60391) );
  INVx1_ASAP7_75t_SL U59952 ( .A(or1200_cpu_or1200_mult_mac_n173), .Y(n63536)
         );
  INVx1_ASAP7_75t_SL U59953 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[4]), .Y(n78334)
         );
  INVxp67_ASAP7_75t_SL U59954 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .Y(
        n70317) );
  INVxp33_ASAP7_75t_SL U59955 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]), .Y(n74050) );
  INVx1_ASAP7_75t_SL U59956 ( .A(or1200_cpu_or1200_mult_mac_n245), .Y(n74114)
         );
  INVxp67_ASAP7_75t_SL U59957 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[26]), .Y(
        n73373) );
  INVx1_ASAP7_75t_SL U59958 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[0]), .Y(n73609)
         );
  INVx1_ASAP7_75t_SL U59959 ( .A(n1356), .Y(n74972) );
  INVx1_ASAP7_75t_SL U59960 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_4_), .Y(n74188) );
  INVx1_ASAP7_75t_SL U59961 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_), .Y(n78433) );
  INVxp67_ASAP7_75t_SL U59962 ( .A(n755), .Y(n59974) );
  INVxp67_ASAP7_75t_SL U59963 ( .A(n3063), .Y(n63742) );
  INVxp67_ASAP7_75t_SL U59964 ( .A(or1200_cpu_or1200_mult_mac_n149), .Y(n63325) );
  INVxp67_ASAP7_75t_SL U59965 ( .A(or1200_cpu_or1200_except_n192), .Y(n63744)
         );
  INVx1_ASAP7_75t_SL U59966 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1[1]), .Y(n78251) );
  INVx1_ASAP7_75t_SL U59967 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[7]), .Y(n70652) );
  INVx1_ASAP7_75t_SL U59968 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[15]), .Y(
        n73150) );
  INVx1_ASAP7_75t_SL U59969 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_1_), .Y(n78250) );
  INVxp67_ASAP7_75t_SL U59970 ( .A(or1200_cpu_or1200_except_n248), .Y(n60005)
         );
  INVx1_ASAP7_75t_SL U59971 ( .A(or1200_cpu_or1200_except_n437), .Y(n77151) );
  INVx1_ASAP7_75t_SL U59972 ( .A(n2739), .Y(n60385) );
  INVx1_ASAP7_75t_SL U59973 ( .A(or1200_cpu_or1200_mult_mac_n393), .Y(n69243)
         );
  INVx1_ASAP7_75t_SL U59974 ( .A(or1200_cpu_or1200_mult_mac_n369), .Y(n69022)
         );
  INVx1_ASAP7_75t_SL U59975 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_3_), .Y(n78333) );
  INVxp33_ASAP7_75t_SL U59976 ( .A(n2798), .Y(n76719) );
  INVxp67_ASAP7_75t_SL U59977 ( .A(n1983), .Y(n60222) );
  INVx1_ASAP7_75t_SL U59978 ( .A(or1200_cpu_or1200_mult_mac_n333), .Y(n65146)
         );
  INVxp33_ASAP7_75t_SL U59979 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .Y(n65613) );
  INVxp67_ASAP7_75t_SL U59980 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[0]), .Y(n28198) );
  INVxp67_ASAP7_75t_SL U59981 ( .A(or1200_cpu_or1200_mult_mac_n257), .Y(n75116) );
  INVxp67_ASAP7_75t_SL U59982 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[1]), .Y(n28199) );
  INVx1_ASAP7_75t_SL U59983 ( .A(n2753), .Y(n60365) );
  INVxp33_ASAP7_75t_SL U59984 ( .A(n783), .Y(n60071) );
  INVxp67_ASAP7_75t_SL U59985 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[2]), .Y(n28200) );
  INVx1_ASAP7_75t_SL U59986 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_15_), .Y(n78353) );
  AND3x1_ASAP7_75t_SL U59987 ( .A(n1533), .B(n1112), .C(n748), .Y(n60236) );
  INVxp67_ASAP7_75t_SL U59988 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[4]), .Y(n28202) );
  INVx1_ASAP7_75t_SL U59989 ( .A(n3000), .Y(n75544) );
  INVxp67_ASAP7_75t_SL U59990 ( .A(n2614), .Y(n77520) );
  INVx1_ASAP7_75t_SL U59991 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[7]), .Y(n78340)
         );
  INVxp67_ASAP7_75t_SL U59992 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[5]), .Y(n28203) );
  INVxp33_ASAP7_75t_SL U59993 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[13]), .Y(n65725) );
  INVx1_ASAP7_75t_SL U59994 ( .A(or1200_cpu_or1200_mult_mac_n323), .Y(n63891)
         );
  AND4x1_ASAP7_75t_SL U59995 ( .A(n1496), .B(n1489), .C(n1519), .D(n1499), .Y(
        n60235) );
  INVxp67_ASAP7_75t_SL U59996 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[6]), .Y(n28204) );
  INVxp33_ASAP7_75t_SL U59997 ( .A(or1200_cpu_or1200_mult_mac_n325), .Y(n61822) );
  INVx1_ASAP7_75t_SL U59998 ( .A(n2499), .Y(n69343) );
  INVxp67_ASAP7_75t_SL U59999 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[44]), .Y(n65855) );
  INVx1_ASAP7_75t_SL U60000 ( .A(or1200_cpu_or1200_except_n679), .Y(n75769) );
  INVxp67_ASAP7_75t_SL U60001 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[7]), .Y(n28161) );
  INVxp33_ASAP7_75t_SL U60002 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .Y(n65583) );
  INVx1_ASAP7_75t_SL U60003 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[0]), .Y(
        n73231) );
  INVxp67_ASAP7_75t_SL U60004 ( .A(or1200_cpu_or1200_mult_mac_n331), .Y(n65124) );
  INVxp33_ASAP7_75t_SL U60005 ( .A(or1200_cpu_or1200_mult_mac_n84), .Y(n64305)
         );
  INVxp67_ASAP7_75t_SL U60006 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[8]), .Y(n28162) );
  INVxp67_ASAP7_75t_SL U60007 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[24]), .Y(n65758) );
  BUFx2_ASAP7_75t_SL U60008 ( .A(n1874), .Y(n59550) );
  INVx1_ASAP7_75t_SL U60009 ( .A(n2691), .Y(n59961) );
  INVxp67_ASAP7_75t_SL U60010 ( .A(or1200_cpu_or1200_mult_mac_n82), .Y(n75579)
         );
  INVxp67_ASAP7_75t_SL U60011 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[9]), .Y(n28163) );
  INVxp67_ASAP7_75t_SL U60012 ( .A(or1200_cpu_or1200_mult_mac_n329), .Y(n65095) );
  INVxp67_ASAP7_75t_SL U60013 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[10]), .Y(n28164)
         );
  INVxp67_ASAP7_75t_SL U60014 ( .A(n1573), .Y(n64865) );
  INVx1_ASAP7_75t_SL U60015 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_38_), .Y(n78391) );
  INVxp67_ASAP7_75t_SL U60016 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[11]), .Y(n28165)
         );
  INVx1_ASAP7_75t_SL U60017 ( .A(n1335), .Y(n77972) );
  INVx1_ASAP7_75t_SL U60018 ( .A(or1200_cpu_or1200_except_n280), .Y(n63764) );
  INVxp67_ASAP7_75t_SL U60019 ( .A(or1200_cpu_or1200_mult_mac_n94), .Y(n75337)
         );
  INVxp67_ASAP7_75t_SL U60020 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[13]), .Y(n28167)
         );
  INVx1_ASAP7_75t_SL U60021 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_47_), .Y(n28256) );
  NAND2xp5_ASAP7_75t_SL U60022 ( .A(or1200_cpu_or1200_mult_mac_n261), .B(
        or1200_cpu_or1200_mult_mac_n407), .Y(n75661) );
  INVxp67_ASAP7_75t_SL U60023 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[14]), .Y(n28168)
         );
  INVx1_ASAP7_75t_SL U60024 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]), .Y(n65805) );
  INVxp67_ASAP7_75t_SL U60025 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[26]), .Y(n78192) );
  INVx1_ASAP7_75t_SL U60026 ( .A(or1200_cpu_or1200_mult_mac_n319), .Y(n63537)
         );
  INVx1_ASAP7_75t_SL U60027 ( .A(or1200_cpu_or1200_except_n476), .Y(n77176) );
  INVx1_ASAP7_75t_SL U60028 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_46_), .Y(n78384) );
  INVxp67_ASAP7_75t_SL U60029 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[15]), .Y(n28169)
         );
  INVxp33_ASAP7_75t_SL U60030 ( .A(n815), .Y(n60090) );
  INVxp67_ASAP7_75t_SL U60031 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[16]), .Y(n28170)
         );
  INVx1_ASAP7_75t_SL U60032 ( .A(n1739), .Y(n78253) );
  INVx1_ASAP7_75t_SL U60033 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[39]), .Y(n65578) );
  INVxp67_ASAP7_75t_SL U60034 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[17]), .Y(n28171)
         );
  INVx1_ASAP7_75t_SL U60035 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[2]), .Y(
        n27721) );
  INVxp67_ASAP7_75t_SL U60036 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_43_), .Y(n78387) );
  INVxp67_ASAP7_75t_SL U60037 ( .A(n1197), .Y(dwb_adr_o[29]) );
  INVx1_ASAP7_75t_SL U60038 ( .A(or1200_cpu_or1200_mult_mac_n305), .Y(n63409)
         );
  INVxp67_ASAP7_75t_SL U60039 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[18]), .Y(n28172)
         );
  INVxp67_ASAP7_75t_SL U60040 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_6_), .Y(n78420) );
  INVx1_ASAP7_75t_SL U60041 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_5_), .Y(n78422) );
  INVxp33_ASAP7_75t_SL U60042 ( .A(or1200_cpu_or1200_mult_mac_n110), .Y(n61348) );
  INVx1_ASAP7_75t_SL U60043 ( .A(or1200_cpu_or1200_except_n544), .Y(n77179) );
  INVxp67_ASAP7_75t_SL U60044 ( .A(n1202), .Y(dwb_adr_o[28]) );
  INVx1_ASAP7_75t_SL U60045 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_17_), .Y(n78430) );
  INVxp33_ASAP7_75t_SL U60046 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[45]), .Y(n65854) );
  INVx1_ASAP7_75t_SL U60047 ( .A(or1200_cpu_or1200_except_n461), .Y(n75619) );
  INVxp33_ASAP7_75t_SL U60048 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .Y(n65856) );
  INVx1_ASAP7_75t_SL U60049 ( .A(n2134), .Y(n76809) );
  NAND2xp5_ASAP7_75t_SL U60050 ( .A(or1200_cpu_or1200_except_n290), .B(
        or1200_cpu_or1200_except_n294), .Y(n77436) );
  INVx1_ASAP7_75t_SL U60051 ( .A(n2747), .Y(n60354) );
  INVx1_ASAP7_75t_SL U60052 ( .A(n829), .Y(iwb_adr_o[3]) );
  INVx1_ASAP7_75t_SL U60053 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_20_), .Y(n78369) );
  INVxp67_ASAP7_75t_SL U60054 ( .A(n1787), .Y(n61741) );
  INVxp67_ASAP7_75t_SL U60055 ( .A(n1004), .Y(iwb_adr_o[29]) );
  INVxp33_ASAP7_75t_SL U60056 ( .A(n917), .Y(n78033) );
  INVx1_ASAP7_75t_SL U60057 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[29]), .Y(n65684) );
  INVx1_ASAP7_75t_SL U60058 ( .A(n1093), .Y(n78062) );
  INVx1_ASAP7_75t_SL U60059 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[31]), .Y(n65681) );
  INVx1_ASAP7_75t_SL U60060 ( .A(or1200_cpu_spr_dat_ppc[26]), .Y(n69367) );
  INVx1_ASAP7_75t_SL U60061 ( .A(n2796), .Y(n61681) );
  INVx1_ASAP7_75t_SL U60062 ( .A(n2749), .Y(n60347) );
  INVx1_ASAP7_75t_SL U60063 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_21_), .Y(n78367) );
  INVxp67_ASAP7_75t_SL U60064 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[25]), .Y(n65761) );
  INVx1_ASAP7_75t_SL U60065 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[6]), .Y(n78338)
         );
  INVx1_ASAP7_75t_SL U60066 ( .A(n1961), .Y(n62237) );
  INVx1_ASAP7_75t_SL U60067 ( .A(or1200_cpu_spr_dat_ppc[27]), .Y(n75795) );
  INVx1_ASAP7_75t_SL U60068 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[27]), .Y(n65831) );
  INVxp67_ASAP7_75t_SL U60069 ( .A(or1200_cpu_or1200_mult_mac_n343), .Y(n75855) );
  INVx1_ASAP7_75t_SL U60070 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), .Y(n65832) );
  INVx1_ASAP7_75t_SL U60071 ( .A(n2751), .Y(n60375) );
  INVx1_ASAP7_75t_SL U60072 ( .A(or1200_cpu_or1200_mult_mac_n341), .Y(n68791)
         );
  INVx1_ASAP7_75t_SL U60073 ( .A(or1200_cpu_or1200_except_n542), .Y(n75798) );
  INVxp67_ASAP7_75t_SL U60074 ( .A(or1200_cpu_or1200_except_n206), .Y(n61271)
         );
  INVxp67_ASAP7_75t_SL U60075 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[17]), .Y(
        n73133) );
  INVxp33_ASAP7_75t_SL U60076 ( .A(n791), .Y(n60060) );
  INVxp67_ASAP7_75t_SL U60077 ( .A(or1200_cpu_except_type_1_), .Y(n77247) );
  INVx1_ASAP7_75t_SL U60078 ( .A(n3006), .Y(n75418) );
  INVx1_ASAP7_75t_SL U60079 ( .A(n2961), .Y(n74034) );
  INVx1_ASAP7_75t_SL U60080 ( .A(n2970), .Y(n59993) );
  OAI21xp33_ASAP7_75t_SL U60081 ( .A1(n2691), .A2(n3123), .B(n2598), .Y(n59957) );
  INVxp67_ASAP7_75t_SL U60082 ( .A(or1200_cpu_or1200_mult_mac_n80), .Y(n61816)
         );
  INVx1_ASAP7_75t_SL U60083 ( .A(or1200_cpu_or1200_mult_mac_n335), .Y(n65140)
         );
  INVxp67_ASAP7_75t_SL U60084 ( .A(n3042), .Y(n61270) );
  INVx1_ASAP7_75t_SL U60085 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[2]), .Y(n73595)
         );
  INVx1_ASAP7_75t_SL U60086 ( .A(or1200_cpu_or1200_mult_mac_n367), .Y(n68985)
         );
  INVx1_ASAP7_75t_SL U60087 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[6]), .Y(
        n27043) );
  NOR2xp33_ASAP7_75t_SRAM U60088 ( .A(n3080), .B(n1832), .Y(n76539) );
  INVx1_ASAP7_75t_SL U60089 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1[0]), .Y(n78248) );
  INVx1_ASAP7_75t_SL U60090 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[9]), .Y(n27516) );
  INVx1_ASAP7_75t_SL U60091 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[5]), .Y(
        n27042) );
  INVx1_ASAP7_75t_SL U60092 ( .A(or1200_cpu_or1200_except_n610), .Y(n76534) );
  NAND2xp5_ASAP7_75t_SL U60093 ( .A(or1200_cpu_or1200_except_n613), .B(n2098), 
        .Y(n63980) );
  INVxp67_ASAP7_75t_SL U60094 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[8]), .Y(n27517) );
  INVxp67_ASAP7_75t_SL U60095 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_31_), .Y(n69602) );
  INVx1_ASAP7_75t_SL U60096 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[4]), .Y(
        n27041) );
  INVx1_ASAP7_75t_SL U60097 ( .A(n3080), .Y(n77460) );
  INVx1_ASAP7_75t_SL U60098 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[7]), .Y(n27518) );
  INVx1_ASAP7_75t_SL U60099 ( .A(or1200_cpu_or1200_mult_mac_n259), .Y(n75126)
         );
  INVxp67_ASAP7_75t_SL U60100 ( .A(n2199), .Y(n60730) );
  INVx1_ASAP7_75t_SL U60101 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[19]), .Y(n78238) );
  INVx1_ASAP7_75t_SL U60102 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_), 
        .Y(n78361) );
  INVx1_ASAP7_75t_SL U60103 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[1]), .Y(n78229) );
  INVx1_ASAP7_75t_SL U60104 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[6]), .Y(n27519) );
  NAND2xp33_ASAP7_75t_SL U60105 ( .A(or1200_cpu_or1200_mult_mac_n147), .B(
        or1200_cpu_or1200_mult_mac_n293), .Y(n63309) );
  INVx1_ASAP7_75t_SL U60106 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[3]), .Y(
        n70152) );
  INVx1_ASAP7_75t_SL U60107 ( .A(or1200_cpu_or1200_except_n664), .Y(n75186) );
  INVx1_ASAP7_75t_SL U60108 ( .A(or1200_cpu_or1200_except_n607), .Y(n63954) );
  INVx1_ASAP7_75t_SL U60109 ( .A(n2122), .Y(n63953) );
  INVxp33_ASAP7_75t_SL U60110 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[7]), .Y(n73710) );
  INVxp33_ASAP7_75t_SL U60111 ( .A(n3088), .Y(n77491) );
  INVxp67_ASAP7_75t_SL U60112 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .Y(
        n70466) );
  INVxp33_ASAP7_75t_SL U60113 ( .A(n1428), .Y(n75691) );
  INVx1_ASAP7_75t_SL U60114 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[5]), .Y(n27520) );
  INVxp67_ASAP7_75t_SL U60115 ( .A(n957), .Y(n65195) );
  NAND2xp33_ASAP7_75t_SL U60116 ( .A(n2134), .B(or1200_cpu_or1200_except_n604), 
        .Y(n63761) );
  INVx1_ASAP7_75t_SL U60117 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_), .Y(
        n74691) );
  INVxp67_ASAP7_75t_SL U60118 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[4]), .Y(n70436) );
  NAND2xp5_ASAP7_75t_SL U60119 ( .A(dbg_stb_i), .B(or1200_du_dbg_ack), .Y(
        n4183) );
  INVxp67_ASAP7_75t_SL U60120 ( .A(or1200_cpu_or1200_mult_mac_n201), .Y(n75692) );
  INVx1_ASAP7_75t_SL U60121 ( .A(n3039), .Y(n63763) );
  INVx1_ASAP7_75t_SL U60122 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_11_), .Y(
        n74657) );
  INVx1_ASAP7_75t_SL U60123 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[3]), .Y(
        n27040) );
  INVx1_ASAP7_75t_SL U60124 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[4]), .Y(n27521) );
  INVx1_ASAP7_75t_SL U60125 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1[1]), .Y(n78249) );
  INVx1_ASAP7_75t_SL U60126 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_23_), .Y(
        n74295) );
  INVx1_ASAP7_75t_SL U60127 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[2]), .Y(
        n27039) );
  INVxp33_ASAP7_75t_SL U60128 ( .A(n1798), .Y(n75764) );
  INVx1_ASAP7_75t_SL U60129 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[3]), .Y(n27522) );
  INVx1_ASAP7_75t_SL U60130 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_25_), .Y(
        n72561) );
  INVx1_ASAP7_75t_SL U60131 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[5]), .Y(n69752) );
  INVxp67_ASAP7_75t_SL U60132 ( .A(n966), .Y(n65221) );
  INVxp67_ASAP7_75t_SL U60133 ( .A(or1200_cpu_or1200_mult_mac_n197), .Y(n75854) );
  INVx1_ASAP7_75t_SL U60134 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[2]), .Y(n27523) );
  INVx1_ASAP7_75t_SL U60135 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_8_), .Y(
        n74660) );
  INVx1_ASAP7_75t_SL U60136 ( .A(or1200_cpu_or1200_except_n667), .Y(n75640) );
  AND4x1_ASAP7_75t_SL U60137 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[24]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[27]), .C(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[28]), .D(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[29]), .Y(n74530) );
  INVx1_ASAP7_75t_SL U60138 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_26_), .Y(
        n74342) );
  NAND2xp33_ASAP7_75t_SL U60139 ( .A(or1200_cpu_or1200_except_n598), .B(n2160), 
        .Y(n63759) );
  INVxp67_ASAP7_75t_SL U60140 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[1]), .Y(n73679) );
  INVx1_ASAP7_75t_SL U60141 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[1]), .Y(n27524) );
  INVx1_ASAP7_75t_SL U60142 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[1]), .Y(
        n27038) );
  AND4x1_ASAP7_75t_SL U60143 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output1_23_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[30]), .C(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[26]), .D(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[25]), .Y(n74529) );
  INVxp67_ASAP7_75t_SL U60144 ( .A(or1200_cpu_or1200_mult_mac_n221), .Y(n69002) );
  INVx1_ASAP7_75t_SL U60145 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[0]), .Y(n27525) );
  INVxp67_ASAP7_75t_SL U60146 ( .A(n975), .Y(n65233) );
  INVx1_ASAP7_75t_SL U60147 ( .A(n2951), .Y(n75455) );
  NAND2xp33_ASAP7_75t_SL U60148 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_), .Y(n71529) );
  INVx1_ASAP7_75t_SL U60149 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_28_), .Y(
        n74356) );
  INVx1_ASAP7_75t_SL U60150 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[12]), .Y(n78235) );
  INVxp67_ASAP7_75t_SL U60151 ( .A(n984), .Y(n75149) );
  INVx1_ASAP7_75t_SL U60152 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_exp_10[6]), .Y(n27033) );
  INVx1_ASAP7_75t_SL U60153 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[2]), .Y(n73833) );
  INVx1_ASAP7_75t_SL U60154 ( .A(or1200_cpu_or1200_except_n670), .Y(n76925) );
  INVx1_ASAP7_75t_SL U60155 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[3]), .Y(n73828) );
  NAND2xp33_ASAP7_75t_SL U60156 ( .A(n2853), .B(n2427), .Y(n74525) );
  INVx1_ASAP7_75t_SL U60157 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_30_), .Y(
        n74314) );
  INVxp33_ASAP7_75t_SL U60158 ( .A(n2119), .Y(n59720) );
  INVx3_ASAP7_75t_SL U60159 ( .A(n3103), .Y(n59706) );
  INVx1_ASAP7_75t_SL U60160 ( .A(n1394), .Y(n76634) );
  INVx1_ASAP7_75t_SL U60161 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_9_), .Y(
        n74655) );
  NAND2xp33_ASAP7_75t_SL U60162 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_29_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_), .Y(n71536) );
  INVxp33_ASAP7_75t_SL U60163 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[14]), .Y(n73697) );
  INVx1_ASAP7_75t_SL U60164 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[0]), .Y(
        n27037) );
  INVx1_ASAP7_75t_SL U60165 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_32_), .Y(
        n74325) );
  NAND2xp5_ASAP7_75t_SL U60166 ( .A(n2450), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_4_), .Y(n70303) );
  INVxp33_ASAP7_75t_SL U60167 ( .A(or1200_cpu_esr[15]), .Y(n77144) );
  INVx1_ASAP7_75t_SL U60168 ( .A(n2577), .Y(n60225) );
  INVxp67_ASAP7_75t_SL U60169 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_30_), .Y(n69598) );
  INVx1_ASAP7_75t_SL U60170 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_1_), 
        .Y(n62046) );
  INVx1_ASAP7_75t_SL U60171 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_34_), .Y(
        n74347) );
  INVxp67_ASAP7_75t_SL U60172 ( .A(n993), .Y(n75163) );
  INVx1_ASAP7_75t_SL U60173 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_1_), .Y(
        n71656) );
  INVx1_ASAP7_75t_SL U60174 ( .A(n3117), .Y(n76558) );
  INVx1_ASAP7_75t_SL U60175 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_11_), .Y(n65245) );
  INVx1_ASAP7_75t_SL U60176 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[23]), .Y(n27502) );
  INVx1_ASAP7_75t_SL U60177 ( .A(n1414), .Y(n76855) );
  NAND2xp5_ASAP7_75t_SL U60178 ( .A(or1200_cpu_or1200_mult_mac_n345), .B(
        or1200_cpu_or1200_mult_mac_n199), .Y(n75008) );
  INVxp33_ASAP7_75t_SL U60179 ( .A(or1200_cpu_or1200_mult_mac_n151), .Y(n63314) );
  INVxp67_ASAP7_75t_SL U60180 ( .A(n3337), .Y(n74733) );
  INVx1_ASAP7_75t_SL U60181 ( .A(or1200_cpu_or1200_except_n586), .Y(n76574) );
  INVx1_ASAP7_75t_SL U60182 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_13_), .Y(n65249) );
  INVx1_ASAP7_75t_SL U60183 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[22]), .Y(n27503) );
  NAND2xp5_ASAP7_75t_SL U60184 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_0_), 
        .Y(n71645) );
  INVxp67_ASAP7_75t_SL U60185 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_), .Y(n78380) );
  NAND2xp33_ASAP7_75t_SL U60186 ( .A(n2685), .B(or1200_cpu_or1200_except_n643), 
        .Y(n75540) );
  INVx1_ASAP7_75t_SL U60187 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[7]), .Y(n69776) );
  INVx1_ASAP7_75t_SL U60188 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_15_), .Y(n65256) );
  INVx1_ASAP7_75t_SL U60189 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[21]), .Y(n27504) );
  INVxp33_ASAP7_75t_SL U60190 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_), .Y(
        n74643) );
  INVxp33_ASAP7_75t_SL U60191 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_7_), .Y(
        n71669) );
  INVx1_ASAP7_75t_SL U60192 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_17_), .Y(n65371) );
  INVx1_ASAP7_75t_SL U60193 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[20]), .Y(n27505) );
  INVx1_ASAP7_75t_SL U60194 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_16_), .Y(
        n74654) );
  INVx1_ASAP7_75t_SL U60195 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_19_), .Y(n65342) );
  INVx1_ASAP7_75t_SL U60196 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[19]), .Y(n27506) );
  INVx1_ASAP7_75t_SL U60197 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_15_), .Y(
        n74664) );
  NAND2xp5_ASAP7_75t_SL U60198 ( .A(n2678), .B(or1200_cpu_or1200_except_n640), 
        .Y(n65201) );
  NAND2xp33_ASAP7_75t_SL U60199 ( .A(or1200_cpu_or1200_mult_mac_n317), .B(
        or1200_cpu_or1200_mult_mac_n171), .Y(n63535) );
  INVx1_ASAP7_75t_SL U60200 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_21_), .Y(n65361) );
  INVx1_ASAP7_75t_SL U60201 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_22_), 
        .Y(n72309) );
  INVx1_ASAP7_75t_SL U60202 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[18]), .Y(n27507) );
  INVxp67_ASAP7_75t_SL U60203 ( .A(n903), .Y(n74969) );
  INVx1_ASAP7_75t_SL U60204 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[17]), .Y(n27508) );
  INVxp67_ASAP7_75t_SL U60205 ( .A(or1200_cpu_or1200_except_n652), .Y(n65222)
         );
  INVxp67_ASAP7_75t_SL U60206 ( .A(n1978), .Y(n61469) );
  INVxp67_ASAP7_75t_SL U60207 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[5]), .Y(
        n73886) );
  INVxp67_ASAP7_75t_SL U60208 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_), 
        .Y(n72348) );
  INVxp33_ASAP7_75t_SL U60209 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_), .Y(
        n74672) );
  INVxp33_ASAP7_75t_SL U60210 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .Y(
        n70297) );
  INVx1_ASAP7_75t_SL U60211 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[6]), .Y(
        n73893) );
  INVx1_ASAP7_75t_SL U60212 ( .A(n1973), .Y(n76870) );
  INVxp67_ASAP7_75t_SL U60213 ( .A(n912), .Y(n64014) );
  INVx1_ASAP7_75t_SL U60214 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[16]), .Y(n27509) );
  NAND2xp5_ASAP7_75t_SL U60215 ( .A(n1582), .B(n1564), .Y(n65261) );
  INVx1_ASAP7_75t_SL U60216 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[7]), .Y(
        n27044) );
  INVx1_ASAP7_75t_SL U60217 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[3]), .Y(n73613)
         );
  INVx1_ASAP7_75t_SL U60218 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_4_), 
        .Y(n74301) );
  INVxp33_ASAP7_75t_SL U60219 ( .A(n1117), .Y(n75531) );
  INVxp67_ASAP7_75t_SL U60220 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_6_), 
        .Y(n73858) );
  INVx1_ASAP7_75t_SL U60221 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_8_), 
        .Y(n74359) );
  INVx1_ASAP7_75t_SL U60222 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[5]), .Y(n73708) );
  INVx1_ASAP7_75t_SL U60223 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_11_), 
        .Y(n74321) );
  INVx1_ASAP7_75t_SL U60224 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[10]), .Y(n27515) );
  INVx1_ASAP7_75t_SL U60225 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_13_), 
        .Y(n74339) );
  INVx1_ASAP7_75t_SL U60226 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[11]), .Y(n27514) );
  INVx1_ASAP7_75t_SL U60227 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[8]), .Y(
        n27045) );
  INVx1_ASAP7_75t_SL U60228 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_15_), 
        .Y(n74386) );
  INVxp67_ASAP7_75t_SL U60229 ( .A(n948), .Y(n75545) );
  INVx1_ASAP7_75t_SL U60230 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_exp_10_o[9]), .Y(
        n27046) );
  INVx1_ASAP7_75t_SL U60231 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_17_), 
        .Y(n74404) );
  NAND2xp5_ASAP7_75t_SL U60232 ( .A(or1200_cpu_or1200_except_n622), .B(n2637), 
        .Y(n64000) );
  INVx1_ASAP7_75t_SL U60233 ( .A(n2193), .Y(n76652) );
  INVx1_ASAP7_75t_SL U60234 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[12]), .Y(n27513) );
  INVx1_ASAP7_75t_SL U60235 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_19_), 
        .Y(n74311) );
  INVxp67_ASAP7_75t_SL U60236 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_output_o_31_), .Y(
        n28158) );
  INVxp67_ASAP7_75t_SL U60237 ( .A(n939), .Y(n64266) );
  INVx1_ASAP7_75t_SL U60238 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_21_), 
        .Y(n74425) );
  INVx1_ASAP7_75t_SL U60239 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[13]), .Y(n27512) );
  INVx1_ASAP7_75t_SL U60240 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_23_), 
        .Y(n74226) );
  INVx1_ASAP7_75t_SL U60241 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_start_i), 
        .Y(n78245) );
  INVx1_ASAP7_75t_SL U60242 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_22_), .Y(
        n74294) );
  INVxp67_ASAP7_75t_SL U60243 ( .A(n930), .Y(n75420) );
  INVx1_ASAP7_75t_SL U60244 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_), 
        .Y(n78379) );
  INVx2_ASAP7_75t_SL U60245 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_1_), .Y(n78437) );
  INVx1_ASAP7_75t_SL U60246 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_), 
        .Y(n78376) );
  INVxp67_ASAP7_75t_SL U60247 ( .A(or1200_cpu_or1200_except_n658), .Y(n75153)
         );
  INVx1_ASAP7_75t_SL U60248 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[11]), .Y(n78234) );
  NAND2xp5_ASAP7_75t_SL U60249 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_1_), .B(
        or1200_cpu_or1200_fpu_fpu_op_r_0_), .Y(n74741) );
  INVxp67_ASAP7_75t_SL U60250 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[3]), .Y(
        n73877) );
  INVx1_ASAP7_75t_SL U60251 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[14]), .Y(n27511) );
  INVx1_ASAP7_75t_SL U60252 ( .A(n2837), .Y(n77285) );
  INVxp67_ASAP7_75t_SL U60253 ( .A(n921), .Y(n64164) );
  INVxp67_ASAP7_75t_SL U60254 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_mul_fract_48[47]), .Y(n28207)
         );
  INVx1_ASAP7_75t_SL U60255 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[15]), .Y(n27510) );
  INVxp67_ASAP7_75t_SL U60256 ( .A(or1200_cpu_or1200_except_n655), .Y(n65234)
         );
  INVxp67_ASAP7_75t_SL U60257 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[28]), .Y(n78196) );
  INVx6_ASAP7_75t_SL U60258 ( .A(n59558), .Y(n57214) );
  INVx1_ASAP7_75t_SL U60259 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_4_), .Y(n74844)
         );
  INVx1_ASAP7_75t_SL U60260 ( .A(or1200_cpu_or1200_mult_mac_n42), .Y(n76045)
         );
  INVx1_ASAP7_75t_SL U60261 ( .A(or1200_cpu_or1200_mult_mac_n40), .Y(n76058)
         );
  INVx1_ASAP7_75t_SL U60262 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[2]), .Y(n27447) );
  INVx1_ASAP7_75t_SL U60263 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[3]), .Y(n69731) );
  INVx1_ASAP7_75t_SL U60264 ( .A(or1200_cpu_or1200_mult_mac_n54), .Y(n76005)
         );
  INVx1_ASAP7_75t_SL U60265 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[1]), .Y(n78330)
         );
  INVxp67_ASAP7_75t_SL U60266 ( .A(or1200_cpu_or1200_mult_mac_n52), .Y(n75928)
         );
  INVxp33_ASAP7_75t_SL U60267 ( .A(n2630), .Y(n62471) );
  INVxp33_ASAP7_75t_SL U60268 ( .A(n1936), .Y(n75532) );
  INVx1_ASAP7_75t_SL U60269 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[13]), .Y(n27477) );
  INVx1_ASAP7_75t_SL U60270 ( .A(or1200_cpu_or1200_mult_mac_n58), .Y(n75991)
         );
  INVxp33_ASAP7_75t_SL U60271 ( .A(n2079), .Y(n77927) );
  INVxp67_ASAP7_75t_SL U60272 ( .A(or1200_cpu_or1200_mult_mac_n303), .Y(n63411) );
  INVx1_ASAP7_75t_SL U60273 ( .A(or1200_cpu_or1200_mult_mac_n62), .Y(n75980)
         );
  INVxp67_ASAP7_75t_SL U60274 ( .A(ex_insn[22]), .Y(n77564) );
  INVxp67_ASAP7_75t_SL U60275 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_6_), .Y(
        n74659) );
  INVx1_ASAP7_75t_SL U60276 ( .A(or1200_cpu_or1200_mult_mac_n36), .Y(n75909)
         );
  INVx1_ASAP7_75t_SL U60277 ( .A(or1200_cpu_or1200_mult_mac_n46), .Y(n75902)
         );
  INVx1_ASAP7_75t_SL U60278 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[5]), .Y(n78336)
         );
  INVx1_ASAP7_75t_SL U60279 ( .A(or1200_cpu_or1200_mult_mac_n8), .Y(n75963) );
  INVx1_ASAP7_75t_SL U60280 ( .A(id_insn_22_), .Y(n62469) );
  INVx1_ASAP7_75t_SL U60281 ( .A(or1200_cpu_or1200_mult_mac_n249), .Y(n69256)
         );
  INVx1_ASAP7_75t_SL U60282 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .Y(n72313) );
  INVx1_ASAP7_75t_SL U60283 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[19]), .Y(n73774) );
  INVx1_ASAP7_75t_SL U60284 ( .A(or1200_cpu_or1200_mult_mac_n2), .Y(n75968) );
  INVx1_ASAP7_75t_SL U60285 ( .A(or1200_cpu_or1200_mult_mac_n4), .Y(n76194) );
  NAND2xp33_ASAP7_75t_SL U60286 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_sign), .Y(n74159) );
  INVxp33_ASAP7_75t_SL U60287 ( .A(or1200_cpu_or1200_except_n292), .Y(n74944)
         );
  INVxp67_ASAP7_75t_SL U60288 ( .A(n2093), .Y(n77554) );
  INVxp33_ASAP7_75t_SL U60289 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_3_), .Y(n69588) );
  INVx1_ASAP7_75t_SL U60290 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[8]), .Y(n78342)
         );
  INVxp67_ASAP7_75t_SL U60291 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_6_), .Y(
        n74794) );
  INVxp67_ASAP7_75t_SL U60292 ( .A(n1826), .Y(n62318) );
  NAND2xp5_ASAP7_75t_SL U60293 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_infa_f_r), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_expa_ff), .Y(n4747) );
  INVxp67_ASAP7_75t_SL U60294 ( .A(n2184), .Y(n77532) );
  INVx1_ASAP7_75t_SL U60295 ( .A(n2397), .Y(n74674) );
  INVx1_ASAP7_75t_SL U60296 ( .A(n2098), .Y(n77381) );
  NOR3xp33_ASAP7_75t_SRAM U60297 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_4_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_7_), .Y(
        n74482) );
  INVxp67_ASAP7_75t_SL U60298 ( .A(n1945), .Y(n62317) );
  INVx1_ASAP7_75t_SL U60299 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_2_), 
        .Y(n72365) );
  INVx1_ASAP7_75t_SL U60300 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .Y(
        n73618) );
  INVxp67_ASAP7_75t_SL U60301 ( .A(n2103), .Y(n77550) );
  INVxp67_ASAP7_75t_SL U60302 ( .A(or1200_cpu_or1200_mult_mac_n261), .Y(n75822) );
  NAND2xp5_ASAP7_75t_SL U60303 ( .A(or1200_cpu_or1200_mult_mac_n331), .B(
        or1200_cpu_or1200_mult_mac_n185), .Y(n65145) );
  INVx1_ASAP7_75t_SL U60304 ( .A(or1200_cpu_or1200_fpu_fpu_conv_shr[0]), .Y(
        n27531) );
  INVx1_ASAP7_75t_SL U60305 ( .A(or1200_cpu_or1200_fpu_fpu_conv_shr[1]), .Y(
        n27532) );
  INVx1_ASAP7_75t_SL U60306 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[9]), .Y(n78344)
         );
  INVx1_ASAP7_75t_SL U60307 ( .A(or1200_cpu_or1200_fpu_fpu_conv_shr[2]), .Y(
        n27533) );
  INVx1_ASAP7_75t_SL U60308 ( .A(or1200_cpu_or1200_fpu_fpu_conv_shr[3]), .Y(
        n27534) );
  INVx1_ASAP7_75t_SL U60309 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[7]), .Y(n78232) );
  INVxp67_ASAP7_75t_SL U60310 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[14]), .Y(n70334) );
  INVx1_ASAP7_75t_SL U60311 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[11]), .Y(n78346) );
  INVxp33_ASAP7_75t_SL U60312 ( .A(or1200_cpu_or1200_mult_mac_n20), .Y(n76146)
         );
  INVx1_ASAP7_75t_SL U60313 ( .A(or1200_cpu_or1200_fpu_fpu_conv_shr[4]), .Y(
        n27535) );
  INVx1_ASAP7_75t_SL U60314 ( .A(or1200_cpu_or1200_fpu_fpu_conv_shr[5]), .Y(
        n27536) );
  INVx1_ASAP7_75t_SL U60315 ( .A(n2172), .Y(n74790) );
  INVx1_ASAP7_75t_SL U60316 ( .A(or1200_cpu_or1200_except_n278), .Y(n76866) );
  INVx1_ASAP7_75t_SL U60317 ( .A(n58422), .Y(n57216) );
  INVx1_ASAP7_75t_SL U60318 ( .A(n2110), .Y(n61161) );
  INVxp67_ASAP7_75t_SL U60319 ( .A(or1200_cpu_or1200_mult_mac_n26), .Y(n76112)
         );
  INVxp67_ASAP7_75t_SL U60320 ( .A(or1200_cpu_or1200_mult_mac_n351), .Y(n68830) );
  INVxp33_ASAP7_75t_SL U60321 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_6_), .Y(
        n74231) );
  INVxp67_ASAP7_75t_SL U60322 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .Y(
        n71899) );
  INVx1_ASAP7_75t_SL U60323 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[21]), .Y(n73753) );
  INVxp67_ASAP7_75t_SL U60324 ( .A(n2115), .Y(n77547) );
  INVx1_ASAP7_75t_SL U60325 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[23]), .Y(n73728) );
  INVxp67_ASAP7_75t_SL U60326 ( .A(n2165), .Y(n77535) );
  INVx1_ASAP7_75t_SL U60327 ( .A(n2552), .Y(n75888) );
  INVx1_ASAP7_75t_SL U60328 ( .A(or1200_cpu_or1200_mult_mac_n353), .Y(n68847)
         );
  INVx1_ASAP7_75t_SL U60329 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[12]), .Y(n78350) );
  INVx1_ASAP7_75t_SL U60330 ( .A(n2160), .Y(n74793) );
  NAND2xp5_ASAP7_75t_SL U60331 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[0]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[1]), .Y(
        n58622) );
  INVxp67_ASAP7_75t_SL U60332 ( .A(n2127), .Y(n77544) );
  INVxp67_ASAP7_75t_SL U60333 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[1]), .Y(
        n73617) );
  INVx1_ASAP7_75t_SL U60334 ( .A(or1200_cpu_or1200_except_n530), .Y(n75433) );
  INVx1_ASAP7_75t_SL U60335 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .Y(
        n73752) );
  INVx1_ASAP7_75t_SL U60336 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[14]), .Y(n78427) );
  INVx1_ASAP7_75t_SL U60337 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]), .Y(n78426) );
  INVx1_ASAP7_75t_SL U60338 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[23]), .Y(n78241) );
  INVxp67_ASAP7_75t_SL U60339 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_5_), .Y(
        n74791) );
  INVx1_ASAP7_75t_SL U60340 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .Y(
        n72241) );
  INVx1_ASAP7_75t_SL U60341 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[15]), .Y(n78236) );
  INVx1_ASAP7_75t_SL U60342 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[17]), .Y(n78424) );
  INVxp67_ASAP7_75t_SL U60343 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[0]), .Y(
        n73641) );
  INVxp33_ASAP7_75t_SL U60344 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .Y(
        n73623) );
  INVx1_ASAP7_75t_SL U60345 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[18]), .Y(n78354) );
  INVxp67_ASAP7_75t_SL U60346 ( .A(n2153), .Y(n77538) );
  INVx1_ASAP7_75t_SL U60347 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[6]), .Y(n78231) );
  INVxp67_ASAP7_75t_SL U60348 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_mul_output[3]), .Y(n74377)
         );
  OAI21xp33_ASAP7_75t_SL U60349 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[7]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[7]), .Y(
        n70192) );
  NAND2xp33_ASAP7_75t_SL U60350 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .Y(
        n72266) );
  INVxp67_ASAP7_75t_SL U60351 ( .A(n2139), .Y(n77541) );
  INVx1_ASAP7_75t_SL U60352 ( .A(n2148), .Y(n74796) );
  INVx1_ASAP7_75t_SL U60353 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .Y(
        n71983) );
  INVx1_ASAP7_75t_SL U60354 ( .A(n58423), .Y(n57217) );
  INVx1_ASAP7_75t_SL U60355 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[20]), .Y(n78368) );
  INVxp67_ASAP7_75t_SL U60356 ( .A(or1200_cpu_or1200_mult_mac_n64), .Y(n75978)
         );
  NAND2xp5_ASAP7_75t_SL U60357 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[7]), .Y(
        n70206) );
  INVxp67_ASAP7_75t_SL U60358 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[7]), .Y(
        n70190) );
  INVxp67_ASAP7_75t_SL U60359 ( .A(n1735), .Y(n65237) );
  INVx1_ASAP7_75t_SL U60360 ( .A(n2517), .Y(n69337) );
  INVxp67_ASAP7_75t_SL U60361 ( .A(or1200_cpu_or1200_except_n258), .Y(n77216)
         );
  INVx1_ASAP7_75t_SL U60362 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_2_), 
        .Y(n62054) );
  INVx1_ASAP7_75t_SL U60363 ( .A(n3419), .Y(n77770) );
  NOR2xp33_ASAP7_75t_SRAM U60364 ( .A(or1200_dc_top_tag_v), .B(n3088), .Y(
        n77478) );
  INVxp67_ASAP7_75t_SL U60365 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[4]), .Y(n69597) );
  INVx1_ASAP7_75t_SL U60366 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_), 
        .Y(n72163) );
  INVx1_ASAP7_75t_SL U60367 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_38_), .Y(
        n74309) );
  INVx1_ASAP7_75t_SL U60368 ( .A(n2410), .Y(n77234) );
  NAND2xp33_ASAP7_75t_SL U60369 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[5]), .Y(
        n70183) );
  NAND2xp5_ASAP7_75t_SL U60370 ( .A(n3309), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .Y(
        n73817) );
  INVx1_ASAP7_75t_SL U60371 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[21]), .Y(n78366) );
  INVx1_ASAP7_75t_SL U60372 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[20]), .Y(n78239) );
  INVx1_ASAP7_75t_SL U60373 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_24_), 
        .Y(n72253) );
  INVx1_ASAP7_75t_SL U60374 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_state), .Y(
        n62047) );
  NAND2xp5_ASAP7_75t_SL U60375 ( .A(or1200_cpu_or1200_mult_mac_n205), .B(
        or1200_cpu_or1200_mult_mac_n351), .Y(n68885) );
  INVx1_ASAP7_75t_SL U60376 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_), 
        .Y(n72212) );
  INVx1_ASAP7_75t_SL U60377 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_25_), 
        .Y(n72234) );
  NAND2xp5_ASAP7_75t_SL U60378 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_0_), .B(or1200_cpu_or1200_fpu_fpu_arith_s_count_1_), .Y(n62053) );
  INVxp67_ASAP7_75t_SL U60379 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[24]), .Y(n78242) );
  INVxp33_ASAP7_75t_SL U60380 ( .A(n2026), .Y(n77924) );
  NAND2xp5_ASAP7_75t_SL U60381 ( .A(n3109), .B(n3107), .Y(n78165) );
  INVx1_ASAP7_75t_SL U60382 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_40_), .Y(
        n74414) );
  NAND2xp5_ASAP7_75t_SL U60383 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .Y(
        n72112) );
  BUFx4f_ASAP7_75t_SL U60384 ( .A(n1802), .Y(n57500) );
  INVxp67_ASAP7_75t_SL U60385 ( .A(n1002), .Y(n75185) );
  NAND2xp33_ASAP7_75t_SL U60386 ( .A(or1200_cpu_or1200_mult_mac_n145), .B(
        or1200_cpu_or1200_mult_mac_n291), .Y(n63308) );
  INVx1_ASAP7_75t_SL U60387 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_42_), .Y(
        n74432) );
  INVx1_ASAP7_75t_SL U60388 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_0_), 
        .Y(n62048) );
  INVxp67_ASAP7_75t_SL U60389 ( .A(n3092), .Y(n78163) );
  INVx1_ASAP7_75t_SL U60390 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .Y(
        n72399) );
  INVx1_ASAP7_75t_SL U60391 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[5]), .Y(n27472) );
  INVx1_ASAP7_75t_SL U60392 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_44_), .Y(
        n74222) );
  INVx1_ASAP7_75t_SL U60393 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_2_), .Y(
        n74685) );
  INVx1_ASAP7_75t_SL U60394 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[2]), .Y(n69724) );
  INVx1_ASAP7_75t_SL U60395 ( .A(n3390), .Y(n62052) );
  INVxp67_ASAP7_75t_SL U60396 ( .A(n1020), .Y(n76917) );
  INVxp67_ASAP7_75t_SL U60397 ( .A(n2031), .Y(n77559) );
  INVx1_ASAP7_75t_SL U60398 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_13_), .Y(n77196)
         );
  INVx1_ASAP7_75t_SL U60399 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[7]), .Y(n73581)
         );
  INVxp67_ASAP7_75t_SL U60400 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_2_), .Y(n69594) );
  INVxp67_ASAP7_75t_SL U60401 ( .A(or1200_cpu_or1200_mult_mac_n165), .Y(n63452) );
  INVxp67_ASAP7_75t_SL U60402 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_3_), .Y(
        n74677) );
  INVx1_ASAP7_75t_SL U60403 ( .A(or1200_cpu_or1200_mult_mac_n38), .Y(n76065)
         );
  INVxp67_ASAP7_75t_SL U60404 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[27]), .Y(n78195) );
  INVx1_ASAP7_75t_SL U60405 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[21]), .Y(n78240) );
  INVxp67_ASAP7_75t_SL U60406 ( .A(n2067), .Y(n77557) );
  INVxp67_ASAP7_75t_SL U60407 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_29_), .Y(n69584) );
  INVx1_ASAP7_75t_SL U60408 ( .A(or1200_cpu_or1200_mult_mac_n34), .Y(n75935)
         );
  INVxp67_ASAP7_75t_SL U60409 ( .A(or1200_cpu_or1200_mult_mac_n269), .Y(n63263) );
  INVxp67_ASAP7_75t_SL U60410 ( .A(n2062), .Y(n77926) );
  INVxp33_ASAP7_75t_SL U60411 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_1_), .Y(n69590) );
  INVx1_ASAP7_75t_SL U60412 ( .A(or1200_cpu_or1200_mult_mac_n28), .Y(n76106)
         );
  INVx1_ASAP7_75t_SL U60413 ( .A(or1200_cpu_or1200_mult_mac_n271), .Y(n63265)
         );
  INVx1_ASAP7_75t_SL U60414 ( .A(or1200_cpu_or1200_mult_mac_n22), .Y(n76129)
         );
  INVxp33_ASAP7_75t_SL U60415 ( .A(n1938), .Y(n62408) );
  INVx1_ASAP7_75t_SL U60416 ( .A(n2054), .Y(n76537) );
  INVx1_ASAP7_75t_SL U60417 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_7_), .Y(n76943)
         );
  INVxp67_ASAP7_75t_SL U60418 ( .A(or1200_cpu_or1200_mult_mac_n233), .Y(n69124) );
  INVxp33_ASAP7_75t_SL U60419 ( .A(or1200_cpu_or1200_except_n286), .Y(n74929)
         );
  INVxp67_ASAP7_75t_SL U60420 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[22]), .Y(n70262) );
  INVx1_ASAP7_75t_SL U60421 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[8]), .Y(n27448) );
  INVx1_ASAP7_75t_SL U60422 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_1_), .Y(
        n74681) );
  INVx1_ASAP7_75t_SL U60423 ( .A(or1200_cpu_or1200_mult_mac_n169), .Y(n63485)
         );
  INVx1_ASAP7_75t_SL U60424 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[6]), .Y(
        n70189) );
  INVx1_ASAP7_75t_SL U60425 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_8_), .Y(n76944)
         );
  INVx1_ASAP7_75t_SL U60426 ( .A(n2440), .Y(n74644) );
  INVx1_ASAP7_75t_SL U60427 ( .A(or1200_cpu_or1200_mult_mac_n10), .Y(n75957)
         );
  INVx1_ASAP7_75t_SL U60428 ( .A(n3321), .Y(n73642) );
  NAND2xp5_ASAP7_75t_SL U60429 ( .A(or1200_cpu_or1200_mult_mac_n329), .B(
        or1200_cpu_or1200_mult_mac_n183), .Y(n65131) );
  INVxp67_ASAP7_75t_SL U60430 ( .A(n2050), .Y(n77562) );
  NAND2xp33_ASAP7_75t_SL U60431 ( .A(or1200_cpu_or1200_mult_mac_n335), .B(
        or1200_cpu_or1200_mult_mac_n189), .Y(n65176) );
  INVxp67_ASAP7_75t_SL U60432 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_9_), .Y(n74880)
         );
  INVxp67_ASAP7_75t_SL U60433 ( .A(or1200_cpu_or1200_mult_mac_n143), .Y(n63272) );
  INVxp67_ASAP7_75t_SL U60434 ( .A(n2045), .Y(n77925) );
  INVx1_ASAP7_75t_SL U60435 ( .A(or1200_cpu_or1200_except_n434), .Y(n77018) );
  INVxp67_ASAP7_75t_SL U60436 ( .A(n3327), .Y(n73695) );
  NAND2xp33_ASAP7_75t_SL U60437 ( .A(or1200_cpu_or1200_mult_mac_n325), .B(
        or1200_cpu_or1200_mult_mac_n179), .Y(n65077) );
  NAND2xp5_ASAP7_75t_SL U60438 ( .A(or1200_cpu_or1200_mult_mac_n207), .B(
        or1200_cpu_or1200_mult_mac_n353), .Y(n68886) );
  INVx1_ASAP7_75t_SL U60439 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[16]), .Y(n27495) );
  NAND2xp33_ASAP7_75t_SL U60440 ( .A(or1200_cpu_or1200_mult_mac_n143), .B(
        or1200_cpu_or1200_mult_mac_n289), .Y(n63276) );
  INVx1_ASAP7_75t_SL U60441 ( .A(n3082), .Y(n61317) );
  INVxp67_ASAP7_75t_SL U60442 ( .A(n2755), .Y(n69332) );
  INVx1_ASAP7_75t_SL U60443 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_36_), .Y(
        n74391) );
  INVx1_ASAP7_75t_SL U60444 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[3]), .Y(n78230) );
  INVxp67_ASAP7_75t_SL U60445 ( .A(or1200_cpu_or1200_except_n640), .Y(n75421)
         );
  INVxp67_ASAP7_75t_SL U60446 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_37_), .Y(n69631) );
  INVx1_ASAP7_75t_SL U60447 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_5_), .Y(
        n74237) );
  INVxp67_ASAP7_75t_SL U60448 ( .A(or1200_cpu_or1200_except_n628), .Y(n64011)
         );
  INVx1_ASAP7_75t_SL U60449 ( .A(n2335), .Y(n70327) );
  NAND2xp33_ASAP7_75t_SL U60450 ( .A(or1200_cpu_or1200_mult_mac_n299), .B(
        or1200_cpu_or1200_mult_mac_n153), .Y(n63376) );
  INVx1_ASAP7_75t_SL U60451 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_), .Y(
        n70552) );
  INVx1_ASAP7_75t_SL U60452 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_), 
        .Y(n72318) );
  INVxp67_ASAP7_75t_SL U60453 ( .A(n1851), .Y(n60286) );
  INVx1_ASAP7_75t_SL U60454 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_), 
        .Y(n72132) );
  INVx1_ASAP7_75t_SL U60455 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_8_), .Y(n69788) );
  INVx1_ASAP7_75t_SL U60456 ( .A(n1123), .Y(n75646) );
  INVxp67_ASAP7_75t_SL U60457 ( .A(n843), .Y(n61587) );
  INVx1_ASAP7_75t_SL U60458 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_12_), .Y(
        n74646) );
  INVx1_ASAP7_75t_SL U60459 ( .A(or1200_cpu_or1200_except_n613), .Y(n63949) );
  NAND2xp33_ASAP7_75t_SL U60460 ( .A(or1200_cpu_or1200_mult_mac_n295), .B(
        or1200_cpu_or1200_mult_mac_n149), .Y(n63339) );
  INVx1_ASAP7_75t_SL U60461 ( .A(or1200_cpu_or1200_mult_mac_n235), .Y(n77042)
         );
  INVxp67_ASAP7_75t_SL U60462 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_5_), .Y(
        n70546) );
  INVxp67_ASAP7_75t_SL U60463 ( .A(n1064), .Y(n63739) );
  INVxp67_ASAP7_75t_SL U60464 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_2_), .Y(
        n71644) );
  INVxp67_ASAP7_75t_SL U60465 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_output_o[29]), .Y(n78209) );
  INVx1_ASAP7_75t_SL U60466 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_37_), 
        .Y(n72054) );
  INVxp67_ASAP7_75t_SL U60467 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_35_), .Y(n69621) );
  INVxp67_ASAP7_75t_SL U60468 ( .A(or1200_cpu_or1200_except_n637), .Y(n64165)
         );
  INVx1_ASAP7_75t_SL U60469 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[0]), .Y(
        n70107) );
  INVx1_ASAP7_75t_SL U60470 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_32_), 
        .Y(n72154) );
  INVxp67_ASAP7_75t_SL U60471 ( .A(n1430), .Y(n75406) );
  INVxp67_ASAP7_75t_SL U60472 ( .A(or1200_cpu_or1200_except_n631), .Y(n74970)
         );
  INVx1_ASAP7_75t_SL U60473 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_), 
        .Y(n71984) );
  INVxp67_ASAP7_75t_SL U60474 ( .A(or1200_cpu_or1200_except_n622), .Y(n63998)
         );
  INVx1_ASAP7_75t_SL U60475 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[8]), .Y(n69787) );
  INVxp67_ASAP7_75t_SL U60476 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[14]), .Y(n69650) );
  NAND2xp33_ASAP7_75t_SL U60477 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_3_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_7_), .Y(
        n72587) );
  INVx1_ASAP7_75t_SL U60478 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[17]), .Y(n78237) );
  INVxp33_ASAP7_75t_SL U60479 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[0]), .Y(
        n70105) );
  INVx1_ASAP7_75t_SL U60480 ( .A(or1200_cpu_or1200_mult_mac_n209), .Y(n68849)
         );
  INVx1_ASAP7_75t_SL U60481 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_36_), 
        .Y(n72079) );
  INVx1_ASAP7_75t_SL U60482 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_7_), .Y(
        n70439) );
  NAND2xp5_ASAP7_75t_SL U60483 ( .A(or1200_cpu_or1200_mult_mac_n315), .B(
        or1200_cpu_or1200_mult_mac_n169), .Y(n63534) );
  INVx1_ASAP7_75t_SL U60484 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .Y(
        n72499) );
  INVxp67_ASAP7_75t_SL U60485 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_0_), .Y(
        n71646) );
  INVxp67_ASAP7_75t_SL U60486 ( .A(n837), .Y(n63748) );
  INVx1_ASAP7_75t_SL U60487 ( .A(or1200_cpu_or1200_except_n272), .Y(n76623) );
  NAND2xp33_ASAP7_75t_SL U60488 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_), .Y(n71525) );
  INVx1_ASAP7_75t_SL U60489 ( .A(or1200_cpu_or1200_mult_mac_n213), .Y(n68892)
         );
  INVxp67_ASAP7_75t_SL U60490 ( .A(or1200_cpu_or1200_mult_mac_n199), .Y(n75219) );
  INVx1_ASAP7_75t_SL U60491 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_), 
        .Y(n72346) );
  INVx1_ASAP7_75t_SL U60492 ( .A(n2963), .Y(n75626) );
  INVxp67_ASAP7_75t_SL U60493 ( .A(n1097), .Y(n63698) );
  INVx1_ASAP7_75t_SL U60494 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_4_), .Y(
        n71692) );
  INVx1_ASAP7_75t_SL U60495 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .Y(n72316) );
  INVxp67_ASAP7_75t_SL U60496 ( .A(n1086), .Y(n61278) );
  INVx1_ASAP7_75t_SL U60497 ( .A(n2850), .Y(n77156) );
  INVx1_ASAP7_75t_SL U60498 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_2_), .Y(
        n71643) );
  INVxp67_ASAP7_75t_SL U60499 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[9]), .Y(n69620) );
  INVx1_ASAP7_75t_SL U60500 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_), 
        .Y(n71993) );
  INVx1_ASAP7_75t_SL U60501 ( .A(n2442), .Y(n74656) );
  INVxp67_ASAP7_75t_SL U60502 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_1_), .Y(
        n71647) );
  INVxp33_ASAP7_75t_SL U60503 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_14_), .Y(n69663) );
  INVx1_ASAP7_75t_SL U60504 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_), 
        .Y(n72263) );
  NAND2xp5_ASAP7_75t_SL U60505 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_6_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_7_), .Y(
        n72590) );
  INVxp67_ASAP7_75t_SL U60506 ( .A(n1510), .Y(n76674) );
  NAND2xp33_ASAP7_75t_SL U60507 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_), .Y(n71513) );
  INVx1_ASAP7_75t_SL U60508 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_13_), 
        .Y(n72351) );
  INVxp67_ASAP7_75t_SL U60509 ( .A(or1200_cpu_or1200_except_n625), .Y(n64006)
         );
  INVx1_ASAP7_75t_SL U60510 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_1_), .Y(
        n74063) );
  INVx1_ASAP7_75t_SL U60511 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n131), .Y(n72565) );
  INVxp67_ASAP7_75t_SL U60512 ( .A(n2974), .Y(n60432) );
  INVxp33_ASAP7_75t_SL U60513 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_3_), .Y(
        n71659) );
  INVx1_ASAP7_75t_SL U60514 ( .A(n1958), .Y(n76626) );
  INVx1_ASAP7_75t_SL U60515 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_35_), 
        .Y(n72080) );
  INVx1_ASAP7_75t_SL U60516 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_4_), .Y(n74809) );
  INVxp67_ASAP7_75t_SL U60517 ( .A(or1200_cpu_or1200_except_n634), .Y(n64015)
         );
  INVx1_ASAP7_75t_SL U60518 ( .A(or1200_cpu_or1200_mult_mac_n215), .Y(n68932)
         );
  INVx1_ASAP7_75t_SL U60519 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .Y(n71863) );
  NAND2xp5_ASAP7_75t_SL U60520 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_5_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_6_), .Y(
        n72574) );
  INVxp67_ASAP7_75t_SL U60521 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[1]), .Y(
        n70125) );
  INVx1_ASAP7_75t_SL U60522 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_17_), 
        .Y(n72317) );
  INVx1_ASAP7_75t_SL U60523 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[12]), .Y(n69840) );
  INVxp33_ASAP7_75t_SL U60524 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[24]), .Y(n70088) );
  INVx1_ASAP7_75t_SL U60525 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_o[0]), .Y(
        n27627) );
  INVx1_ASAP7_75t_SL U60526 ( .A(n2777), .Y(n60281) );
  INVxp67_ASAP7_75t_SL U60527 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[24]), .Y(n27501) );
  INVxp67_ASAP7_75t_SL U60528 ( .A(n885), .Y(n64005) );
  INVx1_ASAP7_75t_SL U60529 ( .A(or1200_cpu_or1200_except_n492), .Y(n76681) );
  INVx1_ASAP7_75t_SL U60530 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[11]), .Y(n69821) );
  INVxp67_ASAP7_75t_SL U60531 ( .A(n1108), .Y(n76533) );
  NAND2xp33_ASAP7_75t_SL U60532 ( .A(or1200_cpu_or1200_mult_mac_n157), .B(
        or1200_cpu_or1200_mult_mac_n303), .Y(n63433) );
  INVxp33_ASAP7_75t_SL U60533 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_15_), .Y(n69665) );
  INVx1_ASAP7_75t_SL U60534 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_24_), .Y(
        n74645) );
  INVxp67_ASAP7_75t_SL U60535 ( .A(n1053), .Y(n76606) );
  INVxp33_ASAP7_75t_SL U60536 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_3_), .Y(
        n72580) );
  NAND2xp5_ASAP7_75t_SL U60537 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_3_), .Y(
        n72572) );
  INVx1_ASAP7_75t_SL U60538 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .Y(n78435) );
  INVx1_ASAP7_75t_SL U60539 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_9_), .Y(n65383) );
  INVx1_ASAP7_75t_SL U60540 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .Y(
        n71894) );
  NAND2xp33_ASAP7_75t_SL U60541 ( .A(or1200_cpu_or1200_mult_mac_n297), .B(
        or1200_cpu_or1200_mult_mac_n151), .Y(n63340) );
  NAND2xp5_ASAP7_75t_SL U60542 ( .A(or1200_cpu_or1200_mult_mac_n201), .B(
        or1200_cpu_or1200_mult_mac_n347), .Y(n68879) );
  INVx1_ASAP7_75t_SL U60543 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[22]), .Y(n73743) );
  INVx1_ASAP7_75t_SL U60544 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_5_), .Y(
        n71667) );
  INVx1_ASAP7_75t_SL U60545 ( .A(or1200_cpu_or1200_except_n260), .Y(n75533) );
  INVxp67_ASAP7_75t_SL U60546 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[25]), .Y(n27500) );
  INVxp67_ASAP7_75t_SL U60547 ( .A(or1200_cpu_or1200_mult_mac_n187), .Y(n75557) );
  INVx1_ASAP7_75t_SL U60548 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_8_), .Y(
        n71677) );
  INVx1_ASAP7_75t_SL U60549 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_), 
        .Y(n71936) );
  INVx1_ASAP7_75t_SL U60550 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_33_), 
        .Y(n72141) );
  INVx1_ASAP7_75t_SL U60551 ( .A(or1200_cpu_or1200_except_n616), .Y(n63960) );
  INVxp67_ASAP7_75t_SL U60552 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[6]), .Y(n73560)
         );
  INVx1_ASAP7_75t_SL U60553 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .Y(n71994) );
  INVx1_ASAP7_75t_SL U60554 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_7_), .Y(n65327) );
  INVx1_ASAP7_75t_SL U60555 ( .A(or1200_cpu_or1200_except_n256), .Y(n75145) );
  INVxp67_ASAP7_75t_SL U60556 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_36_), .Y(n69624) );
  INVx1_ASAP7_75t_SL U60557 ( .A(or1200_cpu_or1200_except_n649), .Y(n65218) );
  INVx1_ASAP7_75t_SL U60558 ( .A(or1200_cpu_or1200_mult_mac_ex_freeze_r), .Y(
        n62011) );
  INVx1_ASAP7_75t_SL U60559 ( .A(n2345), .Y(n70354) );
  INVx1_ASAP7_75t_SL U60560 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[9]), .Y(n78233) );
  INVx1_ASAP7_75t_SL U60561 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_19_), .Y(
        n74662) );
  INVxp67_ASAP7_75t_SL U60562 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_40_), .Y(n69651) );
  INVxp67_ASAP7_75t_SL U60563 ( .A(n876), .Y(n63997) );
  INVx1_ASAP7_75t_SL U60564 ( .A(or1200_cpu_esr[0]), .Y(n76665) );
  NAND2xp5_ASAP7_75t_SL U60565 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_5_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_6_), .Y(
        n71637) );
  INVx1_ASAP7_75t_SL U60566 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .Y(n71950) );
  INVx1_ASAP7_75t_SL U60567 ( .A(n1727), .Y(n76682) );
  INVx1_ASAP7_75t_SL U60568 ( .A(or1200_cpu_or1200_mult_mac_n211), .Y(n68864)
         );
  INVxp33_ASAP7_75t_SL U60569 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[22]), .Y(
        n73338) );
  INVxp67_ASAP7_75t_SL U60570 ( .A(n1031), .Y(n61575) );
  NAND2xp33_ASAP7_75t_SL U60571 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_1_), .Y(
        n72576) );
  INVx1_ASAP7_75t_SL U60572 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[25]), .Y(n27456) );
  INVx1_ASAP7_75t_SL U60573 ( .A(or1200_cpu_or1200_except_n264), .Y(n73959) );
  INVxp67_ASAP7_75t_SL U60574 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_6_), .Y(
        n71664) );
  INVxp67_ASAP7_75t_SL U60575 ( .A(n2761), .Y(n60274) );
  INVxp67_ASAP7_75t_SL U60576 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_0_), 
        .Y(n71835) );
  NAND2xp5_ASAP7_75t_SL U60577 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_1_), .Y(
        n72568) );
  INVxp67_ASAP7_75t_SL U60578 ( .A(or1200_cpu_or1200_mult_mac_n6), .Y(n58665)
         );
  INVx1_ASAP7_75t_SL U60579 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[10]), .Y(n78348) );
  INVx1_ASAP7_75t_SL U60580 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_4_), .Y(
        n72584) );
  INVx1_ASAP7_75t_SL U60581 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_5_), .Y(
        n71724) );
  INVxp33_ASAP7_75t_SL U60582 ( .A(n2826), .Y(n76325) );
  INVx1_ASAP7_75t_SL U60583 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_5_), .Y(n65348) );
  INVx1_ASAP7_75t_SL U60584 ( .A(n1368), .Y(n77140) );
  INVx1_ASAP7_75t_SL U60585 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[13]), .Y(n69855) );
  INVx1_ASAP7_75t_SL U60586 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[26]), .Y(n27499) );
  INVx1_ASAP7_75t_SL U60587 ( .A(or1200_cpu_or1200_except_n268), .Y(n76649) );
  INVxp67_ASAP7_75t_SL U60588 ( .A(n2086), .Y(n76322) );
  INVx1_ASAP7_75t_SL U60589 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_3_), .Y(
        n71733) );
  INVx1_ASAP7_75t_SL U60590 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_1_), 
        .Y(n71869) );
  INVx1_ASAP7_75t_SL U60591 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_2_), .Y(
        n72579) );
  INVx1_ASAP7_75t_SL U60592 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_), 
        .Y(n72005) );
  INVx1_ASAP7_75t_SL U60593 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[2]), .Y(n78331)
         );
  INVx1_ASAP7_75t_SL U60594 ( .A(or1200_cpu_or1200_mult_mac_n263), .Y(n75654)
         );
  INVx1_ASAP7_75t_SL U60595 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_), 
        .Y(n71952) );
  NAND2xp5_ASAP7_75t_SL U60596 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_3_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_4_), .Y(
        n72569) );
  INVx1_ASAP7_75t_SL U60597 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_4_), .Y(
        n71738) );
  INVxp67_ASAP7_75t_SL U60598 ( .A(n2069), .Y(n76321) );
  INVxp33_ASAP7_75t_SL U60599 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .Y(
        n70379) );
  INVxp67_ASAP7_75t_SL U60600 ( .A(n854), .Y(n63945) );
  INVx1_ASAP7_75t_SL U60601 ( .A(n1849), .Y(n60288) );
  INVx1_ASAP7_75t_SL U60602 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_), 
        .Y(n71995) );
  NAND2xp5_ASAP7_75t_SL U60603 ( .A(n78443), .B(n78442), .Y(n78450) );
  NAND2xp5_ASAP7_75t_SL U60604 ( .A(n78445), .B(n78444), .Y(n78449) );
  NAND2xp5_ASAP7_75t_SL U60605 ( .A(n78447), .B(n78446), .Y(n78448) );
  NAND2xp5_ASAP7_75t_SL U60606 ( .A(n59713), .B(dwb_ack_i), .Y(n77414) );
  NAND2xp5_ASAP7_75t_SL U60607 ( .A(iwb_ack_i), .B(n60272), .Y(n77403) );
  INVx1_ASAP7_75t_SL U60608 ( .A(dbg_stall_i), .Y(n77429) );
  INVx1_ASAP7_75t_SL U60609 ( .A(dwb_err_i), .Y(n60208) );
  INVx1_ASAP7_75t_SL U60610 ( .A(dbg_dat_i[2]), .Y(n76570) );
  INVx1_ASAP7_75t_SL U60611 ( .A(dbg_dat_i[10]), .Y(n63695) );
  INVx1_ASAP7_75t_SL U60612 ( .A(dbg_dat_i[4]), .Y(n76591) );
  INVx1_ASAP7_75t_SL U60613 ( .A(dwb_dat_i[5]), .Y(n61079) );
  INVx1_ASAP7_75t_SL U60614 ( .A(pic_ints_i[16]), .Y(n60255) );
  INVx1_ASAP7_75t_SL U60615 ( .A(pic_ints_i[8]), .Y(n60254) );
  INVx1_ASAP7_75t_SL U60616 ( .A(pic_ints_i[6]), .Y(n60253) );
  INVx1_ASAP7_75t_SL U60617 ( .A(pic_ints_i[18]), .Y(n60252) );
  INVx1_ASAP7_75t_SL U60618 ( .A(pic_ints_i[14]), .Y(n60251) );
  INVx1_ASAP7_75t_SL U60619 ( .A(pic_ints_i[4]), .Y(n60250) );
  INVx1_ASAP7_75t_SL U60620 ( .A(pic_ints_i[10]), .Y(n60249) );
  INVx1_ASAP7_75t_SL U60621 ( .A(pic_ints_i[12]), .Y(n60248) );
  INVx1_ASAP7_75t_SL U60622 ( .A(pic_ints_i[13]), .Y(n60247) );
  INVx1_ASAP7_75t_SL U60623 ( .A(pic_ints_i[7]), .Y(n60244) );
  INVx1_ASAP7_75t_SL U60624 ( .A(pic_ints_i[17]), .Y(n60243) );
  INVx1_ASAP7_75t_SL U60625 ( .A(pic_ints_i[9]), .Y(n60242) );
  INVx1_ASAP7_75t_SL U60626 ( .A(pic_ints_i[11]), .Y(n60241) );
  INVx1_ASAP7_75t_SL U60627 ( .A(pic_ints_i[5]), .Y(n60240) );
  INVx1_ASAP7_75t_SL U60628 ( .A(pic_ints_i[2]), .Y(n60239) );
  INVx1_ASAP7_75t_SL U60629 ( .A(pic_ints_i[15]), .Y(n60238) );
  INVx1_ASAP7_75t_SL U60630 ( .A(pic_ints_i[3]), .Y(n60237) );
  INVx1_ASAP7_75t_SL U60631 ( .A(dbg_dat_i[3]), .Y(n61578) );
  INVx1_ASAP7_75t_SL U60632 ( .A(dwb_dat_i[13]), .Y(n61075) );
  INVx1_ASAP7_75t_SL U60633 ( .A(dbg_dat_i[12]), .Y(n63935) );
  INVx1_ASAP7_75t_SL U60634 ( .A(dbg_dat_i[25]), .Y(n60175) );
  INVx1_ASAP7_75t_SL U60635 ( .A(dbg_dat_i[14]), .Y(n60166) );
  INVx1_ASAP7_75t_SL U60636 ( .A(dbg_dat_i[20]), .Y(n60154) );
  INVx1_ASAP7_75t_SL U60637 ( .A(dbg_dat_i[18]), .Y(n60146) );
  INVx1_ASAP7_75t_SL U60638 ( .A(dbg_dat_i[19]), .Y(n60134) );
  INVx1_ASAP7_75t_SL U60639 ( .A(dbg_dat_i[15]), .Y(n60100) );
  INVx1_ASAP7_75t_SL U60640 ( .A(dbg_dat_i[13]), .Y(n60052) );
  INVx1_ASAP7_75t_SL U60641 ( .A(dbg_dat_i[23]), .Y(n60081) );
  INVx1_ASAP7_75t_SL U60642 ( .A(dbg_dat_i[21]), .Y(n60069) );
  INVx1_ASAP7_75t_SL U60643 ( .A(or1200_dc_top_tag_10_), .Y(n59729) );
  INVx1_ASAP7_75t_SL U60644 ( .A(or1200_dc_top_tag_17_), .Y(n59748) );
  INVx1_ASAP7_75t_SL U60645 ( .A(or1200_dc_top_from_dcram_7_), .Y(n60874) );
  INVx1_ASAP7_75t_SL U60646 ( .A(or1200_dc_top_tag_2_), .Y(n59740) );
  INVx1_ASAP7_75t_SL U60647 ( .A(or1200_dc_top_from_dcram_15_), .Y(n60877) );
  INVx1_ASAP7_75t_SL U60648 ( .A(or1200_dc_top_tag_16_), .Y(n59737) );
  INVx1_ASAP7_75t_SL U60649 ( .A(or1200_dc_top_tag_4_), .Y(n59824) );
  INVx1_ASAP7_75t_SL U60650 ( .A(or1200_dc_top_tag_12_), .Y(n59797) );
  INVx1_ASAP7_75t_SL U60651 ( .A(or1200_dc_top_tag_8_), .Y(n59788) );
  INVx1_ASAP7_75t_SL U60652 ( .A(or1200_dc_top_tag_15_), .Y(n59753) );
  INVx1_ASAP7_75t_SL U60653 ( .A(or1200_dc_top_tag_14_), .Y(n59751) );
  INVx1_ASAP7_75t_SL U60654 ( .A(or1200_dc_top_tag_6_), .Y(n59817) );
  INVx1_ASAP7_75t_SL U60655 ( .A(or1200_dc_top_tag_1_), .Y(n59811) );
  INVx1_ASAP7_75t_SL U60656 ( .A(or1200_dc_top_tag_9_), .Y(n59765) );
  INVx1_ASAP7_75t_SL U60657 ( .A(or1200_ic_top_from_icram[17]), .Y(n77948) );
  INVx1_ASAP7_75t_SL U60658 ( .A(or1200_ic_top_from_icram[19]), .Y(n77939) );
  INVx1_ASAP7_75t_SL U60659 ( .A(or1200_ic_top_from_icram[30]), .Y(n60435) );
  INVx1_ASAP7_75t_SL U60660 ( .A(or1200_ic_top_from_icram[31]), .Y(n60448) );
  INVx1_ASAP7_75t_SL U60661 ( .A(or1200_ic_top_from_icram[18]), .Y(n60534) );
  INVx1_ASAP7_75t_SL U60662 ( .A(or1200_ic_top_from_icram[20]), .Y(n60529) );
  XOR2xp5_ASAP7_75t_SL U60663 ( .A(n67766), .B(n57095), .Y(n57249) );
  XNOR2xp5_ASAP7_75t_SL U60664 ( .A(n67656), .B(n59058), .Y(n67766) );
  AOI21x1_ASAP7_75t_SL U60665 ( .A1(n67560), .A2(n59041), .B(n57304), .Y(
        n59040) );
  NAND3xp33_ASAP7_75t_SL U60666 ( .A(n56849), .B(n57569), .C(n57030), .Y(
        n67730) );
  OAI21xp5_ASAP7_75t_SL U60667 ( .A1(n68087), .A2(n59595), .B(n63209), .Y(
        n63636) );
  NAND2x1_ASAP7_75t_SL U60668 ( .A(n64620), .B(n58240), .Y(n64895) );
  NOR2x1p5_ASAP7_75t_SL U60669 ( .A(n59566), .B(n59464), .Y(n57252) );
  XNOR2x1_ASAP7_75t_SL U60670 ( .A(n57543), .B(n57634), .Y(n67795) );
  NAND2x1_ASAP7_75t_SL U60671 ( .A(n67794), .B(n67795), .Y(n67936) );
  NOR2x1_ASAP7_75t_SL U60672 ( .A(n76653), .B(n62646), .Y(n62644) );
  INVx6_ASAP7_75t_SL U60673 ( .A(n58207), .Y(n66258) );
  BUFx12f_ASAP7_75t_SL U60674 ( .A(n75033), .Y(n59518) );
  XNOR2x2_ASAP7_75t_SL U60675 ( .A(n59511), .B(n59640), .Y(n67819) );
  MAJIxp5_ASAP7_75t_SL U60676 ( .A(n63832), .B(n63833), .C(n63834), .Y(n64663)
         );
  OAI22xp5_ASAP7_75t_SL U60677 ( .A1(n63630), .A2(n57360), .B1(n59515), .B2(
        n63823), .Y(n63834) );
  MAJIxp5_ASAP7_75t_SL U60678 ( .A(n68168), .B(n68166), .C(n68167), .Y(n68173)
         );
  XNOR2xp5_ASAP7_75t_SL U60679 ( .A(n68107), .B(n57222), .Y(n68194) );
  XNOR2xp5_ASAP7_75t_SL U60680 ( .A(n68108), .B(n57719), .Y(n57222) );
  XNOR2xp5_ASAP7_75t_SL U60681 ( .A(n63277), .B(n62898), .Y(n63260) );
  NOR2x1_ASAP7_75t_SL U60682 ( .A(n62897), .B(n62896), .Y(n63277) );
  INVx2_ASAP7_75t_SL U60683 ( .A(n59235), .Y(n62808) );
  XNOR2xp5_ASAP7_75t_SL U60684 ( .A(n62756), .B(n58985), .Y(n57473) );
  NAND2x1p5_ASAP7_75t_SL U60685 ( .A(n57716), .B(n58755), .Y(n58757) );
  INVx5_ASAP7_75t_SL U60686 ( .A(n59239), .Y(n59054) );
  NOR2x1p5_ASAP7_75t_SL U60687 ( .A(n57223), .B(n57777), .Y(n68065) );
  INVx4_ASAP7_75t_SL U60688 ( .A(n58336), .Y(n59116) );
  XNOR2x1_ASAP7_75t_SL U60689 ( .A(n68486), .B(n58942), .Y(n68487) );
  AOI21xp5_ASAP7_75t_SL U60690 ( .A1(n68068), .A2(n68070), .B(n68069), .Y(
        n57223) );
  INVx3_ASAP7_75t_SL U60691 ( .A(n59608), .Y(n59611) );
  NAND2xp5_ASAP7_75t_SL U60692 ( .A(n64090), .B(n57226), .Y(n58099) );
  NAND3xp33_ASAP7_75t_SL U60693 ( .A(n64089), .B(n64667), .C(n64665), .Y(
        n57226) );
  OR2x6_ASAP7_75t_SL U60694 ( .A(n67331), .B(n63656), .Y(n59652) );
  XNOR2x1_ASAP7_75t_SL U60695 ( .A(n59652), .B(n59602), .Y(n59332) );
  XOR2x2_ASAP7_75t_SL U60696 ( .A(n57227), .B(n58396), .Y(n67665) );
  AOI21xp5_ASAP7_75t_SL U60697 ( .A1(n67679), .A2(n67672), .B(n67678), .Y(
        n57227) );
  HB1xp67_ASAP7_75t_SL U60698 ( .A(n64957), .Y(n57348) );
  XNOR2xp5_ASAP7_75t_SL U60699 ( .A(n68402), .B(n68399), .Y(n67563) );
  INVx6_ASAP7_75t_SL U60700 ( .A(n66411), .Y(n59239) );
  NOR2x1_ASAP7_75t_SL U60701 ( .A(n68413), .B(n59041), .Y(n67253) );
  MAJIxp5_ASAP7_75t_SL U60702 ( .A(n67407), .B(n67406), .C(n67405), .Y(n67528)
         );
  OAI22xp5_ASAP7_75t_SL U60703 ( .A1(n57076), .A2(n67258), .B1(n67279), .B2(
        n67871), .Y(n67406) );
  INVx1_ASAP7_75t_SL U60704 ( .A(n57900), .Y(n64042) );
  NOR2x1p5_ASAP7_75t_SL U60705 ( .A(n59041), .B(n67562), .Y(n57304) );
  NAND2x1p5_ASAP7_75t_SL U60706 ( .A(n64503), .B(n59144), .Y(n59454) );
  INVx2_ASAP7_75t_SL U60707 ( .A(n67868), .Y(n67967) );
  NAND2xp5_ASAP7_75t_SL U60708 ( .A(n67319), .B(n67967), .Y(n67320) );
  BUFx3_ASAP7_75t_SL U60709 ( .A(n59253), .Y(n57253) );
  OAI21x1_ASAP7_75t_SL U60710 ( .A1(n59456), .A2(n57662), .B(n59359), .Y(
        n68015) );
  INVx4_ASAP7_75t_SL U60711 ( .A(n59418), .Y(n67920) );
  NAND2x1p5_ASAP7_75t_SL U60712 ( .A(n57736), .B(n66988), .Y(n66706) );
  NAND2xp5_ASAP7_75t_SL U60713 ( .A(n59660), .B(n67963), .Y(n67926) );
  INVx2_ASAP7_75t_SL U60714 ( .A(n68111), .Y(n68113) );
  XNOR2x1_ASAP7_75t_SL U60715 ( .A(n67804), .B(n57778), .Y(n68068) );
  NAND2x1_ASAP7_75t_SL U60716 ( .A(n68571), .B(n68570), .Y(n68836) );
  NAND3xp33_ASAP7_75t_SL U60717 ( .A(n68254), .B(n68253), .C(n68836), .Y(
        n68561) );
  NAND2xp33_ASAP7_75t_SRAM U60718 ( .A(n66258), .B(n62609), .Y(n58941) );
  OR2x2_ASAP7_75t_SL U60719 ( .A(n57228), .B(n58343), .Y(n62609) );
  NAND2xp5_ASAP7_75t_SL U60720 ( .A(n57229), .B(n57200), .Y(n57228) );
  INVx1_ASAP7_75t_SL U60721 ( .A(n64896), .Y(n57230) );
  NAND2xp5_ASAP7_75t_SL U60722 ( .A(n59350), .B(n59291), .Y(n64896) );
  OAI21x1_ASAP7_75t_SL U60723 ( .A1(n57122), .A2(n64917), .B(n66296), .Y(
        n68100) );
  AO21x1_ASAP7_75t_SL U60724 ( .A1(n59165), .A2(n57356), .B(n57232), .Y(n64914) );
  OA22x2_ASAP7_75t_SL U60725 ( .A1(n59126), .A2(n60915), .B1(n59538), .B2(
        n64504), .Y(n58906) );
  INVx3_ASAP7_75t_SL U60726 ( .A(n75908), .Y(n75900) );
  BUFx6f_ASAP7_75t_SL U60727 ( .A(n75643), .Y(n59484) );
  INVx1_ASAP7_75t_SL U60728 ( .A(n63482), .Y(n62781) );
  OR2x6_ASAP7_75t_SL U60729 ( .A(n63859), .B(n67308), .Y(n67585) );
  NAND3xp33_ASAP7_75t_SL U60730 ( .A(n59560), .B(n59571), .C(n59542), .Y(
        n59429) );
  NOR2x1_ASAP7_75t_SL U60731 ( .A(n59239), .B(n59455), .Y(n58673) );
  NAND3xp33_ASAP7_75t_SL U60732 ( .A(n62571), .B(n62572), .C(n62570), .Y(
        n59104) );
  OAI21xp5_ASAP7_75t_SL U60733 ( .A1(n59648), .A2(n57108), .B(n58805), .Y(
        n67809) );
  INVx1_ASAP7_75t_SL U60734 ( .A(n57678), .Y(n57233) );
  NAND2x1_ASAP7_75t_SL U60735 ( .A(n57233), .B(n56846), .Y(n67995) );
  BUFx2_ASAP7_75t_SL U60736 ( .A(n64034), .Y(n57234) );
  XNOR2xp5_ASAP7_75t_SL U60737 ( .A(n57150), .B(n64557), .Y(n64495) );
  XNOR2xp5_ASAP7_75t_SL U60738 ( .A(n57401), .B(n64493), .Y(n64557) );
  XOR2x2_ASAP7_75t_SL U60739 ( .A(n68529), .B(n68509), .Y(n68518) );
  XOR2xp5_ASAP7_75t_SL U60740 ( .A(n58358), .B(n68518), .Y(n58435) );
  NAND2xp5_ASAP7_75t_SL U60741 ( .A(n59568), .B(n60751), .Y(n61396) );
  OAI21xp5_ASAP7_75t_SL U60742 ( .A1(n57463), .A2(n53231), .B(n66432), .Y(
        n66434) );
  OAI21xp5_ASAP7_75t_SL U60743 ( .A1(n67891), .A2(n58662), .B(n57236), .Y(
        n67779) );
  NAND2xp5_ASAP7_75t_SL U60744 ( .A(n59223), .B(n67893), .Y(n57236) );
  OAI21xp5_ASAP7_75t_SL U60745 ( .A1(n68235), .A2(n68234), .B(n68231), .Y(
        n68030) );
  INVx5_ASAP7_75t_SL U60746 ( .A(n59509), .Y(n67428) );
  XOR2xp5_ASAP7_75t_SL U60747 ( .A(n57238), .B(n57237), .Y(n64069) );
  INVx1_ASAP7_75t_SL U60748 ( .A(n64086), .Y(n57237) );
  XNOR2xp5_ASAP7_75t_SL U60749 ( .A(n64663), .B(n64085), .Y(n57238) );
  NAND2xp5_ASAP7_75t_SL U60750 ( .A(n75912), .B(n67463), .Y(n57239) );
  NOR2x1_ASAP7_75t_SL U60751 ( .A(n59598), .B(n76028), .Y(n57240) );
  NAND2x1_ASAP7_75t_SL U60752 ( .A(n57164), .B(n57040), .Y(n57440) );
  BUFx6f_ASAP7_75t_SL U60753 ( .A(n1761), .Y(n59707) );
  INVx1_ASAP7_75t_SL U60754 ( .A(n67748), .Y(n58667) );
  AOI22xp33_ASAP7_75t_SL U60755 ( .A1(n64894), .A2(n76653), .B1(n59569), .B2(
        n66258), .Y(n62645) );
  XNOR2x2_ASAP7_75t_SL U60756 ( .A(n66496), .B(n66495), .Y(n67114) );
  INVx8_ASAP7_75t_SL U60757 ( .A(n57637), .Y(n59619) );
  INVx11_ASAP7_75t_SL U60758 ( .A(n59619), .Y(n59012) );
  NOR2x1p5_ASAP7_75t_SL U60759 ( .A(n62562), .B(n59462), .Y(n62555) );
  BUFx2_ASAP7_75t_SL U60760 ( .A(n67836), .Y(n57419) );
  NAND2x1_ASAP7_75t_SL U60761 ( .A(n75904), .B(n67841), .Y(n57282) );
  INVx1_ASAP7_75t_SL U60762 ( .A(n68084), .Y(n59192) );
  XOR2xp5_ASAP7_75t_SL U60763 ( .A(n64415), .B(n64414), .Y(n57760) );
  NOR2x1_ASAP7_75t_SL U60764 ( .A(n64029), .B(n57761), .Y(n64415) );
  NAND2xp5_ASAP7_75t_SL U60765 ( .A(n57113), .B(n67911), .Y(n67224) );
  OAI22xp5_ASAP7_75t_SL U60766 ( .A1(n68383), .A2(n68382), .B1(n53269), .B2(
        n68381), .Y(n68439) );
  INVx3_ASAP7_75t_SL U60767 ( .A(n57104), .Y(n59651) );
  NAND2xp5_ASAP7_75t_SL U60768 ( .A(n2006), .B(n59563), .Y(n66240) );
  INVx1_ASAP7_75t_SL U60769 ( .A(n67599), .Y(n57247) );
  OAI21xp5_ASAP7_75t_SL U60770 ( .A1(n68087), .A2(n59242), .B(n64609), .Y(
        n59009) );
  XNOR2xp5_ASAP7_75t_SL U60771 ( .A(n67768), .B(n57249), .Y(n67769) );
  NAND2xp5_ASAP7_75t_SL U60772 ( .A(n67909), .B(n59604), .Y(n59132) );
  XNOR2xp5_ASAP7_75t_SL U60773 ( .A(n68553), .B(n68554), .Y(n57418) );
  MAJIxp5_ASAP7_75t_SL U60774 ( .A(n68542), .B(n68543), .C(n68544), .Y(n68554)
         );
  NOR2x1p5_ASAP7_75t_SL U60775 ( .A(n57251), .B(n57250), .Y(n62565) );
  INVx2_ASAP7_75t_SL U60776 ( .A(n57252), .Y(n57251) );
  NOR2x1p5_ASAP7_75t_SL U60777 ( .A(n58222), .B(n62613), .Y(n67959) );
  INVx1_ASAP7_75t_SL U60778 ( .A(n63177), .Y(n59128) );
  BUFx6f_ASAP7_75t_SL U60779 ( .A(n2508), .Y(n59462) );
  AND3x2_ASAP7_75t_SL U60780 ( .A(n58205), .B(n57635), .C(n62567), .Y(n58265)
         );
  OR2x2_ASAP7_75t_SL U60781 ( .A(n67898), .B(n66470), .Y(n58859) );
  XNOR2xp5_ASAP7_75t_SL U60782 ( .A(n57456), .B(n57172), .Y(n66470) );
  NOR2x1_ASAP7_75t_SL U60783 ( .A(n67517), .B(n59277), .Y(n57596) );
  AOI22xp5_ASAP7_75t_SL U60784 ( .A1(n67901), .A2(n67561), .B1(n67560), .B2(
        n57101), .Y(n59162) );
  AOI22xp33_ASAP7_75t_SRAM U60785 ( .A1(n67432), .A2(n67948), .B1(n75912), 
        .B2(n67431), .Y(n67433) );
  INVx1_ASAP7_75t_SL U60786 ( .A(n59469), .Y(n67853) );
  INVx1_ASAP7_75t_SL U60787 ( .A(n68147), .Y(n57979) );
  NAND2xp5_ASAP7_75t_SL U60788 ( .A(n57035), .B(n58068), .Y(n68147) );
  NAND2xp5_ASAP7_75t_SL U60789 ( .A(n64609), .B(n57049), .Y(n57671) );
  AOI21xp5_ASAP7_75t_SL U60790 ( .A1(n57108), .A2(n59649), .B(n58806), .Y(
        n58804) );
  NOR2x1p5_ASAP7_75t_SL U60791 ( .A(n58489), .B(n57466), .Y(n58650) );
  XOR2xp5_ASAP7_75t_SL U60792 ( .A(n68506), .B(n68505), .Y(n68507) );
  XOR2xp5_ASAP7_75t_SL U60793 ( .A(n57014), .B(n58133), .Y(n68506) );
  INVx1_ASAP7_75t_SL U60794 ( .A(n57254), .Y(n64355) );
  NOR3xp33_ASAP7_75t_SL U60795 ( .A(n64619), .B(n63174), .C(n58496), .Y(n57254) );
  AO21x2_ASAP7_75t_SL U60796 ( .A1(n57786), .A2(n67603), .B(n57785), .Y(n67814) );
  O2A1O1Ixp5_ASAP7_75t_SL U60797 ( .A1(n57292), .A2(n67244), .B(n67243), .C(
        n58413), .Y(n67245) );
  XNOR2xp5_ASAP7_75t_SL U60798 ( .A(n57169), .B(n57525), .Y(n58413) );
  INVx1_ASAP7_75t_SL U60799 ( .A(n63184), .Y(n63126) );
  NAND2x1_ASAP7_75t_SL U60800 ( .A(n59011), .B(n68694), .Y(n74559) );
  NAND2xp5_ASAP7_75t_SL U60801 ( .A(n76225), .B(n63048), .Y(n58812) );
  NAND2xp5_ASAP7_75t_SL U60802 ( .A(n63047), .B(n63046), .Y(n76225) );
  XNOR2x1_ASAP7_75t_SL U60803 ( .A(n57372), .B(n57255), .Y(n68074) );
  INVx1_ASAP7_75t_SL U60804 ( .A(n57921), .Y(n67938) );
  OR2x2_ASAP7_75t_SL U60805 ( .A(n67804), .B(n67801), .Y(n57921) );
  OAI21xp5_ASAP7_75t_SL U60806 ( .A1(n67867), .A2(n57010), .B(n57256), .Y(
        n68135) );
  OAI21xp5_ASAP7_75t_SL U60807 ( .A1(n67866), .A2(n58015), .B(n67865), .Y(
        n57256) );
  NAND2xp5_ASAP7_75t_SL U60808 ( .A(n57394), .B(n57180), .Y(n64363) );
  XNOR2xp5_ASAP7_75t_SL U60809 ( .A(n63007), .B(n63009), .Y(n62963) );
  NOR2x1_ASAP7_75t_SL U60810 ( .A(n62961), .B(n62962), .Y(n63009) );
  BUFx3_ASAP7_75t_SL U60811 ( .A(n59314), .Y(n58658) );
  INVx2_ASAP7_75t_SL U60812 ( .A(n59613), .Y(n59612) );
  NOR2x1_ASAP7_75t_SL U60813 ( .A(n57094), .B(n67391), .Y(n58910) );
  INVx1_ASAP7_75t_SL U60814 ( .A(n67626), .Y(n67266) );
  XNOR2xp5_ASAP7_75t_SL U60815 ( .A(n65010), .B(n57258), .Y(n65003) );
  XNOR2xp5_ASAP7_75t_SL U60816 ( .A(n65011), .B(n65009), .Y(n57258) );
  OAI21x1_ASAP7_75t_SL U60817 ( .A1(n68024), .A2(n58884), .B(n68023), .Y(
        n58811) );
  BUFx16f_ASAP7_75t_SL U60818 ( .A(n58143), .Y(n59607) );
  INVx4_ASAP7_75t_SL U60819 ( .A(n59607), .Y(n58865) );
  NAND2xp5_ASAP7_75t_SL U60820 ( .A(n56974), .B(n63185), .Y(n63186) );
  NOR2x1p5_ASAP7_75t_SL U60821 ( .A(n57259), .B(n62648), .Y(n57567) );
  NAND2x1_ASAP7_75t_SL U60822 ( .A(n57537), .B(n56979), .Y(n62958) );
  NAND3xp33_ASAP7_75t_SL U60823 ( .A(n57921), .B(n57922), .C(n67936), .Y(
        n57920) );
  INVx3_ASAP7_75t_SL U60824 ( .A(n68012), .Y(n67912) );
  OAI21x1_ASAP7_75t_SL U60825 ( .A1(n67284), .A2(n58113), .B(n57262), .Y(
        n59450) );
  NAND2x1_ASAP7_75t_SL U60826 ( .A(n58675), .B(n56994), .Y(n57262) );
  NAND2x1_ASAP7_75t_SL U60827 ( .A(n64548), .B(n64549), .Y(n64693) );
  AOI21x1_ASAP7_75t_SL U60828 ( .A1(n59620), .A2(n67914), .B(n57176), .Y(
        n67915) );
  NAND2xp5_ASAP7_75t_SL U60829 ( .A(n59523), .B(n71108), .Y(n71112) );
  OAI21x1_ASAP7_75t_SL U60830 ( .A1(n57263), .A2(n57873), .B(n57872), .Y(
        n68184) );
  NAND2xp5_ASAP7_75t_SL U60831 ( .A(n58761), .B(n57025), .Y(n57263) );
  NOR2x1p5_ASAP7_75t_SL U60832 ( .A(n57364), .B(n57363), .Y(n67685) );
  NAND2x1p5_ASAP7_75t_SL U60833 ( .A(n57066), .B(n67419), .Y(n67646) );
  INVx1_ASAP7_75t_SL U60834 ( .A(n59518), .Y(n57264) );
  AND2x2_ASAP7_75t_SL U60835 ( .A(n57264), .B(n58656), .Y(n66322) );
  INVx6_ASAP7_75t_SL U60836 ( .A(n59637), .Y(n59639) );
  OAI21xp5_ASAP7_75t_SL U60837 ( .A1(n68139), .A2(n68137), .B(n68136), .Y(
        n57265) );
  BUFx6f_ASAP7_75t_SL U60838 ( .A(n1683), .Y(n59537) );
  INVx1_ASAP7_75t_SL U60839 ( .A(n64895), .Y(n57340) );
  NAND2xp5_ASAP7_75t_SL U60840 ( .A(n57267), .B(n57266), .Y(n58994) );
  NAND2xp5_ASAP7_75t_SL U60841 ( .A(n64587), .B(n64586), .Y(n57266) );
  OAI21xp5_ASAP7_75t_SL U60842 ( .A1(n64458), .A2(n64457), .B(n57143), .Y(
        n57267) );
  NAND2xp5_ASAP7_75t_SL U60843 ( .A(n59536), .B(n64078), .Y(n58925) );
  XNOR2x1_ASAP7_75t_SL U60844 ( .A(n57268), .B(n57490), .Y(n67888) );
  NAND2xp5_ASAP7_75t_SL U60845 ( .A(n57179), .B(n67920), .Y(n67921) );
  NOR2x1_ASAP7_75t_SL U60846 ( .A(n58933), .B(n67409), .Y(n67477) );
  NAND2x1p5_ASAP7_75t_SL U60847 ( .A(n59093), .B(n59092), .Y(n67765) );
  INVx2_ASAP7_75t_SL U60848 ( .A(n58856), .Y(n58172) );
  NAND2xp5_ASAP7_75t_SL U60849 ( .A(n59605), .B(n67908), .Y(n67910) );
  INVx2_ASAP7_75t_SL U60850 ( .A(n57270), .Y(n64928) );
  NOR2x1_ASAP7_75t_SL U60851 ( .A(n59352), .B(n59291), .Y(n57270) );
  NOR2x1_ASAP7_75t_SL U60852 ( .A(n67595), .B(n67366), .Y(n67905) );
  INVx1_ASAP7_75t_SL U60853 ( .A(n68080), .Y(n57309) );
  XNOR2xp5_ASAP7_75t_SL U60854 ( .A(n59244), .B(n68069), .Y(n68071) );
  OAI21xp5_ASAP7_75t_SL U60855 ( .A1(n57110), .A2(n59470), .B(n62921), .Y(
        n64489) );
  NAND2xp5_ASAP7_75t_SL U60856 ( .A(n67059), .B(n59635), .Y(n58708) );
  OAI21xp5_ASAP7_75t_SL U60857 ( .A1(n57347), .A2(n64949), .B(n57275), .Y(
        n59475) );
  AOI21xp5_ASAP7_75t_SL U60858 ( .A1(n64951), .A2(n57186), .B(n64950), .Y(
        n57275) );
  NOR2xp33_ASAP7_75t_SL U60859 ( .A(n57276), .B(n59460), .Y(n64635) );
  AOI22xp5_ASAP7_75t_SL U60860 ( .A1(n67585), .A2(n59605), .B1(n75906), .B2(
        n57352), .Y(n64634) );
  INVx2_ASAP7_75t_SL U60861 ( .A(n75468), .Y(n59123) );
  AND2x4_ASAP7_75t_SL U60862 ( .A(n57638), .B(n57710), .Y(n57637) );
  NAND2x1_ASAP7_75t_SL U60863 ( .A(n57391), .B(n57390), .Y(n58930) );
  OAI21xp5_ASAP7_75t_SL U60864 ( .A1(n75893), .A2(n59639), .B(n59518), .Y(
        n66923) );
  NOR2x1_ASAP7_75t_SL U60865 ( .A(n76627), .B(n62804), .Y(n59236) );
  MAJIxp5_ASAP7_75t_SL U60866 ( .A(n63054), .B(n57279), .C(n63053), .Y(n63105)
         );
  INVx1_ASAP7_75t_SL U60867 ( .A(n63052), .Y(n57279) );
  XOR2xp5_ASAP7_75t_SL U60868 ( .A(n57280), .B(n62752), .Y(n63052) );
  INVx1_ASAP7_75t_SL U60869 ( .A(n63058), .Y(n57280) );
  OR3x2_ASAP7_75t_SL U60870 ( .A(n58748), .B(n58844), .C(n66291), .Y(n59117)
         );
  INVx2_ASAP7_75t_SL U60871 ( .A(n59117), .Y(n67704) );
  XNOR2x1_ASAP7_75t_SL U60872 ( .A(n59031), .B(n68420), .Y(n67725) );
  INVx2_ASAP7_75t_SL U60873 ( .A(n67725), .Y(n67722) );
  NOR2x1_ASAP7_75t_SL U60874 ( .A(n57281), .B(n67840), .Y(n68176) );
  OAI21xp5_ASAP7_75t_SL U60875 ( .A1(n59067), .A2(n57942), .B(n57282), .Y(
        n57281) );
  AOI31xp67_ASAP7_75t_SL U60876 ( .A1(n63124), .A2(n57118), .A3(n57210), .B(
        n57283), .Y(n59010) );
  INVx1_ASAP7_75t_SL U60877 ( .A(n57665), .Y(n57283) );
  NAND2xp5_ASAP7_75t_SL U60878 ( .A(n68415), .B(n68414), .Y(n68416) );
  NAND2xp5_ASAP7_75t_SL U60879 ( .A(n59599), .B(n67962), .Y(n67252) );
  XNOR2xp5_ASAP7_75t_SL U60880 ( .A(n57054), .B(n67163), .Y(n58355) );
  O2A1O1Ixp5_ASAP7_75t_SL U60881 ( .A1(n71413), .A2(n71412), .B(n57211), .C(
        n28256), .Y(n71416) );
  AO21x2_ASAP7_75t_SL U60882 ( .A1(n67646), .A2(n58475), .B(n67642), .Y(n67776) );
  XNOR2x1_ASAP7_75t_SL U60883 ( .A(n57825), .B(n57824), .Y(n68491) );
  XOR2x1_ASAP7_75t_SL U60884 ( .A(n68491), .B(n68492), .Y(n58987) );
  INVx2_ASAP7_75t_SL U60885 ( .A(n68107), .Y(n58130) );
  XNOR2xp5_ASAP7_75t_SL U60886 ( .A(n57285), .B(n67695), .Y(n58335) );
  AOI21xp5_ASAP7_75t_SL U60887 ( .A1(n57009), .A2(n67549), .B(n67548), .Y(
        n57285) );
  NAND2xp5_ASAP7_75t_SL U60888 ( .A(n57287), .B(n57286), .Y(n52007) );
  AOI21xp5_ASAP7_75t_SL U60889 ( .A1(n58744), .A2(n58839), .B(n68682), .Y(
        n57286) );
  NAND2xp5_ASAP7_75t_SL U60890 ( .A(n57059), .B(n57288), .Y(n57287) );
  NAND2xp5_ASAP7_75t_SL U60891 ( .A(n68686), .B(n58839), .Y(n57288) );
  O2A1O1Ixp5_ASAP7_75t_SL U60892 ( .A1(n67894), .A2(n58706), .B(n58363), .C(
        n67896), .Y(n59136) );
  NAND2xp5_ASAP7_75t_SL U60893 ( .A(n59530), .B(n66258), .Y(n57339) );
  O2A1O1Ixp5_ASAP7_75t_SL U60894 ( .A1(n59647), .A2(n67481), .B(n57291), .C(
        n67480), .Y(n67482) );
  NAND2xp5_ASAP7_75t_SL U60895 ( .A(n53303), .B(n59648), .Y(n57291) );
  NAND2x1p5_ASAP7_75t_SL U60896 ( .A(n57893), .B(n56848), .Y(n67618) );
  INVx8_ASAP7_75t_SL U60897 ( .A(n59505), .Y(n67629) );
  NOR2x1_ASAP7_75t_SL U60898 ( .A(n59609), .B(n62958), .Y(n66716) );
  OAI21xp5_ASAP7_75t_SL U60899 ( .A1(n59227), .A2(n59225), .B(n59224), .Y(
        n63005) );
  AND2x2_ASAP7_75t_SL U60900 ( .A(n57062), .B(n68803), .Y(n68563) );
  OAI21x1_ASAP7_75t_SL U60901 ( .A1(n67906), .A2(n67905), .B(n67904), .Y(
        n67979) );
  XOR2xp5_ASAP7_75t_SL U60902 ( .A(n65004), .B(n58048), .Y(n57293) );
  INVx3_ASAP7_75t_SL U60903 ( .A(n64424), .Y(n67601) );
  A2O1A1Ixp33_ASAP7_75t_SL U60904 ( .A1(n59620), .A2(n64424), .B(n62696), .C(
        n62695), .Y(n62715) );
  NAND2x2_ASAP7_75t_SL U60905 ( .A(n57295), .B(n57294), .Y(n64424) );
  INVx2_ASAP7_75t_SL U60906 ( .A(n62887), .Y(n57294) );
  INVx2_ASAP7_75t_SL U60907 ( .A(n64625), .Y(n57295) );
  NAND2xp5_ASAP7_75t_SL U60908 ( .A(n58786), .B(n57912), .Y(n59327) );
  NOR2x1p5_ASAP7_75t_SL U60909 ( .A(n63206), .B(n58437), .Y(n59180) );
  BUFx6f_ASAP7_75t_SL U60910 ( .A(n1967), .Y(n59556) );
  INVx1_ASAP7_75t_SL U60911 ( .A(n67909), .Y(n57296) );
  NAND2xp5_ASAP7_75t_SL U60912 ( .A(n59602), .B(n57296), .Y(n58517) );
  OAI21xp5_ASAP7_75t_SL U60913 ( .A1(n62735), .A2(n62736), .B(n62734), .Y(
        n57899) );
  MAJIxp5_ASAP7_75t_SL U60914 ( .A(n58878), .B(n62715), .C(n62714), .Y(n62736)
         );
  NAND2x1p5_ASAP7_75t_SL U60915 ( .A(n68348), .B(n68347), .Y(n68754) );
  NAND2x2_ASAP7_75t_SL U60916 ( .A(n56852), .B(n57297), .Y(n66288) );
  INVx2_ASAP7_75t_SL U60917 ( .A(n58927), .Y(n57297) );
  BUFx3_ASAP7_75t_SL U60918 ( .A(n67709), .Y(n57409) );
  NAND2x2_ASAP7_75t_SL U60919 ( .A(n63671), .B(n63670), .Y(n66411) );
  NAND2x1_ASAP7_75t_SL U60920 ( .A(n61920), .B(n58797), .Y(n61918) );
  XOR2xp5_ASAP7_75t_SL U60921 ( .A(n58137), .B(n57147), .Y(n57766) );
  INVx5_ASAP7_75t_SL U60922 ( .A(n58402), .Y(n59057) );
  NAND2xp5_ASAP7_75t_SL U60923 ( .A(n64189), .B(n75552), .Y(n64756) );
  XNOR2xp5_ASAP7_75t_SL U60924 ( .A(n68112), .B(n68113), .Y(n68114) );
  NOR2x1_ASAP7_75t_SL U60925 ( .A(n63188), .B(n57799), .Y(n63250) );
  NAND2x1_ASAP7_75t_SL U60926 ( .A(n75894), .B(n59518), .Y(n66265) );
  NOR2x1p5_ASAP7_75t_SL U60927 ( .A(n58130), .B(n67992), .Y(n67999) );
  MAJIxp5_ASAP7_75t_SL U60928 ( .A(n68521), .B(n68522), .C(n68523), .Y(n68555)
         );
  XOR2xp5_ASAP7_75t_SL U60929 ( .A(n57020), .B(n57298), .Y(n63108) );
  NOR2x1p5_ASAP7_75t_SL U60930 ( .A(n57496), .B(n58046), .Y(n64727) );
  NAND2xp5_ASAP7_75t_SL U60931 ( .A(n62562), .B(n62554), .Y(n57346) );
  XNOR2x1_ASAP7_75t_SL U60932 ( .A(n67496), .B(n67495), .Y(n67763) );
  BUFx6f_ASAP7_75t_SL U60933 ( .A(n3127), .Y(n59581) );
  NAND2xp5_ASAP7_75t_SL U60934 ( .A(n66876), .B(n57610), .Y(n57299) );
  INVx2_ASAP7_75t_SL U60935 ( .A(n67736), .Y(n58015) );
  INVx1_ASAP7_75t_SL U60936 ( .A(n68390), .Y(n68387) );
  NAND2xp5_ASAP7_75t_SL U60937 ( .A(n57301), .B(n57300), .Y(n68390) );
  NAND2xp5_ASAP7_75t_SL U60938 ( .A(n67701), .B(n67700), .Y(n57301) );
  OAI21xp5_ASAP7_75t_SL U60939 ( .A1(n59604), .A2(n67638), .B(n62689), .Y(
        n62699) );
  NAND2xp5_ASAP7_75t_SL U60940 ( .A(n67957), .B(n56830), .Y(n58267) );
  HB1xp67_ASAP7_75t_SL U60941 ( .A(n67407), .Y(n57303) );
  NAND2x2_ASAP7_75t_SL U60942 ( .A(n67914), .B(n66424), .Y(n59253) );
  INVx1_ASAP7_75t_SL U60943 ( .A(n64731), .Y(n64732) );
  INVx1_ASAP7_75t_SL U60944 ( .A(n64528), .Y(n64412) );
  NAND3xp33_ASAP7_75t_SL U60945 ( .A(n57306), .B(n64644), .C(n59298), .Y(
        n64645) );
  NAND3xp33_ASAP7_75t_SL U60946 ( .A(n58668), .B(n57107), .C(n59506), .Y(
        n57306) );
  AOI21xp5_ASAP7_75t_SL U60947 ( .A1(n58397), .A2(n67583), .B(n57307), .Y(
        n57672) );
  NAND3xp33_ASAP7_75t_SL U60948 ( .A(n67589), .B(n58017), .C(n57308), .Y(
        n57307) );
  NAND2xp5_ASAP7_75t_SL U60949 ( .A(n59436), .B(n67584), .Y(n57308) );
  OAI21x1_ASAP7_75t_SL U60950 ( .A1(n57382), .A2(n67468), .B(n57309), .Y(
        n58484) );
  NOR2x1_ASAP7_75t_SL U60951 ( .A(n64382), .B(n64381), .Y(n64438) );
  NAND2xp5_ASAP7_75t_SL U60952 ( .A(n77711), .B(n59589), .Y(n63206) );
  INVx1_ASAP7_75t_SL U60953 ( .A(n64952), .Y(n64628) );
  NAND2x1_ASAP7_75t_SL U60954 ( .A(n64373), .B(n57463), .Y(n64529) );
  NOR2x1_ASAP7_75t_SL U60955 ( .A(n56827), .B(n75958), .Y(n67327) );
  NAND2xp5_ASAP7_75t_SL U60956 ( .A(n59506), .B(n67807), .Y(n67808) );
  INVx2_ASAP7_75t_SL U60957 ( .A(n59588), .Y(n59592) );
  NAND2x1_ASAP7_75t_SL U60958 ( .A(n59464), .B(n59462), .Y(n62553) );
  INVx2_ASAP7_75t_SL U60959 ( .A(n67619), .Y(n57313) );
  INVx2_ASAP7_75t_SL U60960 ( .A(n67463), .Y(n67364) );
  BUFx5_ASAP7_75t_SL U60961 ( .A(n67922), .Y(n57314) );
  MAJx2_ASAP7_75t_SL U60962 ( .A(n68176), .B(n68178), .C(n68177), .Y(n68139)
         );
  AOI22xp5_ASAP7_75t_SL U60963 ( .A1(n67848), .A2(n67847), .B1(n67849), .B2(
        n57501), .Y(n68177) );
  O2A1O1Ixp5_ASAP7_75t_SL U60964 ( .A1(n59459), .A2(n57365), .B(n67060), .C(
        n58001), .Y(n58762) );
  NOR2x1_ASAP7_75t_SL U60965 ( .A(n56999), .B(n58720), .Y(n67329) );
  A2O1A1Ixp33_ASAP7_75t_SL U60966 ( .A1(n67169), .A2(n67178), .B(n67186), .C(
        n67187), .Y(n58635) );
  OAI21x1_ASAP7_75t_SL U60967 ( .A1(n57122), .A2(n62669), .B(n62668), .Y(
        n62672) );
  XNOR2x2_ASAP7_75t_SL U60968 ( .A(n67009), .B(n66866), .Y(n69138) );
  NAND2xp5_ASAP7_75t_SL U60969 ( .A(n64894), .B(n59481), .Y(n64368) );
  NOR2x1_ASAP7_75t_SL U60970 ( .A(n57896), .B(n57895), .Y(n59481) );
  NOR2x1p5_ASAP7_75t_SL U60971 ( .A(n58746), .B(n67917), .Y(n57373) );
  XNOR2x1_ASAP7_75t_SL U60972 ( .A(n59311), .B(n59312), .Y(n68073) );
  NAND3x1_ASAP7_75t_SL U60973 ( .A(n63659), .B(n59477), .C(n59458), .Y(n67947)
         );
  NOR2x1_ASAP7_75t_SL U60974 ( .A(n56993), .B(n68093), .Y(n68105) );
  INVx1_ASAP7_75t_SL U60975 ( .A(n65054), .Y(n64927) );
  NAND2x1_ASAP7_75t_SL U60976 ( .A(n57380), .B(n58492), .Y(n59241) );
  NOR2xp33_ASAP7_75t_SL U60977 ( .A(n53473), .B(n71064), .Y(n57317) );
  BUFx3_ASAP7_75t_SL U60978 ( .A(n67898), .Y(n57410) );
  XNOR2xp5_ASAP7_75t_SL U60979 ( .A(n67773), .B(n67774), .Y(n67775) );
  INVx1_ASAP7_75t_SL U60980 ( .A(n57320), .Y(n57319) );
  NOR2x1_ASAP7_75t_SL U60981 ( .A(n67824), .B(n67434), .Y(n57320) );
  NAND2x1p5_ASAP7_75t_SL U60982 ( .A(n58274), .B(n62575), .Y(n58272) );
  INVx1_ASAP7_75t_SL U60983 ( .A(n59314), .Y(n57323) );
  INVx1_ASAP7_75t_SL U60984 ( .A(n67438), .Y(n57324) );
  AOI21xp5_ASAP7_75t_SL U60985 ( .A1(n57324), .A2(n57323), .B(n57469), .Y(
        n67836) );
  NOR2x1_ASAP7_75t_SL U60986 ( .A(n58508), .B(n59407), .Y(n59135) );
  O2A1O1Ixp5_ASAP7_75t_SL U60987 ( .A1(n57484), .A2(n58901), .B(n56975), .C(
        n53197), .Y(n64077) );
  NAND2xp5_ASAP7_75t_SL U60988 ( .A(n59557), .B(n56861), .Y(n57327) );
  NAND2x1_ASAP7_75t_SL U60989 ( .A(n57328), .B(n56976), .Y(n67480) );
  INVx1_ASAP7_75t_SL U60990 ( .A(n58197), .Y(n57328) );
  OAI21xp5_ASAP7_75t_SL U60991 ( .A1(n59513), .A2(n58439), .B(n62894), .Y(
        n62896) );
  NOR2x1_ASAP7_75t_SL U60992 ( .A(n59581), .B(n59070), .Y(n62658) );
  OAI21x1_ASAP7_75t_SL U60993 ( .A1(n58775), .A2(n67338), .B(n56973), .Y(
        n67344) );
  INVx1_ASAP7_75t_SL U60994 ( .A(n56974), .Y(n63081) );
  NOR2x1_ASAP7_75t_SL U60995 ( .A(n62562), .B(n59336), .Y(n62569) );
  NAND2xp5_ASAP7_75t_SL U60996 ( .A(n59148), .B(n57330), .Y(n59147) );
  NAND3xp33_ASAP7_75t_SL U60997 ( .A(n59149), .B(n58155), .C(n56991), .Y(
        n57330) );
  NAND2x1_ASAP7_75t_SL U60998 ( .A(n59464), .B(n59566), .Y(n62564) );
  NAND2xp5_ASAP7_75t_SL U60999 ( .A(n59614), .B(n67288), .Y(n62628) );
  NAND2x1p5_ASAP7_75t_SL U61000 ( .A(n66411), .B(n57958), .Y(n59436) );
  OAI21xp5_ASAP7_75t_SL U61001 ( .A1(n67802), .A2(n67803), .B(n67776), .Y(
        n58896) );
  XNOR2x1_ASAP7_75t_SL U61002 ( .A(n67065), .B(n67173), .Y(n67199) );
  OAI21xp5_ASAP7_75t_SL U61003 ( .A1(n68106), .A2(n68105), .B(n68151), .Y(
        n57334) );
  NAND2x1_ASAP7_75t_SL U61004 ( .A(n58724), .B(n58725), .Y(n57733) );
  NAND2xp5_ASAP7_75t_SL U61005 ( .A(n62807), .B(n57118), .Y(n59234) );
  OAI21xp5_ASAP7_75t_SL U61006 ( .A1(n62634), .A2(n62593), .B(n76627), .Y(
        n62807) );
  OAI21xp5_ASAP7_75t_SL U61007 ( .A1(n62757), .A2(n59654), .B(n53517), .Y(
        n58057) );
  INVx1_ASAP7_75t_SL U61008 ( .A(n59332), .Y(n68013) );
  NAND2xp5_ASAP7_75t_SL U61009 ( .A(n68581), .B(n68580), .Y(n68915) );
  INVx1_ASAP7_75t_SL U61010 ( .A(n68420), .Y(n68423) );
  INVx1_ASAP7_75t_SL U61011 ( .A(n59186), .Y(n59185) );
  NAND2x1p5_ASAP7_75t_SL U61012 ( .A(n58747), .B(n58138), .Y(n67731) );
  XNOR2xp5_ASAP7_75t_SL U61013 ( .A(n67145), .B(n67143), .Y(n67098) );
  AOI22xp5_ASAP7_75t_SL U61014 ( .A1(n67096), .A2(n67097), .B1(n67095), .B2(
        n56967), .Y(n67145) );
  NAND2xp5_ASAP7_75t_SL U61015 ( .A(n78003), .B(n59589), .Y(n58466) );
  NOR2x1_ASAP7_75t_SL U61016 ( .A(n58466), .B(n62621), .Y(n59419) );
  INVx1_ASAP7_75t_SL U61017 ( .A(n68221), .Y(n65006) );
  XNOR2xp5_ASAP7_75t_SL U61018 ( .A(n57580), .B(n57581), .Y(n68034) );
  NAND2x1_ASAP7_75t_SL U61019 ( .A(n59572), .B(n59394), .Y(n57665) );
  XNOR2x1_ASAP7_75t_SL U61020 ( .A(n68453), .B(n58976), .Y(n68498) );
  NOR2x1_ASAP7_75t_SL U61021 ( .A(n57325), .B(n66479), .Y(n66498) );
  NAND2xp5_ASAP7_75t_SL U61022 ( .A(n66700), .B(n66782), .Y(n68022) );
  NAND2xp5_ASAP7_75t_SL U61023 ( .A(n59508), .B(n59456), .Y(n66700) );
  INVx1_ASAP7_75t_SL U61024 ( .A(n59364), .Y(n64716) );
  OAI21xp5_ASAP7_75t_SL U61025 ( .A1(n58039), .A2(n57337), .B(n64677), .Y(
        n59364) );
  INVx1_ASAP7_75t_SL U61026 ( .A(n64045), .Y(n57337) );
  NAND2xp5_ASAP7_75t_SL U61027 ( .A(n58323), .B(n68213), .Y(n67956) );
  INVx1_ASAP7_75t_SL U61028 ( .A(n68449), .Y(n57338) );
  MAJIxp5_ASAP7_75t_SL U61029 ( .A(n68390), .B(n68389), .C(n68388), .Y(n68449)
         );
  NOR2x1p5_ASAP7_75t_SL U61030 ( .A(n65104), .B(n65101), .Y(n64751) );
  NOR2x1p5_ASAP7_75t_SL U61031 ( .A(n68568), .B(n68569), .Y(n68860) );
  XNOR2x2_ASAP7_75t_SL U61032 ( .A(n67791), .B(n57726), .Y(n68039) );
  NOR2x1_ASAP7_75t_SL U61033 ( .A(n57260), .B(n67640), .Y(n58674) );
  A2O1A1Ixp33_ASAP7_75t_SL U61034 ( .A1(n59518), .A2(n67435), .B(n59504), .C(
        n57342), .Y(n67437) );
  NAND2xp5_ASAP7_75t_SL U61035 ( .A(n59504), .B(n68602), .Y(n57342) );
  INVx11_ASAP7_75t_SL U61036 ( .A(n59598), .Y(n59596) );
  INVx2_ASAP7_75t_SL U61037 ( .A(n58789), .Y(n67244) );
  INVx3_ASAP7_75t_SL U61038 ( .A(n67610), .Y(n67288) );
  BUFx6f_ASAP7_75t_SL U61039 ( .A(n68012), .Y(n59515) );
  INVx1_ASAP7_75t_SL U61040 ( .A(n58997), .Y(n58999) );
  INVx1_ASAP7_75t_SL U61041 ( .A(n63677), .Y(n58002) );
  NAND2x1p5_ASAP7_75t_SL U61042 ( .A(n57994), .B(n58263), .Y(n63669) );
  NAND2x1_ASAP7_75t_SL U61043 ( .A(n63669), .B(n59473), .Y(n63670) );
  NAND3xp33_ASAP7_75t_SL U61044 ( .A(n67910), .B(n59332), .C(n59132), .Y(
        n68001) );
  NAND2xp5_ASAP7_75t_SL U61045 ( .A(n57179), .B(n67444), .Y(n67445) );
  BUFx3_ASAP7_75t_SL U61046 ( .A(n58408), .Y(n57484) );
  XOR2xp5_ASAP7_75t_SL U61047 ( .A(n68530), .B(n68528), .Y(n68509) );
  XNOR2xp5_ASAP7_75t_SL U61048 ( .A(n68508), .B(n68507), .Y(n68530) );
  NAND3x1_ASAP7_75t_SL U61049 ( .A(n57959), .B(n59488), .C(n75378), .Y(n57379)
         );
  NAND2x1_ASAP7_75t_SL U61050 ( .A(n57379), .B(n53624), .Y(n57958) );
  A2O1A1Ixp33_ASAP7_75t_SL U61051 ( .A1(n57414), .A2(n59648), .B(n57344), .C(
        n59596), .Y(n66760) );
  NOR2x1_ASAP7_75t_SL U61052 ( .A(n56978), .B(n57414), .Y(n57344) );
  NOR2x1p5_ASAP7_75t_SL U61053 ( .A(n58084), .B(n62808), .Y(n62806) );
  NOR2x1_ASAP7_75t_SL U61054 ( .A(n57346), .B(n57345), .Y(n58764) );
  INVx5_ASAP7_75t_SL U61055 ( .A(n57781), .Y(n59516) );
  OAI21x1_ASAP7_75t_SL U61056 ( .A1(n57349), .A2(n67253), .B(n58875), .Y(
        n59279) );
  NOR2x1_ASAP7_75t_SL U61057 ( .A(n57315), .B(n67841), .Y(n57349) );
  OAI21xp33_ASAP7_75t_SRAM U61058 ( .A1(n59599), .A2(n59516), .B(n57350), .Y(
        n66797) );
  NAND2xp5_ASAP7_75t_SL U61059 ( .A(n59599), .B(n67741), .Y(n57350) );
  NAND2xp5_ASAP7_75t_SL U61060 ( .A(n67729), .B(n67728), .Y(n67734) );
  INVx1_ASAP7_75t_SL U61061 ( .A(n67734), .Y(n58036) );
  INVx2_ASAP7_75t_SL U61062 ( .A(n63669), .Y(n63667) );
  NAND2x1p5_ASAP7_75t_SL U61063 ( .A(n59533), .B(n63667), .Y(n63671) );
  A2O1A1Ixp33_ASAP7_75t_SL U61064 ( .A1(n67637), .A2(n57221), .B(n67635), .C(
        n68002), .Y(n58749) );
  XNOR2xp5_ASAP7_75t_SL U61065 ( .A(n59601), .B(n57169), .Y(n68002) );
  NOR2x1_ASAP7_75t_SL U61066 ( .A(n64499), .B(n64500), .Y(n65041) );
  NAND2xp5_ASAP7_75t_SL U61067 ( .A(n57351), .B(n57822), .Y(n62695) );
  OAI21xp5_ASAP7_75t_SL U61068 ( .A1(n68097), .A2(n75903), .B(n59503), .Y(
        n57351) );
  BUFx2_ASAP7_75t_SL U61069 ( .A(n62573), .Y(n57353) );
  NAND2xp5_ASAP7_75t_SL U61070 ( .A(n59571), .B(n60595), .Y(n61539) );
  INVx2_ASAP7_75t_SL U61071 ( .A(n58342), .Y(n58343) );
  HB1xp67_ASAP7_75t_SL U61072 ( .A(n66907), .Y(n57354) );
  INVx8_ASAP7_75t_SL U61073 ( .A(n59597), .Y(n59599) );
  AOI22xp5_ASAP7_75t_SL U61074 ( .A1(n68086), .A2(n64956), .B1(n64955), .B2(
        n57478), .Y(n65010) );
  XNOR2x2_ASAP7_75t_SL U61075 ( .A(n59609), .B(n53288), .Y(n67719) );
  NAND2xp5_ASAP7_75t_SL U61076 ( .A(n57355), .B(n58931), .Y(n67358) );
  XNOR2x1_ASAP7_75t_SL U61077 ( .A(n58348), .B(n57357), .Y(n68308) );
  XNOR2x1_ASAP7_75t_SL U61078 ( .A(n57426), .B(n68146), .Y(n57357) );
  OAI22x1_ASAP7_75t_SL U61079 ( .A1(n64374), .A2(n57508), .B1(n58131), .B2(
        n57047), .Y(n63816) );
  INVx4_ASAP7_75t_SL U61080 ( .A(n58273), .Y(n58275) );
  OAI21x1_ASAP7_75t_SL U61081 ( .A1(n57657), .A2(n58953), .B(n67036), .Y(
        n67067) );
  AO21x1_ASAP7_75t_SL U61082 ( .A1(n68101), .A2(n59409), .B(n68095), .Y(n65044) );
  BUFx6f_ASAP7_75t_SL U61083 ( .A(n66418), .Y(n59458) );
  INVx4_ASAP7_75t_SL U61084 ( .A(n57768), .Y(n58788) );
  INVx2_ASAP7_75t_SL U61085 ( .A(n57065), .Y(n68413) );
  NAND2xp5_ASAP7_75t_SL U61086 ( .A(n59124), .B(n59123), .Y(n67884) );
  OAI21xp5_ASAP7_75t_SL U61087 ( .A1(n66384), .A2(n57336), .B(n57078), .Y(
        n66245) );
  NAND2x1_ASAP7_75t_SL U61088 ( .A(n53399), .B(n59243), .Y(n68576) );
  BUFx3_ASAP7_75t_SL U61089 ( .A(n58872), .Y(n58871) );
  NOR2x1_ASAP7_75t_SL U61090 ( .A(n56996), .B(n57361), .Y(n67714) );
  XNOR2x2_ASAP7_75t_SL U61091 ( .A(n59478), .B(n68077), .Y(n58348) );
  NOR2x1_ASAP7_75t_SL U61092 ( .A(n67974), .B(n67478), .Y(n57363) );
  NOR2x1_ASAP7_75t_SL U61093 ( .A(n67719), .B(n57156), .Y(n57364) );
  NOR2x1p5_ASAP7_75t_SL U61094 ( .A(n68575), .B(n58344), .Y(n68850) );
  NAND2x2_ASAP7_75t_SL U61095 ( .A(n3127), .B(n1967), .Y(n61921) );
  NAND2xp5_ASAP7_75t_SL U61096 ( .A(n62993), .B(n57367), .Y(n57383) );
  XOR2xp5_ASAP7_75t_SL U61097 ( .A(n62995), .B(n62994), .Y(n57367) );
  INVx1_ASAP7_75t_SL U61098 ( .A(n67841), .Y(n68418) );
  OAI22xp5_ASAP7_75t_SL U61099 ( .A1(n57801), .A2(n57800), .B1(n67798), .B2(
        n67800), .Y(n67777) );
  NOR2xp33_ASAP7_75t_SL U61100 ( .A(n63173), .B(n63172), .Y(n57995) );
  INVx1_ASAP7_75t_SL U61101 ( .A(n63622), .Y(n63226) );
  A2O1A1Ixp33_ASAP7_75t_SL U61102 ( .A1(n57368), .A2(n63086), .B(n64426), .C(
        n63085), .Y(n63153) );
  NAND2xp5_ASAP7_75t_SL U61103 ( .A(n76028), .B(n63082), .Y(n57368) );
  AND2x4_ASAP7_75t_SL U61104 ( .A(n59286), .B(n59285), .Y(n68146) );
  NAND2xp5_ASAP7_75t_SL U61105 ( .A(n68085), .B(n58025), .Y(n58068) );
  NAND2xp5_ASAP7_75t_SL U61106 ( .A(n59604), .B(n57274), .Y(n63079) );
  HB1xp67_ASAP7_75t_SL U61107 ( .A(n69147), .Y(n57369) );
  BUFx3_ASAP7_75t_SL U61108 ( .A(n67976), .Y(n57371) );
  NAND2x1_ASAP7_75t_SL U61109 ( .A(n58051), .B(n58050), .Y(n58691) );
  AND2x4_ASAP7_75t_SL U61110 ( .A(n65021), .B(n65020), .Y(n58143) );
  NAND2x1_ASAP7_75t_SL U61111 ( .A(n61916), .B(n57838), .Y(n64506) );
  INVx2_ASAP7_75t_SL U61112 ( .A(n61920), .Y(n61925) );
  NOR2x1_ASAP7_75t_SL U61113 ( .A(n61925), .B(n61924), .Y(n63653) );
  NOR2xp33_ASAP7_75t_SL U61114 ( .A(n57257), .B(n58934), .Y(n58933) );
  AOI21x1_ASAP7_75t_SL U61115 ( .A1(n66636), .A2(n74781), .B(n66638), .Y(
        n67410) );
  XNOR2xp5_ASAP7_75t_SL U61116 ( .A(n67761), .B(n57370), .Y(n67762) );
  AOI21xp5_ASAP7_75t_SL U61117 ( .A1(n59177), .A2(n67760), .B(n67759), .Y(
        n57370) );
  NAND2x1p5_ASAP7_75t_SL U61118 ( .A(n57553), .B(n59145), .Y(n68011) );
  NAND2x2_ASAP7_75t_SL U61119 ( .A(n66623), .B(n59204), .Y(n67833) );
  XNOR2x1_ASAP7_75t_SL U61120 ( .A(n67935), .B(n67934), .Y(n57372) );
  AOI21x1_ASAP7_75t_SL U61121 ( .A1(n58746), .A2(n57453), .B(n57373), .Y(
        n58488) );
  NAND2x1_ASAP7_75t_SL U61122 ( .A(n57386), .B(n57440), .Y(n57374) );
  O2A1O1Ixp5_ASAP7_75t_SL U61123 ( .A1(n59654), .A2(n66451), .B(n59578), .C(
        n59044), .Y(n57883) );
  AOI211x1_ASAP7_75t_SL U61124 ( .A1(n64607), .A2(n67608), .B(n58640), .C(
        n56835), .Y(n67816) );
  NOR2x1_ASAP7_75t_SL U61125 ( .A(n62690), .B(n59609), .Y(n62685) );
  AOI21xp5_ASAP7_75t_SL U61126 ( .A1(n68577), .A2(n68578), .B(n68576), .Y(
        n68584) );
  NAND2x1_ASAP7_75t_SL U61127 ( .A(n57181), .B(n62611), .Y(n67909) );
  NOR2x1_ASAP7_75t_SL U61128 ( .A(n66816), .B(n66907), .Y(n67040) );
  MAJIxp5_ASAP7_75t_SL U61129 ( .A(n68547), .B(n68548), .C(n68546), .Y(n66907)
         );
  NAND2x1_ASAP7_75t_SL U61130 ( .A(n74788), .B(n59400), .Y(n59353) );
  OR2x6_ASAP7_75t_SL U61131 ( .A(n67860), .B(n59412), .Y(n67228) );
  XNOR2x1_ASAP7_75t_SL U61132 ( .A(n59330), .B(n68329), .Y(n59329) );
  NAND2xp5_ASAP7_75t_SL U61133 ( .A(n57064), .B(n64891), .Y(n65026) );
  XNOR2xp5_ASAP7_75t_SL U61134 ( .A(n59088), .B(n64640), .Y(n57378) );
  NAND3xp33_ASAP7_75t_SL U61135 ( .A(n59507), .B(n59470), .C(n59608), .Y(
        n66719) );
  AOI21xp5_ASAP7_75t_SL U61136 ( .A1(n59503), .A2(n75906), .B(n63064), .Y(
        n63143) );
  XNOR2x1_ASAP7_75t_SL U61137 ( .A(n67642), .B(n67802), .Y(n58792) );
  AOI21xp5_ASAP7_75t_SL U61138 ( .A1(n59508), .A2(n67920), .B(n63839), .Y(
        n63841) );
  NAND2xp5_ASAP7_75t_SL U61139 ( .A(n75947), .B(n67902), .Y(n67903) );
  INVx1_ASAP7_75t_SL U61140 ( .A(n68480), .Y(n68481) );
  XOR2xp5_ASAP7_75t_SL U61141 ( .A(n57045), .B(n57400), .Y(n68278) );
  XOR2xp5_ASAP7_75t_SL U61142 ( .A(n58363), .B(n67896), .Y(n57381) );
  NOR2x1_ASAP7_75t_SL U61143 ( .A(n59567), .B(n62519), .Y(n60790) );
  NOR2x1_ASAP7_75t_SL U61144 ( .A(n68082), .B(n68083), .Y(n57382) );
  XOR2xp5_ASAP7_75t_SL U61145 ( .A(n68512), .B(n68510), .Y(n57931) );
  XNOR2xp5_ASAP7_75t_SL U61146 ( .A(n68427), .B(n68426), .Y(n68512) );
  XNOR2xp5_ASAP7_75t_SL U61147 ( .A(n63163), .B(n63162), .Y(n57597) );
  NAND2xp5_ASAP7_75t_SL U61148 ( .A(n62994), .B(n62995), .Y(n57384) );
  NAND2xp5_ASAP7_75t_SL U61149 ( .A(n67901), .B(n58499), .Y(n59130) );
  NAND2xp5_ASAP7_75t_SL U61150 ( .A(n57385), .B(n57548), .Y(n58499) );
  NAND2xp5_ASAP7_75t_SL U61151 ( .A(n58402), .B(n67920), .Y(n57385) );
  NAND2xp5_ASAP7_75t_SL U61152 ( .A(n68174), .B(n68169), .Y(n68175) );
  NAND3xp33_ASAP7_75t_SL U61153 ( .A(n58804), .B(n67808), .C(n67810), .Y(
        n57386) );
  XNOR2x1_ASAP7_75t_SL U61154 ( .A(n59511), .B(n58865), .Y(n67968) );
  NAND2xp5_ASAP7_75t_SL U61155 ( .A(n60918), .B(n58251), .Y(n58250) );
  NOR2x1_ASAP7_75t_SL U61156 ( .A(n60599), .B(n57387), .Y(n60918) );
  NAND2xp5_ASAP7_75t_SL U61157 ( .A(n57389), .B(n57388), .Y(n57387) );
  INVx1_ASAP7_75t_SL U61158 ( .A(n58930), .Y(n67498) );
  NAND2xp5_ASAP7_75t_SL U61159 ( .A(n56992), .B(n67462), .Y(n57390) );
  INVx1_ASAP7_75t_SL U61160 ( .A(n67461), .Y(n57391) );
  AOI21xp5_ASAP7_75t_SL U61161 ( .A1(n57392), .A2(n57101), .B(n67330), .Y(
        n59201) );
  INVx1_ASAP7_75t_SL U61162 ( .A(n62581), .Y(n62556) );
  XNOR2xp5_ASAP7_75t_SL U61163 ( .A(n57393), .B(n64910), .Y(n64991) );
  XNOR2xp5_ASAP7_75t_SL U61164 ( .A(n64992), .B(n64993), .Y(n57393) );
  NAND2x1_ASAP7_75t_SL U61165 ( .A(n59034), .B(n63829), .Y(n64048) );
  INVx4_ASAP7_75t_SL U61166 ( .A(n59508), .Y(n67481) );
  INVx1_ASAP7_75t_SL U61167 ( .A(n64875), .Y(n64874) );
  OR2x2_ASAP7_75t_SL U61168 ( .A(n64561), .B(n64560), .Y(n64875) );
  INVx2_ASAP7_75t_SL U61169 ( .A(n58455), .Y(n57834) );
  OAI21x1_ASAP7_75t_SL U61170 ( .A1(n57396), .A2(n57395), .B(n59310), .Y(
        n58897) );
  INVx1_ASAP7_75t_SL U61171 ( .A(n62607), .Y(n57395) );
  NOR2x1_ASAP7_75t_SL U61172 ( .A(n59542), .B(n59400), .Y(n57396) );
  HB1xp67_ASAP7_75t_SL U61173 ( .A(n64509), .Y(n57397) );
  NAND2xp5_ASAP7_75t_SL U61174 ( .A(n57912), .B(n75904), .Y(n58456) );
  INVx1_ASAP7_75t_SL U61175 ( .A(n67519), .Y(n67521) );
  A2O1A1Ixp33_ASAP7_75t_SL U61176 ( .A1(n53288), .A2(n57110), .B(n67417), .C(
        n57399), .Y(n67418) );
  NAND2xp5_ASAP7_75t_SL U61177 ( .A(n67807), .B(n59506), .Y(n57399) );
  AND2x2_ASAP7_75t_SL U61178 ( .A(n59123), .B(n67247), .Y(n67229) );
  OR2x6_ASAP7_75t_SL U61179 ( .A(n58069), .B(n67704), .Y(n58336) );
  NOR2x1_ASAP7_75t_SL U61180 ( .A(n59582), .B(n76679), .Y(n67420) );
  AOI21x1_ASAP7_75t_SL U61181 ( .A1(n67559), .A2(n57163), .B(n59164), .Y(
        n68399) );
  INVx4_ASAP7_75t_SL U61182 ( .A(n59102), .Y(n68119) );
  INVx2_ASAP7_75t_SL U61183 ( .A(n59555), .Y(n76627) );
  MAJIxp5_ASAP7_75t_SL U61184 ( .A(n68135), .B(n68133), .C(n68132), .Y(n68136)
         );
  NOR2x1_ASAP7_75t_SL U61185 ( .A(n59654), .B(n66249), .Y(n58724) );
  XOR2xp5_ASAP7_75t_SL U61186 ( .A(n64494), .B(n57437), .Y(n57401) );
  NOR2x1_ASAP7_75t_SL U61187 ( .A(n58199), .B(n58198), .Y(n57569) );
  NOR2x1_ASAP7_75t_SL U61188 ( .A(n59533), .B(n53615), .Y(n59473) );
  INVx1_ASAP7_75t_SL U61189 ( .A(n67012), .Y(n67013) );
  AND2x2_ASAP7_75t_SL U61190 ( .A(n57797), .B(n58702), .Y(n57795) );
  NOR2x1p5_ASAP7_75t_SL U61191 ( .A(n59548), .B(n66636), .Y(n66286) );
  NAND2x1p5_ASAP7_75t_SL U61192 ( .A(n66258), .B(n78167), .Y(n66269) );
  INVx1_ASAP7_75t_SL U61193 ( .A(n1868), .Y(n75848) );
  XNOR2xp5_ASAP7_75t_SL U61194 ( .A(n57257), .B(n59658), .Y(n58059) );
  AOI21xp5_ASAP7_75t_SL U61195 ( .A1(n58223), .A2(n58746), .B(n57403), .Y(
        n66647) );
  AOI22xp5_ASAP7_75t_SL U61196 ( .A1(n67564), .A2(n59648), .B1(n66623), .B2(
        n59649), .Y(n57403) );
  INVx1_ASAP7_75t_SL U61197 ( .A(n67477), .Y(n67478) );
  XNOR2xp5_ASAP7_75t_SL U61198 ( .A(n68443), .B(n57406), .Y(n57987) );
  MAJIxp5_ASAP7_75t_SL U61199 ( .A(n66936), .B(n66935), .C(n68406), .Y(n68443)
         );
  INVx1_ASAP7_75t_SL U61200 ( .A(n68442), .Y(n57406) );
  O2A1O1Ixp5_ASAP7_75t_SL U61201 ( .A1(n66863), .A2(n66864), .B(n67077), .C(
        n67035), .Y(n58952) );
  INVx4_ASAP7_75t_SL U61202 ( .A(n59445), .Y(n62562) );
  INVxp33_ASAP7_75t_SRAM U61203 ( .A(n66398), .Y(n57408) );
  NAND2x1_ASAP7_75t_SL U61204 ( .A(n65072), .B(n57184), .Y(n66398) );
  NOR2x1p5_ASAP7_75t_SL U61205 ( .A(n58974), .B(n67494), .Y(n67537) );
  XNOR2x1_ASAP7_75t_SL U61206 ( .A(n67491), .B(n67537), .Y(n67291) );
  AO21x2_ASAP7_75t_SL U61207 ( .A1(n68015), .A2(n57709), .B(n67927), .Y(n58454) );
  XOR2x1_ASAP7_75t_SL U61208 ( .A(n57613), .B(n58454), .Y(n57612) );
  INVx2_ASAP7_75t_SL U61209 ( .A(n66810), .Y(n68485) );
  XNOR2x1_ASAP7_75t_SL U61210 ( .A(n58486), .B(n68485), .Y(n58942) );
  INVx1_ASAP7_75t_SL U61211 ( .A(n66296), .Y(n58944) );
  OAI21xp5_ASAP7_75t_SL U61212 ( .A1(n67609), .A2(n62786), .B(n62785), .Y(
        n62787) );
  OAI21xp5_ASAP7_75t_SL U61213 ( .A1(n59513), .A2(n67463), .B(n58523), .Y(
        n62785) );
  NAND2xp5_ASAP7_75t_SL U61214 ( .A(n59514), .B(n59466), .Y(n59072) );
  NAND2xp5_ASAP7_75t_SL U61215 ( .A(n57094), .B(n67391), .Y(n58911) );
  NAND2x1p5_ASAP7_75t_SL U61216 ( .A(n64038), .B(n64037), .Y(n67636) );
  INVx1_ASAP7_75t_SL U61217 ( .A(n57412), .Y(n57411) );
  NAND2xp5_ASAP7_75t_SL U61218 ( .A(n67955), .B(n67948), .Y(n67949) );
  XNOR2xp5_ASAP7_75t_SL U61219 ( .A(n57413), .B(n64903), .Y(n64994) );
  XOR2xp5_ASAP7_75t_SL U61220 ( .A(n65050), .B(n65051), .Y(n57413) );
  NAND2xp5_ASAP7_75t_SL U61221 ( .A(n59664), .B(n68101), .Y(n67600) );
  OAI21xp5_ASAP7_75t_SL U61222 ( .A1(n58015), .A2(n67826), .B(n66929), .Y(
        n66931) );
  XNOR2x1_ASAP7_75t_SL U61223 ( .A(n57415), .B(n64982), .Y(n64986) );
  XNOR2x1_ASAP7_75t_SL U61224 ( .A(n64981), .B(n57416), .Y(n57415) );
  INVx2_ASAP7_75t_SL U61225 ( .A(n64989), .Y(n57416) );
  NOR2x1_ASAP7_75t_SL U61226 ( .A(n59654), .B(n62658), .Y(n58883) );
  NOR2x1_ASAP7_75t_SL U61227 ( .A(n53488), .B(n58883), .Y(n62631) );
  XNOR2xp5_ASAP7_75t_SL U61228 ( .A(n59513), .B(n59616), .Y(n63170) );
  XNOR2xp5_ASAP7_75t_SL U61229 ( .A(n68552), .B(n57418), .Y(n68592) );
  NAND2xp33_ASAP7_75t_SRAM U61230 ( .A(n68086), .B(n64487), .Y(n64460) );
  AOI21xp5_ASAP7_75t_SL U61231 ( .A1(n75900), .A2(n53320), .B(n64459), .Y(
        n64487) );
  OR2x2_ASAP7_75t_SL U61232 ( .A(n59262), .B(n59261), .Y(n66637) );
  O2A1O1Ixp5_ASAP7_75t_SL U61233 ( .A1(n67638), .A2(n56827), .B(n62843), .C(
        n57159), .Y(n62844) );
  NAND2xp5_ASAP7_75t_SL U61234 ( .A(n59470), .B(n59615), .Y(n62921) );
  INVx5_ASAP7_75t_SL U61235 ( .A(n57662), .Y(n67432) );
  NOR2x1_ASAP7_75t_SL U61236 ( .A(n59551), .B(n57116), .Y(n63191) );
  NAND2x1_ASAP7_75t_SL U61237 ( .A(n68349), .B(n68350), .Y(n68737) );
  NAND2xp5_ASAP7_75t_SL U61238 ( .A(n57179), .B(n67610), .Y(n67611) );
  OAI21x1_ASAP7_75t_SL U61239 ( .A1(n53271), .A2(n58431), .B(n67611), .Y(
        n68003) );
  INVx3_ASAP7_75t_SL U61240 ( .A(n57924), .Y(n59508) );
  NOR2x1_ASAP7_75t_SL U61241 ( .A(n64229), .B(n60790), .Y(n62588) );
  AOI22x1_ASAP7_75t_SL U61242 ( .A1(n62588), .A2(n57316), .B1(n78005), .B2(
        n57122), .Y(n62880) );
  NOR2x1_ASAP7_75t_SL U61243 ( .A(n56993), .B(n67367), .Y(n67374) );
  BUFx2_ASAP7_75t_SL U61244 ( .A(n59452), .Y(n57478) );
  OAI21xp5_ASAP7_75t_SL U61245 ( .A1(n59596), .A2(n68087), .B(n67312), .Y(
        n67369) );
  NOR2x1_ASAP7_75t_SL U61246 ( .A(n58732), .B(n58731), .Y(n68722) );
  OAI21xp5_ASAP7_75t_SL U61247 ( .A1(n62730), .A2(n62729), .B(n63058), .Y(
        n62735) );
  NAND2x1p5_ASAP7_75t_SL U61248 ( .A(n67909), .B(n67908), .Y(n68012) );
  NAND2x1p5_ASAP7_75t_SL U61249 ( .A(n67346), .B(n67345), .Y(n67347) );
  NAND2xp5_ASAP7_75t_SL U61250 ( .A(n59464), .B(n59566), .Y(n59322) );
  NAND2xp5_ASAP7_75t_SL U61251 ( .A(n68482), .B(n68481), .Y(n68484) );
  NAND2x1p5_ASAP7_75t_SL U61252 ( .A(n57670), .B(n57998), .Y(n67811) );
  OAI21x1_ASAP7_75t_SL U61253 ( .A1(n58484), .A2(n58653), .B(n58652), .Y(
        n57426) );
  NAND2x1_ASAP7_75t_SL U61254 ( .A(n57427), .B(n57611), .Y(n64037) );
  NOR2x1p5_ASAP7_75t_SL U61255 ( .A(n57480), .B(n57697), .Y(n62579) );
  AOI22x1_ASAP7_75t_SL U61256 ( .A1(n67387), .A2(n68414), .B1(n58746), .B2(
        n67290), .Y(n67491) );
  NOR2x1_ASAP7_75t_SL U61257 ( .A(n67323), .B(n67893), .Y(n58662) );
  NOR2x1p5_ASAP7_75t_SL U61258 ( .A(n61922), .B(n61925), .Y(n59276) );
  INVx2_ASAP7_75t_SL U61259 ( .A(n67635), .Y(n58759) );
  NOR2x1_ASAP7_75t_SL U61260 ( .A(n59578), .B(n59045), .Y(n59044) );
  BUFx3_ASAP7_75t_SL U61261 ( .A(n2186), .Y(n59445) );
  AOI22x1_ASAP7_75t_SL U61262 ( .A1(n59100), .A2(n67556), .B1(n67555), .B2(
        n57067), .Y(n68401) );
  NAND2xp5_ASAP7_75t_SL U61263 ( .A(n59505), .B(n59595), .Y(n67807) );
  INVx1_ASAP7_75t_SL U61264 ( .A(n67594), .Y(n57429) );
  NAND3xp33_ASAP7_75t_SL U61265 ( .A(n75032), .B(n67641), .C(n57429), .Y(
        n57886) );
  NOR2x2_ASAP7_75t_SL U61266 ( .A(n67645), .B(n67303), .Y(n59444) );
  AND2x4_ASAP7_75t_SL U61267 ( .A(n67244), .B(n64928), .Y(n67709) );
  NAND2x2_ASAP7_75t_SL U61268 ( .A(n59054), .B(n67738), .Y(n67914) );
  MAJIxp5_ASAP7_75t_SL U61269 ( .A(n63029), .B(n63027), .C(n63025), .Y(n63044)
         );
  XNOR2xp5_ASAP7_75t_SL U61270 ( .A(n57430), .B(n62697), .Y(n63029) );
  INVx1_ASAP7_75t_SL U61271 ( .A(n58067), .Y(n57430) );
  OAI21xp5_ASAP7_75t_SL U61272 ( .A1(n75947), .A2(n57494), .B(n66400), .Y(
        n66401) );
  NAND2xp5_ASAP7_75t_SL U61273 ( .A(n57431), .B(n68017), .Y(n68020) );
  NOR2x1_ASAP7_75t_SL U61274 ( .A(n59506), .B(n63083), .Y(n68017) );
  NAND2xp5_ASAP7_75t_SL U61275 ( .A(n57433), .B(n57432), .Y(n57431) );
  NAND2xp5_ASAP7_75t_SL U61276 ( .A(n59505), .B(n68019), .Y(n57433) );
  NAND2xp5_ASAP7_75t_SL U61277 ( .A(n59609), .B(n76049), .Y(n58695) );
  NAND2xp5_ASAP7_75t_SL U61278 ( .A(n69231), .B(n69233), .Y(n69232) );
  INVx1_ASAP7_75t_SL U61279 ( .A(n67987), .Y(n67988) );
  NAND3xp33_ASAP7_75t_SL U61280 ( .A(n58692), .B(n58693), .C(n68139), .Y(
        n57861) );
  OA21x2_ASAP7_75t_SL U61281 ( .A1(n66448), .A2(n66447), .B(n57435), .Y(n67112) );
  NAND2x1_ASAP7_75t_SL U61282 ( .A(n74993), .B(n74992), .Y(n65122) );
  AND2x4_ASAP7_75t_SL U61283 ( .A(n59138), .B(n67641), .Y(n67715) );
  AND2x4_ASAP7_75t_SL U61284 ( .A(n59239), .B(n67586), .Y(n59205) );
  NAND2x2_ASAP7_75t_SL U61285 ( .A(n59206), .B(n59205), .Y(n66623) );
  INVx1_ASAP7_75t_SL U61286 ( .A(n64566), .Y(n57437) );
  INVx8_ASAP7_75t_SL U61287 ( .A(n58275), .Y(n76028) );
  OAI21x1_ASAP7_75t_SL U61288 ( .A1(n58431), .A2(n59641), .B(n67342), .Y(
        n67517) );
  AND2x2_ASAP7_75t_SL U61289 ( .A(n64365), .B(n64364), .Y(n57442) );
  NOR2x1_ASAP7_75t_SL U61290 ( .A(n59666), .B(n67231), .Y(n67234) );
  INVx1_ASAP7_75t_SL U61291 ( .A(n62716), .Y(n62698) );
  INVx1_ASAP7_75t_SL U61292 ( .A(n67929), .Y(n58228) );
  NAND2xp5_ASAP7_75t_SL U61293 ( .A(n75098), .B(n75097), .Y(n57444) );
  INVx2_ASAP7_75t_SL U61294 ( .A(n57502), .Y(n67855) );
  BUFx2_ASAP7_75t_SL U61295 ( .A(n57644), .Y(n58882) );
  BUFx6f_ASAP7_75t_SL U61296 ( .A(n59453), .Y(n58903) );
  XNOR2xp5_ASAP7_75t_SL U61297 ( .A(n67085), .B(n57445), .Y(n67046) );
  XNOR2xp5_ASAP7_75t_SL U61298 ( .A(n67083), .B(n67079), .Y(n57445) );
  INVx1_ASAP7_75t_SL U61299 ( .A(n68216), .Y(n68218) );
  XNOR2x2_ASAP7_75t_SL U61300 ( .A(n68218), .B(n68217), .Y(n68219) );
  NAND2x1p5_ASAP7_75t_SL U61301 ( .A(n58078), .B(n58075), .Y(n59266) );
  NOR2x1p5_ASAP7_75t_SL U61302 ( .A(n68346), .B(n68758), .Y(n57870) );
  INVx1_ASAP7_75t_SL U61303 ( .A(n58641), .Y(n58640) );
  NAND2xp5_ASAP7_75t_SL U61304 ( .A(n59154), .B(n64719), .Y(n59153) );
  NOR2x1_ASAP7_75t_SL U61305 ( .A(n58848), .B(n67223), .Y(n67270) );
  HB1xp67_ASAP7_75t_SL U61306 ( .A(n58828), .Y(n57446) );
  NAND2xp5_ASAP7_75t_SL U61307 ( .A(n57447), .B(n58841), .Y(n78172) );
  NAND2xp5_ASAP7_75t_SL U61308 ( .A(n57606), .B(n58773), .Y(n57447) );
  XOR2xp5_ASAP7_75t_SL U61309 ( .A(n57031), .B(n57492), .Y(n66497) );
  XNOR2xp5_ASAP7_75t_SL U61310 ( .A(n58019), .B(n68339), .Y(n57951) );
  AOI22x1_ASAP7_75t_SL U61311 ( .A1(n64384), .A2(n57632), .B1(n64393), .B2(
        n57478), .Y(n64414) );
  INVx1_ASAP7_75t_SL U61312 ( .A(n64527), .Y(n64405) );
  AND2x2_ASAP7_75t_SL U61313 ( .A(n64876), .B(n64877), .Y(n64883) );
  NAND2x1_ASAP7_75t_SL U61314 ( .A(n59591), .B(n57122), .Y(n59197) );
  NOR2x1_ASAP7_75t_SL U61315 ( .A(n59596), .B(n53520), .Y(n67583) );
  NAND2x1_ASAP7_75t_SL U61316 ( .A(n67629), .B(n75761), .Y(n58803) );
  AND2x4_ASAP7_75t_SL U61317 ( .A(n58803), .B(n57166), .Y(n57563) );
  NOR2xp33_ASAP7_75t_SL U61318 ( .A(n65019), .B(n67868), .Y(n65023) );
  OAI22xp5_ASAP7_75t_SL U61319 ( .A1(n67963), .A2(n67971), .B1(n58861), .B2(
        n58536), .Y(n67335) );
  INVx4_ASAP7_75t_SL U61320 ( .A(n57551), .Y(n75927) );
  OAI21xp5_ASAP7_75t_SL U61321 ( .A1(n57486), .A2(n59582), .B(n57969), .Y(
        n67427) );
  OAI21x1_ASAP7_75t_SL U61322 ( .A1(n57858), .A2(n68026), .B(n57857), .Y(
        n68235) );
  OAI21xp5_ASAP7_75t_SL U61323 ( .A1(n67790), .A2(n58370), .B(n67791), .Y(
        n59092) );
  XOR2xp5_ASAP7_75t_SL U61324 ( .A(n57449), .B(n67392), .Y(n67791) );
  INVx1_ASAP7_75t_SL U61325 ( .A(n67400), .Y(n57449) );
  NAND2xp5_ASAP7_75t_SL U61326 ( .A(n57451), .B(n57450), .Y(n58361) );
  OAI21xp5_ASAP7_75t_SL U61327 ( .A1(n62714), .A2(n58878), .B(n62715), .Y(
        n57450) );
  NAND2xp5_ASAP7_75t_SL U61328 ( .A(n62714), .B(n58878), .Y(n57451) );
  OAI22xp5_ASAP7_75t_SL U61329 ( .A1(n62693), .A2(n64489), .B1(n67974), .B2(
        n62694), .Y(n62714) );
  XOR2xp5_ASAP7_75t_SL U61330 ( .A(n57452), .B(n58704), .Y(n67660) );
  XNOR2xp5_ASAP7_75t_SL U61331 ( .A(n67500), .B(n58930), .Y(n57452) );
  NAND2xp5_ASAP7_75t_SL U61332 ( .A(n67850), .B(n59604), .Y(n62689) );
  NAND2xp5_ASAP7_75t_SL U61333 ( .A(n57455), .B(n57454), .Y(n57453) );
  NAND2xp5_ASAP7_75t_SL U61334 ( .A(n59596), .B(n59510), .Y(n57455) );
  NAND4xp75_ASAP7_75t_SL U61335 ( .A(n59559), .B(n59545), .C(n59568), .D(
        n59565), .Y(n57961) );
  NOR2x1p5_ASAP7_75t_SL U61336 ( .A(n57961), .B(n58242), .Y(n58248) );
  INVx2_ASAP7_75t_SL U61337 ( .A(n59450), .Y(n58843) );
  INVx2_ASAP7_75t_SL U61338 ( .A(n63174), .Y(n58342) );
  BUFx3_ASAP7_75t_SL U61339 ( .A(n58208), .Y(n58207) );
  AND2x4_ASAP7_75t_SL U61340 ( .A(n62683), .B(n62684), .Y(n59483) );
  BUFx2_ASAP7_75t_SL U61341 ( .A(n1871), .Y(n59549) );
  INVx1_ASAP7_75t_SL U61342 ( .A(n66471), .Y(n66456) );
  NAND2xp5_ASAP7_75t_SL U61343 ( .A(n57104), .B(n67300), .Y(n67301) );
  OR2x6_ASAP7_75t_SL U61344 ( .A(n59325), .B(n62598), .Y(n58431) );
  XNOR2xp5_ASAP7_75t_SL U61345 ( .A(n67943), .B(n58736), .Y(n68145) );
  XOR2xp5_ASAP7_75t_SL U61346 ( .A(n68116), .B(n59036), .Y(n57862) );
  INVx1_ASAP7_75t_SL U61347 ( .A(n67603), .Y(n57458) );
  INVx1_ASAP7_75t_SL U61348 ( .A(n67905), .Y(n67367) );
  OR2x2_ASAP7_75t_SL U61349 ( .A(n64721), .B(n64709), .Y(n59365) );
  OAI21x1_ASAP7_75t_SL U61350 ( .A1(n67723), .A2(n68425), .B(n67722), .Y(
        n67727) );
  XNOR2xp5_ASAP7_75t_SL U61351 ( .A(n63199), .B(n57459), .Y(n63165) );
  XNOR2xp5_ASAP7_75t_SL U61352 ( .A(n63159), .B(n63201), .Y(n57459) );
  INVx1_ASAP7_75t_SL U61353 ( .A(n64186), .Y(n64197) );
  INVx1_ASAP7_75t_SL U61354 ( .A(n67771), .Y(n57460) );
  INVx1_ASAP7_75t_SL U61355 ( .A(n68035), .Y(n57461) );
  XNOR2xp5_ASAP7_75t_SL U61356 ( .A(n57473), .B(n57464), .Y(n63046) );
  XOR2xp5_ASAP7_75t_SL U61357 ( .A(n63043), .B(n63044), .Y(n57464) );
  INVx1_ASAP7_75t_SL U61358 ( .A(n66692), .Y(n66694) );
  NAND2x1_ASAP7_75t_SL U61359 ( .A(n57558), .B(n57559), .Y(n68032) );
  OR2x2_ASAP7_75t_SL U61360 ( .A(n64471), .B(n64470), .Y(n57467) );
  NOR2x1_ASAP7_75t_SL U61361 ( .A(n59514), .B(n59518), .Y(n67640) );
  OAI21x1_ASAP7_75t_SL U61362 ( .A1(n59639), .A2(n67638), .B(n58893), .Y(
        n67419) );
  NOR2x1_ASAP7_75t_SL U61363 ( .A(n56853), .B(n62691), .Y(n62711) );
  OAI21xp5_ASAP7_75t_SL U61364 ( .A1(n57465), .A2(n62738), .B(n62737), .Y(
        n62740) );
  NOR2x1p5_ASAP7_75t_SL U61365 ( .A(n62740), .B(n62739), .Y(n67839) );
  NAND2xp5_ASAP7_75t_SL U61366 ( .A(n59637), .B(n75904), .Y(n66631) );
  NAND2x1p5_ASAP7_75t_SL U61367 ( .A(n58213), .B(n56831), .Y(n58927) );
  XNOR2xp5_ASAP7_75t_SL U61368 ( .A(n59223), .B(n67891), .Y(n67892) );
  INVx1_ASAP7_75t_SL U61369 ( .A(n62797), .Y(n62856) );
  NOR2x1_ASAP7_75t_SL U61370 ( .A(n67626), .B(n67945), .Y(n57469) );
  INVx2_ASAP7_75t_SL U61371 ( .A(n53627), .Y(n68086) );
  MAJIxp5_ASAP7_75t_SL U61372 ( .A(n57470), .B(n67792), .C(n67793), .Y(n68572)
         );
  XOR2xp5_ASAP7_75t_SL U61373 ( .A(n59176), .B(n68056), .Y(n57470) );
  NAND2xp5_ASAP7_75t_SL U61374 ( .A(n59304), .B(n64929), .Y(n59431) );
  XNOR2xp5_ASAP7_75t_SL U61375 ( .A(n68266), .B(n68267), .Y(n57471) );
  INVx1_ASAP7_75t_SL U61376 ( .A(n68265), .Y(n57472) );
  NOR2x1_ASAP7_75t_SL U61377 ( .A(n67874), .B(n67875), .Y(n68265) );
  INVx1_ASAP7_75t_SL U61378 ( .A(n67561), .Y(n67262) );
  AND2x2_ASAP7_75t_SL U61379 ( .A(n62567), .B(n62565), .Y(n58264) );
  OAI21x1_ASAP7_75t_SL U61380 ( .A1(n58122), .A2(n63127), .B(n63126), .Y(
        n66798) );
  XNOR2x2_ASAP7_75t_SL U61381 ( .A(n64416), .B(n57760), .Y(n64682) );
  XNOR2x1_ASAP7_75t_SL U61382 ( .A(n64660), .B(n64659), .Y(n64661) );
  XNOR2x1_ASAP7_75t_SL U61383 ( .A(n64378), .B(n64377), .Y(n64659) );
  OAI22xp5_ASAP7_75t_SL U61384 ( .A1(n63823), .A2(n59460), .B1(n64022), .B2(
        n59515), .Y(n64049) );
  XNOR2xp5_ASAP7_75t_SL U61385 ( .A(n57476), .B(n75927), .Y(n57818) );
  INVx1_ASAP7_75t_SL U61386 ( .A(n59640), .Y(n57476) );
  NAND2xp5_ASAP7_75t_SL U61387 ( .A(n64035), .B(n67901), .Y(n58697) );
  OAI21x1_ASAP7_75t_SL U61388 ( .A1(n58698), .A2(n58506), .B(n58697), .Y(
        n64346) );
  INVx1_ASAP7_75t_SL U61389 ( .A(n63650), .Y(n63239) );
  INVx2_ASAP7_75t_SL U61390 ( .A(n66258), .Y(n59465) );
  NAND2x1_ASAP7_75t_SL U61391 ( .A(n53502), .B(n57627), .Y(n57626) );
  NAND2xp5_ASAP7_75t_SL U61392 ( .A(n57177), .B(n75761), .Y(n67302) );
  XNOR2xp5_ASAP7_75t_SL U61393 ( .A(n63871), .B(n63872), .Y(n58824) );
  MAJIxp5_ASAP7_75t_SL U61394 ( .A(n63625), .B(n63626), .C(n63624), .Y(n63871)
         );
  NOR2xp33_ASAP7_75t_SL U61395 ( .A(n63182), .B(n63190), .Y(n63234) );
  NAND2xp5_ASAP7_75t_SL U61396 ( .A(n59657), .B(n63826), .Y(n63190) );
  AND3x1_ASAP7_75t_SL U61397 ( .A(n59400), .B(n59563), .C(n74788), .Y(n64515)
         );
  XNOR2x1_ASAP7_75t_SL U61398 ( .A(n64444), .B(n58779), .Y(n64671) );
  NOR2xp33_ASAP7_75t_SL U61399 ( .A(n63144), .B(n63143), .Y(n63145) );
  INVx1_ASAP7_75t_SL U61400 ( .A(n64953), .Y(n63144) );
  OAI21xp5_ASAP7_75t_SL U61401 ( .A1(n68098), .A2(n67598), .B(n67902), .Y(
        n64953) );
  INVx1_ASAP7_75t_SL U61402 ( .A(n64885), .Y(n64637) );
  OAI22xp5_ASAP7_75t_SL U61403 ( .A1(n68124), .A2(n67558), .B1(n59117), .B2(
        n59283), .Y(n59164) );
  NAND2x1_ASAP7_75t_SL U61404 ( .A(n58319), .B(n67733), .Y(n68370) );
  OR3x1_ASAP7_75t_SL U61405 ( .A(n59399), .B(n75032), .C(n67640), .Y(n58629)
         );
  INVx1_ASAP7_75t_SL U61406 ( .A(n62904), .Y(n62902) );
  NOR2x1_ASAP7_75t_SL U61407 ( .A(n64518), .B(n64570), .Y(n64890) );
  INVx1_ASAP7_75t_SL U61408 ( .A(n67747), .Y(n67281) );
  O2A1O1Ixp5_ASAP7_75t_SL U61409 ( .A1(n67569), .A2(n67481), .B(n64939), .C(
        n67480), .Y(n59049) );
  NAND2xp5_ASAP7_75t_SL U61410 ( .A(n67569), .B(n59466), .Y(n64939) );
  AND2x4_ASAP7_75t_SL U61411 ( .A(n59401), .B(n64036), .Y(n58639) );
  XOR2xp5_ASAP7_75t_SL U61412 ( .A(n63625), .B(n57479), .Y(n63227) );
  BUFx2_ASAP7_75t_SL U61413 ( .A(n64353), .Y(n57480) );
  NOR2x1_ASAP7_75t_SL U61414 ( .A(n59579), .B(n59591), .Y(n66266) );
  OAI21xp5_ASAP7_75t_SL U61415 ( .A1(n58227), .A2(n59218), .B(n67981), .Y(
        n67987) );
  NAND2xp5_ASAP7_75t_SL U61416 ( .A(n67137), .B(n67136), .Y(n67195) );
  NAND2x1_ASAP7_75t_SL U61417 ( .A(n57186), .B(n59395), .Y(n59396) );
  INVx1_ASAP7_75t_SL U61418 ( .A(n64481), .Y(n59209) );
  INVx1_ASAP7_75t_SL U61419 ( .A(n68176), .Y(n68179) );
  XNOR2x1_ASAP7_75t_SL U61420 ( .A(n67762), .B(n67763), .Y(n68573) );
  NAND2x1p5_ASAP7_75t_SL U61421 ( .A(n57718), .B(n57937), .Y(n67870) );
  XOR2xp5_ASAP7_75t_SL U61422 ( .A(n68067), .B(n57487), .Y(n68249) );
  XNOR2x1_ASAP7_75t_SL U61423 ( .A(n68344), .B(n57488), .Y(n57950) );
  MAJIxp5_ASAP7_75t_SL U61424 ( .A(n68276), .B(n68277), .C(n68278), .Y(n68343)
         );
  XNOR2xp5_ASAP7_75t_SL U61425 ( .A(n67888), .B(n67890), .Y(n57580) );
  INVx1_ASAP7_75t_SL U61426 ( .A(n67617), .Y(n57490) );
  NOR2x1_ASAP7_75t_SL U61427 ( .A(n66498), .B(n66500), .Y(n57492) );
  NOR2x1_ASAP7_75t_SL U61428 ( .A(n67872), .B(n67871), .Y(n67875) );
  AND2x4_ASAP7_75t_SL U61429 ( .A(n59573), .B(n66301), .Y(n59349) );
  INVx2_ASAP7_75t_SL U61430 ( .A(n59592), .Y(n59045) );
  OAI211xp5_ASAP7_75t_SL U61431 ( .A1(n66800), .A2(n66801), .B(n59475), .C(
        n57359), .Y(n57495) );
  XNOR2x1_ASAP7_75t_SL U61432 ( .A(n57498), .B(n64727), .Y(n57732) );
  INVx1_ASAP7_75t_SL U61433 ( .A(n57497), .Y(n57496) );
  XOR2xp5_ASAP7_75t_SL U61434 ( .A(n64701), .B(n64704), .Y(n57498) );
  NOR2x1p5_ASAP7_75t_SL U61435 ( .A(n57591), .B(n60607), .Y(n63176) );
  INVx1_ASAP7_75t_SL U61436 ( .A(n59567), .Y(n78005) );
  INVx1_ASAP7_75t_SL U61437 ( .A(n63014), .Y(n63015) );
  AND2x2_ASAP7_75t_SL U61438 ( .A(n61930), .B(n61911), .Y(n59371) );
  NOR2x1_ASAP7_75t_SL U61439 ( .A(n57027), .B(n57499), .Y(n64417) );
  OAI21x1_ASAP7_75t_SL U61440 ( .A1(n58793), .A2(n59073), .B(n57042), .Y(
        n67297) );
  AND3x1_ASAP7_75t_SL U61441 ( .A(n66291), .B(n58844), .C(n59485), .Y(n57502)
         );
  XNOR2xp5_ASAP7_75t_SL U61442 ( .A(n67014), .B(n57503), .Y(n66992) );
  XNOR2xp5_ASAP7_75t_SL U61443 ( .A(n67012), .B(n67011), .Y(n57503) );
  NAND2xp5_ASAP7_75t_SL U61444 ( .A(n57117), .B(n62640), .Y(n62641) );
  NAND2xp5_ASAP7_75t_SL U61445 ( .A(n67878), .B(n67879), .Y(n58631) );
  INVx1_ASAP7_75t_SL U61446 ( .A(n66301), .Y(n66300) );
  INVx1_ASAP7_75t_SL U61447 ( .A(n64944), .Y(n64631) );
  AOI22xp5_ASAP7_75t_SL U61448 ( .A1(n75456), .A2(n64353), .B1(n59590), .B2(
        n58655), .Y(n58238) );
  NOR2x1_ASAP7_75t_SL U61449 ( .A(n59466), .B(n59658), .Y(n67223) );
  NOR2x1_ASAP7_75t_SL U61450 ( .A(n68208), .B(n68210), .Y(n68199) );
  INVx1_ASAP7_75t_SL U61451 ( .A(n64539), .Y(n64402) );
  NAND2xp5_ASAP7_75t_SL U61452 ( .A(n67210), .B(n69100), .Y(n59309) );
  INVx1_ASAP7_75t_SL U61453 ( .A(n58776), .Y(n57604) );
  NOR2x1_ASAP7_75t_SL U61454 ( .A(n58762), .B(n66463), .Y(n67140) );
  NAND2xp5_ASAP7_75t_SL U61455 ( .A(n64914), .B(n67833), .Y(n64915) );
  XNOR2x1_ASAP7_75t_SL U61456 ( .A(n68058), .B(n68059), .Y(n58344) );
  INVx1_ASAP7_75t_SL U61457 ( .A(n75900), .Y(n59340) );
  OAI21x1_ASAP7_75t_SL U61458 ( .A1(n67970), .A2(n59440), .B(n67969), .Y(
        n68217) );
  INVx1_ASAP7_75t_SL U61459 ( .A(n64504), .Y(n59471) );
  INVx2_ASAP7_75t_SL U61460 ( .A(n68743), .Y(n58729) );
  NOR2x1p5_ASAP7_75t_SL U61461 ( .A(n67242), .B(n57507), .Y(n59491) );
  INVx2_ASAP7_75t_SL U61462 ( .A(n59268), .Y(n57507) );
  NAND2x1_ASAP7_75t_SL U61463 ( .A(n59113), .B(n59601), .Y(n59268) );
  NAND2xp5_ASAP7_75t_SL U61464 ( .A(n63482), .B(n63481), .Y(n63048) );
  BUFx6f_ASAP7_75t_SL U61465 ( .A(n2001), .Y(n59560) );
  XNOR2xp5_ASAP7_75t_SL U61466 ( .A(n57943), .B(n57853), .Y(n67789) );
  OAI22x1_ASAP7_75t_SL U61467 ( .A1(n59116), .A2(n67003), .B1(n68119), .B2(
        n67002), .Y(n67054) );
  INVx1_ASAP7_75t_SL U61468 ( .A(n58970), .Y(n58966) );
  INVx1_ASAP7_75t_SL U61469 ( .A(n66717), .Y(n66713) );
  AOI21x1_ASAP7_75t_SL U61470 ( .A1(n57157), .A2(n66934), .B(n66713), .Y(
        n68455) );
  INVx2_ASAP7_75t_SL U61471 ( .A(n67151), .Y(n58004) );
  A2O1A1Ixp33_ASAP7_75t_SL U61472 ( .A1(n68414), .A2(n66758), .B(n57509), .C(
        n59599), .Y(n66759) );
  NOR2x1_ASAP7_75t_SL U61473 ( .A(n68104), .B(n57253), .Y(n57509) );
  NOR2xp33_ASAP7_75t_SL U61474 ( .A(n67962), .B(n59517), .Y(n57510) );
  NAND2x2_ASAP7_75t_SL U61475 ( .A(n59538), .B(n59540), .Y(n60599) );
  INVx2_ASAP7_75t_SL U61476 ( .A(n60599), .Y(n60600) );
  OR2x6_ASAP7_75t_SL U61477 ( .A(n59592), .B(n62880), .Y(n67343) );
  AOI22x1_ASAP7_75t_SL U61478 ( .A1(n59100), .A2(n67419), .B1(n67298), .B2(
        n67229), .Y(n67345) );
  NOR2x1_ASAP7_75t_SL U61479 ( .A(n61913), .B(n59254), .Y(n58649) );
  NOR2x1_ASAP7_75t_SL U61480 ( .A(n59284), .B(n68156), .Y(n58653) );
  NOR2x2_ASAP7_75t_SL U61481 ( .A(n58656), .B(n75644), .Y(n67303) );
  NAND2xp5_ASAP7_75t_SL U61482 ( .A(n57182), .B(n75906), .Y(n64938) );
  NAND2xp5_ASAP7_75t_SL U61483 ( .A(n67850), .B(n59639), .Y(n58893) );
  NAND2x1_ASAP7_75t_SL U61484 ( .A(n59537), .B(n66258), .Y(n57799) );
  INVx1_ASAP7_75t_SL U61485 ( .A(n62737), .Y(n62667) );
  INVx2_ASAP7_75t_SL U61486 ( .A(n67870), .Y(n68267) );
  INVx1_ASAP7_75t_SL U61487 ( .A(n66333), .Y(n58648) );
  INVx1_ASAP7_75t_SL U61488 ( .A(n59197), .Y(n62598) );
  NAND2xp5_ASAP7_75t_SL U61489 ( .A(n58481), .B(n64039), .Y(n64041) );
  INVx1_ASAP7_75t_SL U61490 ( .A(n68070), .Y(n59244) );
  A2O1A1Ixp33_ASAP7_75t_SL U61491 ( .A1(n57180), .A2(n57167), .B(n62702), .C(
        n57511), .Y(n62718) );
  NAND2xp5_ASAP7_75t_SL U61492 ( .A(n59510), .B(n67428), .Y(n57511) );
  NOR2x2_ASAP7_75t_SL U61493 ( .A(n63634), .B(n65034), .Y(n67962) );
  NOR2x1_ASAP7_75t_SL U61494 ( .A(n66451), .B(n59654), .Y(n58853) );
  NAND2xp5_ASAP7_75t_SL U61495 ( .A(n58980), .B(n58979), .Y(n58977) );
  INVx1_ASAP7_75t_SL U61496 ( .A(n66772), .Y(n66686) );
  XNOR2xp5_ASAP7_75t_SL U61497 ( .A(n57514), .B(n57513), .Y(n57512) );
  XOR2xp5_ASAP7_75t_SL U61498 ( .A(n68335), .B(n59461), .Y(n57513) );
  INVx1_ASAP7_75t_SL U61499 ( .A(n68334), .Y(n57514) );
  NAND2xp5_ASAP7_75t_SL U61500 ( .A(n58383), .B(n67920), .Y(n58758) );
  INVx1_ASAP7_75t_SL U61501 ( .A(n58803), .Y(n67267) );
  OAI22xp5_ASAP7_75t_SL U61502 ( .A1(n57515), .A2(n57158), .B1(n57410), .B2(
        n67718), .Y(n67405) );
  INVx1_ASAP7_75t_SL U61503 ( .A(n67314), .Y(n57515) );
  XOR2xp5_ASAP7_75t_SL U61504 ( .A(n58874), .B(n57517), .Y(n63041) );
  XOR2xp5_ASAP7_75t_SL U61505 ( .A(n63030), .B(n63032), .Y(n57517) );
  OAI21xp5_ASAP7_75t_SL U61506 ( .A1(n62833), .A2(n57518), .B(n62626), .Y(
        n63030) );
  NAND2x1p5_ASAP7_75t_SL U61507 ( .A(n74776), .B(n57117), .Y(n64622) );
  OAI21x1_ASAP7_75t_SL U61508 ( .A1(n67852), .A2(n59116), .B(n57011), .Y(
        n68107) );
  XNOR2xp5_ASAP7_75t_SL U61509 ( .A(n58702), .B(n68307), .Y(n59362) );
  NOR2x1_ASAP7_75t_SL U61510 ( .A(n64874), .B(n64879), .Y(n64882) );
  NAND3x1_ASAP7_75t_SL U61511 ( .A(n75761), .B(n75762), .C(n59611), .Y(n62647)
         );
  NAND2x1_ASAP7_75t_SL U61512 ( .A(n59535), .B(n59339), .Y(n58014) );
  XNOR2xp5_ASAP7_75t_SL U61513 ( .A(n67055), .B(n58795), .Y(n67050) );
  XNOR2xp5_ASAP7_75t_SL U61514 ( .A(n75922), .B(n59607), .Y(n65019) );
  O2A1O1Ixp5_ASAP7_75t_SL U61515 ( .A1(n56827), .A2(n68104), .B(n68103), .C(
        n68102), .Y(n68106) );
  INVx1_ASAP7_75t_SL U61516 ( .A(n65052), .Y(n64467) );
  NOR2x1_ASAP7_75t_SL U61517 ( .A(n68582), .B(n69004), .Y(n68583) );
  OAI21x1_ASAP7_75t_SL U61518 ( .A1(n68914), .A2(n68584), .B(n68583), .Y(
        n68663) );
  XNOR2x1_ASAP7_75t_SL U61519 ( .A(n68161), .B(n57892), .Y(n57891) );
  BUFx6f_ASAP7_75t_SL U61520 ( .A(n2021), .Y(n59565) );
  NOR2x1p5_ASAP7_75t_SL U61521 ( .A(n68956), .B(n58088), .Y(n68717) );
  NAND2x1p5_ASAP7_75t_SL U61522 ( .A(n68717), .B(n68906), .Y(n68562) );
  INVx1_ASAP7_75t_SL U61523 ( .A(n58738), .Y(n58737) );
  INVx1_ASAP7_75t_SL U61524 ( .A(n68354), .Y(n58781) );
  INVx1_ASAP7_75t_SL U61525 ( .A(n66649), .Y(n66628) );
  XNOR2xp5_ASAP7_75t_SL U61526 ( .A(n75922), .B(n59639), .Y(n67247) );
  NAND3x1_ASAP7_75t_SL U61527 ( .A(n59568), .B(n59565), .C(n59545), .Y(n59186)
         );
  AND2x4_ASAP7_75t_SL U61528 ( .A(n66258), .B(n64895), .Y(n64621) );
  OAI21x1_ASAP7_75t_SL U61529 ( .A1(n57434), .A2(n64621), .B(n59529), .Y(
        n65021) );
  NOR2x1p5_ASAP7_75t_SL U61530 ( .A(n67861), .B(n66625), .Y(n59102) );
  NAND2x1p5_ASAP7_75t_SL U61531 ( .A(n62557), .B(n62558), .Y(n66450) );
  NAND2xp5_ASAP7_75t_SL U61532 ( .A(n58015), .B(n67864), .Y(n67865) );
  XNOR2x1_ASAP7_75t_SL U61533 ( .A(n59028), .B(n68385), .Y(n68420) );
  NOR2x1_ASAP7_75t_SL U61534 ( .A(n62804), .B(n62805), .Y(n64965) );
  NOR2x1_ASAP7_75t_SL U61535 ( .A(n59534), .B(n57186), .Y(n63656) );
  NAND2xp5_ASAP7_75t_SL U61536 ( .A(n67428), .B(n57104), .Y(n64918) );
  NAND2xp5_ASAP7_75t_SL U61537 ( .A(n59711), .B(n59558), .Y(n61910) );
  OAI21x1_ASAP7_75t_SL U61538 ( .A1(n57949), .A2(n57165), .B(n57948), .Y(
        n64891) );
  AND2x4_ASAP7_75t_SL U61539 ( .A(n57783), .B(n57782), .Y(n57781) );
  OAI22x1_ASAP7_75t_SL U61540 ( .A1(n59440), .A2(n57603), .B1(n58398), .B2(
        n59446), .Y(n59223) );
  INVx1_ASAP7_75t_SL U61541 ( .A(n67439), .Y(n67456) );
  INVx1_ASAP7_75t_SL U61542 ( .A(n58969), .Y(n58968) );
  INVx1_ASAP7_75t_SL U61543 ( .A(n67708), .Y(n67710) );
  OAI21x1_ASAP7_75t_SL U61544 ( .A1(n59440), .A2(n67710), .B(n56988), .Y(
        n68388) );
  NOR2x1p5_ASAP7_75t_SL U61545 ( .A(n66332), .B(n59600), .Y(n66864) );
  NAND2x1p5_ASAP7_75t_SL U61546 ( .A(n59488), .B(n64367), .Y(n67634) );
  NOR2x1_ASAP7_75t_SL U61547 ( .A(n68119), .B(n67258), .Y(n59178) );
  AOI21x1_ASAP7_75t_SL U61548 ( .A1(n57603), .A2(n58336), .B(n59178), .Y(
        n67350) );
  INVx2_ASAP7_75t_SL U61549 ( .A(n53615), .Y(n59310) );
  NAND2x1p5_ASAP7_75t_SL U61550 ( .A(n58245), .B(n58047), .Y(n59254) );
  OAI21xp5_ASAP7_75t_SL U61551 ( .A1(n59559), .A2(n62638), .B(n62634), .Y(
        n62635) );
  INVx1_ASAP7_75t_SL U61552 ( .A(n62968), .Y(n62928) );
  OAI21xp5_ASAP7_75t_SL U61553 ( .A1(n57243), .A2(n53280), .B(n63228), .Y(
        n63229) );
  NOR2x1_ASAP7_75t_SL U61554 ( .A(n58907), .B(n63229), .Y(n63230) );
  INVx1_ASAP7_75t_SL U61555 ( .A(n62722), .Y(n58905) );
  NAND2x2_ASAP7_75t_SL U61556 ( .A(n68098), .B(n62580), .Y(n64625) );
  XOR2x2_ASAP7_75t_SL U61557 ( .A(n57050), .B(n68264), .Y(n58702) );
  INVx1_ASAP7_75t_SL U61558 ( .A(n68307), .Y(n57797) );
  NAND2xp5_ASAP7_75t_SL U61559 ( .A(n68307), .B(n57519), .Y(n57796) );
  INVx1_ASAP7_75t_SL U61560 ( .A(n58702), .Y(n57519) );
  INVx1_ASAP7_75t_SL U61561 ( .A(n68128), .Y(n57520) );
  INVx1_ASAP7_75t_SL U61562 ( .A(n68127), .Y(n57521) );
  MAJIxp5_ASAP7_75t_SL U61563 ( .A(n68270), .B(n68269), .C(n68268), .Y(n68307)
         );
  XNOR2xp5_ASAP7_75t_SL U61564 ( .A(n68165), .B(n65055), .Y(n68268) );
  XNOR2x1_ASAP7_75t_SL U61565 ( .A(n57929), .B(n57522), .Y(n57723) );
  MAJIxp5_ASAP7_75t_SL U61566 ( .A(n53495), .B(n67529), .C(n67528), .Y(n67697)
         );
  XNOR2x1_ASAP7_75t_SL U61567 ( .A(n57984), .B(n57767), .Y(n57522) );
  XNOR2x1_ASAP7_75t_SL U61568 ( .A(n57523), .B(n57524), .Y(n67786) );
  INVx1_ASAP7_75t_SL U61569 ( .A(n67510), .Y(n57524) );
  MAJIxp5_ASAP7_75t_SL U61570 ( .A(n67297), .B(n67296), .C(n67295), .Y(n67510)
         );
  BUFx6f_ASAP7_75t_SL U61571 ( .A(n59352), .Y(n57525) );
  NOR2x1_ASAP7_75t_SL U61572 ( .A(n59647), .B(n57179), .Y(n66862) );
  XOR2xp5_ASAP7_75t_SL U61573 ( .A(n57525), .B(n67964), .Y(n67744) );
  XOR2xp5_ASAP7_75t_SL U61574 ( .A(n59620), .B(n57525), .Y(n67440) );
  NOR2x1_ASAP7_75t_SL U61575 ( .A(n57314), .B(n57394), .Y(n66674) );
  NOR2x1_ASAP7_75t_SL U61576 ( .A(n57314), .B(n66758), .Y(n66675) );
  XOR2xp5_ASAP7_75t_SL U61577 ( .A(n57314), .B(n59658), .Y(n66766) );
  NAND2xp5_ASAP7_75t_SL U61578 ( .A(n65005), .B(n65004), .Y(n68220) );
  INVx1_ASAP7_75t_SL U61579 ( .A(n57527), .Y(n57526) );
  AOI21xp5_ASAP7_75t_SL U61580 ( .A1(n57110), .A2(n64933), .B(n58777), .Y(
        n57527) );
  NAND2xp5_ASAP7_75t_SL U61581 ( .A(n57018), .B(n57963), .Y(n57528) );
  XNOR2x1_ASAP7_75t_SL U61582 ( .A(n68532), .B(n68487), .Y(n57529) );
  XOR2xp5_ASAP7_75t_SL U61583 ( .A(n57530), .B(n68521), .Y(n68494) );
  INVx1_ASAP7_75t_SL U61584 ( .A(n68522), .Y(n57530) );
  OAI21xp5_ASAP7_75t_SL U61585 ( .A1(n59531), .A2(n57531), .B(n66244), .Y(
        n59402) );
  XNOR2xp5_ASAP7_75t_SL U61586 ( .A(n57532), .B(n64941), .Y(n64942) );
  XNOR2xp5_ASAP7_75t_SL U61587 ( .A(n57533), .B(n58690), .Y(n57532) );
  INVx1_ASAP7_75t_SL U61588 ( .A(n65013), .Y(n57533) );
  INVx1_ASAP7_75t_SL U61589 ( .A(n57536), .Y(n65066) );
  XNOR2xp5_ASAP7_75t_SL U61590 ( .A(n65058), .B(n57534), .Y(n57536) );
  XNOR2xp5_ASAP7_75t_SL U61591 ( .A(n57535), .B(n65056), .Y(n57534) );
  INVx1_ASAP7_75t_SL U61592 ( .A(n65057), .Y(n57535) );
  MAJx2_ASAP7_75t_SL U61593 ( .A(n57536), .B(n56843), .C(n64942), .Y(n68256)
         );
  NAND2xp5_ASAP7_75t_SL U61594 ( .A(n57005), .B(n64918), .Y(n65057) );
  NOR2x1p5_ASAP7_75t_SL U61595 ( .A(n57019), .B(n58973), .Y(n57537) );
  AOI21x1_ASAP7_75t_SL U61596 ( .A1(n57462), .A2(n76627), .B(n57443), .Y(
        n57538) );
  INVx2_ASAP7_75t_SL U61597 ( .A(n75109), .Y(n57539) );
  AOI31xp67_ASAP7_75t_SL U61598 ( .A1(n57539), .A2(n59427), .A3(n75137), .B(
        n75136), .Y(n58380) );
  NOR2x1_ASAP7_75t_SL U61599 ( .A(n68397), .B(n59090), .Y(n59023) );
  INVx1_ASAP7_75t_SL U61600 ( .A(n68395), .Y(n59090) );
  XNOR2xp5_ASAP7_75t_SL U61601 ( .A(n57540), .B(n68356), .Y(n68395) );
  MAJIxp5_ASAP7_75t_SL U61602 ( .A(n67681), .B(n67682), .C(n67683), .Y(n68356)
         );
  XOR2xp5_ASAP7_75t_SL U61603 ( .A(n56832), .B(n68357), .Y(n57540) );
  MAJIxp5_ASAP7_75t_SL U61604 ( .A(n67692), .B(n67690), .C(n67691), .Y(n68404)
         );
  XOR2xp5_ASAP7_75t_SL U61605 ( .A(n64891), .B(n57064), .Y(n64652) );
  A2O1A1Ixp33_ASAP7_75t_SL U61606 ( .A1(n57180), .A2(n59651), .B(n64650), .C(
        n57542), .Y(n64892) );
  INVx1_ASAP7_75t_SL U61607 ( .A(n67620), .Y(n57543) );
  MAJIxp5_ASAP7_75t_SL U61608 ( .A(n68308), .B(n68309), .C(n68310), .Y(n57544)
         );
  NOR2x1_ASAP7_75t_SL U61609 ( .A(n53483), .B(n57544), .Y(n59216) );
  NAND2xp5_ASAP7_75t_SL U61610 ( .A(n57544), .B(n53483), .Y(n59215) );
  XNOR2xp5_ASAP7_75t_SL U61611 ( .A(n68317), .B(n57544), .Y(n68318) );
  NOR2x1_ASAP7_75t_SL U61612 ( .A(n68263), .B(n68262), .Y(n68306) );
  MAJIxp5_ASAP7_75t_SL U61613 ( .A(n64889), .B(n64887), .C(n64888), .Y(n65028)
         );
  XNOR2x1_ASAP7_75t_SL U61614 ( .A(n59161), .B(n59160), .Y(n67699) );
  XNOR2xp5_ASAP7_75t_SL U61615 ( .A(n57153), .B(n67006), .Y(n66854) );
  INVx1_ASAP7_75t_SL U61616 ( .A(n59447), .Y(n57547) );
  AND2x2_ASAP7_75t_SL U61617 ( .A(n59614), .B(n75927), .Y(n62622) );
  NAND2xp5_ASAP7_75t_SL U61618 ( .A(n57551), .B(n58232), .Y(n57548) );
  NAND2xp5_ASAP7_75t_SL U61619 ( .A(n57912), .B(n57551), .Y(n65040) );
  NAND2xp5_ASAP7_75t_SL U61620 ( .A(n57356), .B(n57178), .Y(n62814) );
  NAND2xp5_ASAP7_75t_SL U61621 ( .A(n57549), .B(n62783), .Y(n62788) );
  OAI21xp5_ASAP7_75t_SL U61622 ( .A1(n57356), .A2(n59618), .B(n57550), .Y(
        n57549) );
  NAND2xp5_ASAP7_75t_SL U61623 ( .A(n57356), .B(n57180), .Y(n57550) );
  INVx1_ASAP7_75t_SL U61624 ( .A(n64678), .Y(n64045) );
  AND2x2_ASAP7_75t_SL U61625 ( .A(n57552), .B(n64678), .Y(n64717) );
  INVx1_ASAP7_75t_SL U61626 ( .A(n64044), .Y(n57552) );
  INVx1_ASAP7_75t_SL U61627 ( .A(n64693), .Y(n64698) );
  OR2x2_ASAP7_75t_SL U61628 ( .A(n64553), .B(n57555), .Y(n64549) );
  NAND2xp5_ASAP7_75t_SL U61629 ( .A(n64553), .B(n57555), .Y(n64548) );
  OR2x2_ASAP7_75t_SL U61630 ( .A(n57215), .B(n57556), .Y(n66254) );
  NOR2x1_ASAP7_75t_SL U61631 ( .A(n57556), .B(n66304), .Y(n66302) );
  INVx1_ASAP7_75t_SL U61632 ( .A(n57557), .Y(n58740) );
  NAND2xp5_ASAP7_75t_SL U61633 ( .A(n57140), .B(n68032), .Y(n57557) );
  NAND3xp33_ASAP7_75t_SL U61634 ( .A(n59220), .B(n59219), .C(n67987), .Y(
        n57558) );
  NAND2xp5_ASAP7_75t_SL U61635 ( .A(n59217), .B(n67990), .Y(n57559) );
  NAND3xp33_ASAP7_75t_SL U61636 ( .A(n75848), .B(n57560), .C(n77732), .Y(
        n74782) );
  AOI21xp5_ASAP7_75t_SL U61637 ( .A1(n66297), .A2(n57561), .B(n59413), .Y(
        n58725) );
  NAND2x2_ASAP7_75t_SL U61638 ( .A(n59242), .B(n59239), .Y(n67837) );
  NAND2xp5_ASAP7_75t_SL U61639 ( .A(n57107), .B(n57065), .Y(n57562) );
  XOR2xp5_ASAP7_75t_SL U61640 ( .A(n68336), .B(n59294), .Y(n59433) );
  XNOR2x1_ASAP7_75t_SL U61641 ( .A(n58687), .B(n68332), .Y(n68330) );
  MAJIxp5_ASAP7_75t_SL U61642 ( .A(n68330), .B(n57420), .C(n58918), .Y(n68336)
         );
  INVx2_ASAP7_75t_SL U61643 ( .A(n57563), .Y(n66915) );
  NOR2x1_ASAP7_75t_SL U61644 ( .A(n57565), .B(n57564), .Y(n57761) );
  NAND2xp5_ASAP7_75t_SL U61645 ( .A(n68079), .B(n66915), .Y(n57564) );
  INVx1_ASAP7_75t_SL U61646 ( .A(n64030), .Y(n57565) );
  NAND2xp5_ASAP7_75t_SL U61647 ( .A(n68087), .B(n59614), .Y(n57566) );
  AND2x2_ASAP7_75t_SL U61648 ( .A(n64971), .B(n57037), .Y(n64973) );
  OAI21xp5_ASAP7_75t_SL U61649 ( .A1(n65052), .A2(n58903), .B(n57022), .Y(
        n64971) );
  OAI21xp5_ASAP7_75t_SL U61650 ( .A1(n64643), .A2(n64642), .B(n57568), .Y(
        n64974) );
  NAND2xp5_ASAP7_75t_SL U61651 ( .A(n68086), .B(n64955), .Y(n57568) );
  XNOR2xp5_ASAP7_75t_SL U61652 ( .A(n53320), .B(n57662), .Y(n64955) );
  NOR2x1_ASAP7_75t_SL U61653 ( .A(n62959), .B(n66716), .Y(n64642) );
  INVx1_ASAP7_75t_SL U61654 ( .A(n66719), .Y(n62959) );
  A2O1A1Ixp33_ASAP7_75t_SL U61655 ( .A1(n57030), .A2(n56849), .B(n57569), .C(
        n57147), .Y(n58136) );
  NAND2xp5_ASAP7_75t_SL U61656 ( .A(n58137), .B(n67487), .Y(n58351) );
  NAND2xp5_ASAP7_75t_SL U61657 ( .A(n56849), .B(n57030), .Y(n67487) );
  INVx1_ASAP7_75t_SL U61658 ( .A(n68143), .Y(n68142) );
  INVx1_ASAP7_75t_SL U61659 ( .A(n65031), .Y(n57572) );
  NAND4xp75_ASAP7_75t_SL U61660 ( .A(n60946), .B(n60600), .C(n56828), .D(
        n57577), .Y(n65031) );
  NOR2x1p5_ASAP7_75t_SL U61661 ( .A(n57578), .B(n59053), .Y(n57577) );
  NAND2x2_ASAP7_75t_SL U61662 ( .A(n59531), .B(n1621), .Y(n64617) );
  XNOR2xp5_ASAP7_75t_SL U61663 ( .A(n58739), .B(n57579), .Y(n68061) );
  XNOR2xp5_ASAP7_75t_SL U61664 ( .A(n68033), .B(n68032), .Y(n57579) );
  INVx1_ASAP7_75t_SL U61665 ( .A(n59008), .Y(n57581) );
  OAI21xp5_ASAP7_75t_SL U61666 ( .A1(n57586), .A2(n64653), .B(n57583), .Y(
        n64878) );
  NAND2xp5_ASAP7_75t_SL U61667 ( .A(n57584), .B(n64580), .Y(n57583) );
  NAND2xp5_ASAP7_75t_SL U61668 ( .A(n64576), .B(n64577), .Y(n64580) );
  NAND2xp5_ASAP7_75t_SL U61669 ( .A(n64512), .B(n64607), .Y(n64577) );
  OAI21xp5_ASAP7_75t_SL U61670 ( .A1(n57585), .A2(n64505), .B(n66860), .Y(
        n64583) );
  OAI21xp5_ASAP7_75t_SL U61671 ( .A1(n64579), .A2(n57587), .B(n64578), .Y(
        n57586) );
  NOR2x1_ASAP7_75t_SL U61672 ( .A(n64574), .B(n64575), .Y(n64893) );
  XNOR2xp5_ASAP7_75t_SL U61673 ( .A(n59614), .B(n59511), .Y(n58509) );
  XOR2xp5_ASAP7_75t_SL U61674 ( .A(n64456), .B(n64455), .Y(n58780) );
  NAND2xp5_ASAP7_75t_SL U61675 ( .A(n59571), .B(n59542), .Y(n57589) );
  NAND2xp5_ASAP7_75t_SL U61676 ( .A(n63125), .B(n59535), .Y(n63172) );
  NOR2x1_ASAP7_75t_SL U61677 ( .A(n57590), .B(n57210), .Y(n63125) );
  INVx1_ASAP7_75t_SL U61678 ( .A(n59537), .Y(n57590) );
  NAND3x1_ASAP7_75t_SL U61679 ( .A(n57199), .B(n58168), .C(n58167), .Y(n61809)
         );
  INVx1_ASAP7_75t_SL U61680 ( .A(n61909), .Y(n57592) );
  NAND2xp5_ASAP7_75t_SL U61681 ( .A(n57595), .B(n58041), .Y(n57594) );
  NAND2xp5_ASAP7_75t_SL U61682 ( .A(n66805), .B(n75899), .Y(n57595) );
  NOR2x1p5_ASAP7_75t_SL U61683 ( .A(n63104), .B(n63103), .Y(n63497) );
  INVxp67_ASAP7_75t_SL U61684 ( .A(n57598), .Y(n57599) );
  O2A1O1Ixp33_ASAP7_75t_SL U61685 ( .A1(n58403), .A2(n58426), .B(n57601), .C(
        n59545), .Y(n57598) );
  NOR2xp67_ASAP7_75t_SL U61686 ( .A(n59482), .B(n62592), .Y(n62634) );
  NOR2x2_ASAP7_75t_SL U61687 ( .A(n58426), .B(n58403), .Y(n59482) );
  INVx1_ASAP7_75t_SL U61688 ( .A(n57817), .Y(n63836) );
  OAI21xp5_ASAP7_75t_SL U61689 ( .A1(n57600), .A2(n59482), .B(n57599), .Y(
        n57817) );
  NAND2xp5_ASAP7_75t_SL U61690 ( .A(n59545), .B(n57601), .Y(n57600) );
  INVx1_ASAP7_75t_SL U61691 ( .A(n62592), .Y(n57601) );
  INVx3_ASAP7_75t_SL U61692 ( .A(n67709), .Y(n59042) );
  NOR2x1_ASAP7_75t_SL U61693 ( .A(n63192), .B(n57347), .Y(n58044) );
  NOR2x1_ASAP7_75t_SL U61694 ( .A(n59551), .B(n63654), .Y(n63192) );
  AND2x2_ASAP7_75t_SL U61695 ( .A(n78327), .B(n66260), .Y(n63654) );
  OAI21xp5_ASAP7_75t_SL U61696 ( .A1(n58688), .A2(n68665), .B(n58677), .Y(
        n69082) );
  NAND2x1_ASAP7_75t_SL U61697 ( .A(n57605), .B(n57604), .Y(n57603) );
  NAND2xp5_ASAP7_75t_SL U61698 ( .A(n75470), .B(n58881), .Y(n58773) );
  NAND2xp5_ASAP7_75t_SL U61699 ( .A(n75463), .B(n57607), .Y(n58842) );
  NAND2xp5_ASAP7_75t_SL U61700 ( .A(n75464), .B(n75465), .Y(n57607) );
  NAND2xp5_ASAP7_75t_SL U61701 ( .A(n75113), .B(n75112), .Y(n75465) );
  A2O1A1Ixp33_ASAP7_75t_SL U61702 ( .A1(n75473), .A2(n58773), .B(n75472), .C(
        n75471), .Y(n78169) );
  XOR2xp5_ASAP7_75t_SL U61703 ( .A(n56843), .B(n65066), .Y(n57608) );
  MAJIxp5_ASAP7_75t_SL U61704 ( .A(n65000), .B(n64999), .C(n64998), .Y(n68276)
         );
  XNOR2xp5_ASAP7_75t_SL U61705 ( .A(n68276), .B(n68277), .Y(n58924) );
  XNOR2xp5_ASAP7_75t_SL U61706 ( .A(n67127), .B(n67128), .Y(n67129) );
  NOR2x1_ASAP7_75t_SL U61707 ( .A(n57609), .B(n57017), .Y(n67127) );
  AOI21xp5_ASAP7_75t_SL U61708 ( .A1(n59639), .A2(n75893), .B(n59518), .Y(
        n66921) );
  NOR2x1_ASAP7_75t_SL U61709 ( .A(n57377), .B(n59591), .Y(n57611) );
  NAND3xp33_ASAP7_75t_SL U61710 ( .A(n59400), .B(n57377), .C(n64036), .Y(
        n64038) );
  INVx2_ASAP7_75t_SL U61711 ( .A(n67977), .Y(n57613) );
  OAI22x1_ASAP7_75t_SL U61712 ( .A1(n57165), .A2(n67923), .B1(n68004), .B2(
        n57099), .Y(n67978) );
  INVx1_ASAP7_75t_SL U61713 ( .A(n57068), .Y(n77730) );
  NOR2x1_ASAP7_75t_SL U61714 ( .A(n57615), .B(n57614), .Y(n67162) );
  XNOR2xp5_ASAP7_75t_SL U61715 ( .A(n67116), .B(n67117), .Y(n57615) );
  OAI21xp5_ASAP7_75t_SL U61716 ( .A1(n57617), .A2(n57616), .B(n68372), .Y(
        n68432) );
  NAND2xp5_ASAP7_75t_SL U61717 ( .A(n68368), .B(n68370), .Y(n57616) );
  INVx1_ASAP7_75t_SL U61718 ( .A(n58783), .Y(n57617) );
  XNOR2x1_ASAP7_75t_SL U61719 ( .A(n57619), .B(n68430), .Y(n68446) );
  NAND2x1_ASAP7_75t_SL U61720 ( .A(n68432), .B(n68431), .Y(n68430) );
  NAND2x1_ASAP7_75t_SL U61721 ( .A(n57618), .B(n68369), .Y(n68431) );
  NAND2x1_ASAP7_75t_SL U61722 ( .A(n68370), .B(n58783), .Y(n68369) );
  XNOR2x1_ASAP7_75t_SL U61723 ( .A(n68434), .B(n68433), .Y(n57619) );
  XNOR2x1_ASAP7_75t_SL U61724 ( .A(n57620), .B(n68447), .Y(n68433) );
  XNOR2x1_ASAP7_75t_SL U61725 ( .A(n57621), .B(n68440), .Y(n68434) );
  XNOR2x2_ASAP7_75t_SL U61726 ( .A(n68074), .B(n57623), .Y(n57894) );
  XNOR2xp5_ASAP7_75t_SL U61727 ( .A(n68047), .B(n68073), .Y(n57623) );
  MAJIxp5_ASAP7_75t_SL U61728 ( .A(n67885), .B(n57863), .C(n68115), .Y(n68047)
         );
  XNOR2xp5_ASAP7_75t_SL U61729 ( .A(n68244), .B(n57894), .Y(n58022) );
  AOI31xp67_ASAP7_75t_SL U61730 ( .A1(n58218), .A2(n57626), .A3(n57625), .B(
        n57624), .Y(n68244) );
  NOR2x1_ASAP7_75t_SL U61731 ( .A(n53502), .B(n57627), .Y(n57624) );
  INVx1_ASAP7_75t_SL U61732 ( .A(n57774), .Y(n57625) );
  OA21x2_ASAP7_75t_SL U61733 ( .A1(n58906), .A2(n57629), .B(n62721), .Y(n57628) );
  NAND2x2_ASAP7_75t_SL U61734 ( .A(n59145), .B(n58463), .Y(n67230) );
  INVx1_ASAP7_75t_SL U61735 ( .A(n63013), .Y(n62985) );
  NAND2xp5_ASAP7_75t_SL U61736 ( .A(n62970), .B(n62971), .Y(n63013) );
  OAI21xp5_ASAP7_75t_SL U61737 ( .A1(n57633), .A2(n53203), .B(n57631), .Y(
        n62971) );
  A2O1A1Ixp33_ASAP7_75t_SL U61738 ( .A1(n58931), .A2(n59514), .B(n58932), .C(
        n57632), .Y(n57631) );
  INVx1_ASAP7_75t_SL U61739 ( .A(n57156), .Y(n57632) );
  INVx1_ASAP7_75t_SL U61740 ( .A(n59308), .Y(n57633) );
  NAND2xp5_ASAP7_75t_SL U61741 ( .A(n66387), .B(n58530), .Y(n66388) );
  AND2x2_ASAP7_75t_SL U61742 ( .A(n66860), .B(n59662), .Y(n66374) );
  OAI22x1_ASAP7_75t_SL U61743 ( .A1(n67439), .A2(n57099), .B1(n57165), .B2(
        n67440), .Y(n67619) );
  INVx1_ASAP7_75t_SL U61744 ( .A(n62563), .Y(n57635) );
  NOR2x1_ASAP7_75t_SL U61745 ( .A(n62561), .B(n2956), .Y(n62567) );
  INVx1_ASAP7_75t_SL U61746 ( .A(n62701), .Y(n57636) );
  INVx1_ASAP7_75t_SL U61747 ( .A(n67322), .Y(n59038) );
  OR2x2_ASAP7_75t_SL U61748 ( .A(n58863), .B(n64928), .Y(n67322) );
  INVx1_ASAP7_75t_SL U61749 ( .A(n61212), .Y(n57639) );
  NAND2xp5_ASAP7_75t_SL U61750 ( .A(n57641), .B(n59541), .Y(n57640) );
  INVx1_ASAP7_75t_SL U61751 ( .A(n59538), .Y(n57641) );
  NAND2xp5_ASAP7_75t_SL U61752 ( .A(n57642), .B(n67332), .Y(n67334) );
  INVx1_ASAP7_75t_SL U61753 ( .A(n67331), .Y(n57642) );
  NOR2x1_ASAP7_75t_SL U61754 ( .A(n63655), .B(n63809), .Y(n67331) );
  NAND2xp5_ASAP7_75t_SL U61755 ( .A(n58518), .B(n57643), .Y(n59218) );
  INVx1_ASAP7_75t_SL U61756 ( .A(n67928), .Y(n57643) );
  NAND2xp5_ASAP7_75t_SL U61757 ( .A(n62582), .B(n62668), .Y(n62560) );
  NOR2x1p5_ASAP7_75t_SL U61758 ( .A(n57082), .B(n57128), .Y(n61212) );
  INVx1_ASAP7_75t_SL U61759 ( .A(n59571), .Y(n77278) );
  OR2x2_ASAP7_75t_SL U61760 ( .A(n57646), .B(n57648), .Y(n60657) );
  NAND2xp5_ASAP7_75t_SL U61761 ( .A(n59565), .B(n59568), .Y(n57646) );
  NOR2x1_ASAP7_75t_SL U61762 ( .A(n57648), .B(n57647), .Y(n57649) );
  NAND4xp25_ASAP7_75t_SL U61763 ( .A(n59555), .B(n59571), .C(n59568), .D(
        n59565), .Y(n57647) );
  NOR2x1_ASAP7_75t_SL U61764 ( .A(n56837), .B(n60915), .Y(n62760) );
  INVx1_ASAP7_75t_SL U61765 ( .A(n63481), .Y(n57650) );
  XOR2xp5_ASAP7_75t_SL U61766 ( .A(n62780), .B(n63049), .Y(n63481) );
  NAND2xp5_ASAP7_75t_SL U61767 ( .A(n58383), .B(n53520), .Y(n57651) );
  NAND2xp5_ASAP7_75t_SL U61768 ( .A(n57912), .B(n57167), .Y(n57652) );
  NAND2x2_ASAP7_75t_SL U61769 ( .A(n57733), .B(n56971), .Y(n59661) );
  XNOR2x1_ASAP7_75t_SL U61770 ( .A(n58175), .B(n62636), .Y(n57653) );
  OAI21x1_ASAP7_75t_SL U61771 ( .A1(n57654), .A2(n63124), .B(n62763), .Y(
        n64957) );
  AOI21xp5_ASAP7_75t_SL U61772 ( .A1(n62760), .A2(n59538), .B(n59560), .Y(
        n57654) );
  NAND2x2_ASAP7_75t_SL U61773 ( .A(n57655), .B(n57182), .Y(n59200) );
  INVx2_ASAP7_75t_SL U61774 ( .A(n57656), .Y(n57655) );
  BUFx6f_ASAP7_75t_SL U61775 ( .A(n64957), .Y(n57656) );
  XNOR2xp5_ASAP7_75t_SL U61776 ( .A(n67068), .B(n67067), .Y(n58237) );
  INVx1_ASAP7_75t_SL U61777 ( .A(n67033), .Y(n57657) );
  OAI22xp5_ASAP7_75t_SL U61778 ( .A1(n67001), .A2(n59612), .B1(n66856), .B2(
        n67627), .Y(n67033) );
  XNOR2xp5_ASAP7_75t_SL U61779 ( .A(n57659), .B(n67158), .Y(n57658) );
  A2O1A1Ixp33_ASAP7_75t_SL U61780 ( .A1(n59551), .A2(n57116), .B(n57122), .C(
        n57661), .Y(n57663) );
  INVxp67_ASAP7_75t_SL U61781 ( .A(n67143), .Y(n57664) );
  O2A1O1Ixp33_ASAP7_75t_SL U61782 ( .A1(n57394), .A2(n67871), .B(n67094), .C(
        n67093), .Y(n67143) );
  NOR2x2_ASAP7_75t_SL U61783 ( .A(n58264), .B(n58265), .Y(n64894) );
  NOR2x1p5_ASAP7_75t_SL U61784 ( .A(n64618), .B(n63173), .Y(n62761) );
  NAND2x2_ASAP7_75t_SL U61785 ( .A(n62557), .B(n62558), .Y(n66244) );
  NAND2xp5_ASAP7_75t_SL U61786 ( .A(n67432), .B(n57941), .Y(n58920) );
  XOR2xp5_ASAP7_75t_SL U61787 ( .A(n64886), .B(n64641), .Y(n64906) );
  MAJIxp5_ASAP7_75t_SL U61788 ( .A(n64640), .B(n64639), .C(n64638), .Y(n64886)
         );
  OAI22xp5_ASAP7_75t_SL U61789 ( .A1(n64501), .A2(n66829), .B1(n57508), .B2(
        n64612), .Y(n64638) );
  OAI22xp5_ASAP7_75t_SL U61790 ( .A1(n64498), .A2(n67627), .B1(n64497), .B2(
        n58658), .Y(n64640) );
  XNOR2x1_ASAP7_75t_SL U61791 ( .A(n67986), .B(n67985), .Y(n58926) );
  XNOR2x1_ASAP7_75t_SL U61792 ( .A(n58453), .B(n57668), .Y(n67985) );
  XNOR2x2_ASAP7_75t_SL U61793 ( .A(n67812), .B(n58787), .Y(n67986) );
  OAI21x1_ASAP7_75t_SL U61794 ( .A1(n67626), .A2(n58658), .B(n57997), .Y(
        n58453) );
  NAND2xp5_ASAP7_75t_SL U61795 ( .A(n57673), .B(n68028), .Y(n68231) );
  NOR2x1_ASAP7_75t_SL U61796 ( .A(n57673), .B(n68028), .Y(n68233) );
  INVx1_ASAP7_75t_SL U61797 ( .A(n68185), .Y(n57673) );
  NAND2xp5_ASAP7_75t_SL U61798 ( .A(n57674), .B(n67591), .Y(n57681) );
  MAJx2_ASAP7_75t_SL U61799 ( .A(n67995), .B(n67996), .C(n58800), .Y(n67813)
         );
  NAND2xp5_ASAP7_75t_SL U61800 ( .A(n58646), .B(n57677), .Y(n58800) );
  NAND2xp5_ASAP7_75t_SL U61801 ( .A(n67609), .B(n67608), .Y(n57677) );
  MAJIxp5_ASAP7_75t_SL U61802 ( .A(n67815), .B(n67814), .C(n67813), .Y(n67890)
         );
  NOR2x1_ASAP7_75t_SL U61803 ( .A(n59440), .B(n57679), .Y(n57678) );
  INVx1_ASAP7_75t_SL U61804 ( .A(n68003), .Y(n57679) );
  NOR2x1_ASAP7_75t_SL U61805 ( .A(n57787), .B(n57680), .Y(n67815) );
  INVx1_ASAP7_75t_SL U61806 ( .A(n57681), .Y(n57680) );
  OR2x2_ASAP7_75t_SL U61807 ( .A(n64556), .B(n64555), .Y(n57682) );
  NOR2x1_ASAP7_75t_SL U61808 ( .A(n64879), .B(n64472), .Y(n64555) );
  NAND2xp5_ASAP7_75t_SL U61809 ( .A(n57683), .B(n57682), .Y(n64908) );
  INVx1_ASAP7_75t_SL U61810 ( .A(n63249), .Y(n63188) );
  OR2x2_ASAP7_75t_SL U61811 ( .A(n60608), .B(n63174), .Y(n63249) );
  NAND2xp5_ASAP7_75t_SL U61812 ( .A(n57696), .B(n57688), .Y(n67466) );
  NAND2xp5_ASAP7_75t_SL U61813 ( .A(n57688), .B(n66333), .Y(n57687) );
  INVx1_ASAP7_75t_SL U61814 ( .A(n67383), .Y(n57688) );
  OAI21xp5_ASAP7_75t_SL U61815 ( .A1(n53271), .A2(n59340), .B(n57689), .Y(
        n67742) );
  NAND2xp5_ASAP7_75t_SL U61816 ( .A(n76077), .B(n67922), .Y(n57689) );
  INVx1_ASAP7_75t_SL U61817 ( .A(n66754), .Y(n66792) );
  OR2x2_ASAP7_75t_SL U61818 ( .A(n57690), .B(n66752), .Y(n66754) );
  INVx1_ASAP7_75t_SL U61819 ( .A(n67615), .Y(n57691) );
  NAND2xp5_ASAP7_75t_SL U61820 ( .A(n57693), .B(n57692), .Y(n67615) );
  A2O1A1Ixp33_ASAP7_75t_SL U61821 ( .A1(n57108), .A2(n75899), .B(n67362), .C(
        n68017), .Y(n57692) );
  NAND2xp5_ASAP7_75t_SL U61822 ( .A(n56390), .B(n57694), .Y(n57693) );
  XOR2xp5_ASAP7_75t_SL U61823 ( .A(n57108), .B(n75947), .Y(n57694) );
  INVx1_ASAP7_75t_SL U61824 ( .A(n68158), .Y(n65062) );
  OAI21xp5_ASAP7_75t_SL U61825 ( .A1(n67569), .A2(n59617), .B(n57695), .Y(
        n68158) );
  NAND2xp5_ASAP7_75t_SL U61826 ( .A(n67846), .B(n57696), .Y(n57695) );
  OR2x2_ASAP7_75t_SL U61827 ( .A(n62574), .B(n62579), .Y(n57698) );
  NOR2x1_ASAP7_75t_SL U61828 ( .A(n58535), .B(n59465), .Y(n57697) );
  NAND2xp5_ASAP7_75t_SL U61829 ( .A(n57699), .B(n58651), .Y(n58368) );
  INVx1_ASAP7_75t_SL U61830 ( .A(n58653), .Y(n57699) );
  NAND2x2_ASAP7_75t_SL U61831 ( .A(n67146), .B(n57700), .Y(n59314) );
  INVx2_ASAP7_75t_SL U61832 ( .A(n58004), .Y(n57700) );
  NAND2x1_ASAP7_75t_SL U61833 ( .A(n59597), .B(n56844), .Y(n67146) );
  OAI21x1_ASAP7_75t_SL U61834 ( .A1(n59601), .A2(n57701), .B(n58456), .Y(
        n67626) );
  NAND2xp5_ASAP7_75t_SL U61835 ( .A(n62727), .B(n63218), .Y(n57704) );
  MAJIxp5_ASAP7_75t_SL U61836 ( .A(n63057), .B(n57708), .C(n63058), .Y(n63140)
         );
  NAND3x1_ASAP7_75t_SL U61837 ( .A(n57705), .B(n57704), .C(n57703), .Y(n62730)
         );
  OAI21x1_ASAP7_75t_SL U61838 ( .A1(n62728), .A2(n57360), .B(n57707), .Y(
        n62729) );
  NOR2x1p5_ASAP7_75t_SL U61839 ( .A(n59619), .B(n57711), .Y(n57709) );
  NAND2xp5_ASAP7_75t_SL U61840 ( .A(n59483), .B(n57924), .Y(n57710) );
  XOR2x2_ASAP7_75t_SL U61841 ( .A(n59456), .B(n59508), .Y(n57711) );
  MAJIxp5_ASAP7_75t_SL U61842 ( .A(n66520), .B(n66519), .C(n66436), .Y(n66443)
         );
  OR2x2_ASAP7_75t_SL U61843 ( .A(n57712), .B(n66449), .Y(n66520) );
  NOR2x1_ASAP7_75t_SL U61844 ( .A(n66445), .B(n66446), .Y(n66449) );
  NOR2x1_ASAP7_75t_SL U61845 ( .A(n57714), .B(n57713), .Y(n59272) );
  NOR2x1_ASAP7_75t_SL U61846 ( .A(n75080), .B(n75104), .Y(n57714) );
  NOR2x1_ASAP7_75t_SL U61847 ( .A(n75111), .B(n57715), .Y(n75104) );
  NOR2x1_ASAP7_75t_SL U61848 ( .A(n75106), .B(n75059), .Y(n57715) );
  INVx1_ASAP7_75t_SL U61849 ( .A(n65061), .Y(n57716) );
  NAND2xp5_ASAP7_75t_SL U61850 ( .A(n59466), .B(n76049), .Y(n57717) );
  NAND2x1_ASAP7_75t_SL U61851 ( .A(n58397), .B(n58743), .Y(n57718) );
  NOR2x1_ASAP7_75t_SL U61852 ( .A(n57155), .B(n57719), .Y(n67992) );
  AND2x2_ASAP7_75t_SL U61853 ( .A(n57155), .B(n57719), .Y(n68000) );
  OAI21x1_ASAP7_75t_SL U61854 ( .A1(n67823), .A2(n59440), .B(n56989), .Y(
        n57719) );
  OR2x2_ASAP7_75t_SL U61855 ( .A(n57181), .B(n58719), .Y(n67328) );
  INVx1_ASAP7_75t_SL U61856 ( .A(n67328), .Y(n57720) );
  XNOR2x1_ASAP7_75t_SL U61857 ( .A(n59319), .B(n57721), .Y(n58847) );
  XNOR2x1_ASAP7_75t_SL U61858 ( .A(n57722), .B(n59318), .Y(n57721) );
  XNOR2x1_ASAP7_75t_SL U61859 ( .A(n67529), .B(n57723), .Y(n59318) );
  AOI21x1_ASAP7_75t_SL U61860 ( .A1(n67400), .A2(n58911), .B(n58910), .Y(
        n57722) );
  O2A1O1Ixp5_ASAP7_75t_SL U61861 ( .A1(n67651), .A2(n67767), .B(n67649), .C(
        n67380), .Y(n67400) );
  XNOR2x1_ASAP7_75t_SL U61862 ( .A(n57765), .B(n57766), .Y(n67529) );
  XNOR2xp5_ASAP7_75t_SL U61863 ( .A(n68039), .B(n57724), .Y(n68053) );
  XNOR2xp5_ASAP7_75t_SL U61864 ( .A(n68040), .B(n68041), .Y(n57724) );
  INVx1_ASAP7_75t_SL U61865 ( .A(n67789), .Y(n57725) );
  XNOR2xp5_ASAP7_75t_SL U61866 ( .A(n67790), .B(n59131), .Y(n57726) );
  AOI21xp5_ASAP7_75t_SL U61867 ( .A1(n67918), .A2(n59651), .B(n59135), .Y(
        n57729) );
  INVx1_ASAP7_75t_SL U61868 ( .A(n58059), .Y(n57730) );
  XNOR2xp5_ASAP7_75t_SL U61869 ( .A(n64715), .B(n64714), .Y(n57731) );
  XNOR2x1_ASAP7_75t_SL U61870 ( .A(n64662), .B(n64661), .Y(n64713) );
  NAND3x1_ASAP7_75t_SL U61871 ( .A(n74992), .B(n74993), .C(n65114), .Y(n64730)
         );
  NAND2x1_ASAP7_75t_SL U61872 ( .A(n64728), .B(n64729), .Y(n65114) );
  NAND2x1_ASAP7_75t_SL U61873 ( .A(n64094), .B(n64093), .Y(n64729) );
  XNOR2x1_ASAP7_75t_SL U61874 ( .A(n64725), .B(n57732), .Y(n64733) );
  NAND2x1_ASAP7_75t_SL U61875 ( .A(n57864), .B(n64736), .Y(n74992) );
  XNOR2x1_ASAP7_75t_SL U61876 ( .A(n64713), .B(n57731), .Y(n64736) );
  XNOR2x1_ASAP7_75t_SL U61877 ( .A(n64708), .B(n57866), .Y(n64725) );
  INVx1_ASAP7_75t_SL U61878 ( .A(n57864), .Y(n64738) );
  XNOR2xp5_ASAP7_75t_SL U61879 ( .A(n64092), .B(n57748), .Y(n64093) );
  OR2x2_ASAP7_75t_SL U61880 ( .A(n57912), .B(n59661), .Y(n66396) );
  OAI22xp33_ASAP7_75t_SL U61881 ( .A1(n59508), .A2(n59072), .B1(n59514), .B2(
        n67826), .Y(n57735) );
  NAND2xp5_ASAP7_75t_SL U61882 ( .A(n59193), .B(n66705), .Y(n57736) );
  OAI21xp5_ASAP7_75t_SL U61883 ( .A1(n66846), .A2(n66987), .B(n57736), .Y(
        n69139) );
  NAND2xp5_ASAP7_75t_SL U61884 ( .A(n59661), .B(n57180), .Y(n67925) );
  INVx1_ASAP7_75t_SL U61885 ( .A(n67899), .Y(n67740) );
  NOR2x1_ASAP7_75t_SL U61886 ( .A(n57446), .B(n63663), .Y(n67899) );
  XNOR2x2_ASAP7_75t_SL U61887 ( .A(n57742), .B(n57737), .Y(n68325) );
  XNOR2xp5_ASAP7_75t_SL U61888 ( .A(n68204), .B(n57738), .Y(n57737) );
  XNOR2xp5_ASAP7_75t_SL U61889 ( .A(n68203), .B(n57739), .Y(n57738) );
  XOR2xp5_ASAP7_75t_SL U61890 ( .A(n68202), .B(n59313), .Y(n57739) );
  XNOR2xp5_ASAP7_75t_SL U61891 ( .A(n57741), .B(n57740), .Y(n68204) );
  INVx1_ASAP7_75t_SL U61892 ( .A(n68139), .Y(n57741) );
  NAND2xp5_ASAP7_75t_SL U61893 ( .A(n68200), .B(n57743), .Y(n57742) );
  NAND2xp5_ASAP7_75t_SL U61894 ( .A(n57744), .B(n68201), .Y(n57743) );
  INVx1_ASAP7_75t_SL U61895 ( .A(n68199), .Y(n57744) );
  XNOR2xp5_ASAP7_75t_SL U61896 ( .A(n57746), .B(n68156), .Y(n57745) );
  NOR2x1_ASAP7_75t_SL U61897 ( .A(n68157), .B(n57747), .Y(n57746) );
  NOR2x1_ASAP7_75t_SL U61898 ( .A(n68158), .B(n58903), .Y(n57747) );
  NOR2x1_ASAP7_75t_SL U61899 ( .A(n64699), .B(n64700), .Y(n65101) );
  NOR2x1_ASAP7_75t_SL U61900 ( .A(n64094), .B(n64093), .Y(n64700) );
  XOR2xp5_ASAP7_75t_SL U61901 ( .A(n64723), .B(n64091), .Y(n57748) );
  OAI21xp5_ASAP7_75t_SL U61902 ( .A1(n59511), .A2(n59641), .B(n57749), .Y(
        n58699) );
  NAND3xp33_ASAP7_75t_SL U61903 ( .A(n57425), .B(n59511), .C(n59485), .Y(
        n57749) );
  INVx1_ASAP7_75t_SL U61904 ( .A(n58927), .Y(n61916) );
  INVx1_ASAP7_75t_SL U61905 ( .A(n66734), .Y(n66913) );
  NAND2xp5_ASAP7_75t_SL U61906 ( .A(n59347), .B(n68483), .Y(n66734) );
  NAND2xp5_ASAP7_75t_SL U61907 ( .A(n68479), .B(n68480), .Y(n68483) );
  NOR3xp33_ASAP7_75t_SL U61908 ( .A(n58276), .B(n59053), .C(n59429), .Y(n57750) );
  NAND2xp5_ASAP7_75t_SL U61909 ( .A(n57753), .B(n57206), .Y(n57754) );
  NAND3x1_ASAP7_75t_SL U61910 ( .A(n57751), .B(n56828), .C(n57750), .Y(n64619)
         );
  NOR2x1p5_ASAP7_75t_SL U61911 ( .A(n60599), .B(n57752), .Y(n57751) );
  NOR2x1_ASAP7_75t_SL U61912 ( .A(n57755), .B(n57754), .Y(n60917) );
  AOI21x1_ASAP7_75t_SL U61913 ( .A1(n57024), .A2(n63819), .B(n57756), .Y(
        n64678) );
  NAND2xp5_ASAP7_75t_SL U61914 ( .A(n57758), .B(n57757), .Y(n57756) );
  NAND2xp5_ASAP7_75t_SL U61915 ( .A(n57148), .B(n57759), .Y(n57757) );
  AOI22xp5_ASAP7_75t_SL U61916 ( .A1(n63819), .A2(n63865), .B1(n63666), .B2(
        n57148), .Y(n57758) );
  NOR2x1_ASAP7_75t_SL U61917 ( .A(n64024), .B(n64023), .Y(n64416) );
  MAJIxp5_ASAP7_75t_SL U61918 ( .A(n66543), .B(n66586), .C(n66588), .Y(n66567)
         );
  NOR2x1_ASAP7_75t_SL U61919 ( .A(n57763), .B(n57762), .Y(n66588) );
  O2A1O1Ixp5_ASAP7_75t_SL U61920 ( .A1(n75947), .A2(n58784), .B(n66538), .C(
        n57764), .Y(n57763) );
  NAND2xp5_ASAP7_75t_SL U61921 ( .A(n67365), .B(n57277), .Y(n57764) );
  NOR2x1_ASAP7_75t_SL U61922 ( .A(n66398), .B(n58143), .Y(n58819) );
  XNOR2xp5_ASAP7_75t_SL U61923 ( .A(n64702), .B(n64703), .Y(n64704) );
  XNOR2xp5_ASAP7_75t_SL U61924 ( .A(n64430), .B(n57769), .Y(n64702) );
  XOR2xp5_ASAP7_75t_SL U61925 ( .A(n64462), .B(n64463), .Y(n57769) );
  OAI21xp5_ASAP7_75t_SL U61926 ( .A1(n68075), .A2(n57772), .B(n57771), .Y(
        n67886) );
  INVx1_ASAP7_75t_SL U61927 ( .A(n68046), .Y(n57771) );
  NOR2x1_ASAP7_75t_SL U61928 ( .A(n68073), .B(n68074), .Y(n68046) );
  INVx1_ASAP7_75t_SL U61929 ( .A(n68048), .Y(n57772) );
  INVx1_ASAP7_75t_SL U61930 ( .A(n66978), .Y(n68553) );
  XOR2xp5_ASAP7_75t_SL U61931 ( .A(n57773), .B(n59005), .Y(n66978) );
  INVx1_ASAP7_75t_SL U61932 ( .A(n66673), .Y(n57773) );
  NOR2x1_ASAP7_75t_SL U61933 ( .A(n53623), .B(n58948), .Y(n57774) );
  MAJIxp5_ASAP7_75t_SL U61934 ( .A(n57776), .B(n57775), .C(n57235), .Y(n68069)
         );
  INVx1_ASAP7_75t_SL U61935 ( .A(n67985), .Y(n57775) );
  XOR2xp5_ASAP7_75t_SL U61936 ( .A(n58715), .B(n57008), .Y(n57776) );
  NOR2x1_ASAP7_75t_SL U61937 ( .A(n68068), .B(n68070), .Y(n57777) );
  XNOR2xp5_ASAP7_75t_SL U61938 ( .A(n58792), .B(n67801), .Y(n57778) );
  A2O1A1Ixp33_ASAP7_75t_SL U61939 ( .A1(n68412), .A2(n59620), .B(n68411), .C(
        n57779), .Y(n68468) );
  AOI22xp5_ASAP7_75t_SL U61940 ( .A1(n57284), .A2(n68409), .B1(n75903), .B2(
        n58784), .Y(n57779) );
  AND2x2_ASAP7_75t_SL U61941 ( .A(n57078), .B(n67639), .Y(n58784) );
  NOR2x1_ASAP7_75t_SL U61942 ( .A(n57322), .B(n56862), .Y(n68409) );
  XNOR2xp5_ASAP7_75t_SL U61943 ( .A(n58734), .B(n64436), .Y(n64056) );
  MAJIxp5_ASAP7_75t_SL U61944 ( .A(n64054), .B(n64053), .C(n64055), .Y(n58734)
         );
  NOR2x1_ASAP7_75t_SL U61945 ( .A(n66422), .B(n63865), .Y(n64053) );
  NOR2x1_ASAP7_75t_SL U61946 ( .A(n57111), .B(n57253), .Y(n63865) );
  NAND2xp5_ASAP7_75t_SL U61947 ( .A(n63862), .B(n57780), .Y(n64054) );
  NAND2xp5_ASAP7_75t_SL U61948 ( .A(n57375), .B(n58767), .Y(n57780) );
  INVx1_ASAP7_75t_SL U61949 ( .A(n69031), .Y(n69043) );
  AO21x1_ASAP7_75t_SL U61950 ( .A1(n57060), .A2(n69030), .B(n69033), .Y(n69031) );
  INVx1_ASAP7_75t_SL U61951 ( .A(n69027), .Y(n69033) );
  NAND2xp5_ASAP7_75t_SL U61952 ( .A(n68589), .B(n68590), .Y(n69027) );
  NAND2xp5_ASAP7_75t_SL U61953 ( .A(n57012), .B(n58898), .Y(n57786) );
  NOR2x1_ASAP7_75t_SL U61954 ( .A(n58787), .B(n57788), .Y(n57787) );
  INVx1_ASAP7_75t_SL U61955 ( .A(n67812), .Y(n57788) );
  NOR2x1_ASAP7_75t_SL U61956 ( .A(n75915), .B(n57791), .Y(n62748) );
  NOR2x1_ASAP7_75t_SL U61957 ( .A(n61809), .B(n61808), .Y(n57791) );
  INVx1_ASAP7_75t_SL U61958 ( .A(n61809), .Y(n57789) );
  INVx1_ASAP7_75t_SL U61959 ( .A(n61808), .Y(n57790) );
  A2O1A1Ixp33_ASAP7_75t_SL U61960 ( .A1(n57791), .A2(n57118), .B(n58433), .C(
        n77701), .Y(n63860) );
  XNOR2xp5_ASAP7_75t_SL U61961 ( .A(n68309), .B(n68310), .Y(n57792) );
  OAI22x1_ASAP7_75t_SL U61962 ( .A1(n68321), .A2(n57794), .B1(n57793), .B2(
        n68322), .Y(n68329) );
  O2A1O1Ixp5_ASAP7_75t_SL U61963 ( .A1(n68319), .A2(n57795), .B(n57796), .C(
        n68320), .Y(n57793) );
  INVx1_ASAP7_75t_SL U61964 ( .A(n68320), .Y(n57794) );
  AOI21x1_ASAP7_75t_SL U61965 ( .A1(n68319), .A2(n57796), .B(n57795), .Y(
        n68321) );
  INVx1_ASAP7_75t_SL U61966 ( .A(n57798), .Y(n63127) );
  OAI21xp5_ASAP7_75t_SL U61967 ( .A1(n63184), .A2(n57798), .B(n57665), .Y(
        n63187) );
  INVx3_ASAP7_75t_SL U61968 ( .A(n59452), .Y(n67974) );
  NAND4xp25_ASAP7_75t_SL U61969 ( .A(n57802), .B(n65020), .C(n58810), .D(
        n65021), .Y(n58809) );
  INVx2_ASAP7_75t_SL U61970 ( .A(n58809), .Y(n67861) );
  NAND2xp5_ASAP7_75t_SL U61971 ( .A(n65021), .B(n65020), .Y(n66291) );
  AND2x2_ASAP7_75t_SL U61972 ( .A(n58844), .B(n66291), .Y(n66625) );
  XNOR2xp5_ASAP7_75t_SL U61973 ( .A(n68042), .B(n68043), .Y(n68044) );
  MAJIxp5_ASAP7_75t_SL U61974 ( .A(n67770), .B(n67658), .C(n57803), .Y(n68042)
         );
  XNOR2xp5_ASAP7_75t_SL U61975 ( .A(n57095), .B(n67768), .Y(n57803) );
  XNOR2xp5_ASAP7_75t_SL U61976 ( .A(n57805), .B(n57804), .Y(n68043) );
  XOR2xp5_ASAP7_75t_SL U61977 ( .A(n58703), .B(n67660), .Y(n57804) );
  INVx1_ASAP7_75t_SL U61978 ( .A(n67661), .Y(n57805) );
  OR2x2_ASAP7_75t_SL U61979 ( .A(n57806), .B(n64621), .Y(n65020) );
  NAND2xp5_ASAP7_75t_SL U61980 ( .A(n57807), .B(n59590), .Y(n57806) );
  NAND2xp5_ASAP7_75t_SL U61981 ( .A(n57810), .B(n57809), .Y(n58959) );
  NAND3xp33_ASAP7_75t_SL U61982 ( .A(n65035), .B(n59606), .C(n56854), .Y(
        n57809) );
  INVx1_ASAP7_75t_SL U61983 ( .A(n67820), .Y(n57810) );
  NOR2x1_ASAP7_75t_SL U61984 ( .A(n59467), .B(n67962), .Y(n67820) );
  NAND2x1_ASAP7_75t_SL U61985 ( .A(n59397), .B(n62675), .Y(n57811) );
  INVx3_ASAP7_75t_SL U61986 ( .A(n75915), .Y(n59655) );
  NAND2xp5_ASAP7_75t_SL U61987 ( .A(n66641), .B(n66971), .Y(n66644) );
  NOR2x1_ASAP7_75t_SL U61988 ( .A(n66941), .B(n66939), .Y(n66971) );
  INVx1_ASAP7_75t_SL U61989 ( .A(n66940), .Y(n66939) );
  NAND2xp5_ASAP7_75t_SL U61990 ( .A(n56850), .B(n56997), .Y(n66940) );
  AOI22xp5_ASAP7_75t_SL U61991 ( .A1(n57067), .A2(n66749), .B1(n66953), .B2(
        n59100), .Y(n66941) );
  OAI21xp5_ASAP7_75t_SL U61992 ( .A1(n75903), .A2(n59637), .B(n66630), .Y(
        n66953) );
  NAND2xp5_ASAP7_75t_SL U61993 ( .A(n66969), .B(n57812), .Y(n66641) );
  OAI21xp5_ASAP7_75t_SL U61994 ( .A1(n57158), .A2(n66793), .B(n66633), .Y(
        n66970) );
  NAND2xp33_ASAP7_75t_SL U61995 ( .A(n66330), .B(n66329), .Y(n57813) );
  NAND2xp5_ASAP7_75t_SL U61996 ( .A(n57813), .B(n57814), .Y(n66340) );
  OR2x2_ASAP7_75t_SL U61997 ( .A(n66330), .B(n66329), .Y(n57814) );
  INVx1_ASAP7_75t_SL U61998 ( .A(n57814), .Y(n66556) );
  INVxp67_ASAP7_75t_SL U61999 ( .A(n66329), .Y(n66335) );
  NAND2xp5_ASAP7_75t_SL U62000 ( .A(n67901), .B(n57815), .Y(n67260) );
  AO21x1_ASAP7_75t_SL U62001 ( .A1(n53315), .A2(n57662), .B(n57816), .Y(n67825) );
  NAND2xp5_ASAP7_75t_SL U62002 ( .A(n59117), .B(n57111), .Y(n67857) );
  OR2x2_ASAP7_75t_SL U62003 ( .A(n67326), .B(n68078), .Y(n67749) );
  NAND2xp5_ASAP7_75t_SL U62004 ( .A(n59590), .B(n57817), .Y(n67326) );
  XNOR2x1_ASAP7_75t_SL U62005 ( .A(n58120), .B(n58121), .Y(n68309) );
  MAJIxp5_ASAP7_75t_SL U62006 ( .A(n58726), .B(n68288), .C(n68289), .Y(n68310)
         );
  XNOR2xp5_ASAP7_75t_SL U62007 ( .A(n57819), .B(n64076), .Y(n58100) );
  INVx1_ASAP7_75t_SL U62008 ( .A(n64347), .Y(n57819) );
  NAND2xp5_ASAP7_75t_SL U62009 ( .A(n59656), .B(n57422), .Y(n57820) );
  OAI21xp5_ASAP7_75t_SL U62010 ( .A1(n75947), .A2(n57821), .B(n67903), .Y(
        n67904) );
  INVx1_ASAP7_75t_SL U62011 ( .A(n67864), .Y(n57821) );
  OAI21xp5_ASAP7_75t_SL U62012 ( .A1(n57173), .A2(n57422), .B(n57178), .Y(
        n57822) );
  NAND2xp5_ASAP7_75t_SL U62013 ( .A(n57823), .B(n64421), .Y(n64422) );
  OAI21xp5_ASAP7_75t_SL U62014 ( .A1(n57422), .A2(n57107), .B(n57178), .Y(
        n57823) );
  XOR2xp5_ASAP7_75t_SL U62015 ( .A(n68489), .B(n68444), .Y(n57824) );
  INVx1_ASAP7_75t_SL U62016 ( .A(n68490), .Y(n57825) );
  MAJIxp5_ASAP7_75t_SL U62017 ( .A(n68437), .B(n68435), .C(n68436), .Y(n68490)
         );
  AOI22xp5_ASAP7_75t_SL U62018 ( .A1(n58152), .A2(n58153), .B1(n68404), .B2(
        n58149), .Y(n68437) );
  INVx1_ASAP7_75t_SL U62019 ( .A(n67821), .Y(n67442) );
  INVx1_ASAP7_75t_SL U62020 ( .A(n67447), .Y(n67622) );
  OAI21xp5_ASAP7_75t_SL U62021 ( .A1(n53258), .A2(n58919), .B(n57827), .Y(
        n57826) );
  NOR2x1_ASAP7_75t_SL U62022 ( .A(n67441), .B(n63097), .Y(n67821) );
  OAI21xp5_ASAP7_75t_SL U62023 ( .A1(n57171), .A2(n57829), .B(n57023), .Y(
        n57828) );
  NAND2xp5_ASAP7_75t_SL U62024 ( .A(n59200), .B(n63120), .Y(n57829) );
  AOI21xp5_ASAP7_75t_SL U62025 ( .A1(n68048), .A2(n58354), .B(n68046), .Y(
        n68066) );
  INVx1_ASAP7_75t_SL U62026 ( .A(n68065), .Y(n57830) );
  XNOR2xp5_ASAP7_75t_SL U62027 ( .A(n57832), .B(n57831), .Y(n67940) );
  XOR2xp5_ASAP7_75t_SL U62028 ( .A(n67579), .B(n67578), .Y(n57831) );
  NOR2x1_ASAP7_75t_SL U62029 ( .A(n67771), .B(n57833), .Y(n67394) );
  NOR2x1_ASAP7_75t_SL U62030 ( .A(n67772), .B(n57834), .Y(n57833) );
  NOR2x1_ASAP7_75t_SL U62031 ( .A(n67349), .B(n67348), .Y(n67771) );
  AND2x2_ASAP7_75t_SL U62032 ( .A(n57834), .B(n67772), .Y(n67395) );
  INVx1_ASAP7_75t_SL U62033 ( .A(n67107), .Y(n67106) );
  NAND2xp5_ASAP7_75t_SL U62034 ( .A(n69140), .B(n57835), .Y(n67107) );
  NAND2xp5_ASAP7_75t_SL U62035 ( .A(n57836), .B(n67104), .Y(n57835) );
  INVx1_ASAP7_75t_SL U62036 ( .A(n69142), .Y(n57836) );
  NOR2x1_ASAP7_75t_SL U62037 ( .A(n57837), .B(n67105), .Y(n69142) );
  NAND2xp5_ASAP7_75t_SL U62038 ( .A(n57837), .B(n67105), .Y(n69140) );
  INVx1_ASAP7_75t_SL U62039 ( .A(n67103), .Y(n57837) );
  INVx1_ASAP7_75t_SL U62040 ( .A(n59333), .Y(n57838) );
  NAND2xp5_ASAP7_75t_SL U62041 ( .A(n59547), .B(n61915), .Y(n59333) );
  NOR2x1_ASAP7_75t_SL U62042 ( .A(n59095), .B(n61912), .Y(n61915) );
  INVx1_ASAP7_75t_SL U62043 ( .A(n63019), .Y(n63024) );
  XNOR2xp5_ASAP7_75t_SL U62044 ( .A(n57840), .B(n57839), .Y(n63019) );
  XOR2xp5_ASAP7_75t_SL U62045 ( .A(n63035), .B(n63034), .Y(n57839) );
  INVx1_ASAP7_75t_SL U62046 ( .A(n63033), .Y(n57840) );
  XOR2xp5_ASAP7_75t_SL U62047 ( .A(n63017), .B(n57841), .Y(n63033) );
  INVx1_ASAP7_75t_SL U62048 ( .A(n63018), .Y(n57841) );
  NAND2xp5_ASAP7_75t_SL U62049 ( .A(n75058), .B(n57843), .Y(n68614) );
  NAND2xp5_ASAP7_75t_SL U62050 ( .A(n57845), .B(n57844), .Y(n57843) );
  NAND2xp5_ASAP7_75t_SL U62051 ( .A(n68955), .B(n68730), .Y(n69032) );
  NOR2x1_ASAP7_75t_SL U62052 ( .A(n59383), .B(n57847), .Y(n68730) );
  INVx1_ASAP7_75t_SL U62053 ( .A(n69006), .Y(n57847) );
  INVx1_ASAP7_75t_SL U62054 ( .A(n69012), .Y(n59383) );
  AND2x2_ASAP7_75t_SL U62055 ( .A(n59094), .B(n67398), .Y(n58427) );
  AOI21x1_ASAP7_75t_SL U62056 ( .A1(n57851), .A2(n53486), .B(n57850), .Y(
        n67398) );
  NOR2xp67_ASAP7_75t_SL U62057 ( .A(n57852), .B(n67786), .Y(n57850) );
  NAND2x1_ASAP7_75t_SL U62058 ( .A(n57852), .B(n67786), .Y(n57851) );
  INVx1_ASAP7_75t_SL U62059 ( .A(n67787), .Y(n57852) );
  XNOR2xp5_ASAP7_75t_SL U62060 ( .A(n57855), .B(n57048), .Y(n59094) );
  XOR2xp5_ASAP7_75t_SL U62061 ( .A(n67485), .B(n67486), .Y(n57855) );
  INVx1_ASAP7_75t_SL U62062 ( .A(n59232), .Y(n57856) );
  NAND2xp5_ASAP7_75t_SL U62063 ( .A(n68188), .B(n57859), .Y(n57857) );
  NOR3xp33_ASAP7_75t_SL U62064 ( .A(n67997), .B(n57860), .C(n57859), .Y(n57858) );
  INVx1_ASAP7_75t_SL U62065 ( .A(n68187), .Y(n57859) );
  XOR2xp5_ASAP7_75t_SL U62066 ( .A(n58800), .B(n57955), .Y(n68187) );
  INVx1_ASAP7_75t_SL U62067 ( .A(n68027), .Y(n57860) );
  AND2x2_ASAP7_75t_SL U62068 ( .A(n57036), .B(n62793), .Y(n59308) );
  INVx1_ASAP7_75t_SL U62069 ( .A(n68116), .Y(n57863) );
  XOR2xp5_ASAP7_75t_SL U62070 ( .A(n64707), .B(n64706), .Y(n57866) );
  NOR2x1_ASAP7_75t_SL U62071 ( .A(n57865), .B(n64731), .Y(n57864) );
  AOI21x1_ASAP7_75t_SL U62072 ( .A1(n64725), .A2(n64726), .B(n64727), .Y(
        n64731) );
  NOR2x1_ASAP7_75t_SL U62073 ( .A(n64726), .B(n64725), .Y(n57865) );
  INVx1_ASAP7_75t_SL U62074 ( .A(n68471), .Y(n57867) );
  INVx1_ASAP7_75t_SL U62075 ( .A(n68391), .Y(n57868) );
  NAND2x1_ASAP7_75t_SL U62076 ( .A(n65070), .B(n65069), .Y(n68756) );
  NOR2x1_ASAP7_75t_SL U62077 ( .A(n65069), .B(n65070), .Y(n68346) );
  INVx2_ASAP7_75t_SL U62078 ( .A(n68753), .Y(n58731) );
  OR2x2_ASAP7_75t_SL U62079 ( .A(n68348), .B(n68347), .Y(n68753) );
  NAND2xp5_ASAP7_75t_SL U62080 ( .A(n59664), .B(n57243), .Y(n67376) );
  OAI21xp5_ASAP7_75t_SL U62081 ( .A1(n67933), .A2(n67932), .B(n67931), .Y(
        n58253) );
  NAND2xp5_ASAP7_75t_SL U62082 ( .A(n57871), .B(n58254), .Y(n67931) );
  INVx1_ASAP7_75t_SL U62083 ( .A(n67993), .Y(n57871) );
  AOI22xp5_ASAP7_75t_SL U62084 ( .A1(n67842), .A2(n67824), .B1(n57380), .B2(
        n67825), .Y(n67993) );
  OAI22xp5_ASAP7_75t_SL U62085 ( .A1(n68003), .A2(n57099), .B1(n68004), .B2(
        n59454), .Y(n68182) );
  INVx1_ASAP7_75t_SL U62086 ( .A(n67629), .Y(n58990) );
  NAND3xp33_ASAP7_75t_SL U62087 ( .A(n67416), .B(n57166), .C(n58803), .Y(
        n67810) );
  OR2x2_ASAP7_75t_SL U62088 ( .A(n59593), .B(n67629), .Y(n67416) );
  A2O1A1Ixp33_ASAP7_75t_SL U62089 ( .A1(n57877), .A2(n64675), .B(n63803), .C(
        n63804), .Y(n64680) );
  NAND2xp5_ASAP7_75t_SL U62090 ( .A(n57006), .B(n63657), .Y(n63804) );
  OAI21xp5_ASAP7_75t_SL U62091 ( .A1(n57875), .A2(n57158), .B(n57874), .Y(
        n63803) );
  INVx1_ASAP7_75t_SL U62092 ( .A(n63801), .Y(n57875) );
  OAI21xp5_ASAP7_75t_SL U62093 ( .A1(n67850), .A2(n59616), .B(n57876), .Y(
        n63801) );
  NAND2xp5_ASAP7_75t_SL U62094 ( .A(n58402), .B(n67638), .Y(n57876) );
  OAI22xp5_ASAP7_75t_SL U62095 ( .A1(n64035), .A2(n68383), .B1(n59453), .B2(
        n63170), .Y(n64675) );
  NOR2x1_ASAP7_75t_SL U62096 ( .A(n57878), .B(n63189), .Y(n58904) );
  OAI21xp5_ASAP7_75t_SL U62097 ( .A1(n67850), .A2(n67898), .B(n53613), .Y(
        n57878) );
  NAND2x2_ASAP7_75t_SL U62098 ( .A(n59448), .B(n57912), .Y(n66332) );
  NOR2x1p5_ASAP7_75t_SL U62099 ( .A(n53289), .B(n57179), .Y(n59245) );
  NAND2xp5_ASAP7_75t_SRAM U62100 ( .A(n59448), .B(n57184), .Y(n67071) );
  INVx1_ASAP7_75t_SL U62101 ( .A(n62580), .Y(n67596) );
  NAND2x2_ASAP7_75t_SL U62102 ( .A(n62580), .B(n67598), .Y(n67906) );
  NAND2x2_ASAP7_75t_SL U62103 ( .A(n57881), .B(n57880), .Y(n62580) );
  INVx1_ASAP7_75t_SL U62104 ( .A(n58784), .Y(n58785) );
  OAI21xp5_ASAP7_75t_SL U62105 ( .A1(n76057), .A2(n58784), .B(n57882), .Y(
        n66742) );
  NAND2xp5_ASAP7_75t_SL U62106 ( .A(n76057), .B(n75045), .Y(n57882) );
  NAND2xp5_ASAP7_75t_SL U62107 ( .A(n59518), .B(n67532), .Y(n75045) );
  NAND2x1_ASAP7_75t_SL U62108 ( .A(n57884), .B(n57465), .Y(n59043) );
  NOR2x1_ASAP7_75t_SL U62109 ( .A(n59578), .B(n66451), .Y(n57884) );
  XNOR2xp5_ASAP7_75t_SL U62110 ( .A(n66476), .B(n66475), .Y(n66468) );
  AO21x1_ASAP7_75t_SL U62111 ( .A1(n57161), .A2(n66467), .B(n57885), .Y(n66476) );
  NAND2x2_ASAP7_75t_SL U62112 ( .A(n56862), .B(n58711), .Y(n67641) );
  A2O1A1Ixp33_ASAP7_75t_SL U62113 ( .A1(n57274), .A2(n57277), .B(n67239), .C(
        n57886), .Y(n67294) );
  XOR2x1_ASAP7_75t_SL U62114 ( .A(n59644), .B(n59504), .Y(n67594) );
  OAI21xp5_ASAP7_75t_SL U62115 ( .A1(n63475), .A2(n57888), .B(n57887), .Y(
        n58818) );
  NAND2xp5_ASAP7_75t_SL U62116 ( .A(n63476), .B(n63477), .Y(n57888) );
  NAND3xp33_ASAP7_75t_SL U62117 ( .A(n57890), .B(n63882), .C(n58813), .Y(
        n63880) );
  OAI21xp5_ASAP7_75t_SL U62118 ( .A1(n63361), .A2(n58817), .B(n57889), .Y(
        n58813) );
  AOI211x1_ASAP7_75t_SL U62119 ( .A1(n63045), .A2(n63444), .B(n63475), .C(
        n58814), .Y(n57889) );
  NOR2x1_ASAP7_75t_SL U62120 ( .A(n63877), .B(n63878), .Y(n63882) );
  NOR2x1_ASAP7_75t_SL U62121 ( .A(n63686), .B(n63685), .Y(n63877) );
  AO21x2_ASAP7_75t_SL U62122 ( .A1(n58495), .A2(n59215), .B(n59216), .Y(n59461) );
  NOR2x1_ASAP7_75t_SL U62123 ( .A(n58943), .B(n57894), .Y(n68245) );
  NOR2x1_ASAP7_75t_SL U62124 ( .A(n64504), .B(n59481), .Y(n66271) );
  NAND2xp5_ASAP7_75t_SL U62125 ( .A(n59104), .B(n59108), .Y(n57895) );
  NAND2xp5_ASAP7_75t_SL U62126 ( .A(n59107), .B(n62573), .Y(n57896) );
  NAND3xp33_ASAP7_75t_SL U62127 ( .A(n62553), .B(n62554), .C(n62562), .Y(
        n62573) );
  XNOR2xp5_ASAP7_75t_SL U62128 ( .A(n63106), .B(n63105), .Y(n57897) );
  NOR2x1_ASAP7_75t_SL U62129 ( .A(n57898), .B(n62733), .Y(n63054) );
  INVx1_ASAP7_75t_SL U62130 ( .A(n57899), .Y(n57898) );
  AND2x2_ASAP7_75t_SL U62131 ( .A(n57284), .B(n67601), .Y(n62587) );
  INVx1_ASAP7_75t_SL U62132 ( .A(n69227), .Y(n68628) );
  AOI21xp5_ASAP7_75t_SL U62133 ( .A1(n57903), .A2(n57902), .B(n57901), .Y(
        n75105) );
  AO21x1_ASAP7_75t_SL U62134 ( .A1(n68666), .A2(n68678), .B(n59195), .Y(n59274) );
  OR2x2_ASAP7_75t_SL U62135 ( .A(n57087), .B(n69227), .Y(n68678) );
  NOR2x1_ASAP7_75t_SL U62136 ( .A(n57132), .B(n59271), .Y(n57902) );
  AND2x2_ASAP7_75t_SL U62137 ( .A(n74112), .B(n68684), .Y(n59271) );
  NAND2xp5_ASAP7_75t_SL U62138 ( .A(n68624), .B(n68623), .Y(n68685) );
  INVx1_ASAP7_75t_SL U62139 ( .A(n59275), .Y(n57903) );
  XOR2xp5_ASAP7_75t_SL U62140 ( .A(n62995), .B(n62988), .Y(n63363) );
  NOR2x1_ASAP7_75t_SL U62141 ( .A(n59227), .B(n59228), .Y(n63004) );
  OAI21xp5_ASAP7_75t_SL U62142 ( .A1(n56985), .A2(n75036), .B(n57905), .Y(
        n66688) );
  NAND2xp5_ASAP7_75t_SL U62143 ( .A(n66666), .B(n59100), .Y(n57905) );
  INVx1_ASAP7_75t_SL U62144 ( .A(n59370), .Y(n64710) );
  OR2x2_ASAP7_75t_SL U62145 ( .A(n64046), .B(n64044), .Y(n59370) );
  OAI21xp5_ASAP7_75t_SL U62146 ( .A1(n63805), .A2(n57906), .B(n64680), .Y(
        n64044) );
  INVx1_ASAP7_75t_SL U62147 ( .A(n64676), .Y(n57906) );
  INVx1_ASAP7_75t_SL U62148 ( .A(n64677), .Y(n64046) );
  INVx1_ASAP7_75t_SL U62149 ( .A(n59226), .Y(n59228) );
  OR2x2_ASAP7_75t_SL U62150 ( .A(n62964), .B(n62963), .Y(n59226) );
  O2A1O1Ixp33_ASAP7_75t_SL U62151 ( .A1(n57292), .A2(n67244), .B(n67243), .C(
        n65022), .Y(n59374) );
  NOR2x1_ASAP7_75t_SL U62152 ( .A(n56982), .B(n59335), .Y(n65022) );
  NAND2xp5_ASAP7_75t_SL U62153 ( .A(n63853), .B(n63852), .Y(n64059) );
  OA21x2_ASAP7_75t_SL U62154 ( .A1(n59073), .A2(n63843), .B(n57907), .Y(n63852) );
  NAND2xp5_ASAP7_75t_SL U62155 ( .A(n57478), .B(n63613), .Y(n57907) );
  OAI21xp5_ASAP7_75t_SL U62156 ( .A1(n59620), .A2(n58931), .B(n58936), .Y(
        n63843) );
  NAND2xp5_ASAP7_75t_SL U62157 ( .A(n58384), .B(n58786), .Y(n64503) );
  OA21x2_ASAP7_75t_SL U62158 ( .A1(n64356), .A2(n58210), .B(n58209), .Y(n58384) );
  XNOR2xp5_ASAP7_75t_SL U62159 ( .A(n59594), .B(n59652), .Y(n64406) );
  OAI21xp5_ASAP7_75t_SL U62160 ( .A1(n68243), .A2(n57423), .B(n68141), .Y(
        n57908) );
  NAND2xp5_ASAP7_75t_SL U62161 ( .A(n57423), .B(n68243), .Y(n57909) );
  XNOR2xp5_ASAP7_75t_SL U62162 ( .A(n68064), .B(n68063), .Y(n68243) );
  INVx1_ASAP7_75t_SL U62163 ( .A(n68827), .Y(n68571) );
  NAND2xp5_ASAP7_75t_SL U62164 ( .A(n68828), .B(n68827), .Y(n68718) );
  XNOR2xp5_ASAP7_75t_SL U62165 ( .A(n64888), .B(n64887), .Y(n64613) );
  OAI21x1_ASAP7_75t_SL U62166 ( .A1(n59067), .A2(n64612), .B(n57910), .Y(
        n64887) );
  OAI21x1_ASAP7_75t_SL U62167 ( .A1(n65042), .A2(n67434), .B(n64610), .Y(
        n64888) );
  AOI22xp5_ASAP7_75t_SL U62168 ( .A1(n67401), .A2(n66764), .B1(n57463), .B2(
        n66830), .Y(n66826) );
  INVx1_ASAP7_75t_SL U62169 ( .A(n67467), .Y(n67360) );
  MAJIxp5_ASAP7_75t_SL U62170 ( .A(n66825), .B(n66824), .C(n66826), .Y(n66849)
         );
  NOR2x1_ASAP7_75t_SL U62171 ( .A(n74781), .B(n61912), .Y(n57913) );
  INVx1_ASAP7_75t_SL U62172 ( .A(n67155), .Y(n67154) );
  NAND2xp5_ASAP7_75t_SL U62173 ( .A(n57916), .B(n57914), .Y(n67155) );
  NAND2xp5_ASAP7_75t_SL U62174 ( .A(n57260), .B(n57915), .Y(n57914) );
  OAI21xp5_ASAP7_75t_SL U62175 ( .A1(n58861), .A2(n75644), .B(n67060), .Y(
        n57915) );
  NAND2xp5_ASAP7_75t_SL U62176 ( .A(n67061), .B(n67715), .Y(n57916) );
  XNOR2xp5_ASAP7_75t_SL U62177 ( .A(n67942), .B(n57919), .Y(n59428) );
  MAJIxp5_ASAP7_75t_SL U62178 ( .A(n67890), .B(n67889), .C(n67888), .Y(n67942)
         );
  XNOR2xp5_ASAP7_75t_SL U62179 ( .A(n67614), .B(n57917), .Y(n67889) );
  XOR2xp5_ASAP7_75t_SL U62180 ( .A(n67613), .B(n57918), .Y(n57917) );
  INVx1_ASAP7_75t_SL U62181 ( .A(n67612), .Y(n57918) );
  NAND2xp5_ASAP7_75t_SL U62182 ( .A(n57923), .B(n57920), .Y(n57919) );
  INVx1_ASAP7_75t_SL U62183 ( .A(n67939), .Y(n57922) );
  INVx1_ASAP7_75t_SL U62184 ( .A(n67937), .Y(n57923) );
  NOR2x1_ASAP7_75t_SL U62185 ( .A(n67794), .B(n67795), .Y(n67937) );
  OAI22xp5_ASAP7_75t_SL U62186 ( .A1(n57926), .A2(n67340), .B1(n58711), .B2(
        n57925), .Y(n67894) );
  INVx1_ASAP7_75t_SL U62187 ( .A(n67344), .Y(n57925) );
  INVx1_ASAP7_75t_SL U62188 ( .A(n56862), .Y(n57927) );
  OAI21xp5_ASAP7_75t_SL U62189 ( .A1(n56862), .A2(n67340), .B(n58711), .Y(
        n67531) );
  XNOR2xp5_ASAP7_75t_SL U62190 ( .A(n58701), .B(n59518), .Y(n67454) );
  XNOR2xp5_ASAP7_75t_SL U62191 ( .A(n68130), .B(n68129), .Y(n57928) );
  AOI22xp5_ASAP7_75t_SL U62192 ( .A1(n56972), .A2(n58916), .B1(n58913), .B2(
        n58914), .Y(n68129) );
  INVx1_ASAP7_75t_SL U62193 ( .A(n68208), .Y(n68209) );
  OAI22xp5_ASAP7_75t_SL U62194 ( .A1(n67415), .A2(n67414), .B1(n67413), .B2(
        n59042), .Y(n67488) );
  INVx1_ASAP7_75t_SL U62195 ( .A(n67836), .Y(n57930) );
  XNOR2xp5_ASAP7_75t_SL U62196 ( .A(n57931), .B(n68513), .Y(n58997) );
  XOR2xp5_ASAP7_75t_SL U62197 ( .A(n57932), .B(n57933), .Y(n68513) );
  INVx1_ASAP7_75t_SL U62198 ( .A(n59202), .Y(n57932) );
  XNOR2xp5_ASAP7_75t_SL U62199 ( .A(n68445), .B(n68446), .Y(n57933) );
  MAJIxp5_ASAP7_75t_SL U62200 ( .A(n59000), .B(n68393), .C(n68394), .Y(n68510)
         );
  INVx1_ASAP7_75t_SL U62201 ( .A(n66812), .Y(n57934) );
  AOI22xp5_ASAP7_75t_SL U62202 ( .A1(n75048), .A2(n66748), .B1(n66749), .B2(
        n59100), .Y(n66812) );
  INVx1_ASAP7_75t_SL U62203 ( .A(n63133), .Y(n63134) );
  NOR2x1_ASAP7_75t_SL U62204 ( .A(n57021), .B(n57935), .Y(n63133) );
  INVx1_ASAP7_75t_SL U62205 ( .A(n62890), .Y(n62889) );
  OR2x2_ASAP7_75t_SL U62206 ( .A(n57938), .B(n62875), .Y(n62890) );
  NAND2xp5_ASAP7_75t_SL U62207 ( .A(n57111), .B(n67902), .Y(n57939) );
  O2A1O1Ixp5_ASAP7_75t_SL U62208 ( .A1(n59594), .A2(n57940), .B(n57310), .C(
        n64335), .Y(n64339) );
  NAND2x1_ASAP7_75t_SL U62209 ( .A(n58971), .B(n58032), .Y(n67668) );
  XNOR2x1_ASAP7_75t_SL U62210 ( .A(n58035), .B(n58049), .Y(n67669) );
  INVx2_ASAP7_75t_SL U62211 ( .A(n58073), .Y(n67758) );
  OAI21x1_ASAP7_75t_SL U62212 ( .A1(n57945), .A2(n53485), .B(n57944), .Y(
        n67275) );
  NAND2xp5_ASAP7_75t_SL U62213 ( .A(n57946), .B(n67350), .Y(n57944) );
  INVx1_ASAP7_75t_SL U62214 ( .A(n56990), .Y(n57946) );
  NAND2xp5_ASAP7_75t_SL U62215 ( .A(n57947), .B(n59620), .Y(n62677) );
  INVx1_ASAP7_75t_SL U62216 ( .A(n67250), .Y(n57947) );
  AND2x2_ASAP7_75t_SL U62217 ( .A(n57698), .B(n58173), .Y(n67250) );
  NOR2x1_ASAP7_75t_SL U62218 ( .A(n57064), .B(n64891), .Y(n65025) );
  NAND2xp5_ASAP7_75t_SL U62219 ( .A(n65022), .B(n58070), .Y(n57948) );
  INVx1_ASAP7_75t_SL U62220 ( .A(n67970), .Y(n57949) );
  NAND2xp5_ASAP7_75t_SL U62221 ( .A(n64571), .B(n64890), .Y(n65027) );
  AOI22xp5_ASAP7_75t_SL U62222 ( .A1(n58336), .A2(n67004), .B1(n57163), .B2(
        n66461), .Y(n67141) );
  NOR2x1_ASAP7_75t_SL U62223 ( .A(n56977), .B(n66454), .Y(n66461) );
  XNOR2xp5_ASAP7_75t_SL U62224 ( .A(n59607), .B(n75895), .Y(n67004) );
  XNOR2x1_ASAP7_75t_SL U62225 ( .A(n57952), .B(n57950), .Y(n68347) );
  XNOR2x1_ASAP7_75t_SL U62226 ( .A(n68340), .B(n57951), .Y(n65069) );
  XNOR2x1_ASAP7_75t_SL U62227 ( .A(n68341), .B(n68342), .Y(n57952) );
  NAND2xp5_ASAP7_75t_SL U62228 ( .A(n75071), .B(n75056), .Y(n75078) );
  OR2x2_ASAP7_75t_SL U62229 ( .A(n57149), .B(n75055), .Y(n75056) );
  XNOR2x1_ASAP7_75t_SL U62230 ( .A(n68187), .B(n68188), .Y(n68189) );
  NAND2x1_ASAP7_75t_SL U62231 ( .A(n68027), .B(n68025), .Y(n68188) );
  OAI21xp5_ASAP7_75t_SL U62232 ( .A1(n68000), .A2(n67999), .B(n67998), .Y(
        n68027) );
  XNOR2xp5_ASAP7_75t_SL U62233 ( .A(n67996), .B(n67995), .Y(n57955) );
  MAJIxp5_ASAP7_75t_SL U62234 ( .A(n68223), .B(n68224), .C(n68279), .Y(n68271)
         );
  MAJIxp5_ASAP7_75t_SL U62235 ( .A(n65010), .B(n65009), .C(n65011), .Y(n68224)
         );
  NOR2x1_ASAP7_75t_SL U62236 ( .A(n64961), .B(n57956), .Y(n65009) );
  NOR2x1_ASAP7_75t_SL U62237 ( .A(n67849), .B(n68383), .Y(n57956) );
  OAI21xp5_ASAP7_75t_SL U62238 ( .A1(n59456), .A2(n59668), .B(n57957), .Y(
        n66701) );
  NAND2xp5_ASAP7_75t_SL U62239 ( .A(n58536), .B(n59668), .Y(n57957) );
  INVx1_ASAP7_75t_SL U62240 ( .A(n63672), .Y(n57959) );
  BUFx6f_ASAP7_75t_SL U62241 ( .A(n58248), .Y(n57960) );
  INVx1_ASAP7_75t_SL U62242 ( .A(n58248), .Y(n64618) );
  INVx2_ASAP7_75t_SL U62243 ( .A(n75277), .Y(n57962) );
  NOR2x1p5_ASAP7_75t_SL U62244 ( .A(n75275), .B(n75274), .Y(n75277) );
  AND2x2_ASAP7_75t_SL U62245 ( .A(n67217), .B(n67218), .Y(n75278) );
  INVx1_ASAP7_75t_SL U62246 ( .A(n68694), .Y(n67219) );
  NAND2xp5_ASAP7_75t_SL U62247 ( .A(n59653), .B(n67302), .Y(n57963) );
  NAND2xp5_ASAP7_75t_SL U62248 ( .A(n57964), .B(n68617), .Y(n68639) );
  NAND2xp5_ASAP7_75t_SL U62249 ( .A(n57966), .B(n57965), .Y(n68617) );
  NAND2xp5_ASAP7_75t_SL U62250 ( .A(n57968), .B(n57967), .Y(n57966) );
  NAND2xp5_ASAP7_75t_SL U62251 ( .A(n66586), .B(n66567), .Y(n57968) );
  NAND2xp5_ASAP7_75t_SL U62252 ( .A(n57970), .B(n57486), .Y(n57969) );
  NAND2xp5_ASAP7_75t_SL U62253 ( .A(n57122), .B(n67420), .Y(n57970) );
  NAND2xp5_ASAP7_75t_SL U62254 ( .A(n62864), .B(n57971), .Y(n62909) );
  NAND2xp5_ASAP7_75t_SL U62255 ( .A(n62863), .B(n57972), .Y(n57971) );
  NAND2xp5_ASAP7_75t_SL U62256 ( .A(n62862), .B(n57973), .Y(n62864) );
  XNOR2xp5_ASAP7_75t_SL U62257 ( .A(n62788), .B(n62787), .Y(n57973) );
  NAND2xp5_ASAP7_75t_SL U62258 ( .A(n53490), .B(n57974), .Y(n58954) );
  INVx1_ASAP7_75t_SL U62259 ( .A(n57371), .Y(n57974) );
  NAND2xp5_ASAP7_75t_SL U62260 ( .A(n57979), .B(n57975), .Y(n68159) );
  NAND2xp5_ASAP7_75t_SL U62261 ( .A(n57371), .B(n68148), .Y(n57975) );
  OAI22xp5_ASAP7_75t_SL U62262 ( .A1(n67976), .A2(n57977), .B1(n68148), .B2(
        n57976), .Y(n57978) );
  INVx1_ASAP7_75t_SL U62263 ( .A(n57979), .Y(n57976) );
  MAJIxp5_ASAP7_75t_SL U62264 ( .A(n57978), .B(n68160), .C(n68161), .Y(n68232)
         );
  XNOR2x1_ASAP7_75t_SL U62265 ( .A(n57980), .B(n53274), .Y(n68161) );
  MAJx2_ASAP7_75t_SL U62266 ( .A(n68216), .B(n58170), .C(n68217), .Y(n67976)
         );
  NAND2xp5_ASAP7_75t_SL U62267 ( .A(n75092), .B(n57981), .Y(n75093) );
  NAND2xp5_ASAP7_75t_SL U62268 ( .A(n75286), .B(n57983), .Y(n75288) );
  INVx1_ASAP7_75t_SL U62269 ( .A(n58691), .Y(n57984) );
  OAI21xp5_ASAP7_75t_SL U62270 ( .A1(n58495), .A2(n59216), .B(n59215), .Y(
        n57986) );
  INVx1_ASAP7_75t_SL U62271 ( .A(n68444), .Y(n68488) );
  XOR2xp5_ASAP7_75t_SL U62272 ( .A(n57988), .B(n57987), .Y(n68444) );
  INVx1_ASAP7_75t_SL U62273 ( .A(n68441), .Y(n57988) );
  XNOR2xp5_ASAP7_75t_SL U62274 ( .A(n68387), .B(n68388), .Y(n59029) );
  NOR2x1_ASAP7_75t_SL U62275 ( .A(n62910), .B(n62909), .Y(n63292) );
  XNOR2xp5_ASAP7_75t_SL U62276 ( .A(n62867), .B(n57989), .Y(n62910) );
  XNOR2xp5_ASAP7_75t_SL U62277 ( .A(n62866), .B(n62865), .Y(n57989) );
  OAI21xp5_ASAP7_75t_SL U62278 ( .A1(n57990), .A2(n62865), .B(n62855), .Y(
        n62867) );
  NOR2x1_ASAP7_75t_SL U62279 ( .A(n62870), .B(n62849), .Y(n62865) );
  NOR2x1_ASAP7_75t_SL U62280 ( .A(n57991), .B(n67474), .Y(n67700) );
  O2A1O1Ixp5_ASAP7_75t_SL U62281 ( .A1(n57991), .A2(n66786), .B(n66785), .C(
        n66784), .Y(n68464) );
  NOR2x1_ASAP7_75t_SL U62282 ( .A(n59603), .B(n75947), .Y(n57991) );
  XOR2xp5_ASAP7_75t_SL U62283 ( .A(n66848), .B(n66847), .Y(n66832) );
  OAI21xp5_ASAP7_75t_SL U62284 ( .A1(n59491), .A2(n66831), .B(n57992), .Y(
        n66847) );
  NAND2xp5_ASAP7_75t_SL U62285 ( .A(n57463), .B(n57993), .Y(n57992) );
  NAND2xp5_ASAP7_75t_SL U62286 ( .A(n67393), .B(n58627), .Y(n58429) );
  NAND2xp5_ASAP7_75t_SL U62287 ( .A(n67578), .B(n67579), .Y(n67393) );
  NAND2xp5_ASAP7_75t_SL U62288 ( .A(n57067), .B(n66666), .Y(n58798) );
  AOI22xp5_ASAP7_75t_SL U62289 ( .A1(n57067), .A2(n66954), .B1(n66923), .B2(
        n66922), .Y(n68360) );
  NAND2xp5_ASAP7_75t_SL U62290 ( .A(n58342), .B(n57995), .Y(n57994) );
  NOR2x1_ASAP7_75t_SL U62291 ( .A(n59535), .B(n63184), .Y(n63661) );
  AND2x2_ASAP7_75t_SL U62292 ( .A(n57996), .B(n58342), .Y(n63184) );
  NOR2xp33_ASAP7_75t_SL U62293 ( .A(n57201), .B(n63173), .Y(n57996) );
  AND2x2_ASAP7_75t_SL U62294 ( .A(n59539), .B(n62748), .Y(n63859) );
  MAJIxp5_ASAP7_75t_SL U62295 ( .A(n67633), .B(n67811), .C(n58453), .Y(n67801)
         );
  NAND2xp5_ASAP7_75t_SL U62296 ( .A(n57999), .B(n58649), .Y(n63673) );
  NAND2xp5_ASAP7_75t_SL U62297 ( .A(n59551), .B(n58650), .Y(n58000) );
  NAND2xp5_ASAP7_75t_SL U62298 ( .A(n75031), .B(n75032), .Y(n58001) );
  OR2x2_ASAP7_75t_SL U62299 ( .A(n57365), .B(n59518), .Y(n75031) );
  O2A1O1Ixp5_ASAP7_75t_SL U62300 ( .A1(n53221), .A2(n58658), .B(n58005), .C(
        n67152), .Y(n67138) );
  NOR2xp33_ASAP7_75t_SL U62301 ( .A(n53310), .B(n59314), .Y(n58003) );
  NAND2xp5_ASAP7_75t_SL U62302 ( .A(n59596), .B(n75947), .Y(n67062) );
  NAND3xp33_ASAP7_75t_SL U62303 ( .A(n68805), .B(n59489), .C(n58006), .Y(
        n58727) );
  NAND2xp5_ASAP7_75t_SL U62304 ( .A(n53622), .B(n59294), .Y(n58006) );
  INVx1_ASAP7_75t_SL U62305 ( .A(n67272), .Y(n67509) );
  NAND2xp5_ASAP7_75t_SL U62306 ( .A(n58009), .B(n58007), .Y(n67272) );
  NAND2xp5_ASAP7_75t_SL U62307 ( .A(n57358), .B(n58008), .Y(n58007) );
  XNOR2xp5_ASAP7_75t_SL U62308 ( .A(n59603), .B(n57104), .Y(n67404) );
  NAND2xp5_ASAP7_75t_SL U62309 ( .A(n67363), .B(n57273), .Y(n58009) );
  OAI21xp5_ASAP7_75t_SL U62310 ( .A1(n67569), .A2(n57112), .B(n58010), .Y(
        n63210) );
  NAND2xp5_ASAP7_75t_SL U62311 ( .A(n67846), .B(n57112), .Y(n58010) );
  OAI21xp5_ASAP7_75t_SL U62312 ( .A1(n75644), .A2(n57484), .B(n58012), .Y(
        n67282) );
  NAND2xp5_ASAP7_75t_SL U62313 ( .A(n67444), .B(n75644), .Y(n58012) );
  AOI21xp5_ASAP7_75t_SL U62314 ( .A1(n63672), .A2(n53624), .B(n58013), .Y(
        n66418) );
  NAND2xp5_ASAP7_75t_SL U62315 ( .A(n64368), .B(n58014), .Y(n58013) );
  NAND2xp5_ASAP7_75t_SL U62316 ( .A(n59668), .B(n59600), .Y(n66285) );
  XNOR2xp5_ASAP7_75t_SL U62317 ( .A(n59670), .B(n57314), .Y(n66535) );
  INVx1_ASAP7_75t_SL U62318 ( .A(n75962), .Y(n58016) );
  INVx2_ASAP7_75t_SL U62319 ( .A(n67914), .Y(n59055) );
  OAI21xp5_ASAP7_75t_SL U62320 ( .A1(n59596), .A2(n58892), .B(n58696), .Y(
        n58017) );
  MAJIxp5_ASAP7_75t_SL U62321 ( .A(n66893), .B(n66891), .C(n66892), .Y(n66990)
         );
  XNOR2xp5_ASAP7_75t_SL U62322 ( .A(n58018), .B(n66680), .Y(n66893) );
  INVx1_ASAP7_75t_SL U62323 ( .A(n66873), .Y(n58018) );
  AOI22xp5_ASAP7_75t_SL U62324 ( .A1(n67077), .A2(n67306), .B1(n66677), .B2(
        n57161), .Y(n66873) );
  MAJIxp5_ASAP7_75t_SL U62325 ( .A(n64993), .B(n64992), .C(n64994), .Y(n68339)
         );
  XOR2xp5_ASAP7_75t_SL U62326 ( .A(n65067), .B(n65068), .Y(n58019) );
  XOR2xp5_ASAP7_75t_SL U62327 ( .A(n68256), .B(n68257), .Y(n65067) );
  INVx1_ASAP7_75t_SL U62328 ( .A(n67074), .Y(n66863) );
  OR2x2_ASAP7_75t_SL U62329 ( .A(n58020), .B(n53271), .Y(n67074) );
  NAND2xp5_ASAP7_75t_SL U62330 ( .A(n58021), .B(n58384), .Y(n58020) );
  XNOR2x2_ASAP7_75t_SL U62331 ( .A(n58832), .B(n58022), .Y(n68241) );
  XNOR2x1_ASAP7_75t_SL U62332 ( .A(n68241), .B(n58023), .Y(n68803) );
  XNOR2x1_ASAP7_75t_SL U62333 ( .A(n68242), .B(n58024), .Y(n58023) );
  NAND2x1_ASAP7_75t_SL U62334 ( .A(n68230), .B(n68229), .Y(n58024) );
  XNOR2x2_ASAP7_75t_SL U62335 ( .A(n68237), .B(n68236), .Y(n68242) );
  BUFx6f_ASAP7_75t_SL U62336 ( .A(n59452), .Y(n58025) );
  AOI22x1_ASAP7_75t_SL U62337 ( .A1(n58025), .A2(n68084), .B1(n59171), .B2(
        n68085), .Y(n68156) );
  NOR2x1p5_ASAP7_75t_SL U62338 ( .A(n67973), .B(n58026), .Y(n68085) );
  NAND2x1p5_ASAP7_75t_SL U62339 ( .A(n62647), .B(n66719), .Y(n59452) );
  OAI21xp5_ASAP7_75t_SL U62340 ( .A1(n64604), .A2(n58027), .B(n64603), .Y(
        n64996) );
  NOR2x1_ASAP7_75t_SL U62341 ( .A(n64600), .B(n64599), .Y(n64597) );
  NAND3xp33_ASAP7_75t_SL U62342 ( .A(n58030), .B(n64596), .C(n64595), .Y(
        n58029) );
  NAND2xp5_ASAP7_75t_SL U62343 ( .A(n64540), .B(n64541), .Y(n64595) );
  OAI21xp5_ASAP7_75t_SL U62344 ( .A1(n64540), .A2(n64541), .B(n64539), .Y(
        n64596) );
  NAND2xp5_ASAP7_75t_SL U62345 ( .A(n64600), .B(n64599), .Y(n58030) );
  INVx1_ASAP7_75t_SL U62346 ( .A(n68286), .Y(n58031) );
  XNOR2xp5_ASAP7_75t_SL U62347 ( .A(n68174), .B(n68173), .Y(n68284) );
  OAI211xp5_ASAP7_75t_SL U62348 ( .A1(n67485), .A2(n67486), .B(n58034), .C(
        n58033), .Y(n58032) );
  NAND2xp5_ASAP7_75t_SL U62349 ( .A(n67273), .B(n67275), .Y(n58033) );
  OAI21xp5_ASAP7_75t_SL U62350 ( .A1(n67275), .A2(n67273), .B(n67274), .Y(
        n58034) );
  XNOR2x1_ASAP7_75t_SL U62351 ( .A(n58036), .B(n67732), .Y(n58035) );
  NAND2xp5_ASAP7_75t_SL U62352 ( .A(n67275), .B(n67274), .Y(n67483) );
  OAI21xp5_ASAP7_75t_SL U62353 ( .A1(n67275), .A2(n67274), .B(n67273), .Y(
        n67484) );
  INVx1_ASAP7_75t_SL U62354 ( .A(n57331), .Y(n76237) );
  INVx1_ASAP7_75t_SL U62355 ( .A(n58037), .Y(n76678) );
  NAND2xp5_ASAP7_75t_SL U62356 ( .A(n1770), .B(n1686), .Y(n58037) );
  NAND2xp5_ASAP7_75t_SL U62357 ( .A(n1571), .B(n1588), .Y(n59258) );
  XNOR2xp5_ASAP7_75t_SL U62358 ( .A(n58038), .B(n64069), .Y(n63847) );
  INVx1_ASAP7_75t_SL U62359 ( .A(n64067), .Y(n58038) );
  XNOR2xp5_ASAP7_75t_SL U62360 ( .A(n58039), .B(n63821), .Y(n64067) );
  INVx1_ASAP7_75t_SL U62361 ( .A(n64044), .Y(n58039) );
  AOI22xp5_ASAP7_75t_SL U62362 ( .A1(n62801), .A2(n57007), .B1(n67251), .B2(
        n62813), .Y(n62823) );
  NAND2xp5_ASAP7_75t_SL U62363 ( .A(n58040), .B(n62800), .Y(n62813) );
  INVx1_ASAP7_75t_SL U62364 ( .A(n68486), .Y(n66809) );
  MAJIxp5_ASAP7_75t_SL U62365 ( .A(n68466), .B(n58042), .C(n57058), .Y(n68486)
         );
  INVx1_ASAP7_75t_SL U62366 ( .A(n68465), .Y(n58042) );
  AOI22xp5_ASAP7_75t_SL U62367 ( .A1(n66795), .A2(n57380), .B1(n66793), .B2(
        n66794), .Y(n68465) );
  NAND2x2_ASAP7_75t_SL U62368 ( .A(n64394), .B(n64395), .Y(n67964) );
  NAND2x1_ASAP7_75t_SL U62369 ( .A(n58043), .B(n63191), .Y(n64395) );
  NOR2x1p5_ASAP7_75t_SL U62370 ( .A(n58045), .B(n58044), .Y(n64394) );
  INVx2_ASAP7_75t_SL U62371 ( .A(n60747), .Y(n58047) );
  INVx1_ASAP7_75t_SL U62372 ( .A(n68371), .Y(n58049) );
  OR2x2_ASAP7_75t_SL U62373 ( .A(n64088), .B(n64087), .Y(n64667) );
  INVx1_ASAP7_75t_SL U62374 ( .A(n64419), .Y(n64532) );
  OR2x2_ASAP7_75t_SL U62375 ( .A(n64418), .B(n64417), .Y(n64419) );
  NAND2xp5_ASAP7_75t_SL U62376 ( .A(n67810), .B(n58052), .Y(n58051) );
  OAI21xp5_ASAP7_75t_SL U62377 ( .A1(n67257), .A2(n57038), .B(n67256), .Y(
        n67407) );
  OAI21xp5_ASAP7_75t_SL U62378 ( .A1(n59460), .A2(n67361), .B(n58053), .Y(
        n67617) );
  NAND3xp33_ASAP7_75t_SL U62379 ( .A(n67912), .B(n59048), .C(n58054), .Y(
        n58053) );
  XNOR2xp5_ASAP7_75t_SL U62380 ( .A(n63797), .B(n63799), .Y(n63681) );
  XNOR2xp5_ASAP7_75t_SL U62381 ( .A(n63665), .B(n58055), .Y(n63799) );
  XNOR2xp5_ASAP7_75t_SL U62382 ( .A(n63804), .B(n63803), .Y(n58055) );
  AND2x2_ASAP7_75t_SL U62383 ( .A(n61932), .B(n59371), .Y(n58797) );
  AND2x2_ASAP7_75t_SL U62384 ( .A(n57213), .B(n63063), .Y(n62757) );
  INVx1_ASAP7_75t_SL U62385 ( .A(n63063), .Y(n67311) );
  NAND2x1_ASAP7_75t_SL U62386 ( .A(n59019), .B(n61923), .Y(n63063) );
  XNOR2xp5_ASAP7_75t_SL U62387 ( .A(n57078), .B(n59620), .Y(n67559) );
  NOR2x1_ASAP7_75t_SL U62388 ( .A(n59348), .B(n59349), .Y(n59485) );
  INVx1_ASAP7_75t_SL U62389 ( .A(n67326), .Y(n58058) );
  NAND2xp5_ASAP7_75t_SL U62390 ( .A(n58060), .B(n68001), .Y(n67919) );
  OAI21xp5_ASAP7_75t_SL U62391 ( .A1(n58490), .A2(n67913), .B(n67912), .Y(
        n58060) );
  NAND2xp5_ASAP7_75t_SL U62392 ( .A(n67536), .B(n58061), .Y(n62868) );
  XOR2xp5_ASAP7_75t_SL U62393 ( .A(n62908), .B(n62907), .Y(n62884) );
  NOR2x1_ASAP7_75t_SL U62394 ( .A(n58062), .B(n57162), .Y(n62908) );
  NAND2xp5_ASAP7_75t_SL U62395 ( .A(n59657), .B(n67230), .Y(n58062) );
  NAND2xp5_ASAP7_75t_SL U62396 ( .A(n66819), .B(n58063), .Y(n66901) );
  NAND3xp33_ASAP7_75t_SL U62397 ( .A(n66818), .B(n66821), .C(n58064), .Y(
        n58063) );
  OR2x2_ASAP7_75t_SL U62398 ( .A(n66821), .B(n66822), .Y(n66902) );
  INVx1_ASAP7_75t_SL U62399 ( .A(n68589), .Y(n68588) );
  XNOR2xp5_ASAP7_75t_SL U62400 ( .A(n69035), .B(n58065), .Y(n68589) );
  XNOR2xp5_ASAP7_75t_SL U62401 ( .A(n58066), .B(n69036), .Y(n58065) );
  AOI21xp5_ASAP7_75t_SL U62402 ( .A1(n59015), .A2(n68551), .B(n59014), .Y(
        n58066) );
  INVx1_ASAP7_75t_SL U62403 ( .A(n58878), .Y(n58067) );
  NOR2x1_ASAP7_75t_SL U62404 ( .A(n62710), .B(n62711), .Y(n58878) );
  AOI22xp5_ASAP7_75t_SL U62405 ( .A1(n62692), .A2(n59171), .B1(n62956), .B2(
        n57157), .Y(n62710) );
  INVx1_ASAP7_75t_SL U62406 ( .A(n68147), .Y(n58171) );
  INVx1_ASAP7_75t_SL U62407 ( .A(n67855), .Y(n58069) );
  OA21x2_ASAP7_75t_SL U62408 ( .A1(n56841), .A2(n59328), .B(n59327), .Y(n58070) );
  AOI22xp33_ASAP7_75t_SL U62409 ( .A1(n57161), .A2(n67076), .B1(n67306), .B2(
        n66467), .Y(n67142) );
  NAND4xp75_ASAP7_75t_SL U62410 ( .A(n57457), .B(n57353), .C(n53492), .D(
        n59107), .Y(n58071) );
  INVx3_ASAP7_75t_SL U62411 ( .A(n59474), .Y(n64353) );
  INVx1_ASAP7_75t_SL U62412 ( .A(n59220), .Y(n67989) );
  OR2x2_ASAP7_75t_SL U62413 ( .A(n67983), .B(n58072), .Y(n59220) );
  MAJIxp5_ASAP7_75t_SL U62414 ( .A(n58488), .B(n59490), .C(n67979), .Y(n67980)
         );
  NAND2xp5_ASAP7_75t_SL U62415 ( .A(n58073), .B(n58074), .Y(n58077) );
  NOR2x1p5_ASAP7_75t_SL U62416 ( .A(n58427), .B(n67765), .Y(n58076) );
  NAND2x1_ASAP7_75t_SL U62417 ( .A(n67758), .B(n59334), .Y(n58078) );
  XNOR2xp5_ASAP7_75t_SL U62418 ( .A(n56990), .B(n67350), .Y(n58921) );
  AOI22xp5_ASAP7_75t_SL U62419 ( .A1(n75048), .A2(n67016), .B1(n58079), .B2(
        n59635), .Y(n67079) );
  INVx1_ASAP7_75t_SL U62420 ( .A(n66696), .Y(n58079) );
  INVx1_ASAP7_75t_SL U62421 ( .A(n75644), .Y(n58080) );
  NOR3xp33_ASAP7_75t_SL U62422 ( .A(n61188), .B(n61189), .C(n58082), .Y(n61195) );
  A2O1A1Ixp33_ASAP7_75t_SL U62423 ( .A1(n77097), .A2(n58084), .B(n75736), .C(
        n78004), .Y(n61653) );
  XNOR2xp5_ASAP7_75t_SL U62424 ( .A(n58084), .B(n60767), .Y(n61619) );
  INVx1_ASAP7_75t_SL U62425 ( .A(n59545), .Y(n58084) );
  NAND2xp5_ASAP7_75t_SL U62426 ( .A(n58087), .B(n58086), .Y(n58085) );
  INVx1_ASAP7_75t_SL U62427 ( .A(n58088), .Y(n68907) );
  INVx1_ASAP7_75t_SL U62428 ( .A(n68907), .Y(n68960) );
  INVx1_ASAP7_75t_SL U62429 ( .A(n74565), .Y(n68692) );
  OR2x2_ASAP7_75t_SL U62430 ( .A(n67216), .B(n67215), .Y(n74565) );
  OAI21xp5_ASAP7_75t_SL U62431 ( .A1(n67182), .A2(n67181), .B(n67180), .Y(
        n67215) );
  MAJIxp5_ASAP7_75t_SL U62432 ( .A(n67205), .B(n67206), .C(n67208), .Y(n67216)
         );
  INVx1_ASAP7_75t_SL U62433 ( .A(n67164), .Y(n58089) );
  NAND2xp5_ASAP7_75t_SL U62434 ( .A(n68868), .B(n58090), .Y(n68870) );
  NAND2xp5_ASAP7_75t_SL U62435 ( .A(n57129), .B(n68867), .Y(n58090) );
  NAND2xp5_ASAP7_75t_SL U62436 ( .A(n57061), .B(n58091), .Y(n68867) );
  NAND3xp33_ASAP7_75t_SL U62437 ( .A(n59345), .B(n59341), .C(n68809), .Y(
        n58091) );
  XOR2xp5_ASAP7_75t_SL U62438 ( .A(n56860), .B(n58092), .Y(n52008) );
  OAI21xp5_ASAP7_75t_SL U62439 ( .A1(n74567), .A2(n58881), .B(n74566), .Y(
        n58092) );
  INVx1_ASAP7_75t_SL U62440 ( .A(n68093), .Y(n58093) );
  INVx1_ASAP7_75t_SL U62441 ( .A(n58094), .Y(n67214) );
  NAND2xp5_ASAP7_75t_SL U62442 ( .A(n58095), .B(n67180), .Y(n58094) );
  INVx1_ASAP7_75t_SL U62443 ( .A(n67162), .Y(n58095) );
  XNOR2xp5_ASAP7_75t_SL U62444 ( .A(n58097), .B(n58096), .Y(n67108) );
  XOR2xp5_ASAP7_75t_SL U62445 ( .A(n67184), .B(n67185), .Y(n58096) );
  XNOR2xp5_ASAP7_75t_SL U62446 ( .A(n58752), .B(n58751), .Y(n67184) );
  INVx1_ASAP7_75t_SL U62447 ( .A(n67186), .Y(n58752) );
  INVx1_ASAP7_75t_SL U62448 ( .A(n67183), .Y(n58097) );
  MAJIxp5_ASAP7_75t_SL U62449 ( .A(n67102), .B(n67101), .C(n58098), .Y(n67183)
         );
  INVx1_ASAP7_75t_SL U62450 ( .A(n67100), .Y(n58098) );
  INVxp33_ASAP7_75t_SL U62451 ( .A(n64088), .Y(n64086) );
  INVx1_ASAP7_75t_SL U62452 ( .A(n64087), .Y(n64085) );
  O2A1O1Ixp5_ASAP7_75t_SL U62453 ( .A1(n58102), .A2(n58101), .B(n57141), .C(
        n58099), .Y(n64669) );
  XNOR2xp5_ASAP7_75t_SL U62454 ( .A(n64075), .B(n58100), .Y(n64090) );
  INVx1_ASAP7_75t_SL U62455 ( .A(n64089), .Y(n58101) );
  INVx1_ASAP7_75t_SL U62456 ( .A(n64667), .Y(n58102) );
  INVx1_ASAP7_75t_SL U62457 ( .A(n67951), .Y(n68380) );
  NAND2xp5_ASAP7_75t_SL U62458 ( .A(n57173), .B(n67951), .Y(n58104) );
  INVx1_ASAP7_75t_SL U62459 ( .A(n62721), .Y(n62723) );
  OR2x2_ASAP7_75t_SL U62460 ( .A(n58106), .B(n62760), .Y(n62721) );
  NAND2xp5_ASAP7_75t_SL U62461 ( .A(n59538), .B(n64504), .Y(n58106) );
  NAND2xp5_ASAP7_75t_SL U62462 ( .A(n58108), .B(n58107), .Y(n58783) );
  INVx1_ASAP7_75t_SL U62463 ( .A(n68371), .Y(n58107) );
  NAND4xp25_ASAP7_75t_SL U62464 ( .A(n67728), .B(n58351), .C(n67729), .D(
        n58109), .Y(n58108) );
  NAND2xp5_ASAP7_75t_SL U62465 ( .A(n67731), .B(n67730), .Y(n58109) );
  INVx1_ASAP7_75t_SL U62466 ( .A(n63103), .Y(n63101) );
  XOR2xp5_ASAP7_75t_SL U62467 ( .A(n58110), .B(n58888), .Y(n63106) );
  INVx1_ASAP7_75t_SL U62468 ( .A(n63139), .Y(n58110) );
  XOR2xp5_ASAP7_75t_SL U62469 ( .A(n58112), .B(n63108), .Y(n58111) );
  INVx1_ASAP7_75t_SL U62470 ( .A(n58502), .Y(n58112) );
  NAND2xp5_ASAP7_75t_SL U62471 ( .A(n58114), .B(n58674), .Y(n58113) );
  INVx1_ASAP7_75t_SL U62472 ( .A(n59399), .Y(n58114) );
  XNOR2xp5_ASAP7_75t_SL U62473 ( .A(n68471), .B(n68391), .Y(n67754) );
  NOR2x1_ASAP7_75t_SL U62474 ( .A(n57039), .B(n58115), .Y(n68471) );
  O2A1O1Ixp5_ASAP7_75t_SL U62475 ( .A1(n59670), .A2(n58668), .B(n58667), .C(
        n58116), .Y(n58115) );
  INVx1_ASAP7_75t_SL U62476 ( .A(n57108), .Y(n58668) );
  XNOR2x1_ASAP7_75t_SL U62477 ( .A(n67758), .B(n59334), .Y(n67495) );
  NAND2x1_ASAP7_75t_SL U62478 ( .A(n58118), .B(n58117), .Y(n59334) );
  NAND2xp5_ASAP7_75t_SL U62479 ( .A(n59656), .B(n67855), .Y(n67856) );
  XNOR2x1_ASAP7_75t_SL U62480 ( .A(n67976), .B(n58119), .Y(n58120) );
  INVx2_ASAP7_75t_SL U62481 ( .A(n58171), .Y(n58119) );
  INVx1_ASAP7_75t_SL U62482 ( .A(n68148), .Y(n58121) );
  OAI22xp5_ASAP7_75t_SL U62483 ( .A1(n63857), .A2(n63858), .B1(n64408), .B2(
        n57362), .Y(n64055) );
  NAND2xp5_ASAP7_75t_SL U62484 ( .A(n57900), .B(n58481), .Y(n63857) );
  OR2x2_ASAP7_75t_SL U62485 ( .A(n59435), .B(n68098), .Y(n58481) );
  INVx1_ASAP7_75t_SL U62486 ( .A(n63826), .Y(n63171) );
  INVx1_ASAP7_75t_SL U62487 ( .A(n63185), .Y(n58122) );
  INVx1_ASAP7_75t_SL U62488 ( .A(n66911), .Y(n66733) );
  MAJx2_ASAP7_75t_SL U62489 ( .A(n58125), .B(n66949), .C(n66952), .Y(n66911)
         );
  NOR2x1_ASAP7_75t_SL U62490 ( .A(n58123), .B(n66723), .Y(n66952) );
  INVx1_ASAP7_75t_SL U62491 ( .A(n58124), .Y(n58123) );
  AOI22xp5_ASAP7_75t_SL U62492 ( .A1(n66755), .A2(n59447), .B1(n67744), .B2(
        n67446), .Y(n66949) );
  O2A1O1Ixp5_ASAP7_75t_SL U62493 ( .A1(n64340), .A2(n64339), .B(n58127), .C(
        n58126), .Y(n59410) );
  OAI21xp5_ASAP7_75t_SL U62494 ( .A1(n64338), .A2(n64340), .B(n64337), .Y(
        n58126) );
  INVx1_ASAP7_75t_SL U62495 ( .A(n64338), .Y(n64336) );
  NOR2x1_ASAP7_75t_SL U62496 ( .A(n58128), .B(n64082), .Y(n64338) );
  INVx1_ASAP7_75t_SL U62497 ( .A(n58129), .Y(n58128) );
  NAND2xp5_ASAP7_75t_SL U62498 ( .A(n76078), .B(n64083), .Y(n58129) );
  AOI21xp5_ASAP7_75t_SL U62499 ( .A1(n58536), .A2(n67227), .B(n62724), .Y(
        n63122) );
  INVx1_ASAP7_75t_SL U62500 ( .A(n63816), .Y(n64350) );
  MAJIxp5_ASAP7_75t_SL U62501 ( .A(n68508), .B(n58132), .C(n66942), .Y(n68525)
         );
  INVx1_ASAP7_75t_SL U62502 ( .A(n68506), .Y(n58132) );
  XNOR2xp5_ASAP7_75t_SL U62503 ( .A(n66938), .B(n66937), .Y(n58133) );
  MAJIxp5_ASAP7_75t_SL U62504 ( .A(n68441), .B(n68443), .C(n57220), .Y(n68508)
         );
  NOR2x1_ASAP7_75t_SL U62505 ( .A(n66927), .B(n68365), .Y(n68441) );
  NOR2x1_ASAP7_75t_SL U62506 ( .A(n66926), .B(n68360), .Y(n68365) );
  NAND2xp5_ASAP7_75t_SL U62507 ( .A(n58135), .B(n67252), .Y(n67368) );
  NAND2xp33_ASAP7_75t_SL U62508 ( .A(n59596), .B(n75908), .Y(n58135) );
  INVx1_ASAP7_75t_SL U62509 ( .A(n67732), .Y(n67733) );
  NAND2xp5_ASAP7_75t_SL U62510 ( .A(n67465), .B(n59613), .Y(n58138) );
  NAND2xp5_ASAP7_75t_SL U62511 ( .A(n58139), .B(n66325), .Y(n66328) );
  INVx1_ASAP7_75t_SL U62512 ( .A(n58140), .Y(n58139) );
  NOR2x1_ASAP7_75t_SL U62513 ( .A(n58962), .B(n66356), .Y(n58140) );
  NOR2x1_ASAP7_75t_SL U62514 ( .A(n58863), .B(n59446), .Y(n66356) );
  INVx1_ASAP7_75t_SL U62515 ( .A(n68011), .Y(n64083) );
  XNOR2xp5_ASAP7_75t_SL U62516 ( .A(n57003), .B(n66932), .Y(n68358) );
  OAI21xp5_ASAP7_75t_SL U62517 ( .A1(n67465), .A2(n57099), .B(n58142), .Y(
        n66932) );
  NAND2xp5_ASAP7_75t_SL U62518 ( .A(n66928), .B(n67306), .Y(n58142) );
  OAI21xp5_ASAP7_75t_SL U62519 ( .A1(n64566), .A2(n64565), .B(n64564), .Y(
        n64877) );
  NAND2xp5_ASAP7_75t_SL U62520 ( .A(n64566), .B(n64565), .Y(n64876) );
  OAI21xp5_ASAP7_75t_SL U62521 ( .A1(n64489), .A2(n64643), .B(n64488), .Y(
        n64565) );
  INVx1_ASAP7_75t_SL U62522 ( .A(n62877), .Y(n68094) );
  NOR2x1_ASAP7_75t_SL U62523 ( .A(n58144), .B(n67519), .Y(n67523) );
  INVx1_ASAP7_75t_SL U62524 ( .A(n58145), .Y(n58144) );
  NAND3xp33_ASAP7_75t_SL U62525 ( .A(n67641), .B(n75032), .C(n67517), .Y(
        n58145) );
  INVx1_ASAP7_75t_SL U62526 ( .A(or1200_cpu_or1200_except_n681), .Y(n58146) );
  INVx1_ASAP7_75t_SL U62527 ( .A(n66944), .Y(n66945) );
  XNOR2xp5_ASAP7_75t_SL U62528 ( .A(n66736), .B(n58147), .Y(n66944) );
  XNOR2xp5_ASAP7_75t_SL U62529 ( .A(n59237), .B(n66735), .Y(n58147) );
  AOI22xp5_ASAP7_75t_SL U62530 ( .A1(n67306), .A2(n66611), .B1(n66751), .B2(
        n57161), .Y(n66735) );
  OAI22xp5_ASAP7_75t_SL U62531 ( .A1(n66756), .A2(n59440), .B1(n66857), .B2(
        n59042), .Y(n59237) );
  AOI21xp5_ASAP7_75t_SL U62532 ( .A1(n57311), .A2(n58148), .B(n68377), .Y(
        n68378) );
  INVx1_ASAP7_75t_SL U62533 ( .A(n67739), .Y(n58148) );
  AOI21xp5_ASAP7_75t_SL U62534 ( .A1(n68400), .A2(n68401), .B(n58152), .Y(
        n58150) );
  INVx1_ASAP7_75t_SL U62535 ( .A(n68399), .Y(n58151) );
  INVx1_ASAP7_75t_SL U62536 ( .A(n68398), .Y(n58152) );
  NAND2xp33_ASAP7_75t_SL U62537 ( .A(n59637), .B(n75900), .Y(n58154) );
  AOI22xp33_ASAP7_75t_SL U62538 ( .A1(n57067), .A2(n66850), .B1(n66851), .B2(
        n59100), .Y(n67007) );
  NAND2xp5_ASAP7_75t_SL U62539 ( .A(n58156), .B(n67358), .Y(n59074) );
  O2A1O1Ixp5_ASAP7_75t_SL U62540 ( .A1(n77730), .A2(n57109), .B(n57428), .C(
        n58158), .Y(n58157) );
  NOR2x1_ASAP7_75t_SL U62541 ( .A(n57428), .B(n57109), .Y(n58158) );
  INVx1_ASAP7_75t_SL U62542 ( .A(n68456), .Y(n68497) );
  NOR2x1_ASAP7_75t_SL U62543 ( .A(n59289), .B(n59287), .Y(n58160) );
  NOR2x1_ASAP7_75t_SL U62544 ( .A(n59288), .B(n75076), .Y(n59287) );
  INVx1_ASAP7_75t_SL U62545 ( .A(n68450), .Y(n58161) );
  NAND2xp5_ASAP7_75t_SL U62546 ( .A(n64675), .B(n57877), .Y(n63805) );
  INVx1_ASAP7_75t_SL U62547 ( .A(n67883), .Y(n58162) );
  NOR3xp33_ASAP7_75t_SL U62548 ( .A(n64492), .B(n64491), .C(n58163), .Y(n64493) );
  INVx1_ASAP7_75t_SL U62549 ( .A(n67056), .Y(n67057) );
  NAND2xp5_ASAP7_75t_SL U62550 ( .A(n58164), .B(n66995), .Y(n67056) );
  OAI21xp5_ASAP7_75t_SL U62551 ( .A1(n66993), .A2(n58165), .B(n56839), .Y(
        n58164) );
  INVx1_ASAP7_75t_SL U62552 ( .A(n59664), .Y(n58165) );
  NOR2x1_ASAP7_75t_SL U62553 ( .A(n59598), .B(n57253), .Y(n66993) );
  INVx1_ASAP7_75t_SL U62554 ( .A(n68687), .Y(n74112) );
  NOR2x1p5_ASAP7_75t_SL U62555 ( .A(n57214), .B(n61909), .Y(n58166) );
  NAND3x2_ASAP7_75t_SL U62556 ( .A(n59442), .B(n59567), .C(n59544), .Y(n61909)
         );
  NAND3x2_ASAP7_75t_SL U62557 ( .A(n58166), .B(n57199), .C(n58168), .Y(n62629)
         );
  INVx1_ASAP7_75t_SL U62558 ( .A(n57214), .Y(n58167) );
  INVx2_ASAP7_75t_SL U62559 ( .A(n59711), .Y(n58169) );
  INVx1_ASAP7_75t_SL U62560 ( .A(n61921), .Y(n58707) );
  OR2x2_ASAP7_75t_SL U62561 ( .A(n58174), .B(n58172), .Y(n67902) );
  NAND2xp5_ASAP7_75t_SL U62562 ( .A(n58173), .B(n62649), .Y(n58174) );
  XNOR2x1_ASAP7_75t_SL U62563 ( .A(n59081), .B(n58177), .Y(n68580) );
  XNOR2x1_ASAP7_75t_SL U62564 ( .A(n68351), .B(n59266), .Y(n58177) );
  XNOR2x1_ASAP7_75t_SL U62565 ( .A(n68353), .B(n58178), .Y(n68351) );
  XNOR2x2_ASAP7_75t_SL U62566 ( .A(n68355), .B(n68354), .Y(n58178) );
  MAJIxp5_ASAP7_75t_SL U62567 ( .A(n66834), .B(n58529), .C(n66835), .Y(n66897)
         );
  XNOR2xp5_ASAP7_75t_SL U62568 ( .A(n58180), .B(n59296), .Y(n66835) );
  XOR2xp5_ASAP7_75t_SL U62569 ( .A(n57151), .B(n66688), .Y(n58180) );
  AO21x1_ASAP7_75t_SL U62570 ( .A1(n57041), .A2(n58181), .B(n58182), .Y(n63161) );
  NAND2xp5_ASAP7_75t_SL U62571 ( .A(n58183), .B(n63107), .Y(n58181) );
  NOR2x1_ASAP7_75t_SL U62572 ( .A(n58183), .B(n63107), .Y(n58182) );
  NAND2xp5_ASAP7_75t_SL U62573 ( .A(n58186), .B(n57380), .Y(n64429) );
  OAI21xp5_ASAP7_75t_SL U62574 ( .A1(n67944), .A2(n59617), .B(n58187), .Y(
        n64428) );
  NAND2xp5_ASAP7_75t_SL U62575 ( .A(n59617), .B(n75930), .Y(n58187) );
  OAI21xp5_ASAP7_75t_SL U62576 ( .A1(n57257), .A2(n76071), .B(n58188), .Y(
        n64461) );
  NAND2xp5_ASAP7_75t_SL U62577 ( .A(n67585), .B(n57257), .Y(n58188) );
  NOR2xp33_ASAP7_75t_SL U62578 ( .A(n57477), .B(n53314), .Y(n68959) );
  NOR3xp33_ASAP7_75t_SL U62579 ( .A(n53314), .B(n57477), .C(n68960), .Y(n68962) );
  NOR2x1_ASAP7_75t_SL U62580 ( .A(n68581), .B(n68580), .Y(n68956) );
  NOR2x1p5_ASAP7_75t_SL U62581 ( .A(n69117), .B(n58688), .Y(n58830) );
  AND2x2_ASAP7_75t_SL U62582 ( .A(n68919), .B(n68649), .Y(n58190) );
  AOI21x1_ASAP7_75t_SL U62583 ( .A1(n68920), .A2(n68919), .B(n68663), .Y(
        n58677) );
  O2A1O1Ixp5_ASAP7_75t_SL U62584 ( .A1(n67655), .A2(n67547), .B(n58195), .C(
        n67546), .Y(n67548) );
  NAND2xp5_ASAP7_75t_SL U62585 ( .A(n67544), .B(n67545), .Y(n58195) );
  OR2x2_ASAP7_75t_SL U62586 ( .A(n57140), .B(n68032), .Y(n58738) );
  NOR2x1_ASAP7_75t_SL U62587 ( .A(n67404), .B(n59460), .Y(n58198) );
  NOR2x1_ASAP7_75t_SL U62588 ( .A(n67473), .B(n59515), .Y(n58199) );
  OAI21xp5_ASAP7_75t_SL U62589 ( .A1(n59601), .A2(n75912), .B(n58200), .Y(
        n67751) );
  NAND2xp5_ASAP7_75t_SL U62590 ( .A(n59601), .B(n57662), .Y(n58200) );
  INVx1_ASAP7_75t_SL U62591 ( .A(n58201), .Y(n58204) );
  BUFx6f_ASAP7_75t_SL U62592 ( .A(n68010), .Y(n58202) );
  INVx1_ASAP7_75t_SL U62593 ( .A(n68010), .Y(n68008) );
  NAND2x2_ASAP7_75t_SL U62594 ( .A(n56840), .B(n59437), .Y(n68010) );
  NAND2xp5_ASAP7_75t_SL U62595 ( .A(n58203), .B(n62639), .Y(n58201) );
  INVx1_ASAP7_75t_SL U62596 ( .A(n62564), .Y(n58205) );
  OAI21xp33_ASAP7_75t_SL U62597 ( .A1(n62566), .A2(n62565), .B(n62567), .Y(
        n58208) );
  NAND2xp5_ASAP7_75t_SL U62598 ( .A(n64355), .B(n66258), .Y(n58210) );
  NOR2xp67_ASAP7_75t_SL U62599 ( .A(n57214), .B(n61909), .Y(n58214) );
  INVx1_ASAP7_75t_SL U62600 ( .A(n57466), .Y(n58213) );
  INVx2_ASAP7_75t_SL U62601 ( .A(n60747), .Y(n58215) );
  OAI21xp5_ASAP7_75t_SL U62602 ( .A1(n58216), .A2(n59380), .B(n67906), .Y(
        n67516) );
  NOR2x1_ASAP7_75t_SL U62603 ( .A(n58672), .B(n67250), .Y(n59380) );
  NAND2xp5_ASAP7_75t_SL U62604 ( .A(n57321), .B(n67248), .Y(n67249) );
  NAND2xp5_ASAP7_75t_SL U62605 ( .A(n58172), .B(n57112), .Y(n67248) );
  MAJIxp5_ASAP7_75t_SL U62606 ( .A(n63158), .B(n58217), .C(n63157), .Y(n63199)
         );
  OAI21xp5_ASAP7_75t_SL U62607 ( .A1(n75927), .A2(n58931), .B(n58935), .Y(
        n63066) );
  OAI21xp5_ASAP7_75t_SL U62608 ( .A1(n63070), .A2(n57159), .B(n63069), .Y(
        n58217) );
  OAI21xp5_ASAP7_75t_SL U62609 ( .A1(n63067), .A2(n56851), .B(n57159), .Y(
        n63069) );
  OAI21xp5_ASAP7_75t_SL U62610 ( .A1(n68834), .A2(n58219), .B(n68721), .Y(
        n58866) );
  INVx1_ASAP7_75t_SL U62611 ( .A(n62684), .Y(n58222) );
  OAI21xp5_ASAP7_75t_SL U62612 ( .A1(n59540), .A2(n62612), .B(n59479), .Y(
        n62684) );
  OA21x2_ASAP7_75t_SL U62613 ( .A1(n59378), .A2(n60915), .B(n64504), .Y(n59479) );
  NOR2x1_ASAP7_75t_SL U62614 ( .A(n60915), .B(n60596), .Y(n62612) );
  NAND2xp5_ASAP7_75t_SL U62615 ( .A(n67530), .B(n59179), .Y(n67258) );
  OR2x2_ASAP7_75t_SL U62616 ( .A(n57176), .B(n57104), .Y(n66658) );
  MAJIxp5_ASAP7_75t_SL U62617 ( .A(n66361), .B(n58224), .C(n66362), .Y(n66366)
         );
  INVx1_ASAP7_75t_SL U62618 ( .A(n66408), .Y(n58224) );
  O2A1O1Ixp5_ASAP7_75t_SL U62619 ( .A1(n53221), .A2(n66356), .B(n66355), .C(
        n66354), .Y(n66408) );
  NOR2x1_ASAP7_75t_SL U62620 ( .A(n57466), .B(n59264), .Y(n59263) );
  INVx1_ASAP7_75t_SL U62621 ( .A(n61964), .Y(n59264) );
  NOR2x1_ASAP7_75t_SL U62622 ( .A(n58226), .B(n58225), .Y(n61964) );
  NAND2xp5_ASAP7_75t_SL U62623 ( .A(n59546), .B(n59578), .Y(n58225) );
  NAND2xp5_ASAP7_75t_SL U62624 ( .A(n57068), .B(n59547), .Y(n58226) );
  OAI21xp33_ASAP7_75t_SL U62625 ( .A1(n53274), .A2(n67979), .B(n58228), .Y(
        n58227) );
  XNOR2xp5_ASAP7_75t_SL U62626 ( .A(n63154), .B(n63153), .Y(n63087) );
  NOR2x1_ASAP7_75t_SL U62627 ( .A(n58229), .B(n58632), .Y(n61931) );
  NAND2xp5_ASAP7_75t_SL U62628 ( .A(n1690), .B(n1929), .Y(n58229) );
  INVx1_ASAP7_75t_SL U62629 ( .A(n64516), .Y(n67851) );
  NOR2x1_ASAP7_75t_SL U62630 ( .A(n58231), .B(n58230), .Y(n64516) );
  NOR2x1_ASAP7_75t_SL U62631 ( .A(n63571), .B(n59654), .Y(n58230) );
  AOI21xp5_ASAP7_75t_SL U62632 ( .A1(n58353), .A2(n59712), .B(n59443), .Y(
        n58231) );
  NOR2x1p5_ASAP7_75t_SL U62633 ( .A(n63128), .B(n66798), .Y(n63182) );
  XNOR2xp5_ASAP7_75t_SL U62634 ( .A(n66972), .B(n66941), .Y(n58233) );
  OAI21xp5_ASAP7_75t_SL U62635 ( .A1(n57478), .A2(n59171), .B(n66712), .Y(
        n66972) );
  INVx1_ASAP7_75t_SL U62636 ( .A(n58460), .Y(n58234) );
  NAND2xp5_ASAP7_75t_SL U62637 ( .A(n58236), .B(n58941), .Y(n58235) );
  XNOR2xp5_ASAP7_75t_SL U62638 ( .A(n67070), .B(n58237), .Y(n67049) );
  XNOR2xp5_ASAP7_75t_SL U62639 ( .A(n68501), .B(n68502), .Y(n68503) );
  MAJIxp5_ASAP7_75t_SL U62640 ( .A(n58160), .B(n68450), .C(n68451), .Y(n68502)
         );
  NOR2xp67_ASAP7_75t_SL U62641 ( .A(n58239), .B(n58343), .Y(n58655) );
  NAND2xp33_ASAP7_75t_SL U62642 ( .A(n67623), .B(n67622), .Y(n58970) );
  INVx1_ASAP7_75t_SL U62643 ( .A(n59557), .Y(n59079) );
  NAND2xp5_ASAP7_75t_SL U62644 ( .A(n56861), .B(n59557), .Y(n58242) );
  OR2x2_ASAP7_75t_SL U62645 ( .A(n68566), .B(n68565), .Y(n68837) );
  XOR2xp5_ASAP7_75t_SL U62646 ( .A(n58243), .B(n68243), .Y(n68565) );
  NAND2xp5_ASAP7_75t_SL U62647 ( .A(n68250), .B(n68251), .Y(n68566) );
  XNOR2xp5_ASAP7_75t_SL U62648 ( .A(n58638), .B(n68249), .Y(n58243) );
  OAI21xp5_ASAP7_75t_SL U62649 ( .A1(n57119), .A2(n66270), .B(n58244), .Y(
        n58656) );
  NAND2xp5_ASAP7_75t_SL U62650 ( .A(n59576), .B(n66269), .Y(n58244) );
  INVx1_ASAP7_75t_SL U62651 ( .A(n59254), .Y(n59423) );
  INVx1_ASAP7_75t_SL U62652 ( .A(n57214), .Y(n58245) );
  MAJIxp5_ASAP7_75t_SL U62653 ( .A(n66875), .B(n59439), .C(n66874), .Y(n67012)
         );
  OAI22xp5_ASAP7_75t_SL U62654 ( .A1(n59165), .A2(n58246), .B1(n67586), .B2(
        n59666), .Y(n67097) );
  INVx1_ASAP7_75t_SL U62655 ( .A(n59666), .Y(n58246) );
  OAI22xp5_ASAP7_75t_SL U62656 ( .A1(n67738), .A2(n58934), .B1(n57172), .B2(
        n67408), .Y(n66768) );
  NAND2xp5_ASAP7_75t_SL U62657 ( .A(n58247), .B(n57000), .Y(n59439) );
  OAI21xp5_ASAP7_75t_SL U62658 ( .A1(n58669), .A2(n66617), .B(n67829), .Y(
        n58247) );
  NOR2x1_ASAP7_75t_SL U62659 ( .A(n58250), .B(n58249), .Y(n64357) );
  NAND2xp5_ASAP7_75t_SL U62660 ( .A(n60917), .B(n57960), .Y(n58249) );
  INVx1_ASAP7_75t_SL U62661 ( .A(n57424), .Y(n58251) );
  MAJx2_ASAP7_75t_SL U62662 ( .A(n59172), .B(n58252), .C(n68461), .Y(n66810)
         );
  INVx1_ASAP7_75t_SL U62663 ( .A(n68464), .Y(n58252) );
  MAJIxp5_ASAP7_75t_SL U62664 ( .A(n67934), .B(n67935), .C(n58253), .Y(n68033)
         );
  INVx1_ASAP7_75t_SL U62665 ( .A(n67994), .Y(n58254) );
  AOI22xp5_ASAP7_75t_SL U62666 ( .A1(n57161), .A2(n58413), .B1(n67456), .B2(
        n67306), .Y(n67835) );
  INVx1_ASAP7_75t_SL U62667 ( .A(n66938), .Y(n66732) );
  OAI21xp5_ASAP7_75t_SL U62668 ( .A1(n57158), .A2(n66731), .B(n58256), .Y(
        n66938) );
  OAI21xp5_ASAP7_75t_SL U62669 ( .A1(n59651), .A2(n68380), .B(n58257), .Y(
        n58256) );
  OAI21xp5_ASAP7_75t_SL U62670 ( .A1(n68900), .A2(n57481), .B(n76881), .Y(
        n58260) );
  OAI21xp5_ASAP7_75t_SL U62671 ( .A1(n68964), .A2(n68965), .B(n68963), .Y(
        n68978) );
  AOI21xp5_ASAP7_75t_SL U62672 ( .A1(n68962), .A2(n68961), .B(n57475), .Y(
        n68963) );
  INVx1_ASAP7_75t_SL U62673 ( .A(n68962), .Y(n68965) );
  XNOR2xp5_ASAP7_75t_SL U62674 ( .A(n68407), .B(n68405), .Y(n59150) );
  AOI22xp5_ASAP7_75t_SL U62675 ( .A1(n67702), .A2(n59229), .B1(n67912), .B2(
        n66964), .Y(n68407) );
  NOR2x1_ASAP7_75t_SL U62676 ( .A(n58261), .B(n56855), .Y(n67702) );
  NAND2xp5_ASAP7_75t_SL U62677 ( .A(n56847), .B(n59425), .Y(n58262) );
  INVx1_ASAP7_75t_SL U62678 ( .A(n64894), .Y(n58263) );
  INVx1_ASAP7_75t_SL U62679 ( .A(n67956), .Y(n58266) );
  NOR2xp33_ASAP7_75t_SL U62680 ( .A(n58808), .B(n74776), .Y(n58268) );
  XNOR2xp5_ASAP7_75t_SL U62681 ( .A(n58271), .B(n67683), .Y(n59159) );
  NAND2xp5_ASAP7_75t_SL U62682 ( .A(n58270), .B(n58269), .Y(n67683) );
  NAND2xp5_ASAP7_75t_SL U62683 ( .A(n67465), .B(n67464), .Y(n58269) );
  NAND2xp5_ASAP7_75t_SL U62684 ( .A(n67751), .B(n59613), .Y(n58270) );
  OAI21x1_ASAP7_75t_SL U62685 ( .A1(n62575), .A2(n56954), .B(n58272), .Y(
        n58273) );
  AND2x2_ASAP7_75t_SL U62686 ( .A(n56954), .B(n59588), .Y(n58274) );
  NAND2xp5_ASAP7_75t_SL U62687 ( .A(n58273), .B(n59644), .Y(n67711) );
  NAND2xp5_ASAP7_75t_SL U62688 ( .A(n59569), .B(n59570), .Y(n58276) );
  INVxp33_ASAP7_75t_SL U62689 ( .A(n62615), .Y(n62617) );
  NAND2xp5_ASAP7_75t_SL U62690 ( .A(n59555), .B(n64894), .Y(n58277) );
  NAND2xp5_ASAP7_75t_SL U62691 ( .A(or1200_ic_top_from_icram[27]), .B(n58387), 
        .Y(n60440) );
  OAI21xp5_ASAP7_75t_SL U62692 ( .A1(n73291), .A2(n73410), .B(n73290), .Y(
        n58278) );
  AO21x1_ASAP7_75t_SL U62693 ( .A1(n59678), .A2(n77870), .B(n58279), .Y(n9614)
         );
  AO211x2_ASAP7_75t_SL U62694 ( .A1(or1200_cpu_rf_datab[25]), .A2(n57091), .B(
        n77184), .C(n64257), .Y(n58279) );
  NAND2xp5_ASAP7_75t_SL U62695 ( .A(n61672), .B(n61671), .Y(n60776) );
  AOI21xp5_ASAP7_75t_SL U62696 ( .A1(n76275), .A2(n59499), .B(n75359), .Y(
        n75382) );
  NAND2xp5_ASAP7_75t_SL U62697 ( .A(n73235), .B(n73230), .Y(n73236) );
  NOR2x1_ASAP7_75t_SL U62698 ( .A(n63995), .B(n63996), .Y(n64001) );
  NOR2x1_ASAP7_75t_SL U62699 ( .A(n63994), .B(n63993), .Y(n63996) );
  NAND2xp5_ASAP7_75t_SL U62700 ( .A(n68879), .B(n68891), .Y(n76887) );
  NAND2xp5_ASAP7_75t_SL U62701 ( .A(n77958), .B(n77960), .Y(n77959) );
  NOR2x1_ASAP7_75t_SL U62702 ( .A(n74301), .B(n74304), .Y(n74333) );
  NAND2xp5_ASAP7_75t_SL U62703 ( .A(n62456), .B(n62455), .Y(n62454) );
  NAND2xp5_ASAP7_75t_SL U62704 ( .A(n61054), .B(n61053), .Y(n9675) );
  OAI21xp5_ASAP7_75t_SL U62705 ( .A1(n76117), .A2(n76116), .B(n76115), .Y(
        n76118) );
  INVx1_ASAP7_75t_SL U62706 ( .A(n76117), .Y(n76110) );
  XNOR2xp5_ASAP7_75t_SL U62707 ( .A(n76106), .B(n57107), .Y(n76117) );
  NOR2x1_ASAP7_75t_SL U62708 ( .A(n74057), .B(n74056), .Y(n74201) );
  NOR2x1_ASAP7_75t_SL U62709 ( .A(n66211), .B(n74875), .Y(n74056) );
  NAND2xp5_ASAP7_75t_SL U62710 ( .A(n74877), .B(n77195), .Y(n74905) );
  NOR2x1_ASAP7_75t_SL U62711 ( .A(n53290), .B(n57483), .Y(n60644) );
  NAND2xp5_ASAP7_75t_SL U62712 ( .A(n62096), .B(n75360), .Y(n63562) );
  NAND2xp5_ASAP7_75t_SL U62713 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[0]), .B(n57193), .Y(
        n66081) );
  NAND2xp5_ASAP7_75t_SL U62714 ( .A(n69407), .B(n69406), .Y(n69408) );
  INVx1_ASAP7_75t_SL U62715 ( .A(n60872), .Y(n60791) );
  NAND2xp5_ASAP7_75t_SL U62716 ( .A(n60618), .B(n60617), .Y(n61649) );
  NAND2xp5_ASAP7_75t_SL U62717 ( .A(n77351), .B(n77350), .Y(n77505) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U62718 ( .A1(n77623), .A2(n77622), .B(n77621), 
        .C(n77620), .Y(n77625) );
  NAND2xp5_ASAP7_75t_SL U62719 ( .A(n76906), .B(n76897), .Y(n63269) );
  NAND2xp5_ASAP7_75t_SL U62720 ( .A(n69182), .B(n68813), .Y(n76909) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U62721 ( .A1(n71512), .A2(n78368), .B(n78364), 
        .C(n70104), .Y(n70056) );
  INVx1_ASAP7_75t_SL U62722 ( .A(n72393), .Y(n72415) );
  AND2x2_ASAP7_75t_SL U62723 ( .A(n60440), .B(n60439), .Y(n58282) );
  AOI21xp5_ASAP7_75t_SL U62724 ( .A1(or1200_ic_top_from_icram[27]), .A2(n58387), .B(n60438), .Y(n61045) );
  NAND2xp5_ASAP7_75t_SL U62725 ( .A(n64808), .B(n64807), .Y(n9615) );
  AOI21xp5_ASAP7_75t_SL U62726 ( .A1(n63527), .A2(n63524), .B(n63523), .Y(
        n63528) );
  NAND3xp33_ASAP7_75t_SL U62727 ( .A(n74358), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_10_), 
        .C(or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_9_), .Y(n58283) );
  NAND2xp5_ASAP7_75t_SL U62728 ( .A(n70501), .B(n70099), .Y(n70101) );
  INVx1_ASAP7_75t_SL U62729 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[25]), .Y(n73690) );
  NAND2xp5_ASAP7_75t_SL U62730 ( .A(n60165), .B(n57100), .Y(n4130) );
  NAND2xp5_ASAP7_75t_SL U62731 ( .A(n63257), .B(n63256), .Y(n63258) );
  NOR2x1_ASAP7_75t_SL U62732 ( .A(n74750), .B(n74204), .Y(n74058) );
  NOR2x1_ASAP7_75t_SL U62733 ( .A(n74061), .B(n74060), .Y(n78199) );
  AOI21xp5_ASAP7_75t_SL U62734 ( .A1(n75901), .A2(n59230), .B(n63822), .Y(
        n64022) );
  NAND2xp5_ASAP7_75t_SL U62735 ( .A(n76040), .B(n75931), .Y(n76061) );
  NAND2x1p5_ASAP7_75t_SL U62736 ( .A(n78327), .B(n66260), .Y(n75915) );
  NAND2xp5_ASAP7_75t_SL U62737 ( .A(n66227), .B(n66226), .Y(n66231) );
  NAND2xp5_ASAP7_75t_SL U62738 ( .A(n75646), .B(n75647), .Y(n76891) );
  NAND2xp5_ASAP7_75t_SL U62739 ( .A(n74049), .B(n74048), .Y(
        or1200_cpu_or1200_except_n1706) );
  NAND2xp5_ASAP7_75t_SL U62740 ( .A(n77023), .B(n77022), .Y(
        or1200_cpu_or1200_except_n1716) );
  NOR2x1_ASAP7_75t_SL U62741 ( .A(n63704), .B(n77209), .Y(n63713) );
  NAND2xp5_ASAP7_75t_SL U62742 ( .A(n63362), .B(n63361), .Y(n63447) );
  NAND2xp5_ASAP7_75t_SL U62743 ( .A(n72318), .B(n71556), .Y(n71635) );
  NAND2xp5_ASAP7_75t_SL U62744 ( .A(n71548), .B(n71622), .Y(n71547) );
  OR2x2_ASAP7_75t_SL U62745 ( .A(n64217), .B(n64216), .Y(n58286) );
  NAND2xp5_ASAP7_75t_SL U62746 ( .A(n2843), .B(n77770), .Y(n62254) );
  OAI21xp5_ASAP7_75t_SL U62747 ( .A1(n74039), .A2(n74038), .B(n74037), .Y(
        or1200_cpu_to_sr[10]) );
  NOR2x1_ASAP7_75t_SL U62748 ( .A(n71218), .B(n71217), .Y(n71226) );
  XOR2xp5_ASAP7_75t_SL U62749 ( .A(n62946), .B(n62991), .Y(n62952) );
  NAND2xp5_ASAP7_75t_SL U62750 ( .A(n75929), .B(n76014), .Y(n76026) );
  NOR2x1_ASAP7_75t_SL U62751 ( .A(n64003), .B(n64004), .Y(n64008) );
  NOR2x1_ASAP7_75t_SL U62752 ( .A(n64002), .B(n64001), .Y(n64004) );
  NOR2x1_ASAP7_75t_SL U62753 ( .A(n74404), .B(n74405), .Y(n74403) );
  NAND2xp5_ASAP7_75t_SL U62754 ( .A(or1200_cpu_or1200_mult_mac_n145), .B(
        n63282), .Y(n63302) );
  INVx1_ASAP7_75t_SL U62755 ( .A(or1200_cpu_or1200_mult_mac_n291), .Y(n63282)
         );
  OAI21xp5_ASAP7_75t_SL U62756 ( .A1(n63781), .A2(n63782), .B(n63780), .Y(
        n63532) );
  NAND2xp5_ASAP7_75t_SL U62757 ( .A(n60068), .B(n57100), .Y(n4116) );
  NAND2xp5_ASAP7_75t_SL U62758 ( .A(n72597), .B(n74239), .Y(n74275) );
  NOR2x1_ASAP7_75t_SL U62759 ( .A(n74072), .B(n74739), .Y(n74250) );
  NAND2xp5_ASAP7_75t_SL U62760 ( .A(n76209), .B(n76208), .Y(
        or1200_cpu_or1200_except_n1725) );
  OAI21xp5_ASAP7_75t_SL U62761 ( .A1(n2991), .A2(n74953), .B(n60033), .Y(
        n60034) );
  INVx1_ASAP7_75t_SL U62762 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[2]), .Y(n74093) );
  NAND2xp5_ASAP7_75t_SL U62763 ( .A(n75800), .B(n75799), .Y(
        or1200_cpu_or1200_except_n1703) );
  NAND2xp5_ASAP7_75t_SL U62764 ( .A(n75435), .B(n75434), .Y(
        or1200_cpu_or1200_except_n1709) );
  NAND2xp5_ASAP7_75t_SL U62765 ( .A(n74988), .B(n74987), .Y(
        or1200_cpu_or1200_except_n1712) );
  NAND2xp5_ASAP7_75t_SL U62766 ( .A(n75785), .B(n75784), .Y(
        or1200_cpu_or1200_except_n1720) );
  NAND2xp5_ASAP7_75t_SL U62767 ( .A(n62205), .B(n62319), .Y(n60549) );
  NAND2xp5_ASAP7_75t_SL U62768 ( .A(n76248), .B(n76247), .Y(
        or1200_cpu_or1200_except_n1721) );
  NAND2xp5_ASAP7_75t_SL U62769 ( .A(n75624), .B(n75623), .Y(
        or1200_cpu_or1200_except_n1707) );
  NAND2xp5_ASAP7_75t_SL U62770 ( .A(n75451), .B(n75450), .Y(
        or1200_cpu_or1200_except_n1708) );
  NAND2xp5_ASAP7_75t_SL U62771 ( .A(n74597), .B(n74596), .Y(n74595) );
  OAI22xp5_ASAP7_75t_SL U62772 ( .A1(n60435), .A2(n77954), .B1(n2974), .B2(
        n78009), .Y(n60436) );
  NOR2x1_ASAP7_75t_SL U62773 ( .A(n74325), .B(n74326), .Y(n74338) );
  NAND2xp5_ASAP7_75t_SL U62774 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_31_), .B(
        n74320), .Y(n74326) );
  NAND2xp5_ASAP7_75t_SL U62775 ( .A(n65245), .B(n65244), .Y(n65246) );
  INVx1_ASAP7_75t_SL U62776 ( .A(n59531), .Y(n76874) );
  BUFx6f_ASAP7_75t_SL U62777 ( .A(n1636), .Y(n59531) );
  AOI22xp5_ASAP7_75t_SL U62778 ( .A1(n59531), .A2(n59711), .B1(n57377), .B2(
        n59712), .Y(n61492) );
  NAND2xp5_ASAP7_75t_SL U62779 ( .A(n59531), .B(n61946), .Y(n62073) );
  NAND2xp5_ASAP7_75t_SL U62780 ( .A(n59531), .B(n77715), .Y(n74598) );
  OAI21xp5_ASAP7_75t_SL U62781 ( .A1(n71182), .A2(n71205), .B(n71181), .Y(
        n71185) );
  NAND2xp5_ASAP7_75t_SL U62782 ( .A(n60228), .B(n77663), .Y(n58287) );
  NAND2xp5_ASAP7_75t_SL U62783 ( .A(n60228), .B(n77663), .Y(n60231) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U62784 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .A2(
        n72313), .B(n57125), .C(n72312), .Y(n72314) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U62785 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .A2(
        n72341), .B(n57127), .C(n72342), .Y(n72258) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U62786 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .A2(
        n72351), .B(n57125), .C(n72349), .Y(n72260) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U62787 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .A2(
        n72309), .B(n57127), .C(n72293), .Y(n72254) );
  INVx1_ASAP7_75t_SL U62788 ( .A(n60438), .Y(n60439) );
  NAND2xp5_ASAP7_75t_SL U62789 ( .A(n61429), .B(n61215), .Y(n61514) );
  NOR2x1_ASAP7_75t_SL U62790 ( .A(n58592), .B(n64008), .Y(n64010) );
  NOR2x1_ASAP7_75t_SL U62791 ( .A(n59526), .B(n70686), .Y(n70674) );
  NAND2xp5_ASAP7_75t_SL U62792 ( .A(or1200_dc_top_tag_v), .B(n59768), .Y(
        n59769) );
  NAND2xp5_ASAP7_75t_SL U62793 ( .A(n71254), .B(n71258), .Y(n71240) );
  OR2x2_ASAP7_75t_SL U62794 ( .A(n70841), .B(n70840), .Y(n58288) );
  OR2x2_ASAP7_75t_SL U62795 ( .A(dbg_adr_i[11]), .B(n78439), .Y(n58289) );
  OR2x2_ASAP7_75t_SL U62796 ( .A(dbg_stb_i), .B(n76547), .Y(n58290) );
  NAND2xp5_ASAP7_75t_SL U62797 ( .A(n60099), .B(n57100), .Y(n4128) );
  NAND2xp5_ASAP7_75t_SL U62798 ( .A(n59755), .B(n59754), .Y(n59756) );
  INVx1_ASAP7_75t_SL U62799 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .Y(n78373) );
  NOR2x1_ASAP7_75t_SL U62800 ( .A(n74495), .B(n69977), .Y(n70081) );
  NAND2xp5_ASAP7_75t_SL U62801 ( .A(n74499), .B(n70081), .Y(n70166) );
  NAND2xp5_ASAP7_75t_SL U62802 ( .A(n59736), .B(n59735), .Y(n59745) );
  NOR2x1_ASAP7_75t_SL U62803 ( .A(n77678), .B(n60229), .Y(n73960) );
  NAND2xp5_ASAP7_75t_SL U62804 ( .A(n74580), .B(n74579), .Y(
        or1200_cpu_or1200_except_n1711) );
  NAND2xp5_ASAP7_75t_SL U62805 ( .A(n76234), .B(n76233), .Y(
        or1200_cpu_or1200_except_n1714) );
  NAND2xp5_ASAP7_75t_SL U62806 ( .A(n75305), .B(n75304), .Y(
        or1200_cpu_or1200_except_n1713) );
  NAND2xp5_ASAP7_75t_SL U62807 ( .A(n75202), .B(n75201), .Y(
        or1200_cpu_or1200_except_n1701) );
  INVx1_ASAP7_75t_SL U62808 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[5]), .Y(
        n73221) );
  NAND2xp5_ASAP7_75t_SL U62809 ( .A(n4122), .B(n78257), .Y(icqmem_adr_qmem[18]) );
  NAND2xp5_ASAP7_75t_SL U62810 ( .A(n75678), .B(n75677), .Y(
        or1200_cpu_or1200_except_n1700) );
  OAI21xp5_ASAP7_75t_SL U62811 ( .A1(or1200_cpu_or1200_mult_mac_n52), .A2(
        n76158), .B(n76017), .Y(or1200_cpu_or1200_mult_mac_n1520) );
  OAI21xp5_ASAP7_75t_SL U62812 ( .A1(or1200_cpu_or1200_mult_mac_n22), .A2(
        n76158), .B(n76142), .Y(or1200_cpu_or1200_mult_mac_n1505) );
  OAI21xp5_ASAP7_75t_SL U62813 ( .A1(or1200_cpu_or1200_mult_mac_n18), .A2(
        n76158), .B(n76157), .Y(or1200_cpu_or1200_mult_mac_n1503) );
  AOI21xp5_ASAP7_75t_SL U62814 ( .A1(n71258), .A2(n71257), .B(n71256), .Y(
        n71259) );
  NAND2xp5_ASAP7_75t_SL U62815 ( .A(n76072), .B(n57133), .Y(n76073) );
  NAND2xp5_ASAP7_75t_SL U62816 ( .A(n76055), .B(n57133), .Y(n76056) );
  NAND2xp5_ASAP7_75t_SL U62817 ( .A(n76029), .B(n57133), .Y(n76030) );
  NAND2xp5_ASAP7_75t_SL U62818 ( .A(n75992), .B(n57133), .Y(n75993) );
  NAND2xp5_ASAP7_75t_SL U62819 ( .A(n75982), .B(n75981), .Y(
        or1200_cpu_or1200_mult_mac_n1526) );
  AOI21xp5_ASAP7_75t_SL U62820 ( .A1(n71785), .A2(n71709), .B(n71720), .Y(
        n71686) );
  INVx6_ASAP7_75t_SL U62821 ( .A(n56827), .Y(n59594) );
  XNOR2xp5_ASAP7_75t_SL U62822 ( .A(n56827), .B(n59510), .Y(n63070) );
  OAI21xp5_ASAP7_75t_SL U62823 ( .A1(n69780), .A2(n69785), .B(n69781), .Y(
        n69789) );
  NAND2xp5_ASAP7_75t_SL U62824 ( .A(n69601), .B(n69786), .Y(n69781) );
  NAND2xp5_ASAP7_75t_SL U62825 ( .A(n76182), .B(n57133), .Y(n76183) );
  NAND2xp5_ASAP7_75t_SL U62826 ( .A(n76119), .B(n57133), .Y(n76120) );
  NAND2xp5_ASAP7_75t_SL U62827 ( .A(n76168), .B(n57133), .Y(n76169) );
  NAND2xp5_ASAP7_75t_SL U62828 ( .A(n76178), .B(n57133), .Y(n76179) );
  AOI22xp5_ASAP7_75t_SL U62829 ( .A1(n60805), .A2(n57121), .B1(n59498), .B2(
        n60965), .Y(n60936) );
  NOR2x1_ASAP7_75t_SL U62830 ( .A(n53429), .B(n78182), .Y(n61827) );
  AOI22xp5_ASAP7_75t_SL U62831 ( .A1(n63422), .A2(n57121), .B1(n61827), .B2(
        n61764), .Y(n61830) );
  AOI22xp5_ASAP7_75t_SL U62832 ( .A1(n63483), .A2(n57121), .B1(n53430), .B2(
        n60811), .Y(n61829) );
  AOI22xp5_ASAP7_75t_SL U62833 ( .A1(n75341), .A2(n57121), .B1(n61827), .B2(
        n75337), .Y(n62096) );
  AOI22xp5_ASAP7_75t_SL U62834 ( .A1(n61822), .A2(n57121), .B1(n61827), .B2(
        n74609), .Y(n74597) );
  NAND2xp5_ASAP7_75t_SL U62835 ( .A(n72990), .B(n72769), .Y(n73032) );
  OAI21xp5_ASAP7_75t_SL U62836 ( .A1(n59627), .A2(n78337), .B(n72820), .Y(
        n72938) );
  NAND2xp5_ASAP7_75t_SL U62837 ( .A(n63705), .B(n63726), .Y(n76931) );
  NAND2xp5_ASAP7_75t_SL U62838 ( .A(n76173), .B(n57133), .Y(n76174) );
  NOR2xp33_ASAP7_75t_SL U62839 ( .A(n58295), .B(n71205), .Y(n58292) );
  OR2x2_ASAP7_75t_SL U62840 ( .A(n58292), .B(n58293), .Y(n71217) );
  AND2x2_ASAP7_75t_SL U62841 ( .A(n58294), .B(n71238), .Y(n58293) );
  OR2x2_ASAP7_75t_SL U62842 ( .A(n71206), .B(n71214), .Y(n58295) );
  NAND2xp5_ASAP7_75t_SL U62843 ( .A(n70855), .B(n70856), .Y(n71026) );
  NAND2xp5_ASAP7_75t_SL U62844 ( .A(n70854), .B(n70853), .Y(n70856) );
  OAI21xp5_ASAP7_75t_SL U62845 ( .A1(or1200_cpu_or1200_mult_mac_n44), .A2(
        n76158), .B(n76046), .Y(or1200_cpu_or1200_mult_mac_n1516) );
  OAI21xp5_ASAP7_75t_SL U62846 ( .A1(or1200_cpu_or1200_mult_mac_n40), .A2(
        n76158), .B(n76066), .Y(or1200_cpu_or1200_mult_mac_n1514) );
  OAI21xp5_ASAP7_75t_SL U62847 ( .A1(or1200_cpu_or1200_mult_mac_n56), .A2(
        n76158), .B(n76000), .Y(or1200_cpu_or1200_mult_mac_n1522) );
  OAI21xp5_ASAP7_75t_SL U62848 ( .A1(or1200_cpu_or1200_mult_mac_n50), .A2(
        n76158), .B(n76024), .Y(or1200_cpu_or1200_mult_mac_n1519) );
  OAI21xp5_ASAP7_75t_SL U62849 ( .A1(or1200_cpu_or1200_mult_mac_n28), .A2(
        n76158), .B(n76113), .Y(or1200_cpu_or1200_mult_mac_n1508) );
  NOR2x1_ASAP7_75t_SL U62850 ( .A(n64009), .B(n64010), .Y(n64012) );
  NAND2xp5_ASAP7_75t_SL U62851 ( .A(n71434), .B(n71470), .Y(n71494) );
  NAND2xp5_ASAP7_75t_SL U62852 ( .A(n60120), .B(n57100), .Y(n4126) );
  OAI21xp5_ASAP7_75t_SL U62853 ( .A1(or1200_cpu_or1200_mult_mac_n411), .A2(
        n76894), .B(n76893), .Y(n76916) );
  OAI21xp5_ASAP7_75t_SL U62854 ( .A1(n77846), .A2(n77845), .B(n77844), .Y(
        or1200_cpu_or1200_rf_N36) );
  OAI22xp5_ASAP7_75t_SL U62855 ( .A1(n57115), .A2(n70735), .B1(n70722), .B2(
        n59524), .Y(n71064) );
  NAND2xp5_ASAP7_75t_SL U62856 ( .A(n76058), .B(n76057), .Y(n76067) );
  OAI21xp5_ASAP7_75t_SL U62857 ( .A1(n71365), .A2(n70828), .B(n70827), .Y(
        n70830) );
  AOI21xp5_ASAP7_75t_SL U62858 ( .A1(n77012), .A2(n59945), .B(n59727), .Y(
        n59838) );
  NAND2xp5_ASAP7_75t_SL U62859 ( .A(n60113), .B(n57100), .Y(n4124) );
  NOR2x1_ASAP7_75t_SL U62860 ( .A(n74361), .B(n74418), .Y(n74258) );
  AOI21xp5_ASAP7_75t_SL U62861 ( .A1(n71180), .A2(n71179), .B(n71178), .Y(
        n71201) );
  NAND2xp5_ASAP7_75t_SL U62862 ( .A(n71168), .B(n71167), .Y(n71180) );
  INVx1_ASAP7_75t_SL U62863 ( .A(n70986), .Y(n71117) );
  OR2x2_ASAP7_75t_SL U62864 ( .A(n74361), .B(n74736), .Y(n58298) );
  INVx1_ASAP7_75t_SL U62865 ( .A(n74418), .Y(n74736) );
  NAND2xp5_ASAP7_75t_SL U62866 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[8]), .B(
        n73382), .Y(n73207) );
  NOR2x1_ASAP7_75t_SL U62867 ( .A(n70935), .B(n70936), .Y(n70970) );
  OR2x2_ASAP7_75t_SL U62868 ( .A(n76503), .B(n58287), .Y(n58299) );
  NAND2xp5_ASAP7_75t_SL U62869 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[23]), .B(n71013), 
        .Y(n58301) );
  NOR2xp33_ASAP7_75t_SL U62870 ( .A(n60834), .B(n60833), .Y(n61060) );
  INVx1_ASAP7_75t_SL U62871 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_2_), .Y(n76946)
         );
  NAND2xp5_ASAP7_75t_SL U62872 ( .A(n57100), .B(n65192), .Y(n4108) );
  NAND2xp5_ASAP7_75t_SL U62873 ( .A(n77506), .B(n77343), .Y(n77399) );
  AOI21xp5_ASAP7_75t_SL U62874 ( .A1(n78090), .A2(n78092), .B(n69362), .Y(
        n69364) );
  OR3x1_ASAP7_75t_SL U62875 ( .A(n78100), .B(n69362), .C(n75188), .Y(n75794)
         );
  INVx1_ASAP7_75t_SL U62876 ( .A(n59798), .Y(n69362) );
  NAND2xp5_ASAP7_75t_SL U62877 ( .A(n60133), .B(n57100), .Y(n4120) );
  NAND2xp5_ASAP7_75t_SL U62878 ( .A(n70153), .B(n69899), .Y(n69877) );
  NAND2xp5_ASAP7_75t_SL U62879 ( .A(n70153), .B(n70135), .Y(n69878) );
  NOR2x1_ASAP7_75t_SL U62880 ( .A(n62582), .B(n62675), .Y(n67625) );
  NOR2x1_ASAP7_75t_SL U62881 ( .A(or1200_cpu_or1200_mult_mac_n46), .B(n53261), 
        .Y(n76042) );
  NAND2xp5_ASAP7_75t_SL U62882 ( .A(or1200_cpu_or1200_mult_mac_n26), .B(n59459), .Y(n75938) );
  NOR2x1_ASAP7_75t_SL U62883 ( .A(n60216), .B(n76542), .Y(n74925) );
  NAND2xp5_ASAP7_75t_SL U62884 ( .A(n70673), .B(n70672), .Y(n70681) );
  OAI21xp5_ASAP7_75t_SL U62885 ( .A1(n63877), .A2(n63687), .B(n64746), .Y(
        n63885) );
  OAI22xp5_ASAP7_75t_SL U62886 ( .A1(n70704), .A2(n70703), .B1(n70702), .B2(
        n70701), .Y(n70714) );
  INVx1_ASAP7_75t_SL U62887 ( .A(or1200_cpu_or1200_mult_mac_n321), .Y(n75341)
         );
  AOI21xp5_ASAP7_75t_SL U62888 ( .A1(n73576), .A2(n73544), .B(n73543), .Y(
        n73549) );
  NAND2xp5_ASAP7_75t_SL U62889 ( .A(n73578), .B(n73577), .Y(n73576) );
  NOR2x1_ASAP7_75t_SL U62890 ( .A(n58601), .B(n64012), .Y(n74968) );
  NAND2xp5_ASAP7_75t_SL U62891 ( .A(n59854), .B(n74122), .Y(n74982) );
  NAND2xp5_ASAP7_75t_SL U62892 ( .A(n75299), .B(n59854), .Y(n74123) );
  INVx3_ASAP7_75t_SL U62893 ( .A(n75841), .Y(n59646) );
  NAND2x1_ASAP7_75t_SL U62894 ( .A(n59711), .B(n59442), .Y(n75841) );
  NAND2xp5_ASAP7_75t_SL U62895 ( .A(n73437), .B(n58278), .Y(n73442) );
  NOR2xp33_ASAP7_75t_SL U62896 ( .A(n70921), .B(n70920), .Y(n70973) );
  INVx1_ASAP7_75t_SL U62897 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[21]), .Y(
        n73119) );
  OAI21xp5_ASAP7_75t_SL U62898 ( .A1(n53288), .A2(n76181), .B(n75963), .Y(
        n75969) );
  NAND2xp5_ASAP7_75t_SL U62899 ( .A(n59954), .B(n77304), .Y(n60325) );
  NOR2x1_ASAP7_75t_SL U62900 ( .A(n60191), .B(n77356), .Y(n60202) );
  NOR2x1_ASAP7_75t_SL U62901 ( .A(n60421), .B(n60401), .Y(n77356) );
  OR2x2_ASAP7_75t_SL U62902 ( .A(n73581), .B(n73562), .Y(n58304) );
  NAND2xp5_ASAP7_75t_SL U62903 ( .A(n71263), .B(n71140), .Y(n70957) );
  NAND2xp5_ASAP7_75t_SL U62904 ( .A(n70953), .B(n70952), .Y(n71140) );
  NAND2xp5_ASAP7_75t_SL U62905 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_29_), .B(n71121), 
        .Y(n71127) );
  AND2x2_ASAP7_75t_SL U62906 ( .A(n61201), .B(n60748), .Y(n58305) );
  OAI21xp5_ASAP7_75t_SL U62907 ( .A1(n59443), .A2(n60747), .B(n57214), .Y(
        n61201) );
  INVx1_ASAP7_75t_SL U62908 ( .A(n62519), .Y(n60748) );
  NOR2x1_ASAP7_75t_SL U62909 ( .A(n61855), .B(n60626), .Y(n76782) );
  INVx1_ASAP7_75t_SL U62910 ( .A(n75453), .Y(n60834) );
  AOI21xp5_ASAP7_75t_SL U62911 ( .A1(n76298), .A2(n59499), .B(n62390), .Y(
        n76654) );
  OAI21xp5_ASAP7_75t_SL U62912 ( .A1(n71281), .A2(n71103), .B(n71102), .Y(
        n71248) );
  OAI21xp5_ASAP7_75t_SL U62913 ( .A1(n71281), .A2(n71221), .B(n71220), .Y(
        n71393) );
  NAND2xp5_ASAP7_75t_SL U62914 ( .A(n61944), .B(n62094), .Y(n64146) );
  INVx1_ASAP7_75t_SL U62915 ( .A(n64208), .Y(n60552) );
  INVx1_ASAP7_75t_SL U62916 ( .A(n58287), .Y(n60229) );
  NOR2x1p5_ASAP7_75t_SL U62917 ( .A(n59596), .B(n67837), .Y(n67566) );
  NAND2xp5_ASAP7_75t_SL U62918 ( .A(n65249), .B(n65248), .Y(n65250) );
  NOR2x1_ASAP7_75t_SL U62919 ( .A(n76529), .B(n76528), .Y(n63981) );
  OAI21xp5_ASAP7_75t_SL U62920 ( .A1(or1200_cpu_or1200_mult_mac_n34), .A2(
        n76158), .B(n76086), .Y(or1200_cpu_or1200_mult_mac_n1511) );
  INVx1_ASAP7_75t_SL U62921 ( .A(n75940), .Y(n76165) );
  NAND2xp5_ASAP7_75t_SL U62922 ( .A(n71731), .B(n71687), .Y(n71690) );
  OAI21xp5_ASAP7_75t_SL U62923 ( .A1(n71719), .A2(n71718), .B(n71800), .Y(
        n71717) );
  INVx1_ASAP7_75t_SL U62924 ( .A(n71679), .Y(n71718) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U62925 ( .A1(n74713), .A2(n74712), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .C(
        n74711), .Y(n74714) );
  NAND2xp5_ASAP7_75t_SL U62926 ( .A(n70566), .B(n74285), .Y(n74711) );
  OAI22xp5_ASAP7_75t_SL U62927 ( .A1(n76057), .A2(n58517), .B1(n67328), .B2(
        n57167), .Y(n59129) );
  NAND2xp5_ASAP7_75t_SL U62928 ( .A(n63686), .B(n63685), .Y(n64746) );
  INVx1_ASAP7_75t_SL U62929 ( .A(n58281), .Y(n58306) );
  NAND2xp5_ASAP7_75t_SL U62930 ( .A(n68747), .B(n68746), .Y(n52061) );
  NAND2xp5_ASAP7_75t_SL U62931 ( .A(n69355), .B(n59764), .Y(n75440) );
  FAx1_ASAP7_75t_SL U62932 ( .A(or1200_dc_top_tag_10_), .B(n59767), .CI(n59766), .CON(), .SN(n59768) );
  NAND2xp5_ASAP7_75t_SL U62933 ( .A(n61838), .B(n74593), .Y(n64107) );
  NAND2xp5_ASAP7_75t_SL U62934 ( .A(n69373), .B(n64814), .Y(n73905) );
  NAND2xp5_ASAP7_75t_SL U62935 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_25_), .B(n71062), 
        .Y(n71080) );
  AOI22xp5_ASAP7_75t_SL U62936 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[5]), .A2(n70668), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[13]), .B2(
        n58300), .Y(n70670) );
  AOI22xp5_ASAP7_75t_SL U62937 ( .A1(n70668), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[4]), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[12]), .B2(n58300), 
        .Y(n70663) );
  AOI22xp5_ASAP7_75t_SL U62938 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[6]), .A2(n70668), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[14]), .B2(
        n58300), .Y(n70660) );
  NAND2xp5_ASAP7_75t_SL U62939 ( .A(n71350), .B(n58311), .Y(n58308) );
  AND2x2_ASAP7_75t_SL U62940 ( .A(n58308), .B(n58309), .Y(n71388) );
  OR2x2_ASAP7_75t_SL U62941 ( .A(n58310), .B(n71344), .Y(n58309) );
  AND2x2_ASAP7_75t_SL U62942 ( .A(n71309), .B(n71327), .Y(n58311) );
  NAND2xp5_ASAP7_75t_SL U62943 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_0_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_1_), .Y(n74840)
         );
  OAI22xp5_ASAP7_75t_SL U62944 ( .A1(dbg_stb_i), .A2(n76199), .B1(dbg_adr_i[5]), .B2(n78439), .Y(n60573) );
  OAI21xp5_ASAP7_75t_SL U62945 ( .A1(n60874), .A2(n61078), .B(n60873), .Y(
        n77087) );
  INVx1_ASAP7_75t_SL U62946 ( .A(n61547), .Y(n61078) );
  OAI22xp5_ASAP7_75t_SL U62947 ( .A1(n72993), .A2(n72900), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), 
        .B2(n72886), .Y(n72723) );
  NOR2x1_ASAP7_75t_SL U62948 ( .A(n2589), .B(n57072), .Y(n61155) );
  NAND2xp5_ASAP7_75t_SL U62949 ( .A(n77425), .B(n60360), .Y(n61160) );
  INVx1_ASAP7_75t_SL U62950 ( .A(n60756), .Y(n60979) );
  NAND2xp5_ASAP7_75t_SL U62951 ( .A(n75265), .B(n75264), .Y(n75270) );
  NAND2xp5_ASAP7_75t_SL U62952 ( .A(n71327), .B(n71326), .Y(n58312) );
  NAND2xp5_ASAP7_75t_SL U62953 ( .A(n73448), .B(n73447), .Y(n73446) );
  NAND2xp5_ASAP7_75t_SL U62954 ( .A(n73364), .B(n73446), .Y(n73365) );
  NAND2xp5_ASAP7_75t_SL U62955 ( .A(n58416), .B(n77163), .Y(n77239) );
  AND2x2_ASAP7_75t_SL U62956 ( .A(n68723), .B(n68722), .Y(n58313) );
  AOI21xp5_ASAP7_75t_SL U62957 ( .A1(n76299), .A2(n59499), .B(n61376), .Y(
        n77907) );
  NAND2xp5_ASAP7_75t_SL U62958 ( .A(n53468), .B(n76108), .Y(n76116) );
  NAND2xp5_ASAP7_75t_SL U62959 ( .A(n60549), .B(n60548), .Y(n73907) );
  NAND2xp5_ASAP7_75t_SL U62960 ( .A(n77621), .B(n60559), .Y(n60548) );
  OAI21xp5_ASAP7_75t_SL U62961 ( .A1(n76075), .A2(n75911), .B(n75910), .Y(
        n76087) );
  NAND2xp5_ASAP7_75t_SL U62962 ( .A(n76079), .B(n76074), .Y(n75911) );
  INVx1_ASAP7_75t_SL U62963 ( .A(n76089), .Y(n76125) );
  INVx1_ASAP7_75t_SL U62964 ( .A(n58307), .Y(n58314) );
  OAI21xp5_ASAP7_75t_SL U62965 ( .A1(n63954), .A2(n63953), .B(n63952), .Y(
        n76528) );
  INVx1_ASAP7_75t_SL U62966 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_), 
        .Y(n72350) );
  NAND2xp5_ASAP7_75t_SL U62967 ( .A(n72234), .B(n71424), .Y(n71481) );
  AOI21xp5_ASAP7_75t_SL U62968 ( .A1(n61560), .A2(n61399), .B(n61400), .Y(
        n60764) );
  NAND2xp5_ASAP7_75t_SL U62969 ( .A(n3327), .B(n73633), .Y(n73523) );
  INVx1_ASAP7_75t_SL U62970 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[9]), .Y(n73633) );
  NOR2x1_ASAP7_75t_SL U62971 ( .A(n68745), .B(n68744), .Y(n76882) );
  XNOR2x2_ASAP7_75t_SL U62972 ( .A(n27420), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n254), .Y(n73379) );
  NOR2x1_ASAP7_75t_SL U62973 ( .A(n66205), .B(n76954), .Y(n74884) );
  NAND2xp5_ASAP7_75t_SL U62974 ( .A(n57318), .B(n60645), .Y(n62012) );
  NAND2xp5_ASAP7_75t_SL U62975 ( .A(n57353), .B(n62012), .Y(n76751) );
  NOR2x1_ASAP7_75t_SL U62976 ( .A(n73899), .B(n73898), .Y(n74739) );
  NAND2xp5_ASAP7_75t_SL U62977 ( .A(n66213), .B(n74161), .Y(n74205) );
  INVx1_ASAP7_75t_SL U62978 ( .A(n74203), .Y(n74161) );
  AOI22xp5_ASAP7_75t_SL U62979 ( .A1(dwb_dat_i[23]), .A2(n61548), .B1(n75569), 
        .B2(dwb_dat_i[31]), .Y(n60881) );
  NOR2x1_ASAP7_75t_SL U62980 ( .A(n62254), .B(n61547), .Y(n61548) );
  NAND2xp5_ASAP7_75t_SL U62981 ( .A(n76138), .B(n76123), .Y(n76145) );
  OAI21xp5_ASAP7_75t_SL U62982 ( .A1(or1200_cpu_or1200_mult_mac_n46), .A2(
        n76158), .B(n76039), .Y(or1200_cpu_or1200_mult_mac_n1517) );
  OAI21xp5_ASAP7_75t_SL U62983 ( .A1(or1200_cpu_or1200_mult_mac_n30), .A2(
        n76158), .B(n76107), .Y(or1200_cpu_or1200_mult_mac_n1509) );
  INVx1_ASAP7_75t_SL U62984 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[16]), .Y(
        n73128) );
  NAND2xp5_ASAP7_75t_SL U62985 ( .A(n71005), .B(n71006), .Y(n71027) );
  NAND2xp5_ASAP7_75t_SL U62986 ( .A(n60145), .B(n57100), .Y(n4122) );
  NAND2xp5_ASAP7_75t_SL U62987 ( .A(n60220), .B(n76538), .Y(n76541) );
  NAND2x1_ASAP7_75t_SL U62988 ( .A(n66634), .B(n65017), .Y(n66376) );
  AOI21xp5_ASAP7_75t_SL U62989 ( .A1(n76270), .A2(n59499), .B(n75756), .Y(
        n77857) );
  BUFx10_ASAP7_75t_SL U62990 ( .A(n75923), .Y(n59511) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U62991 ( .A1(n77998), .A2(n77470), .B(n58570), 
        .C(n3418), .Y(n77762) );
  NAND2xp5_ASAP7_75t_SL U62992 ( .A(n58684), .B(n76879), .Y(n58683) );
  XNOR2xp5_ASAP7_75t_SL U62993 ( .A(n63038), .B(n58461), .Y(n63444) );
  INVx1_ASAP7_75t_SL U62994 ( .A(n63038), .Y(n63039) );
  NAND2xp5_ASAP7_75t_SL U62995 ( .A(n59694), .B(n77897), .Y(n77024) );
  AO21x2_ASAP7_75t_SL U62996 ( .A1(n72611), .A2(n72610), .B(n72609), .Y(n73047) );
  OAI21xp5_ASAP7_75t_SL U62997 ( .A1(n59631), .A2(n73239), .B(n73237), .Y(
        n73247) );
  NAND2xp5_ASAP7_75t_SL U62998 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[3]), .B(
        n59630), .Y(n73237) );
  AOI21xp5_ASAP7_75t_SL U62999 ( .A1(n57316), .A2(n62656), .B(n78002), .Y(
        n62632) );
  INVx1_ASAP7_75t_SL U63000 ( .A(n59867), .Y(n75190) );
  NAND2x1_ASAP7_75t_SL U63001 ( .A(n2145), .B(n59555), .Y(n59935) );
  AND2x4_ASAP7_75t_SL U63002 ( .A(n59655), .B(n66637), .Y(n66634) );
  NOR2x1_ASAP7_75t_SL U63003 ( .A(n59526), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_0_), .Y(n70676) );
  NOR2x1_ASAP7_75t_SL U63004 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_0_), .B(n71365), .Y(
        n70675) );
  NAND2xp5_ASAP7_75t_SL U63005 ( .A(n74629), .B(n74628), .Y(n74627) );
  OAI21xp5_ASAP7_75t_SL U63006 ( .A1(n62085), .A2(n75306), .B(n62084), .Y(
        n74628) );
  OAI22xp5_ASAP7_75t_SL U63007 ( .A1(n68798), .A2(n74998), .B1(n68797), .B2(
        n75016), .Y(n68818) );
  NAND2xp5_ASAP7_75t_SL U63008 ( .A(n60320), .B(n77839), .Y(n60458) );
  NAND2xp5_ASAP7_75t_SL U63009 ( .A(n78009), .B(n61043), .Y(n60320) );
  NAND2xp5_ASAP7_75t_SL U63010 ( .A(n77841), .B(n60458), .Y(n61046) );
  NAND2xp5_ASAP7_75t_SL U63011 ( .A(n77229), .B(n77228), .Y(
        or1200_cpu_or1200_except_n1717) );
  NAND2xp5_ASAP7_75t_SL U63012 ( .A(n62313), .B(n60774), .Y(n62077) );
  NAND2xp5_ASAP7_75t_SL U63013 ( .A(n69281), .B(n69288), .Y(n69161) );
  OAI21xp5_ASAP7_75t_SL U63014 ( .A1(n69127), .A2(n69126), .B(n69125), .Y(
        n69288) );
  INVx1_ASAP7_75t_SL U63015 ( .A(n59388), .Y(n69114) );
  INVx2_ASAP7_75t_SL U63016 ( .A(n59634), .Y(n59636) );
  AOI22xp5_ASAP7_75t_SL U63017 ( .A1(n59634), .A2(n68594), .B1(n75073), .B2(
        n75048), .Y(n68601) );
  NAND2xp5_ASAP7_75t_SL U63018 ( .A(n60153), .B(n57100), .Y(n4118) );
  NOR2x1p5_ASAP7_75t_SL U63019 ( .A(n58870), .B(n53608), .Y(n69160) );
  AOI22xp5_ASAP7_75t_SL U63020 ( .A1(n75133), .A2(n75132), .B1(n75131), .B2(
        n75130), .Y(n75658) );
  AOI21xp5_ASAP7_75t_SL U63021 ( .A1(n76916), .A2(n76899), .B(n76898), .Y(
        n76914) );
  NOR2x1_ASAP7_75t_SL U63022 ( .A(n807), .B(n60114), .Y(n60142) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63023 ( .A1(n771), .A2(n59703), .B(n60173), .C(
        n76821), .Y(n60035) );
  INVx1_ASAP7_75t_SL U63024 ( .A(n76882), .Y(n68746) );
  NAND2xp5_ASAP7_75t_SL U63025 ( .A(n63912), .B(n75387), .Y(n62218) );
  NAND2xp5_ASAP7_75t_SL U63026 ( .A(n62404), .B(n62403), .Y(n62407) );
  NAND2xp5_ASAP7_75t_SL U63027 ( .A(n67210), .B(n59388), .Y(n59392) );
  INVx1_ASAP7_75t_SL U63028 ( .A(n61753), .Y(n76729) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63029 ( .A1(n61753), .A2(n60568), .B(n77582), 
        .C(n60567), .Y(n60569) );
  NAND2xp5_ASAP7_75t_SL U63030 ( .A(n73406), .B(n73405), .Y(n73407) );
  NAND2xp5_ASAP7_75t_SL U63031 ( .A(n73358), .B(n73357), .Y(n73405) );
  OAI22xp5_ASAP7_75t_SL U63032 ( .A1(dbg_stb_i), .A2(n59935), .B1(dbg_adr_i[6]), .B2(n78439), .Y(n60572) );
  NAND2xp5_ASAP7_75t_SL U63033 ( .A(n73586), .B(n73567), .Y(n3275) );
  INVx3_ASAP7_75t_SL U63034 ( .A(n59586), .Y(n59584) );
  INVx1_ASAP7_75t_SL U63035 ( .A(n64351), .Y(n63817) );
  NAND2xp5_ASAP7_75t_SL U63036 ( .A(n64351), .B(n64350), .Y(n64043) );
  O2A1O1Ixp5_ASAP7_75t_SL U63037 ( .A1(n65106), .A2(n65105), .B(n65103), .C(
        n65104), .Y(n75790) );
  INVx1_ASAP7_75t_SL U63038 ( .A(n64728), .Y(n65106) );
  NOR2xp33_ASAP7_75t_SL U63039 ( .A(n68664), .B(n69117), .Y(n58831) );
  INVx1_ASAP7_75t_SL U63040 ( .A(n76542), .Y(n75768) );
  INVx1_ASAP7_75t_SL U63041 ( .A(n60454), .Y(n77407) );
  NAND2xp5_ASAP7_75t_SL U63042 ( .A(n70118), .B(n70077), .Y(n69944) );
  AOI21xp5_ASAP7_75t_SL U63043 ( .A1(n69505), .A2(n70118), .B(n69462), .Y(
        n69573) );
  NAND2xp5_ASAP7_75t_SL U63044 ( .A(n77115), .B(n77114), .Y(n77113) );
  OAI21xp5_ASAP7_75t_SL U63045 ( .A1(n67039), .A2(n66839), .B(n67043), .Y(
        n66905) );
  AOI21xp5_ASAP7_75t_SL U63046 ( .A1(n64187), .A2(n64196), .B(n61970), .Y(
        n64193) );
  OAI21xp5_ASAP7_75t_SL U63047 ( .A1(n64269), .A2(n64270), .B(n64271), .Y(
        n64187) );
  AND2x2_ASAP7_75t_SL U63048 ( .A(n59280), .B(n75085), .Y(n75464) );
  NAND2xp5_ASAP7_75t_SL U63049 ( .A(n71953), .B(n71561), .Y(n71551) );
  INVx1_ASAP7_75t_SL U63050 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), 
        .Y(n71953) );
  NAND2xp5_ASAP7_75t_SL U63051 ( .A(n71435), .B(n71616), .Y(n71619) );
  AOI21xp5_ASAP7_75t_SL U63052 ( .A1(n76320), .A2(n77031), .B(n62139), .Y(
        n77878) );
  OAI21xp5_ASAP7_75t_SL U63053 ( .A1(n75882), .A2(n62138), .B(n62137), .Y(
        n62139) );
  NOR2x1p5_ASAP7_75t_SL U63054 ( .A(n53608), .B(n58325), .Y(n75095) );
  AOI21xp5_ASAP7_75t_SL U63055 ( .A1(n68761), .A2(n68755), .B(n64988), .Y(
        n65071) );
  XNOR2x1_ASAP7_75t_SL U63056 ( .A(n58988), .B(n58987), .Y(n58317) );
  NOR2xp33_ASAP7_75t_SL U63057 ( .A(n74558), .B(n57474), .Y(n58318) );
  INVx1_ASAP7_75t_SL U63058 ( .A(n68736), .Y(n68727) );
  NAND2xp5_ASAP7_75t_SL U63059 ( .A(n74753), .B(n74934), .Y(n74808) );
  HB1xp67_ASAP7_75t_SL U63060 ( .A(n67734), .Y(n58319) );
  XNOR2xp5_ASAP7_75t_SL U63061 ( .A(n57051), .B(n66838), .Y(n58320) );
  NAND2xp5_ASAP7_75t_SL U63062 ( .A(n67306), .B(n67571), .Y(n67265) );
  NAND2xp5_ASAP7_75t_SL U63063 ( .A(n73202), .B(n73460), .Y(n73465) );
  OAI22xp5_ASAP7_75t_SL U63064 ( .A1(n63636), .A2(n57097), .B1(n63838), .B2(
        n57159), .Y(n63832) );
  OAI21xp5_ASAP7_75t_SL U63065 ( .A1(n75900), .A2(n59594), .B(n63635), .Y(
        n63838) );
  XNOR2xp5_ASAP7_75t_SL U63066 ( .A(n68312), .B(n68311), .Y(n68315) );
  INVx1_ASAP7_75t_SL U63067 ( .A(n67340), .Y(n59138) );
  NAND2xp5_ASAP7_75t_SL U63068 ( .A(n71026), .B(n71033), .Y(n71051) );
  INVx1_ASAP7_75t_SL U63069 ( .A(n68419), .Y(n67723) );
  NOR2xp33_ASAP7_75t_SL U63070 ( .A(n66671), .B(n66690), .Y(n58321) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63071 ( .A1(n59591), .A2(n66637), .B(n57186), 
        .C(n59548), .Y(n66639) );
  INVx1_ASAP7_75t_SL U63072 ( .A(n58957), .Y(n58322) );
  NAND2xp5_ASAP7_75t_SL U63073 ( .A(n59326), .B(n62600), .Y(n59325) );
  AOI31xp33_ASAP7_75t_SL U63074 ( .A1(n59613), .A2(n58761), .A3(n57025), .B(
        n58760), .Y(n58323) );
  A2O1A1Ixp33_ASAP7_75t_SL U63075 ( .A1(n56830), .A2(n67957), .B(n68214), .C(
        n67956), .Y(n58324) );
  O2A1O1Ixp5_ASAP7_75t_SL U63076 ( .A1(n67863), .A2(n59642), .B(n67862), .C(
        n58917), .Y(n58916) );
  INVx1_ASAP7_75t_SL U63077 ( .A(n75642), .Y(n59642) );
  XNOR2xp5_ASAP7_75t_SL U63078 ( .A(n67670), .B(n67671), .Y(n58396) );
  XNOR2x2_ASAP7_75t_SL U63079 ( .A(n68401), .B(n67563), .Y(n67670) );
  INVx1_ASAP7_75t_SL U63080 ( .A(n57269), .Y(n59063) );
  NAND2xp5_ASAP7_75t_SL U63081 ( .A(n58885), .B(n68809), .Y(n59207) );
  NAND2x1_ASAP7_75t_SL U63082 ( .A(n59344), .B(n68808), .Y(n68809) );
  NOR2x1_ASAP7_75t_SL U63083 ( .A(n64669), .B(n64670), .Y(n64708) );
  NAND2xp5_ASAP7_75t_SL U63084 ( .A(n66782), .B(n66781), .Y(n66785) );
  INVx1_ASAP7_75t_SL U63085 ( .A(n68724), .Y(n59403) );
  INVx1_ASAP7_75t_SL U63086 ( .A(n64055), .Y(n63868) );
  NAND2xp5_ASAP7_75t_SL U63087 ( .A(n59596), .B(n57104), .Y(n66624) );
  NAND2xp5_ASAP7_75t_SL U63088 ( .A(n58353), .B(n76430), .Y(n58909) );
  NAND2xp5_ASAP7_75t_SL U63089 ( .A(n67281), .B(n75032), .Y(n67283) );
  XNOR2x1_ASAP7_75t_SL U63090 ( .A(n67471), .B(n67285), .Y(n67485) );
  AOI22xp5_ASAP7_75t_SL U63091 ( .A1(n64535), .A2(n64534), .B1(n64533), .B2(
        n64532), .Y(n64604) );
  INVx1_ASAP7_75t_SL U63092 ( .A(n62858), .Y(n62810) );
  INVx1_ASAP7_75t_SL U63093 ( .A(n68279), .Y(n68281) );
  INVx1_ASAP7_75t_SL U63094 ( .A(n63137), .Y(n63100) );
  OAI21xp5_ASAP7_75t_SL U63095 ( .A1(n75947), .A2(n57176), .B(n67062), .Y(
        n66884) );
  XNOR2x2_ASAP7_75t_SL U63096 ( .A(n62777), .B(n62680), .Y(n62754) );
  INVx1_ASAP7_75t_SL U63097 ( .A(n57277), .Y(n68603) );
  AOI21xp5_ASAP7_75t_SL U63098 ( .A1(n57277), .A2(n59475), .B(n66357), .Y(
        n66358) );
  AOI21xp5_ASAP7_75t_SL U63099 ( .A1(n57277), .A2(n76049), .B(n66959), .Y(
        n59289) );
  XNOR2x1_ASAP7_75t_SL U63100 ( .A(n68295), .B(n68294), .Y(n68344) );
  NAND2xp5_ASAP7_75t_SL U63101 ( .A(n57260), .B(n67876), .Y(n67877) );
  OAI21xp5_ASAP7_75t_SL U63102 ( .A1(n70879), .A2(n70878), .B(n70877), .Y(
        n58326) );
  AOI21xp5_ASAP7_75t_SL U63103 ( .A1(n70876), .A2(n70875), .B(n70874), .Y(
        n70877) );
  INVx1_ASAP7_75t_SL U63104 ( .A(n67598), .Y(n62887) );
  MAJIxp5_ASAP7_75t_SL U63105 ( .A(n67070), .B(n67069), .C(n67068), .Y(n58327)
         );
  NAND2xp5_ASAP7_75t_SL U63106 ( .A(or1200_cpu_or1200_except_n586), .B(n2517), 
        .Y(n63752) );
  NOR2x1_ASAP7_75t_SL U63107 ( .A(n63129), .B(n64079), .Y(n63677) );
  NOR2x1_ASAP7_75t_SL U63108 ( .A(n62888), .B(n62889), .Y(n62893) );
  NAND2xp5_ASAP7_75t_SL U63109 ( .A(n62893), .B(n62885), .Y(n62899) );
  OAI22xp5_ASAP7_75t_SL U63110 ( .A1(n60331), .A2(n78006), .B1(n2705), .B2(
        n78009), .Y(n60438) );
  NAND2x1p5_ASAP7_75t_SL U63111 ( .A(n59252), .B(n59457), .Y(n58839) );
  OAI22xp5_ASAP7_75t_SL U63112 ( .A1(n59446), .A2(n58794), .B1(n67004), .B2(
        n59440), .Y(n67053) );
  AOI22xp5_ASAP7_75t_SL U63113 ( .A1(n57323), .A2(n67402), .B1(n67386), .B2(
        n67401), .Y(n67503) );
  INVx1_ASAP7_75t_SL U63114 ( .A(n68326), .Y(n59066) );
  INVx1_ASAP7_75t_SL U63115 ( .A(n68258), .Y(n65046) );
  INVx1_ASAP7_75t_SL U63116 ( .A(n68748), .Y(n58329) );
  INVx1_ASAP7_75t_SL U63117 ( .A(n68737), .Y(n68748) );
  NAND2xp5_ASAP7_75t_SL U63118 ( .A(n61399), .B(n61396), .Y(n60765) );
  INVx1_ASAP7_75t_SL U63119 ( .A(n64604), .Y(n64544) );
  INVx1_ASAP7_75t_SL U63120 ( .A(n63231), .Y(n63117) );
  XNOR2x1_ASAP7_75t_SL U63121 ( .A(n59013), .B(n68545), .Y(n69035) );
  OAI21xp5_ASAP7_75t_SL U63122 ( .A1(n1145), .A2(n75391), .B(n74979), .Y(n9257) );
  OAI21xp5_ASAP7_75t_SL U63123 ( .A1(n63010), .A2(n63009), .B(n63008), .Y(
        n63035) );
  NAND2xp5_ASAP7_75t_SL U63124 ( .A(n71295), .B(n71294), .Y(n71306) );
  AOI22xp5_ASAP7_75t_SL U63125 ( .A1(n66957), .A2(n57463), .B1(n67401), .B2(
        n66956), .Y(n68454) );
  AOI22xp5_ASAP7_75t_SL U63126 ( .A1(n75048), .A2(n66953), .B1(n59100), .B2(
        n66954), .Y(n68453) );
  AO22x1_ASAP7_75t_SL U63127 ( .A1(n71087), .A2(n71085), .B1(n70996), .B2(
        n71086), .Y(n58330) );
  NAND2xp5_ASAP7_75t_SL U63128 ( .A(n70935), .B(n70936), .Y(n58331) );
  XNOR2xp5_ASAP7_75t_SL U63129 ( .A(n67295), .B(n58661), .Y(n67784) );
  INVx1_ASAP7_75t_SL U63130 ( .A(n67698), .Y(n58332) );
  NOR2x1_ASAP7_75t_SL U63131 ( .A(n66556), .B(n66555), .Y(n66591) );
  NAND2xp5_ASAP7_75t_SL U63132 ( .A(n69804), .B(n69803), .Y(n69835) );
  OAI21xp5_ASAP7_75t_SL U63133 ( .A1(n69802), .A2(n69801), .B(n69800), .Y(
        n69803) );
  NAND2xp5_ASAP7_75t_SL U63134 ( .A(n71203), .B(n71270), .Y(n71198) );
  INVx1_ASAP7_75t_SL U63135 ( .A(n67017), .Y(n63097) );
  HB1xp67_ASAP7_75t_SL U63136 ( .A(n68034), .Y(n58334) );
  XOR2xp5_ASAP7_75t_SL U63137 ( .A(n68428), .B(n68429), .Y(n68426) );
  AOI21xp5_ASAP7_75t_SL U63138 ( .A1(n68621), .A2(n68622), .B(n66607), .Y(
        n68627) );
  NOR2x1_ASAP7_75t_SL U63139 ( .A(n68634), .B(n68633), .Y(n69300) );
  AOI21xp5_ASAP7_75t_SL U63140 ( .A1(n67434), .A2(n57410), .B(n66470), .Y(
        n67126) );
  NAND2xp5_ASAP7_75t_SL U63141 ( .A(n66696), .B(n75032), .Y(n66698) );
  XNOR2xp5_ASAP7_75t_SL U63142 ( .A(n70525), .B(n70101), .Y(n70102) );
  INVx1_ASAP7_75t_SL U63143 ( .A(n68678), .Y(n69225) );
  INVx1_ASAP7_75t_SL U63144 ( .A(n59279), .Y(n67254) );
  NAND2xp5_ASAP7_75t_SL U63145 ( .A(n57376), .B(n68666), .Y(n68675) );
  XNOR2xp5_ASAP7_75t_SL U63146 ( .A(n66592), .B(n66593), .Y(n66605) );
  OAI21xp5_ASAP7_75t_SL U63147 ( .A1(n73952), .A2(n73951), .B(n75813), .Y(
        n76266) );
  NAND2xp5_ASAP7_75t_SL U63148 ( .A(n73951), .B(n73952), .Y(n75813) );
  OAI21xp5_ASAP7_75t_SL U63149 ( .A1(n66596), .A2(n66597), .B(n66343), .Y(
        n66593) );
  OAI21xp5_ASAP7_75t_SL U63150 ( .A1(n59630), .A2(n73159), .B(n73155), .Y(
        n73457) );
  NAND2xp5_ASAP7_75t_SL U63151 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[9]), .B(
        n59630), .Y(n73155) );
  NAND2xp5_ASAP7_75t_SL U63152 ( .A(n73289), .B(n73409), .Y(n73291) );
  INVx1_ASAP7_75t_SL U63153 ( .A(n66691), .Y(n66690) );
  NOR2x1p5_ASAP7_75t_SL U63154 ( .A(n68711), .B(n75277), .Y(n74557) );
  NOR2x1_ASAP7_75t_SL U63155 ( .A(n66203), .B(n74900), .Y(n74846) );
  NAND2xp5_ASAP7_75t_SL U63156 ( .A(n76956), .B(n74218), .Y(n58820) );
  OAI22xp5_ASAP7_75t_SL U63157 ( .A1(n59537), .A2(n66271), .B1(n63251), .B2(
        n63250), .Y(n59115) );
  NAND2x1_ASAP7_75t_SL U63158 ( .A(n64034), .B(n67586), .Y(n64897) );
  INVx1_ASAP7_75t_SL U63159 ( .A(n64053), .Y(n63866) );
  XOR2xp5_ASAP7_75t_SL U63160 ( .A(n67697), .B(n58335), .Y(n67667) );
  INVx1_ASAP7_75t_SL U63161 ( .A(n59243), .Y(n68961) );
  NOR2x1_ASAP7_75t_SL U63162 ( .A(or1200_cpu_or1200_mult_mac_n12), .B(n76171), 
        .Y(n75959) );
  OAI21xp5_ASAP7_75t_SL U63163 ( .A1(n75951), .A2(n53471), .B(n75950), .Y(
        n75952) );
  AOI21xp5_ASAP7_75t_SL U63164 ( .A1(n76171), .A2(
        or1200_cpu_or1200_mult_mac_n12), .B(n57336), .Y(n75960) );
  NAND2xp5_ASAP7_75t_SL U63165 ( .A(n59666), .B(n76181), .Y(n75970) );
  NAND2xp5_ASAP7_75t_SL U63166 ( .A(n75969), .B(n75970), .Y(n76185) );
  INVx1_ASAP7_75t_SL U63167 ( .A(n68180), .Y(n68181) );
  NAND2xp5_ASAP7_75t_SL U63168 ( .A(n59316), .B(n59315), .Y(n68180) );
  XNOR2x1_ASAP7_75t_SL U63169 ( .A(n68182), .B(n68181), .Y(n68183) );
  OAI22xp5_ASAP7_75t_SL U63170 ( .A1(n67001), .A2(n59491), .B1(n67000), .B2(
        n59612), .Y(n67055) );
  INVx1_ASAP7_75t_SL U63171 ( .A(n67170), .Y(n67172) );
  INVx1_ASAP7_75t_SL U63172 ( .A(n75077), .Y(n75034) );
  INVx2_ASAP7_75t_SL U63173 ( .A(n69008), .Y(n59382) );
  INVx2_ASAP7_75t_SL U63174 ( .A(n59542), .Y(n62604) );
  NOR2x1_ASAP7_75t_SL U63175 ( .A(n77278), .B(n63174), .Y(n62606) );
  NAND2xp5_ASAP7_75t_SL U63176 ( .A(n77338), .B(n77307), .Y(n77500) );
  INVx1_ASAP7_75t_SL U63177 ( .A(n60456), .Y(n61044) );
  NOR2x1_ASAP7_75t_SL U63178 ( .A(n60324), .B(n77840), .Y(n60456) );
  XNOR2x1_ASAP7_75t_SL U63179 ( .A(n67780), .B(n67781), .Y(n59082) );
  INVx1_ASAP7_75t_SL U63180 ( .A(n67778), .Y(n67781) );
  NAND2xp5_ASAP7_75t_SL U63181 ( .A(n1770), .B(n1686), .Y(n59106) );
  INVx1_ASAP7_75t_SL U63182 ( .A(n68389), .Y(n59030) );
  NAND2xp5_ASAP7_75t_SL U63183 ( .A(n67707), .B(n59293), .Y(n68389) );
  INVx1_ASAP7_75t_SL U63184 ( .A(n58819), .Y(n67243) );
  NAND2xp5_ASAP7_75t_SL U63185 ( .A(n75899), .B(n66803), .Y(n66632) );
  INVx1_ASAP7_75t_SL U63186 ( .A(n67560), .Y(n66803) );
  NOR2x1_ASAP7_75t_SL U63187 ( .A(n69226), .B(n68628), .Y(n68650) );
  OAI21xp5_ASAP7_75t_SL U63188 ( .A1(n67569), .A2(n59642), .B(n66916), .Y(
        n66962) );
  INVx1_ASAP7_75t_SL U63189 ( .A(n67270), .Y(n67226) );
  INVx1_ASAP7_75t_SL U63190 ( .A(n68462), .Y(n59172) );
  NAND2xp5_ASAP7_75t_SL U63191 ( .A(n69065), .B(n69068), .Y(n68831) );
  OAI21xp5_ASAP7_75t_SL U63192 ( .A1(n68819), .A2(n68818), .B(n68817), .Y(
        n69068) );
  AOI21xp5_ASAP7_75t_SL U63193 ( .A1(n68993), .A2(n69051), .B(n69058), .Y(
        n69017) );
  OAI21xp5_ASAP7_75t_SL U63194 ( .A1(n70592), .A2(n70591), .B(n70601), .Y(
        n70594) );
  OAI21xp5_ASAP7_75t_SL U63195 ( .A1(n70585), .A2(n70608), .B(n70584), .Y(
        n70592) );
  INVx11_ASAP7_75t_SL U63196 ( .A(n58402), .Y(n59617) );
  NAND2xp5_ASAP7_75t_SL U63197 ( .A(n59616), .B(n76049), .Y(n64960) );
  INVx3_ASAP7_75t_SL U63198 ( .A(n59646), .Y(n59645) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63199 ( .A1(n59577), .A2(n59645), .B(n64231), 
        .C(n61507), .Y(n60937) );
  AOI21xp5_ASAP7_75t_SL U63200 ( .A1(n76352), .A2(n59645), .B(n61183), .Y(
        n75701) );
  INVx1_ASAP7_75t_SL U63201 ( .A(n67198), .Y(n67201) );
  NOR2x1_ASAP7_75t_SL U63202 ( .A(n64518), .B(n64517), .Y(n64579) );
  INVx1_ASAP7_75t_SL U63203 ( .A(n59281), .Y(n58338) );
  XNOR2x1_ASAP7_75t_SL U63204 ( .A(n58394), .B(n64909), .Y(n64591) );
  INVx1_ASAP7_75t_SL U63205 ( .A(n68487), .Y(n68531) );
  INVx1_ASAP7_75t_SL U63206 ( .A(n68698), .Y(n58957) );
  OAI21xp5_ASAP7_75t_SL U63207 ( .A1(n58490), .A2(n67913), .B(n67912), .Y(
        n59133) );
  NAND2xp5_ASAP7_75t_SL U63208 ( .A(n57180), .B(n75962), .Y(n68092) );
  NAND2xp5_ASAP7_75t_SL U63209 ( .A(n65256), .B(n65255), .Y(n65298) );
  NOR2x1_ASAP7_75t_SL U63210 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_14_), .B(n65250), .Y(
        n65255) );
  NOR2x1_ASAP7_75t_SL U63211 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_20_), .B(n65344), .Y(
        n65353) );
  AO21x2_ASAP7_75t_SL U63212 ( .A1(n60303), .A2(n62150), .B(n60302), .Y(n77459) );
  NAND2xp5_ASAP7_75t_SL U63213 ( .A(n57160), .B(n76817), .Y(n77249) );
  INVx1_ASAP7_75t_SL U63214 ( .A(n64018), .Y(n64019) );
  INVx8_ASAP7_75t_SL U63215 ( .A(n59709), .Y(n59708) );
  AOI21x1_ASAP7_75t_SL U63216 ( .A1(n58882), .A2(n59709), .B(n67860), .Y(
        n59513) );
  AOI21x1_ASAP7_75t_SL U63217 ( .A1(n58882), .A2(n59709), .B(n67860), .Y(
        n59512) );
  INVx1_ASAP7_75t_SL U63218 ( .A(n68245), .Y(n68247) );
  XOR2x2_ASAP7_75t_SL U63219 ( .A(n68055), .B(n59176), .Y(n68059) );
  OAI21xp5_ASAP7_75t_SL U63220 ( .A1(n62977), .A2(n63144), .B(n57362), .Y(
        n62978) );
  INVx1_ASAP7_75t_SL U63221 ( .A(n66475), .Y(n66477) );
  INVx1_ASAP7_75t_SL U63222 ( .A(n64445), .Y(n63824) );
  AOI22xp5_ASAP7_75t_SL U63223 ( .A1(n71209), .A2(n71115), .B1(n71245), .B2(
        n71172), .Y(n71262) );
  OAI22xp5_ASAP7_75t_SL U63224 ( .A1(n57115), .A2(n70786), .B1(n70776), .B2(
        n59524), .Y(n71115) );
  XOR2xp5_ASAP7_75t_SL U63225 ( .A(n66981), .B(n58340), .Y(n67212) );
  INVx1_ASAP7_75t_SL U63226 ( .A(n64581), .Y(n64458) );
  INVx1_ASAP7_75t_SL U63227 ( .A(n67918), .Y(n67231) );
  NOR2x1_ASAP7_75t_SL U63228 ( .A(n58432), .B(n59594), .Y(n67918) );
  INVx1_ASAP7_75t_SL U63229 ( .A(n70758), .Y(n70725) );
  XOR2x2_ASAP7_75t_SL U63230 ( .A(n68056), .B(n68057), .Y(n68058) );
  OAI21xp5_ASAP7_75t_SL U63231 ( .A1(n69327), .A2(n69326), .B(n69325), .Y(
        n75130) );
  NAND2x1p5_ASAP7_75t_SL U63232 ( .A(n58202), .B(n67607), .Y(n67237) );
  XNOR2x2_ASAP7_75t_SL U63233 ( .A(n68259), .B(n65046), .Y(n65047) );
  NAND2xp5_ASAP7_75t_SL U63234 ( .A(n67923), .B(n67446), .Y(n67449) );
  HB1xp67_ASAP7_75t_SL U63235 ( .A(n67761), .Y(n58346) );
  NAND2x1_ASAP7_75t_SL U63236 ( .A(n68575), .B(n68574), .Y(n59243) );
  OAI31xp33_ASAP7_75t_SL U63237 ( .A1(n76269), .A2(n76268), .A3(n73953), .B(
        n64801), .Y(n64804) );
  AOI22xp5_ASAP7_75t_SL U63238 ( .A1(n59100), .A2(n67454), .B1(n67453), .B2(
        n75048), .Y(n67500) );
  AOI21xp5_ASAP7_75t_SL U63239 ( .A1(n59637), .A2(n67343), .B(n67286), .Y(
        n67453) );
  INVx1_ASAP7_75t_SL U63240 ( .A(n66909), .Y(n59085) );
  MAJx2_ASAP7_75t_SL U63241 ( .A(n68520), .B(n58388), .C(n68518), .Y(n58347)
         );
  OAI21xp5_ASAP7_75t_SL U63242 ( .A1(n67620), .A2(n58968), .B(n57033), .Y(
        n67653) );
  INVx1_ASAP7_75t_SL U63243 ( .A(n59596), .Y(n59206) );
  NOR2x1_ASAP7_75t_SL U63244 ( .A(n64350), .B(n64351), .Y(n58735) );
  INVx1_ASAP7_75t_SL U63245 ( .A(n67659), .Y(n58703) );
  OAI22xp5_ASAP7_75t_SL U63246 ( .A1(n57115), .A2(n70910), .B1(n70893), .B2(
        n59524), .Y(n71171) );
  NAND2xp5_ASAP7_75t_SL U63247 ( .A(n71052), .B(n71053), .Y(n71056) );
  OAI21xp5_ASAP7_75t_SL U63248 ( .A1(n62699), .A2(n57360), .B(n62698), .Y(
        n62720) );
  NAND2xp5_ASAP7_75t_SL U63249 ( .A(n60452), .B(n60453), .Y(n77843) );
  NAND2xp5_ASAP7_75t_SL U63250 ( .A(n59657), .B(n59605), .Y(n62767) );
  OA21x2_ASAP7_75t_SL U63251 ( .A1(n63070), .A2(n57159), .B(n63069), .Y(n58350) );
  NAND2x2_ASAP7_75t_SL U63252 ( .A(n58202), .B(n67230), .Y(n68102) );
  INVx1_ASAP7_75t_SL U63253 ( .A(n64964), .Y(n64629) );
  INVx1_ASAP7_75t_SL U63254 ( .A(n66307), .Y(n66312) );
  OAI22xp5_ASAP7_75t_SL U63255 ( .A1(n66828), .A2(n66829), .B1(n57508), .B2(
        n66884), .Y(n66848) );
  XNOR2xp5_ASAP7_75t_SL U63256 ( .A(n68462), .B(n68461), .Y(n68463) );
  INVx1_ASAP7_75t_SL U63257 ( .A(n63041), .Y(n63036) );
  OAI22xp5_ASAP7_75t_SL U63258 ( .A1(n66464), .A2(n59491), .B1(n66397), .B2(
        n59612), .Y(n66493) );
  NAND2xp5_ASAP7_75t_SL U63259 ( .A(n70745), .B(n70744), .Y(n70752) );
  XNOR2x1_ASAP7_75t_SL U63260 ( .A(n58366), .B(n67694), .Y(n59081) );
  INVx1_ASAP7_75t_SL U63261 ( .A(n66898), .Y(n66837) );
  XNOR2xp5_ASAP7_75t_SL U63262 ( .A(n59660), .B(n57109), .Y(n65053) );
  XNOR2x1_ASAP7_75t_SL U63263 ( .A(n68212), .B(n68211), .Y(n68298) );
  NAND2x1p5_ASAP7_75t_SL U63264 ( .A(n58347), .B(n68541), .Y(n69029) );
  INVx1_ASAP7_75t_SL U63265 ( .A(n66560), .Y(n68604) );
  OAI22xp5_ASAP7_75t_SL U63266 ( .A1(n68119), .A2(n66560), .B1(n66561), .B2(
        n59116), .Y(n66590) );
  XNOR2x2_ASAP7_75t_SL U63267 ( .A(n57078), .B(n53275), .Y(n66560) );
  OAI21xp5_ASAP7_75t_SL U63268 ( .A1(n75947), .A2(n57172), .B(n66650), .Y(
        n66767) );
  NAND2xp5_ASAP7_75t_SL U63269 ( .A(n76067), .B(n76059), .Y(n76076) );
  NAND2xp5_ASAP7_75t_SL U63270 ( .A(n76045), .B(n59510), .Y(n76059) );
  OAI21x1_ASAP7_75t_SL U63271 ( .A1(n68094), .A2(n64486), .B(n64485), .Y(
        n64566) );
  NAND2xp5_ASAP7_75t_SL U63272 ( .A(n64480), .B(n64479), .Y(n64486) );
  XNOR2x1_ASAP7_75t_SL U63273 ( .A(n58317), .B(n58986), .Y(n68537) );
  XNOR2x1_ASAP7_75t_SL U63274 ( .A(n68514), .B(n68515), .Y(n58986) );
  NAND2xp5_ASAP7_75t_SL U63275 ( .A(n59499), .B(n76256), .Y(n61988) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63276 ( .A1(n59656), .A2(n57827), .B(n67441), 
        .C(n59119), .Y(n59118) );
  AND2x4_ASAP7_75t_SL U63277 ( .A(n78327), .B(n66260), .Y(n58353) );
  HB1xp67_ASAP7_75t_SL U63278 ( .A(n68047), .Y(n58354) );
  INVx1_ASAP7_75t_SL U63279 ( .A(n68500), .Y(n68504) );
  NAND2xp5_ASAP7_75t_SL U63280 ( .A(n78207), .B(n4106), .Y(icqmem_adr_qmem[26]) );
  INVx1_ASAP7_75t_SL U63281 ( .A(n77398), .Y(n59156) );
  AOI211xp5_ASAP7_75t_SL U63282 ( .A1(iwb_dat_i[22]), .A2(n77373), .B(n58540), 
        .C(n60409), .Y(n2087) );
  OAI21xp5_ASAP7_75t_SL U63283 ( .A1(n71229), .A2(n70985), .B(n70984), .Y(
        n71146) );
  XNOR2x1_ASAP7_75t_SL U63284 ( .A(n67177), .B(n67176), .Y(n67190) );
  INVx1_ASAP7_75t_SL U63285 ( .A(n67157), .Y(n67177) );
  INVx1_ASAP7_75t_SL U63286 ( .A(n66775), .Y(n66653) );
  INVx1_ASAP7_75t_SL U63287 ( .A(n76661), .Y(n77218) );
  NAND2xp5_ASAP7_75t_SL U63288 ( .A(n77048), .B(n77163), .Y(n76661) );
  NAND2xp5_ASAP7_75t_SL U63289 ( .A(n77732), .B(n58433), .Y(n66296) );
  XOR2xp5_ASAP7_75t_SL U63290 ( .A(n68321), .B(n68320), .Y(n68311) );
  AOI21xp5_ASAP7_75t_SL U63291 ( .A1(n68380), .A2(n75901), .B(n65015), .Y(
        n59004) );
  NAND2xp5_ASAP7_75t_SL U63292 ( .A(n59534), .B(n1626), .Y(n61806) );
  NAND2xp5_ASAP7_75t_SL U63293 ( .A(n75670), .B(n75669), .Y(
        or1200_cpu_or1200_mult_mac_n1594) );
  NOR2x1_ASAP7_75t_SL U63294 ( .A(n58696), .B(n59596), .Y(n66421) );
  INVx1_ASAP7_75t_SL U63295 ( .A(n64943), .Y(n64630) );
  NAND2x1p5_ASAP7_75t_SL U63296 ( .A(n59269), .B(n59268), .Y(n67401) );
  OAI21xp5_ASAP7_75t_SL U63297 ( .A1(n57213), .A2(n57465), .B(n64026), .Y(
        n63634) );
  OAI21x1_ASAP7_75t_SL U63298 ( .A1(n75893), .A2(n66265), .B(n66264), .Y(
        n59634) );
  XNOR2x1_ASAP7_75t_SL U63299 ( .A(n66707), .B(n66706), .Y(n66840) );
  INVx1_ASAP7_75t_SL U63300 ( .A(n62935), .Y(n62838) );
  NAND2xp5_ASAP7_75t_SL U63301 ( .A(n59657), .B(n59171), .Y(n62935) );
  NAND2xp5_ASAP7_75t_SL U63302 ( .A(n70730), .B(n70731), .Y(n70715) );
  NAND2xp5_ASAP7_75t_SL U63303 ( .A(n70714), .B(n70713), .Y(n70731) );
  NAND2xp5_ASAP7_75t_SL U63304 ( .A(n67947), .B(n59620), .Y(n58857) );
  NAND2xp5_ASAP7_75t_SL U63305 ( .A(n68626), .B(n68625), .Y(n68687) );
  NAND2xp5_ASAP7_75t_SL U63306 ( .A(n70889), .B(n70888), .Y(n70908) );
  OAI22xp5_ASAP7_75t_SL U63307 ( .A1(n66465), .A2(n67627), .B1(n59612), .B2(
        n66464), .Y(n66478) );
  INVx2_ASAP7_75t_SL U63308 ( .A(n67464), .Y(n67627) );
  INVx1_ASAP7_75t_SL U63309 ( .A(n57335), .Y(n68925) );
  AOI21x1_ASAP7_75t_SL U63310 ( .A1(n68917), .A2(n68915), .B(n58686), .Y(
        n69004) );
  NAND2xp5_ASAP7_75t_SL U63311 ( .A(n68208), .B(n68210), .Y(n68200) );
  NOR2x1_ASAP7_75t_SL U63312 ( .A(n59598), .B(n66882), .Y(n66656) );
  NOR3x1_ASAP7_75t_SL U63313 ( .A(n59477), .B(n57348), .C(n59467), .Y(n63169)
         );
  INVx1_ASAP7_75t_SL U63314 ( .A(n68524), .Y(n66943) );
  INVx1_ASAP7_75t_SL U63315 ( .A(n68505), .Y(n66942) );
  NAND2xp5_ASAP7_75t_SL U63316 ( .A(n66288), .B(n58487), .Y(n58950) );
  NOR2x2_ASAP7_75t_SL U63317 ( .A(n75468), .B(n66322), .Y(n75048) );
  NAND2xp5_ASAP7_75t_SL U63318 ( .A(n59638), .B(n75468), .Y(n75046) );
  OA21x2_ASAP7_75t_SL U63319 ( .A1(n57352), .A2(n62687), .B(n62686), .Y(n58356) );
  INVx1_ASAP7_75t_SL U63320 ( .A(n58889), .Y(n62687) );
  NAND2x1_ASAP7_75t_SL U63321 ( .A(n57352), .B(n62685), .Y(n62686) );
  INVx1_ASAP7_75t_SL U63322 ( .A(n64534), .Y(n64375) );
  XNOR2x2_ASAP7_75t_SL U63323 ( .A(n64524), .B(n64525), .Y(n64377) );
  INVx1_ASAP7_75t_SL U63324 ( .A(n63674), .Y(n58938) );
  NAND2xp5_ASAP7_75t_SL U63325 ( .A(n63569), .B(n57120), .Y(n60749) );
  NAND2xp5_ASAP7_75t_SL U63326 ( .A(n61201), .B(n60748), .Y(n63569) );
  NOR2x1_ASAP7_75t_SL U63327 ( .A(n61620), .B(n61619), .Y(n62308) );
  NAND2xp5_ASAP7_75t_SL U63328 ( .A(n70815), .B(n70814), .Y(n70835) );
  AOI21xp5_ASAP7_75t_SL U63329 ( .A1(n58326), .A2(n71035), .B(n71034), .Y(
        n71036) );
  INVx1_ASAP7_75t_SL U63330 ( .A(n68721), .Y(n59426) );
  AOI211xp5_ASAP7_75t_SL U63331 ( .A1(n62619), .A2(n59020), .B(n64358), .C(
        n62618), .Y(n68016) );
  OR2x2_ASAP7_75t_SL U63332 ( .A(n63683), .B(n63684), .Y(n65102) );
  NAND2xp5_ASAP7_75t_SL U63333 ( .A(n70990), .B(n70991), .Y(n71023) );
  AOI22xp5_ASAP7_75t_SL U63334 ( .A1(n58746), .A2(n66473), .B1(n67095), .B2(
        n67096), .Y(n67123) );
  AOI21xp5_ASAP7_75t_SL U63335 ( .A1(n67096), .A2(n64616), .B(n64474), .Y(
        n64477) );
  OAI22xp5_ASAP7_75t_SL U63336 ( .A1(n62751), .A2(n59460), .B1(n63080), .B2(
        n64920), .Y(n63056) );
  NAND2xp5_ASAP7_75t_SL U63337 ( .A(n59455), .B(n75947), .Y(n66650) );
  OAI21xp5_ASAP7_75t_SL U63338 ( .A1(n64880), .A2(n64879), .B(n64878), .Y(
        n64881) );
  XNOR2x1_ASAP7_75t_SL U63339 ( .A(n59188), .B(n58452), .Y(n68335) );
  XNOR2x2_ASAP7_75t_SL U63340 ( .A(n58754), .B(n68186), .Y(n59188) );
  INVx1_ASAP7_75t_SL U63341 ( .A(n61037), .Y(n77840) );
  NAND2xp5_ASAP7_75t_SL U63342 ( .A(n71058), .B(n71154), .Y(n71063) );
  INVx1_ASAP7_75t_SL U63343 ( .A(n68523), .Y(n58357) );
  INVx1_ASAP7_75t_SL U63344 ( .A(n67045), .Y(n67048) );
  INVx1_ASAP7_75t_SL U63345 ( .A(n71087), .Y(n71076) );
  NOR2x1_ASAP7_75t_SL U63346 ( .A(n73963), .B(n76662), .Y(n77217) );
  AOI21xp5_ASAP7_75t_SL U63347 ( .A1(n70978), .A2(n70977), .B(n70976), .Y(
        n71024) );
  INVx1_ASAP7_75t_SL U63348 ( .A(n63011), .Y(n62987) );
  INVx1_ASAP7_75t_SL U63349 ( .A(n63363), .Y(n63446) );
  INVx5_ASAP7_75t_SL U63350 ( .A(n59530), .Y(n74776) );
  NAND2xp5_ASAP7_75t_SL U63351 ( .A(n57078), .B(n57163), .Y(n66479) );
  INVx1_ASAP7_75t_SL U63352 ( .A(n66530), .Y(n66531) );
  AOI22xp5_ASAP7_75t_SL U63353 ( .A1(n59100), .A2(n67247), .B1(n75048), .B2(
        n67246), .Y(n67656) );
  NOR2x1_ASAP7_75t_SL U63354 ( .A(n68366), .B(n68365), .Y(n68459) );
  XNOR2x1_ASAP7_75t_SL U63355 ( .A(n68475), .B(n68474), .Y(n68514) );
  HB1xp67_ASAP7_75t_SL U63356 ( .A(n64594), .Y(n58359) );
  AOI22xp5_ASAP7_75t_SL U63357 ( .A1(n59635), .A2(n66542), .B1(n66550), .B2(
        n75048), .Y(n66585) );
  AO21x2_ASAP7_75t_SL U63358 ( .A1(n67901), .A2(n68158), .B(n67900), .Y(n59490) );
  OAI21xp5_ASAP7_75t_SL U63359 ( .A1(n67972), .A2(n59615), .B(n59506), .Y(
        n58777) );
  NAND2xp5_ASAP7_75t_SL U63360 ( .A(n60454), .B(n77455), .Y(n61038) );
  INVx1_ASAP7_75t_SL U63361 ( .A(n63090), .Y(n62764) );
  AOI21xp5_ASAP7_75t_SL U63362 ( .A1(n63090), .A2(n63089), .B(n63088), .Y(
        n63091) );
  XNOR2x2_ASAP7_75t_SL U63363 ( .A(n63078), .B(n62779), .Y(n63051) );
  INVx1_ASAP7_75t_SL U63364 ( .A(or1200_cpu_rf_rdb), .Y(n77455) );
  AOI22xp5_ASAP7_75t_SL U63365 ( .A1(n67251), .A2(n62848), .B1(n62879), .B2(
        n62847), .Y(n62870) );
  NOR2x1_ASAP7_75t_SL U63366 ( .A(n59065), .B(n67566), .Y(n59067) );
  OAI21xp5_ASAP7_75t_SL U63367 ( .A1(n67566), .A2(n59660), .B(n67565), .Y(
        n67687) );
  NAND2xp5_ASAP7_75t_SL U63368 ( .A(n65016), .B(n59004), .Y(n59003) );
  HB1xp67_ASAP7_75t_SL U63369 ( .A(n68339), .Y(n58360) );
  NAND2xp5_ASAP7_75t_SL U63370 ( .A(n57180), .B(n59664), .Y(n67859) );
  NAND2x1p5_ASAP7_75t_SL U63371 ( .A(n59057), .B(n67441), .Y(n67511) );
  OAI21xp5_ASAP7_75t_SL U63372 ( .A1(n58931), .A2(n58431), .B(n58937), .Y(
        n62741) );
  NAND2xp5_ASAP7_75t_SL U63373 ( .A(n58931), .B(n57274), .Y(n58937) );
  OAI21xp5_ASAP7_75t_SL U63374 ( .A1(n63075), .A2(n62773), .B(n63073), .Y(
        n62778) );
  NAND2xp5_ASAP7_75t_SL U63375 ( .A(n75125), .B(n75664), .Y(n75141) );
  OAI21xp5_ASAP7_75t_SL U63376 ( .A1(n75124), .A2(n75123), .B(n75122), .Y(
        n75664) );
  NAND2xp5_ASAP7_75t_SL U63377 ( .A(n64078), .B(n57120), .Y(n61933) );
  NAND2x1_ASAP7_75t_SL U63378 ( .A(n59018), .B(n59017), .Y(n64078) );
  BUFx3_ASAP7_75t_SL U63379 ( .A(n59660), .Y(n59381) );
  NAND2xp5_ASAP7_75t_SL U63380 ( .A(n77701), .B(n59589), .Y(n58647) );
  BUFx3_ASAP7_75t_SL U63381 ( .A(n66450), .Y(n59589) );
  AOI21xp5_ASAP7_75t_SL U63382 ( .A1(n67076), .A2(n67306), .B(n67075), .Y(
        n67133) );
  OAI21xp5_ASAP7_75t_SL U63383 ( .A1(n67074), .A2(n59651), .B(n67073), .Y(
        n67075) );
  HB1xp67_ASAP7_75t_SL U63384 ( .A(n58170), .Y(n58362) );
  AOI22xp5_ASAP7_75t_SL U63385 ( .A1(n57463), .A2(n66472), .B1(n66883), .B2(
        n53231), .Y(n67121) );
  NAND2xp5_ASAP7_75t_SL U63386 ( .A(n57108), .B(n58531), .Y(n59298) );
  NAND2xp5_ASAP7_75t_SL U63387 ( .A(n57108), .B(n64396), .Y(n64400) );
  NAND2xp5_ASAP7_75t_SL U63388 ( .A(n74363), .B(n74362), .Y(n74505) );
  NOR2x1_ASAP7_75t_SL U63389 ( .A(n74224), .B(n74739), .Y(n74362) );
  OAI21xp5_ASAP7_75t_SL U63390 ( .A1(n67844), .A2(n57158), .B(n59040), .Y(
        n58363) );
  NAND2xp5_ASAP7_75t_SL U63391 ( .A(n78262), .B(n4101), .Y(icqmem_adr_qmem[28]) );
  NAND2xp5_ASAP7_75t_SL U63392 ( .A(n66338), .B(n66337), .Y(n66554) );
  HB1xp67_ASAP7_75t_SL U63393 ( .A(n68433), .Y(n58364) );
  NAND2xp5_ASAP7_75t_SL U63394 ( .A(n64420), .B(n64419), .Y(n64448) );
  XNOR2xp5_ASAP7_75t_SL U63395 ( .A(n68059), .B(n68058), .Y(n68574) );
  INVx1_ASAP7_75t_SL U63396 ( .A(n63196), .Y(n58877) );
  NOR2x1_ASAP7_75t_SL U63397 ( .A(n53193), .B(n58313), .Y(n68749) );
  OAI21xp5_ASAP7_75t_SL U63398 ( .A1(n76162), .A2(n75940), .B(
        or1200_cpu_or1200_mult_mac_n14), .Y(n75946) );
  NAND2xp5_ASAP7_75t_SL U63399 ( .A(n53505), .B(n68851), .Y(n68858) );
  NAND2xp5_ASAP7_75t_SL U63400 ( .A(n58931), .B(n67920), .Y(n58935) );
  OAI22xp5_ASAP7_75t_SL U63401 ( .A1(n57115), .A2(n70850), .B1(n70843), .B2(
        n59524), .Y(n71172) );
  OAI22xp5_ASAP7_75t_SL U63402 ( .A1(n75157), .A2(n75156), .B1(n2054), .B2(
        or1200_cpu_or1200_except_n655), .Y(n75159) );
  INVx1_ASAP7_75t_SL U63403 ( .A(n72490), .Y(n72503) );
  NOR2x1_ASAP7_75t_SL U63404 ( .A(n73581), .B(n73562), .Y(n73661) );
  NAND2xp5_ASAP7_75t_SL U63405 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[6]), .B(n73585), 
        .Y(n73562) );
  OAI21xp5_ASAP7_75t_SL U63406 ( .A1(n68079), .A2(n58509), .B(n59307), .Y(
        n62970) );
  NAND2xp5_ASAP7_75t_SL U63407 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[20]), .B(
        n73123), .Y(n73089) );
  OAI21xp5_ASAP7_75t_SL U63408 ( .A1(n73279), .A2(n73154), .B(n73153), .Y(
        n73440) );
  NOR2x1_ASAP7_75t_SL U63409 ( .A(n61438), .B(n64116), .Y(n62682) );
  NAND2xp5_ASAP7_75t_SL U63410 ( .A(n59513), .B(n67713), .Y(n58675) );
  NOR2x1_ASAP7_75t_SL U63411 ( .A(n59598), .B(n59436), .Y(n59065) );
  INVx2_ASAP7_75t_SL U63412 ( .A(n63825), .Y(n64032) );
  INVx1_ASAP7_75t_SL U63413 ( .A(n64639), .Y(n59088) );
  XNOR2x1_ASAP7_75t_SL U63414 ( .A(n64496), .B(n64495), .Y(n64552) );
  INVx1_ASAP7_75t_SL U63415 ( .A(n64555), .Y(n64496) );
  AOI31xp33_ASAP7_75t_SL U63416 ( .A1(n67551), .A2(n67549), .A3(n67550), .B(
        n67548), .Y(n58365) );
  NAND2xp5_ASAP7_75t_SL U63417 ( .A(n62302), .B(n62303), .Y(n62397) );
  NAND2xp5_ASAP7_75t_SL U63418 ( .A(n57100), .B(n53439), .Y(n76817) );
  NAND2xp5_ASAP7_75t_SL U63419 ( .A(n68086), .B(n66712), .Y(n66717) );
  XNOR2xp5_ASAP7_75t_SL U63420 ( .A(n65068), .B(n57290), .Y(n58367) );
  INVx1_ASAP7_75t_SL U63421 ( .A(n66985), .Y(n66903) );
  NAND2xp5_ASAP7_75t_SL U63422 ( .A(n59617), .B(n53258), .Y(n67084) );
  INVx2_ASAP7_75t_SL U63423 ( .A(n64355), .Y(n66241) );
  NAND2xp5_ASAP7_75t_SL U63424 ( .A(n57335), .B(n68899), .Y(n68923) );
  NAND2xp5_ASAP7_75t_SL U63425 ( .A(n62964), .B(n62963), .Y(n63008) );
  NOR2x1_ASAP7_75t_SL U63426 ( .A(n67028), .B(n67027), .Y(n67070) );
  NAND2x1_ASAP7_75t_SL U63427 ( .A(n67222), .B(n75112), .Y(n75096) );
  INVx1_ASAP7_75t_SL U63428 ( .A(n67503), .Y(n67506) );
  OAI21xp5_ASAP7_75t_SL U63429 ( .A1(n69160), .A2(n69159), .B(n69158), .Y(
        n52011) );
  INVx1_ASAP7_75t_SL U63430 ( .A(n62989), .Y(n62933) );
  XNOR2xp5_ASAP7_75t_SL U63431 ( .A(n67689), .B(n59068), .Y(n67572) );
  OAI22xp5_ASAP7_75t_SL U63432 ( .A1(n57494), .A2(n67570), .B1(n59440), .B2(
        n67571), .Y(n59068) );
  INVx1_ASAP7_75t_SL U63433 ( .A(n75906), .Y(n76071) );
  INVx1_ASAP7_75t_SL U63434 ( .A(n68469), .Y(n68470) );
  INVx1_ASAP7_75t_SL U63435 ( .A(n65014), .Y(n64941) );
  XNOR2xp5_ASAP7_75t_SL U63436 ( .A(n66704), .B(n66703), .Y(n66705) );
  INVx1_ASAP7_75t_SL U63437 ( .A(n66870), .Y(n66704) );
  OAI22xp5_ASAP7_75t_SL U63438 ( .A1(n67744), .A2(n67743), .B1(n57099), .B2(
        n67742), .Y(n68373) );
  NOR2x1_ASAP7_75t_SL U63439 ( .A(n67616), .B(n67617), .Y(n67378) );
  INVx1_ASAP7_75t_SL U63440 ( .A(n67009), .Y(n58964) );
  INVx1_ASAP7_75t_SL U63441 ( .A(n67108), .Y(n69141) );
  INVx1_ASAP7_75t_SL U63442 ( .A(n66700), .Y(n66786) );
  INVx1_ASAP7_75t_SL U63443 ( .A(n64049), .Y(n63831) );
  AOI22xp5_ASAP7_75t_SL U63444 ( .A1(n67609), .A2(n62655), .B1(n62654), .B2(
        n64607), .Y(n62777) );
  INVx1_ASAP7_75t_SL U63445 ( .A(n67777), .Y(n67782) );
  HB1xp67_ASAP7_75t_SL U63446 ( .A(n68232), .Y(n58369) );
  MAJIxp5_ASAP7_75t_SL U63447 ( .A(n67783), .B(n67325), .C(n67324), .Y(n58370)
         );
  NAND2xp5_ASAP7_75t_SL U63448 ( .A(n75652), .B(n75135), .Y(n75139) );
  NAND2xp5_ASAP7_75t_SL U63449 ( .A(n75134), .B(n75658), .Y(n75135) );
  NAND2xp5_ASAP7_75t_SL U63450 ( .A(n58999), .B(n68579), .Y(n68917) );
  NAND2xp5_ASAP7_75t_SL U63451 ( .A(n66345), .B(n66349), .Y(n66347) );
  INVx1_ASAP7_75t_SL U63452 ( .A(n59330), .Y(n58918) );
  INVx3_ASAP7_75t_SL U63453 ( .A(n59581), .Y(n78002) );
  OAI21xp5_ASAP7_75t_SL U63454 ( .A1(n78002), .A2(n57347), .B(n62629), .Y(
        n62630) );
  NAND2xp5_ASAP7_75t_SL U63455 ( .A(n59571), .B(n78002), .Y(n73981) );
  OAI22xp5_ASAP7_75t_SL U63456 ( .A1(n57115), .A2(n70767), .B1(n70759), .B2(
        n59524), .Y(n71085) );
  NAND2xp5_ASAP7_75t_SL U63457 ( .A(n64602), .B(n64601), .Y(n64603) );
  INVx1_ASAP7_75t_SL U63458 ( .A(n59451), .Y(n76880) );
  INVx1_ASAP7_75t_SL U63459 ( .A(n59346), .Y(n59343) );
  INVx1_ASAP7_75t_SL U63460 ( .A(n62620), .Y(n62621) );
  NAND2xp5_ASAP7_75t_SL U63461 ( .A(n62614), .B(n59655), .Y(n62620) );
  INVx1_ASAP7_75t_SL U63462 ( .A(n59396), .Y(n62739) );
  NOR2x1_ASAP7_75t_SL U63463 ( .A(n61913), .B(n61912), .Y(n61920) );
  AOI22xp5_ASAP7_75t_SL U63464 ( .A1(n59100), .A2(n66414), .B1(n66351), .B2(
        n75048), .Y(n66407) );
  NOR2x1p5_ASAP7_75t_SL U63465 ( .A(n68561), .B(n68562), .Y(n68919) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63466 ( .A1(n61043), .A2(n57090), .B(n61042), 
        .C(n77840), .Y(n61052) );
  NAND2xp5_ASAP7_75t_SL U63467 ( .A(n75246), .B(n57120), .Y(n60755) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63468 ( .A1(n75246), .A2(n62682), .B(n61635), 
        .C(n61634), .Y(n61636) );
  INVx1_ASAP7_75t_SL U63469 ( .A(n62688), .Y(n75246) );
  INVx2_ASAP7_75t_SL U63470 ( .A(n66322), .Y(n67298) );
  NAND2xp5_ASAP7_75t_SL U63471 ( .A(n57436), .B(n75467), .Y(n66417) );
  INVx1_ASAP7_75t_SL U63472 ( .A(n63796), .Y(n63682) );
  INVx1_ASAP7_75t_SL U63473 ( .A(n64742), .Y(n64745) );
  NAND2xp5_ASAP7_75t_SL U63474 ( .A(n63683), .B(n63684), .Y(n64742) );
  NAND2x1_ASAP7_75t_SL U63475 ( .A(n62738), .B(n62581), .Y(n62676) );
  NAND2xp5_ASAP7_75t_SL U63476 ( .A(n66571), .B(n66570), .Y(n68594) );
  NAND2xp5_ASAP7_75t_SL U63477 ( .A(n68601), .B(n68600), .Y(n75058) );
  NAND2xp5_ASAP7_75t_SL U63478 ( .A(n68599), .B(n68598), .Y(n68600) );
  INVx1_ASAP7_75t_SL U63479 ( .A(n59566), .Y(n59336) );
  AOI31xp33_ASAP7_75t_SL U63480 ( .A1(n70685), .A2(n70684), .A3(n70683), .B(
        n70682), .Y(n58372) );
  AOI31xp33_ASAP7_75t_SL U63481 ( .A1(n70685), .A2(n70684), .A3(n70683), .B(
        n70682), .Y(n58373) );
  AOI31xp33_ASAP7_75t_SL U63482 ( .A1(n70685), .A2(n70683), .A3(n70684), .B(
        n70682), .Y(n70721) );
  NAND2xp5_ASAP7_75t_SL U63483 ( .A(n76851), .B(n76795), .Y(n62333) );
  AOI21xp5_ASAP7_75t_SL U63484 ( .A1(n77112), .A2(n61902), .B(n61901), .Y(
        n61989) );
  XNOR2xp5_ASAP7_75t_SL U63485 ( .A(n68362), .B(n66925), .Y(n66926) );
  AOI22xp5_ASAP7_75t_SL U63486 ( .A1(n67912), .A2(n65060), .B1(n65059), .B2(
        n67701), .Y(n68153) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63487 ( .A1(n67475), .A2(n67701), .B(n66667), 
        .C(n66739), .Y(n66671) );
  INVx1_ASAP7_75t_SL U63488 ( .A(n62736), .Y(n58984) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63489 ( .A1(n76963), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_17_), .B(n76962), 
        .C(n76961), .Y(n76964) );
  NAND2xp5_ASAP7_75t_SL U63490 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_18_), .B(n76963), 
        .Y(n76962) );
  OAI21xp5_ASAP7_75t_SL U63491 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_7_), .A2(n74849), 
        .B(n74848), .Y(n52494) );
  AOI22xp5_ASAP7_75t_SL U63492 ( .A1(n71087), .A2(n71016), .B1(n59522), .B2(
        n71085), .Y(n70867) );
  OAI22xp5_ASAP7_75t_SL U63493 ( .A1(n57115), .A2(n70717), .B1(n70709), .B2(
        n59524), .Y(n71016) );
  NAND2xp5_ASAP7_75t_SL U63494 ( .A(n59493), .B(n61064), .Y(n60818) );
  INVx1_ASAP7_75t_SL U63495 ( .A(n64721), .Y(n64065) );
  XNOR2x2_ASAP7_75t_SL U63496 ( .A(n64437), .B(n64056), .Y(n64721) );
  AOI22xp5_ASAP7_75t_SL U63497 ( .A1(n59171), .A2(n66934), .B1(n58025), .B2(
        n67720), .Y(n68405) );
  INVx1_ASAP7_75t_SL U63498 ( .A(n68405), .Y(n66935) );
  INVx1_ASAP7_75t_SL U63499 ( .A(n64091), .Y(n58374) );
  OAI22xp5_ASAP7_75t_SL U63500 ( .A1(n67442), .A2(n67021), .B1(n53269), .B2(
        n66682), .Y(n66770) );
  NAND2xp5_ASAP7_75t_SL U63501 ( .A(n62762), .B(n66271), .Y(n62763) );
  INVx2_ASAP7_75t_SL U63502 ( .A(n59560), .Y(n62762) );
  OAI21xp5_ASAP7_75t_SL U63503 ( .A1(n59659), .A2(n68124), .B(n59641), .Y(
        n67092) );
  INVx1_ASAP7_75t_SL U63504 ( .A(n64694), .Y(n64695) );
  XOR2x1_ASAP7_75t_SL U63505 ( .A(n64698), .B(n64697), .Y(n65108) );
  OAI22xp5_ASAP7_75t_SL U63506 ( .A1(n59603), .A2(n67432), .B1(n59605), .B2(
        n75912), .Y(n65060) );
  NAND2xp5_ASAP7_75t_SL U63507 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[7]), .B(
        n73191), .Y(n73053) );
  INVx1_ASAP7_75t_SL U63508 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[7]), .Y(
        n73191) );
  OAI21xp5_ASAP7_75t_SL U63509 ( .A1(n59630), .A2(n73161), .B(n73160), .Y(
        n73164) );
  AOI21xp5_ASAP7_75t_SL U63510 ( .A1(n71690), .A2(n71689), .B(n71735), .Y(
        n71688) );
  NAND2xp5_ASAP7_75t_SL U63511 ( .A(n71723), .B(n71652), .Y(n71735) );
  INVx1_ASAP7_75t_SL U63512 ( .A(n64906), .Y(n64656) );
  AOI22xp5_ASAP7_75t_SL U63513 ( .A1(n57380), .A2(n66726), .B1(n66795), .B2(
        n66794), .Y(n66937) );
  INVx1_ASAP7_75t_SL U63514 ( .A(n59470), .Y(n75762) );
  OAI22xp5_ASAP7_75t_SL U63515 ( .A1(n63838), .A2(n57097), .B1(n63837), .B2(
        n57159), .Y(n64052) );
  INVx1_ASAP7_75t_SL U63516 ( .A(n64052), .Y(n63846) );
  BUFx6f_ASAP7_75t_SL U63517 ( .A(n1766), .Y(n59538) );
  BUFx6f_ASAP7_75t_SL U63518 ( .A(n1785), .Y(n59540) );
  NAND2xp5_ASAP7_75t_SL U63519 ( .A(n66341), .B(n66340), .Y(n66342) );
  NAND2xp5_ASAP7_75t_SL U63520 ( .A(n64984), .B(n64983), .Y(n68345) );
  AOI22xp5_ASAP7_75t_SL U63521 ( .A1(n66683), .A2(n57163), .B1(n66740), .B2(
        n53616), .Y(n66646) );
  NAND2x1p5_ASAP7_75t_SL U63522 ( .A(n59117), .B(n67855), .Y(n59300) );
  NAND2xp5_ASAP7_75t_SL U63523 ( .A(n78185), .B(n4097), .Y(icqmem_adr_qmem[30]) );
  INVx1_ASAP7_75t_SL U63524 ( .A(n68308), .Y(n58955) );
  NAND2xp5_ASAP7_75t_SL U63525 ( .A(n77363), .B(n61038), .Y(n60468) );
  INVx1_ASAP7_75t_SL U63526 ( .A(n68126), .Y(n68266) );
  NAND2xp5_ASAP7_75t_SL U63527 ( .A(n77722), .B(n57644), .Y(n64948) );
  AOI21xp5_ASAP7_75t_SL U63528 ( .A1(n57195), .A2(n59554), .B(n59543), .Y(
        n62582) );
  AOI21x1_ASAP7_75t_SL U63529 ( .A1(n74204), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]), .B(n74200), .Y(
        n74190) );
  NOR2x1_ASAP7_75t_SL U63530 ( .A(n66219), .B(n74875), .Y(n74200) );
  INVx1_ASAP7_75t_SL U63531 ( .A(n59436), .Y(n66882) );
  NAND2xp5_ASAP7_75t_SL U63532 ( .A(n68674), .B(n68673), .Y(n69238) );
  INVx1_ASAP7_75t_SL U63533 ( .A(n66841), .Y(n66708) );
  XNOR2x2_ASAP7_75t_SL U63534 ( .A(n64912), .B(n64911), .Y(n64871) );
  NAND2xp5_ASAP7_75t_SL U63535 ( .A(n59278), .B(n62923), .Y(n62966) );
  NAND2xp5_ASAP7_75t_SL U63536 ( .A(n68608), .B(n68607), .Y(n75072) );
  NAND2xp5_ASAP7_75t_SL U63537 ( .A(n68514), .B(n68515), .Y(n59122) );
  INVx1_ASAP7_75t_SL U63538 ( .A(n67121), .Y(n67125) );
  XNOR2xp5_ASAP7_75t_SL U63539 ( .A(n67204), .B(n58375), .Y(n67218) );
  XNOR2x1_ASAP7_75t_SL U63540 ( .A(n58709), .B(n67064), .Y(n67173) );
  INVx1_ASAP7_75t_SL U63541 ( .A(n58710), .Y(n58709) );
  NAND4xp25_ASAP7_75t_SL U63542 ( .A(n58322), .B(n68699), .C(n68700), .D(
        n69102), .Y(n58376) );
  NAND2x1_ASAP7_75t_SL U63543 ( .A(n69025), .B(n69027), .Y(n68698) );
  OR2x2_ASAP7_75t_SL U63544 ( .A(n68564), .B(n68563), .Y(n58377) );
  OAI22xp5_ASAP7_75t_SL U63545 ( .A1(n64922), .A2(n59460), .B1(n64920), .B2(
        n64921), .Y(n65056) );
  NAND2x1p5_ASAP7_75t_SL U63546 ( .A(n59408), .B(n57106), .Y(n68101) );
  INVx1_ASAP7_75t_SL U63547 ( .A(n67539), .Y(n67551) );
  OAI21x1_ASAP7_75t_SL U63548 ( .A1(n63120), .A2(n59617), .B(n67511), .Y(
        n67842) );
  NAND2xp5_ASAP7_75t_SL U63549 ( .A(n71315), .B(n70851), .Y(n70738) );
  OAI21xp5_ASAP7_75t_SL U63550 ( .A1(n71076), .A2(n70882), .B(n70718), .Y(
        n70851) );
  AOI21xp5_ASAP7_75t_SL U63551 ( .A1(n70753), .A2(n70752), .B(n70751), .Y(
        n70799) );
  INVx1_ASAP7_75t_SL U63552 ( .A(n68902), .Y(n68728) );
  INVx1_ASAP7_75t_SL U63553 ( .A(n71745), .Y(n71744) );
  INVx1_ASAP7_75t_SL U63554 ( .A(n68342), .Y(n58378) );
  INVx1_ASAP7_75t_SL U63555 ( .A(n58378), .Y(n58379) );
  NOR2x1_ASAP7_75t_SL U63556 ( .A(n66779), .B(n66778), .Y(n66817) );
  AOI22xp5_ASAP7_75t_SL U63557 ( .A1(n76653), .A2(n59720), .B1(n76639), .B2(
        n76696), .Y(n75778) );
  INVx1_ASAP7_75t_SL U63558 ( .A(n63163), .Y(n58381) );
  INVx1_ASAP7_75t_SL U63559 ( .A(n58381), .Y(n58382) );
  AOI21xp5_ASAP7_75t_SL U63560 ( .A1(n66283), .A2(n59573), .B(n59574), .Y(
        n66304) );
  INVx1_ASAP7_75t_SL U63561 ( .A(n68648), .Y(n59389) );
  NOR2x1_ASAP7_75t_SL U63562 ( .A(n78003), .B(n62614), .Y(n59070) );
  INVx2_ASAP7_75t_SL U63563 ( .A(n59556), .Y(n78003) );
  INVx1_ASAP7_75t_SL U63564 ( .A(n62710), .Y(n62996) );
  INVx1_ASAP7_75t_SL U63565 ( .A(n63022), .Y(n63006) );
  OAI21xp5_ASAP7_75t_SL U63566 ( .A1(n1737), .A2(n77214), .B(n60232), .Y(
        or1200_cpu_to_sr[1]) );
  OAI22xp5_ASAP7_75t_SL U63567 ( .A1(n66482), .A2(n67743), .B1(n57099), .B2(
        n66481), .Y(n66501) );
  INVx1_ASAP7_75t_SL U63568 ( .A(n64966), .Y(n67748) );
  NOR2x1_ASAP7_75t_SL U63569 ( .A(n63148), .B(n59337), .Y(n63237) );
  XNOR2xp5_ASAP7_75t_SL U63570 ( .A(n59222), .B(n67765), .Y(n68055) );
  BUFx6f_ASAP7_75t_SL U63571 ( .A(n58384), .Y(n58383) );
  NAND2x1_ASAP7_75t_SL U63572 ( .A(n68569), .B(n68568), .Y(n68853) );
  NAND2xp5_ASAP7_75t_SL U63573 ( .A(n61131), .B(n75687), .Y(n60550) );
  OAI22xp5_ASAP7_75t_SL U63574 ( .A1(n67952), .A2(n59460), .B1(n68014), .B2(
        n59515), .Y(n68214) );
  INVx1_ASAP7_75t_SL U63575 ( .A(n64061), .Y(n63869) );
  NOR2x1_ASAP7_75t_SL U63576 ( .A(n58532), .B(n62629), .Y(n62671) );
  XOR2x2_ASAP7_75t_SL U63577 ( .A(n68327), .B(n53481), .Y(n68743) );
  NAND2x1_ASAP7_75t_SL U63578 ( .A(n58830), .B(n58829), .Y(n59252) );
  OAI21xp5_ASAP7_75t_SL U63579 ( .A1(n72544), .A2(n72547), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .Y(
        n72545) );
  OAI21xp5_ASAP7_75t_SL U63580 ( .A1(n72547), .A2(n72546), .B(n72545), .Y(
        n72558) );
  NAND2xp5_ASAP7_75t_SL U63581 ( .A(n72544), .B(n72433), .Y(n72508) );
  MAJIxp5_ASAP7_75t_SL U63582 ( .A(n58348), .B(n68146), .C(n58368), .Y(n58385)
         );
  INVx1_ASAP7_75t_SL U63583 ( .A(n67126), .Y(n67128) );
  INVx1_ASAP7_75t_SL U63584 ( .A(n67873), .Y(n67874) );
  XNOR2x1_ASAP7_75t_SL U63585 ( .A(n58628), .B(n67818), .Y(n67935) );
  AOI22xp5_ASAP7_75t_SL U63586 ( .A1(n68086), .A2(n63613), .B1(n63224), .B2(
        n57478), .Y(n63621) );
  HB1xp67_ASAP7_75t_SL U63587 ( .A(n68343), .Y(n58386) );
  INVx1_ASAP7_75t_SL U63588 ( .A(n67784), .Y(n67325) );
  AND2x2_ASAP7_75t_SL U63589 ( .A(n22057), .B(n60330), .Y(n58387) );
  OAI21xp5_ASAP7_75t_SL U63590 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .A2(n71316), .B(
        n71017), .Y(n71175) );
  OAI21xp5_ASAP7_75t_SL U63591 ( .A1(n71015), .A2(n71207), .B(n71014), .Y(
        n71316) );
  NAND2xp5_ASAP7_75t_SL U63592 ( .A(n71203), .B(n71202), .Y(n71238) );
  NOR2x1_ASAP7_75t_SL U63593 ( .A(n53429), .B(n78182), .Y(n59498) );
  AOI22xp5_ASAP7_75t_SL U63594 ( .A1(n60647), .A2(n57121), .B1(n59498), .B2(
        n60631), .Y(n60935) );
  XNOR2x1_ASAP7_75t_SL U63595 ( .A(n65048), .B(n65047), .Y(n68277) );
  OAI21xp5_ASAP7_75t_SL U63596 ( .A1(n66915), .A2(n59506), .B(n67750), .Y(
        n68362) );
  AOI21xp5_ASAP7_75t_SL U63597 ( .A1(n59594), .A2(n75901), .B(n62653), .Y(
        n63156) );
  INVx1_ASAP7_75t_SL U63598 ( .A(n63200), .Y(n63159) );
  OA21x2_ASAP7_75t_SL U63599 ( .A1(n65031), .A2(n61208), .B(n64504), .Y(n66301) );
  NAND2xp5_ASAP7_75t_SL U63600 ( .A(n60929), .B(n62761), .Y(n63660) );
  AOI21xp5_ASAP7_75t_SL U63601 ( .A1(n57210), .A2(n63124), .B(n63123), .Y(
        n63128) );
  INVx1_ASAP7_75t_SL U63602 ( .A(n57665), .Y(n63123) );
  HB1xp67_ASAP7_75t_SL U63603 ( .A(n68519), .Y(n58388) );
  INVx1_ASAP7_75t_SL U63604 ( .A(n67686), .Y(n59161) );
  OAI21xp5_ASAP7_75t_SL U63605 ( .A1(n68098), .A2(n59510), .B(n62674), .Y(
        n63114) );
  NAND2xp5_ASAP7_75t_SL U63606 ( .A(n68098), .B(n76049), .Y(n62674) );
  INVx1_ASAP7_75t_SL U63607 ( .A(n62754), .Y(n62755) );
  INVx1_ASAP7_75t_SL U63608 ( .A(n64889), .Y(n64614) );
  NAND2xp5_ASAP7_75t_SL U63609 ( .A(n58520), .B(n61911), .Y(n59095) );
  INVx1_ASAP7_75t_SL U63610 ( .A(n68301), .Y(n68292) );
  OAI21xp5_ASAP7_75t_SL U63611 ( .A1(n75977), .A2(n76190), .B(n75976), .Y(
        n76187) );
  NAND2xp5_ASAP7_75t_SL U63612 ( .A(n76092), .B(n57133), .Y(n76093) );
  NAND2xp5_ASAP7_75t_SL U63613 ( .A(n61915), .B(n61914), .Y(n74787) );
  AO22x1_ASAP7_75t_SL U63614 ( .A1(n76631), .A2(n58390), .B1(n75909), .B2(
        n58600), .Y(or1200_cpu_or1200_mult_mac_n1513) );
  XOR2xp5_ASAP7_75t_SL U63615 ( .A(or1200_cpu_or1200_mult_mac_n38), .B(n76073), 
        .Y(n58390) );
  AO22x1_ASAP7_75t_SL U63616 ( .A1(n76631), .A2(n58391), .B1(n75902), .B2(
        n58600), .Y(or1200_cpu_or1200_mult_mac_n1518) );
  XOR2xp5_ASAP7_75t_SL U63617 ( .A(or1200_cpu_or1200_mult_mac_n48), .B(n76030), 
        .Y(n58391) );
  AO22x1_ASAP7_75t_SL U63618 ( .A1(n76631), .A2(n58392), .B1(n75924), .B2(
        n58600), .Y(or1200_cpu_or1200_mult_mac_n1523) );
  XOR2xp5_ASAP7_75t_SL U63619 ( .A(or1200_cpu_or1200_mult_mac_n58), .B(n75993), 
        .Y(n58392) );
  INVx1_ASAP7_75t_SL U63620 ( .A(or1200_cpu_or1200_mult_mac_n56), .Y(n75924)
         );
  OAI21xp5_ASAP7_75t_SL U63621 ( .A1(n59485), .A2(n75643), .B(n59487), .Y(
        n67881) );
  NAND2xp5_ASAP7_75t_SL U63622 ( .A(n75906), .B(n57277), .Y(n59112) );
  NOR2x1_ASAP7_75t_SL U63623 ( .A(n67881), .B(n68133), .Y(n68109) );
  NAND2xp5_ASAP7_75t_SL U63624 ( .A(n66806), .B(n57277), .Y(n66404) );
  AOI21xp5_ASAP7_75t_SL U63625 ( .A1(n57277), .A2(n76077), .B(n66620), .Y(
        n66621) );
  AOI21xp5_ASAP7_75t_SL U63626 ( .A1(n71132), .A2(n71129), .B(n71128), .Y(
        n71134) );
  OAI21xp5_ASAP7_75t_SL U63627 ( .A1(n71097), .A2(n71096), .B(n71111), .Y(
        n71129) );
  NAND2xp5_ASAP7_75t_SL U63628 ( .A(n67845), .B(n67262), .Y(n67263) );
  OAI21xp5_ASAP7_75t_SL U63629 ( .A1(n59631), .A2(n73244), .B(n73240), .Y(
        n73246) );
  OAI22xp5_ASAP7_75t_SL U63630 ( .A1(n57115), .A2(n70881), .B1(n70863), .B2(
        n59524), .Y(n71208) );
  INVx1_ASAP7_75t_SL U63631 ( .A(n71176), .Y(n71318) );
  INVx2_ASAP7_75t_SL U63632 ( .A(n2547), .Y(n62561) );
  AOI22xp5_ASAP7_75t_SL U63633 ( .A1(n66466), .A2(n59635), .B1(n66281), .B2(
        n75048), .Y(n66433) );
  AOI21xp5_ASAP7_75t_SL U63634 ( .A1(n67741), .A2(n75644), .B(n66255), .Y(
        n66466) );
  NAND2xp5_ASAP7_75t_SL U63635 ( .A(n58758), .B(n65040), .Y(n67946) );
  NAND2xp5_ASAP7_75t_SL U63636 ( .A(n75102), .B(n75098), .Y(n75111) );
  NAND2xp5_ASAP7_75t_SL U63637 ( .A(n68620), .B(n68619), .Y(n75098) );
  NOR2x1_ASAP7_75t_SL U63638 ( .A(n59147), .B(n59146), .Y(n68375) );
  OAI22xp5_ASAP7_75t_SL U63639 ( .A1(n66754), .A2(n59491), .B1(n66753), .B2(
        n59612), .Y(n66813) );
  INVx1_ASAP7_75t_SL U63640 ( .A(n66815), .Y(n66761) );
  NAND2x1p5_ASAP7_75t_SL U63641 ( .A(n64511), .B(n63808), .Y(n67972) );
  NAND2xp5_ASAP7_75t_SL U63642 ( .A(n63806), .B(n63809), .Y(n64511) );
  NAND2xp5_ASAP7_75t_SL U63643 ( .A(n57100), .B(n60058), .Y(n4114) );
  OAI21xp5_ASAP7_75t_SL U63644 ( .A1(n65008), .A2(n65007), .B(n65006), .Y(
        n65012) );
  NAND2xp5_ASAP7_75t_SL U63645 ( .A(n57122), .B(n64481), .Y(n64923) );
  NAND2xp5_ASAP7_75t_SL U63646 ( .A(n59210), .B(n59310), .Y(n64481) );
  AOI22xp5_ASAP7_75t_SL U63647 ( .A1(n67609), .A2(n64927), .B1(n64926), .B2(
        n64925), .Y(n68222) );
  OAI22xp5_ASAP7_75t_SL U63648 ( .A1(n63679), .A2(n67452), .B1(n63858), .B2(
        n67906), .Y(n63819) );
  OAI21xp5_ASAP7_75t_SL U63649 ( .A1(n59609), .A2(n59510), .B(n58695), .Y(
        n63842) );
  INVx1_ASAP7_75t_SL U63650 ( .A(n64540), .Y(n64404) );
  OAI22xp5_ASAP7_75t_SL U63651 ( .A1(n59440), .A2(n56984), .B1(n59446), .B2(
        n66933), .Y(n68406) );
  INVx1_ASAP7_75t_SL U63652 ( .A(n66981), .Y(n66839) );
  BUFx6f_ASAP7_75t_SL U63653 ( .A(n2835), .Y(n59570) );
  OAI21xp5_ASAP7_75t_SL U63654 ( .A1(n76190), .A2(n75975), .B(n76193), .Y(
        n75976) );
  NAND2xp5_ASAP7_75t_SL U63655 ( .A(n75985), .B(n57133), .Y(n75986) );
  INVx1_ASAP7_75t_SL U63656 ( .A(n59065), .Y(n67564) );
  INVx1_ASAP7_75t_SL U63657 ( .A(n66647), .Y(n66627) );
  OAI21xp5_ASAP7_75t_SL U63658 ( .A1(n59472), .A2(n64365), .B(n64364), .Y(
        n64651) );
  OAI21xp5_ASAP7_75t_SL U63659 ( .A1(n69071), .A2(n69070), .B(n69069), .Y(
        n69085) );
  INVx1_ASAP7_75t_SL U63660 ( .A(n67880), .Y(n68110) );
  INVx1_ASAP7_75t_SL U63661 ( .A(n59407), .Y(n68095) );
  OAI22xp5_ASAP7_75t_SL U63662 ( .A1(or1200_cpu_or1200_except_n661), .A2(
        n77388), .B1(n2037), .B2(n75180), .Y(n77389) );
  INVx1_ASAP7_75t_SL U63663 ( .A(n67390), .Y(n67571) );
  INVx1_ASAP7_75t_SL U63664 ( .A(n66814), .Y(n59071) );
  INVx1_ASAP7_75t_SL U63665 ( .A(n65041), .Y(n64612) );
  INVx1_ASAP7_75t_SL U63666 ( .A(n56993), .Y(n58802) );
  INVx1_ASAP7_75t_SL U63667 ( .A(n68421), .Y(n68422) );
  OAI21xp5_ASAP7_75t_SL U63668 ( .A1(n75947), .A2(n57242), .B(n58384), .Y(
        n67063) );
  INVx1_ASAP7_75t_SL U63669 ( .A(n68627), .Y(n69226) );
  OAI21xp5_ASAP7_75t_SL U63670 ( .A1(n64041), .A2(n64042), .B(n58491), .Y(
        n64344) );
  OAI21xp5_ASAP7_75t_SL U63671 ( .A1(n67288), .A2(n59637), .B(n67287), .Y(
        n67556) );
  AOI22xp5_ASAP7_75t_SL U63672 ( .A1(n67251), .A2(n62879), .B1(n62878), .B2(
        n62877), .Y(n62906) );
  OAI21xp5_ASAP7_75t_SL U63673 ( .A1(n62901), .A2(n63299), .B(n62900), .Y(
        n62904) );
  NAND2x1_ASAP7_75t_SL U63674 ( .A(n59557), .B(n59559), .Y(n62590) );
  INVx1_ASAP7_75t_SL U63675 ( .A(n66554), .Y(n66555) );
  OAI21xp5_ASAP7_75t_SL U63676 ( .A1(n63450), .A2(n63449), .B(n63448), .Y(
        n63480) );
  AOI21xp5_ASAP7_75t_SL U63677 ( .A1(n63447), .A2(n63446), .B(n63445), .Y(
        n63449) );
  INVx1_ASAP7_75t_SL U63678 ( .A(n67889), .Y(n59008) );
  NAND2xp5_ASAP7_75t_SL U63679 ( .A(n59512), .B(n59641), .Y(n67338) );
  XNOR2xp5_ASAP7_75t_SL U63680 ( .A(n68052), .B(n68051), .Y(n59355) );
  INVx1_ASAP7_75t_SL U63681 ( .A(n63835), .Y(n63130) );
  INVx1_ASAP7_75t_SL U63682 ( .A(n63108), .Y(n58947) );
  INVx2_ASAP7_75t_SL U63683 ( .A(n64990), .Y(n64981) );
  XNOR2x1_ASAP7_75t_SL U63684 ( .A(n57489), .B(n64980), .Y(n64990) );
  NAND2xp5_ASAP7_75t_SL U63685 ( .A(n59438), .B(n60644), .Y(n75478) );
  NAND2xp5_ASAP7_75t_SL U63686 ( .A(n62075), .B(n62084), .Y(n61956) );
  NAND2xp5_ASAP7_75t_SL U63687 ( .A(n66311), .B(n66307), .Y(n66308) );
  NOR2x1_ASAP7_75t_SL U63688 ( .A(n59574), .B(n59020), .Y(n66307) );
  XNOR2xp5_ASAP7_75t_SL U63689 ( .A(n66950), .B(n66949), .Y(n66951) );
  INVx1_ASAP7_75t_SL U63690 ( .A(n69026), .Y(n69038) );
  OAI22xp5_ASAP7_75t_SL U63691 ( .A1(n67974), .A2(n62741), .B1(n57156), .B2(
        n63066), .Y(n63059) );
  OAI21xp5_ASAP7_75t_SL U63692 ( .A1(n67971), .A2(n59641), .B(n66858), .Y(
        n67003) );
  AOI21xp5_ASAP7_75t_SL U63693 ( .A1(n66487), .A2(n66486), .B(n66485), .Y(
        n66489) );
  NOR2x1_ASAP7_75t_SL U63694 ( .A(n59358), .B(n58436), .Y(n68371) );
  XNOR2xp5_ASAP7_75t_SL U63695 ( .A(n59006), .B(n57354), .Y(n68552) );
  OAI21xp5_ASAP7_75t_SL U63696 ( .A1(n66692), .A2(n58321), .B(n66843), .Y(
        n66977) );
  XOR2xp5_ASAP7_75t_SL U63697 ( .A(n64869), .B(n58338), .Y(n64753) );
  NAND2xp5_ASAP7_75t_SL U63698 ( .A(n57111), .B(n63171), .Y(n63183) );
  NAND2xp5_ASAP7_75t_SL U63699 ( .A(n57111), .B(n64366), .Y(n64370) );
  OAI22xp5_ASAP7_75t_SL U63700 ( .A1(n57172), .A2(n63183), .B1(n57111), .B2(
        n66805), .Y(n63189) );
  OAI21xp5_ASAP7_75t_SL U63701 ( .A1(n67748), .A2(n57111), .B(n67749), .Y(
        n62822) );
  INVx1_ASAP7_75t_SL U63702 ( .A(n67199), .Y(n67200) );
  OAI22xp5_ASAP7_75t_SL U63703 ( .A1(n67752), .A2(n59491), .B1(n58658), .B2(
        n66955), .Y(n68359) );
  NAND2xp5_ASAP7_75t_SL U63704 ( .A(n57491), .B(n59664), .Y(n66482) );
  O2A1O1Ixp5_ASAP7_75t_SL U63705 ( .A1(n67232), .A2(n64441), .B(n59660), .C(
        n64387), .Y(n64388) );
  O2A1O1Ixp5_ASAP7_75t_SL U63706 ( .A1(n67232), .A2(n53280), .B(n63115), .C(
        n58907), .Y(n63116) );
  INVx1_ASAP7_75t_SL U63707 ( .A(n62990), .Y(n62932) );
  OAI22xp5_ASAP7_75t_SL U63708 ( .A1(n64042), .A2(n62816), .B1(n57362), .B2(
        n62815), .Y(n62929) );
  OAI21xp5_ASAP7_75t_SL U63709 ( .A1(n53197), .A2(n68022), .B(n66702), .Y(
        n66869) );
  NAND2xp5_ASAP7_75t_SL U63710 ( .A(n59012), .B(n68022), .Y(n68117) );
  NAND2xp5_ASAP7_75t_SL U63711 ( .A(n75974), .B(n75973), .Y(n75977) );
  AND2x4_ASAP7_75t_SL U63712 ( .A(n76631), .B(n57133), .Y(n76195) );
  NAND2xp5_ASAP7_75t_SL U63713 ( .A(n59573), .B(n66301), .Y(n66305) );
  INVx1_ASAP7_75t_SL U63714 ( .A(n64904), .Y(n64654) );
  OAI22xp5_ASAP7_75t_SL U63715 ( .A1(n57253), .A2(n66883), .B1(n66885), .B2(
        n66884), .Y(n67024) );
  INVx1_ASAP7_75t_SL U63716 ( .A(n66994), .Y(n66883) );
  OAI22xp5_ASAP7_75t_SL U63717 ( .A1(n68119), .A2(n66480), .B1(n59116), .B2(
        n67078), .Y(n66500) );
  NAND2xp5_ASAP7_75t_SL U63718 ( .A(n59641), .B(n59651), .Y(n66480) );
  XNOR2x2_ASAP7_75t_SL U63719 ( .A(n66347), .B(n66346), .Y(n66506) );
  INVx1_ASAP7_75t_SL U63720 ( .A(n66687), .Y(n59296) );
  OAI21xp5_ASAP7_75t_SL U63721 ( .A1(n59670), .A2(n57172), .B(n58666), .Y(
        n67020) );
  NOR2x1_ASAP7_75t_SL U63722 ( .A(n67082), .B(n67081), .Y(n67085) );
  NOR2x1_ASAP7_75t_SL U63723 ( .A(n57158), .B(n67022), .Y(n67081) );
  NOR2x1_ASAP7_75t_SL U63724 ( .A(n53242), .B(n67020), .Y(n67082) );
  NAND2xp5_ASAP7_75t_SL U63725 ( .A(n65371), .B(n65289), .Y(n65375) );
  NAND2xp5_ASAP7_75t_SL U63726 ( .A(n2854), .B(n65271), .Y(n65263) );
  AOI21xp5_ASAP7_75t_SL U63727 ( .A1(n63135), .A2(n63134), .B(n63150), .Y(
        n63138) );
  NAND2xp5_ASAP7_75t_SL U63728 ( .A(n57082), .B(n64353), .Y(n62683) );
  INVx1_ASAP7_75t_SL U63729 ( .A(n64589), .Y(n64520) );
  OAI21xp5_ASAP7_75t_SL U63730 ( .A1(n57099), .A2(n67923), .B(n58801), .Y(
        n67996) );
  NAND2xp5_ASAP7_75t_SL U63731 ( .A(n67306), .B(n58413), .Y(n58801) );
  NAND2xp5_ASAP7_75t_SL U63732 ( .A(n75832), .B(n66244), .Y(n58676) );
  NAND2xp5_ASAP7_75t_SL U63733 ( .A(n74557), .B(n68702), .Y(n68709) );
  OAI22xp5_ASAP7_75t_SL U63734 ( .A1(n67974), .A2(n63843), .B1(n57156), .B2(
        n63842), .Y(n64050) );
  NAND2xp5_ASAP7_75t_SL U63735 ( .A(n57312), .B(n58353), .Y(n64079) );
  NOR2x1_ASAP7_75t_SL U63736 ( .A(n66817), .B(n66820), .Y(n66822) );
  AOI22xp5_ASAP7_75t_SL U63737 ( .A1(n66507), .A2(n66273), .B1(n66272), .B2(
        n66433), .Y(n66276) );
  NOR2x1_ASAP7_75t_SL U63738 ( .A(n66250), .B(n66252), .Y(n66507) );
  AOI21xp5_ASAP7_75t_SL U63739 ( .A1(n66394), .A2(n66395), .B(n66282), .Y(
        n66606) );
  INVx1_ASAP7_75t_SL U63740 ( .A(n67785), .Y(n67324) );
  XNOR2x1_ASAP7_75t_SL U63741 ( .A(n67624), .B(n58694), .Y(n67794) );
  OAI21xp5_ASAP7_75t_SL U63742 ( .A1(n59599), .A2(n67276), .B(n66790), .Y(
        n68415) );
  NAND2xp5_ASAP7_75t_SL U63743 ( .A(n59598), .B(n67911), .Y(n66790) );
  NAND2xp5_ASAP7_75t_SL U63744 ( .A(n2779), .B(n60281), .Y(n77349) );
  AOI31xp67_ASAP7_75t_SL U63745 ( .A1(n62150), .A2(n60309), .A3(n62148), .B(
        n60308), .Y(or1200_cpu_or1200_if_if_bypass) );
  OAI21xp5_ASAP7_75t_SL U63746 ( .A1(n67489), .A2(n53619), .B(n58691), .Y(
        n67728) );
  OAI22xp5_ASAP7_75t_SL U63747 ( .A1(n57115), .A2(n70759), .B1(n70735), .B2(
        n70993), .Y(n71074) );
  NAND2xp5_ASAP7_75t_SL U63748 ( .A(n67963), .B(n59651), .Y(n67479) );
  INVx1_ASAP7_75t_SL U63749 ( .A(n68322), .Y(n68312) );
  INVx1_ASAP7_75t_SL U63750 ( .A(n64017), .Y(n64020) );
  INVx1_ASAP7_75t_SL U63751 ( .A(n63005), .Y(n63023) );
  NOR2x1_ASAP7_75t_SL U63752 ( .A(n53615), .B(n58906), .Y(n62722) );
  NOR2x1_ASAP7_75t_SL U63753 ( .A(n62857), .B(n62797), .Y(n62931) );
  OAI22x1_ASAP7_75t_SL U63754 ( .A1(n68425), .A2(n68424), .B1(n68423), .B2(
        n68422), .Y(n68429) );
  OAI21xp5_ASAP7_75t_SL U63755 ( .A1(n68420), .A2(n68421), .B(n68419), .Y(
        n68424) );
  OAI21xp5_ASAP7_75t_SL U63756 ( .A1(n64428), .A2(n59453), .B(n59241), .Y(
        n64600) );
  INVx1_ASAP7_75t_SL U63757 ( .A(n59297), .Y(n67632) );
  NAND2xp5_ASAP7_75t_SL U63758 ( .A(n64718), .B(n59370), .Y(n59368) );
  NOR2x1_ASAP7_75t_SL U63759 ( .A(n64709), .B(n59368), .Y(n59366) );
  BUFx3_ASAP7_75t_SL U63760 ( .A(n67972), .Y(n58861) );
  INVx1_ASAP7_75t_SL U63761 ( .A(n67815), .Y(n59312) );
  AOI21xp5_ASAP7_75t_SL U63762 ( .A1(n66258), .A2(n57448), .B(n53316), .Y(
        n62576) );
  NAND2xp5_ASAP7_75t_SL U63763 ( .A(n62808), .B(n62807), .Y(n68078) );
  OAI22xp5_ASAP7_75t_SL U63764 ( .A1(n64538), .A2(n53269), .B1(n58499), .B2(
        n68383), .Y(n64337) );
  NAND2xp5_ASAP7_75t_SL U63765 ( .A(n58699), .B(n67531), .Y(n67436) );
  OAI21xp5_ASAP7_75t_SL U63766 ( .A1(n57179), .A2(n75927), .B(n67921), .Y(
        n68004) );
  INVx1_ASAP7_75t_SL U63767 ( .A(n68190), .Y(n68026) );
  OAI22xp5_ASAP7_75t_SL U63768 ( .A1(n58903), .A2(n67021), .B1(n67442), .B2(
        n66853), .Y(n66868) );
  NOR2x1_ASAP7_75t_SL U63769 ( .A(n67212), .B(n67211), .Y(n69100) );
  INVx1_ASAP7_75t_SL U63770 ( .A(n67497), .Y(n67499) );
  INVx1_ASAP7_75t_SL U63771 ( .A(n67499), .Y(n58704) );
  NAND2xp5_ASAP7_75t_SL U63772 ( .A(n64374), .B(n67464), .Y(n64531) );
  OAI21xp5_ASAP7_75t_SL U63773 ( .A1(n59598), .A2(n59514), .B(n63815), .Y(
        n64374) );
  INVx1_ASAP7_75t_SL U63774 ( .A(n64352), .Y(n64075) );
  NAND2xp5_ASAP7_75t_SL U63775 ( .A(n64074), .B(n64073), .Y(n64352) );
  NAND2xp5_ASAP7_75t_SL U63776 ( .A(n59513), .B(n67740), .Y(n63664) );
  AOI22xp5_ASAP7_75t_SL U63777 ( .A1(n63799), .A2(n63798), .B1(n63797), .B2(
        n63796), .Y(n64068) );
  INVx1_ASAP7_75t_SL U63778 ( .A(n64068), .Y(n63848) );
  HB1xp67_ASAP7_75t_SL U63779 ( .A(n64714), .Y(n58395) );
  INVx1_ASAP7_75t_SL U63780 ( .A(n64060), .Y(n63855) );
  XNOR2x1_ASAP7_75t_SL U63781 ( .A(n63623), .B(n63855), .Y(n63872) );
  BUFx2_ASAP7_75t_SL U63782 ( .A(n66450), .Y(n59590) );
  INVx1_ASAP7_75t_SL U63783 ( .A(n64051), .Y(n63844) );
  NAND2xp5_ASAP7_75t_SL U63784 ( .A(n53617), .B(n57195), .Y(n62737) );
  NAND2xp5_ASAP7_75t_SL U63785 ( .A(n57377), .B(n61943), .Y(n62094) );
  INVx1_ASAP7_75t_SL U63786 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_), .Y(
        n74265) );
  OAI22xp5_ASAP7_75t_SL U63787 ( .A1(n64064), .A2(n64063), .B1(n64062), .B2(
        n64061), .Y(n64712) );
  INVx1_ASAP7_75t_SL U63788 ( .A(n64057), .Y(n64062) );
  NAND2xp5_ASAP7_75t_SL U63789 ( .A(n67083), .B(n67085), .Y(n67088) );
  AOI22xp5_ASAP7_75t_SL U63790 ( .A1(n57161), .A2(n66750), .B1(n66751), .B2(
        n67306), .Y(n66811) );
  OAI21xp5_ASAP7_75t_SL U63791 ( .A1(n59600), .A2(n67276), .B(n66610), .Y(
        n66751) );
  OAI21xp5_ASAP7_75t_SL U63792 ( .A1(n59668), .A2(n67144), .B(n58858), .Y(
        n67130) );
  INVx1_ASAP7_75t_SL U63793 ( .A(n68278), .Y(n58880) );
  OAI21xp5_ASAP7_75t_SL U63794 ( .A1(n63072), .A2(n62772), .B(n62771), .Y(
        n63073) );
  OAI22xp5_ASAP7_75t_SL U63795 ( .A1(n53203), .A2(n62693), .B1(n57156), .B2(
        n62741), .Y(n62771) );
  AO21x2_ASAP7_75t_SL U63796 ( .A1(n64510), .A2(n64511), .B(n57397), .Y(n67276) );
  INVx1_ASAP7_75t_SL U63797 ( .A(n64509), .Y(n58979) );
  INVx1_ASAP7_75t_SL U63798 ( .A(n64994), .Y(n64910) );
  NAND2xp5_ASAP7_75t_SL U63799 ( .A(n71153), .B(n71154), .Y(n71137) );
  OAI22xp5_ASAP7_75t_SL U63800 ( .A1(n58878), .A2(n59051), .B1(n62712), .B2(
        n62713), .Y(n63025) );
  OAI22xp5_ASAP7_75t_SL U63801 ( .A1(n62996), .A2(n62999), .B1(n62997), .B2(
        n62998), .Y(n59051) );
  NAND2xp5_ASAP7_75t_SL U63802 ( .A(n4132), .B(n78264), .Y(icqmem_adr_qmem[13]) );
  NAND2xp5_ASAP7_75t_SL U63803 ( .A(n57126), .B(n75589), .Y(n75338) );
  NAND2xp5_ASAP7_75t_SL U63804 ( .A(n57126), .B(n75847), .Y(n75722) );
  NAND2xp5_ASAP7_75t_SL U63805 ( .A(n57126), .B(n61494), .Y(n77105) );
  INVx1_ASAP7_75t_SL U63806 ( .A(n75338), .Y(n75741) );
  OAI21xp5_ASAP7_75t_SL U63807 ( .A1(n59612), .A2(n66613), .B(n66612), .Y(
        n66736) );
  NAND2xp5_ASAP7_75t_SL U63808 ( .A(n58981), .B(n67687), .Y(n67688) );
  OAI21xp5_ASAP7_75t_SL U63809 ( .A1(n72640), .A2(n72636), .B(n72638), .Y(
        n72632) );
  NAND2xp5_ASAP7_75t_SL U63810 ( .A(n72625), .B(n72624), .Y(n72638) );
  NAND2xp5_ASAP7_75t_SL U63811 ( .A(n75628), .B(n59589), .Y(n64514) );
  NOR2x1_ASAP7_75t_SL U63812 ( .A(n74336), .B(n74337), .Y(n74346) );
  OAI21xp5_ASAP7_75t_SL U63813 ( .A1(n66860), .A2(n67736), .B(n56981), .Y(
        n67076) );
  OAI21xp5_ASAP7_75t_SL U63814 ( .A1(n66860), .A2(n59668), .B(n66285), .Y(
        n66334) );
  INVx1_ASAP7_75t_SL U63815 ( .A(n68306), .Y(n65048) );
  INVx1_ASAP7_75t_SL U63816 ( .A(n57184), .Y(n66860) );
  INVx1_ASAP7_75t_SL U63817 ( .A(n63842), .Y(n64393) );
  AOI21xp5_ASAP7_75t_SL U63818 ( .A1(n57167), .A2(n53320), .B(n64031), .Y(
        n64384) );
  NAND2xp5_ASAP7_75t_SL U63819 ( .A(n59601), .B(n67146), .Y(n67150) );
  NAND2xp5_ASAP7_75t_SL U63820 ( .A(n64742), .B(n65102), .Y(n63881) );
  AOI21xp5_ASAP7_75t_SL U63821 ( .A1(n57332), .A2(n65105), .B(n65106), .Y(
        n64095) );
  INVx1_ASAP7_75t_SL U63822 ( .A(n60945), .Y(n59405) );
  NAND2x1p5_ASAP7_75t_SL U63823 ( .A(n59528), .B(n59529), .Y(n60945) );
  NAND2xp5_ASAP7_75t_SL U63824 ( .A(n58383), .B(n67444), .Y(n58761) );
  INVx1_ASAP7_75t_SL U63825 ( .A(n62611), .Y(n58720) );
  INVx1_ASAP7_75t_SL U63826 ( .A(n68355), .Y(n58782) );
  OAI21xp5_ASAP7_75t_SL U63827 ( .A1(n68306), .A2(n68305), .B(n68304), .Y(
        n68319) );
  NAND2xp5_ASAP7_75t_SL U63828 ( .A(n68259), .B(n68258), .Y(n68304) );
  INVx1_ASAP7_75t_SL U63829 ( .A(n68057), .Y(n67792) );
  INVx1_ASAP7_75t_SL U63830 ( .A(n70661), .Y(n70685) );
  OAI21xp5_ASAP7_75t_SL U63831 ( .A1(n71015), .A2(n70864), .B(n70710), .Y(
        n70931) );
  NAND2xp5_ASAP7_75t_SL U63832 ( .A(n71015), .B(n71016), .Y(n70710) );
  NOR2x1_ASAP7_75t_SL U63833 ( .A(n59709), .B(n61921), .Y(n61930) );
  AOI22xp5_ASAP7_75t_SL U63834 ( .A1(n75895), .A2(n57112), .B1(n64923), .B2(
        n64484), .Y(n64626) );
  NAND2xp5_ASAP7_75t_SL U63835 ( .A(n59655), .B(n62676), .Y(n59395) );
  INVx1_ASAP7_75t_SL U63836 ( .A(n64592), .Y(n64545) );
  INVx1_ASAP7_75t_SL U63837 ( .A(n64593), .Y(n64546) );
  INVx1_ASAP7_75t_SL U63838 ( .A(n68017), .Y(n64426) );
  NAND2xp5_ASAP7_75t_SL U63839 ( .A(n63700), .B(n62150), .Y(n63712) );
  NAND2xp5_ASAP7_75t_SL U63840 ( .A(n68649), .B(n68919), .Y(n68665) );
  NOR2x1p5_ASAP7_75t_SL U63841 ( .A(n75710), .B(n59645), .Y(n64229) );
  XNOR2xp5_ASAP7_75t_SL U63842 ( .A(n64705), .B(n64704), .Y(n64726) );
  NAND2xp5_ASAP7_75t_SL U63843 ( .A(n59379), .B(n60914), .Y(n59378) );
  NAND2x1_ASAP7_75t_SL U63844 ( .A(n71308), .B(n71307), .Y(n71350) );
  OAI21xp5_ASAP7_75t_SL U63845 ( .A1(n70907), .A2(n70906), .B(n70908), .Y(
        n70978) );
  OAI22xp5_ASAP7_75t_SL U63846 ( .A1(n58315), .A2(n71018), .B1(n70844), .B2(
        n58328), .Y(n70869) );
  NAND2xp5_ASAP7_75t_SL U63847 ( .A(n71229), .B(n71263), .Y(n70708) );
  NAND2xp5_ASAP7_75t_SL U63848 ( .A(n1924), .B(n59572), .Y(n59922) );
  BUFx6f_ASAP7_75t_SL U63849 ( .A(n2848), .Y(n59572) );
  NAND2xp5_ASAP7_75t_SL U63850 ( .A(n68922), .B(n68921), .Y(n68930) );
  INVx1_ASAP7_75t_SL U63851 ( .A(n58901), .Y(n64401) );
  NAND2xp5_ASAP7_75t_SL U63852 ( .A(n67481), .B(n57182), .Y(n58901) );
  INVx1_ASAP7_75t_SL U63853 ( .A(n67042), .Y(n59007) );
  INVx1_ASAP7_75t_SL U63854 ( .A(n63008), .Y(n59227) );
  NAND2xp5_ASAP7_75t_SL U63855 ( .A(n67211), .B(n67212), .Y(n59388) );
  OAI21xp5_ASAP7_75t_SL U63856 ( .A1(n63674), .A2(n57315), .B(n58879), .Y(
        n63679) );
  NAND2xp5_ASAP7_75t_SL U63857 ( .A(n57112), .B(n76078), .Y(n58879) );
  INVx1_ASAP7_75t_SL U63858 ( .A(n63795), .Y(n63797) );
  INVx1_ASAP7_75t_SL U63859 ( .A(n67398), .Y(n59221) );
  NAND2xp5_ASAP7_75t_SL U63860 ( .A(n68149), .B(n68152), .Y(n59286) );
  NOR2x1_ASAP7_75t_SL U63861 ( .A(n68106), .B(n68105), .Y(n68152) );
  AOI21xp5_ASAP7_75t_SL U63862 ( .A1(n73413), .A2(n73289), .B(n73288), .Y(
        n73290) );
  NAND2xp5_ASAP7_75t_SL U63863 ( .A(n58461), .B(n63039), .Y(n63448) );
  INVx1_ASAP7_75t_SL U63864 ( .A(n62683), .Y(n62613) );
  NOR2x1_ASAP7_75t_SL U63865 ( .A(n62587), .B(n62586), .Y(n63018) );
  INVx1_ASAP7_75t_SL U63866 ( .A(n63166), .Y(n58946) );
  OAI21xp5_ASAP7_75t_SL U63867 ( .A1(n67279), .A2(n57076), .B(n67278), .Y(
        n67470) );
  NAND2xp5_ASAP7_75t_SL U63868 ( .A(n67920), .B(n75644), .Y(n67280) );
  O2A1O1Ixp5_ASAP7_75t_SL U63869 ( .A1(n59333), .A2(n58927), .B(n59655), .C(
        n59591), .Y(n67354) );
  INVx1_ASAP7_75t_SL U63870 ( .A(n59402), .Y(n59401) );
  NAND2xp5_ASAP7_75t_SL U63871 ( .A(n59360), .B(n58714), .Y(n58713) );
  OAI22xp5_ASAP7_75t_SL U63872 ( .A1(n59515), .A2(n63110), .B1(n63080), .B2(
        n58356), .Y(n63155) );
  NAND2xp5_ASAP7_75t_SL U63873 ( .A(n71023), .B(n70992), .Y(n71009) );
  AOI21xp5_ASAP7_75t_SL U63874 ( .A1(n70982), .A2(n70981), .B(n70980), .Y(
        n70992) );
  AOI21xp5_ASAP7_75t_SL U63875 ( .A1(n58730), .A2(n58902), .B(n68901), .Y(
        n68649) );
  NAND2x1_ASAP7_75t_SL U63876 ( .A(n58902), .B(n68559), .Y(n68726) );
  OAI21xp5_ASAP7_75t_SL U63877 ( .A1(n57253), .A2(n59469), .B(n59415), .Y(
        n68170) );
  NAND2xp5_ASAP7_75t_SL U63878 ( .A(n65042), .B(n67096), .Y(n59415) );
  NOR2x1_ASAP7_75t_SL U63879 ( .A(n63187), .B(n63186), .Y(n63825) );
  XNOR2xp5_ASAP7_75t_SL U63880 ( .A(n63844), .B(n64050), .Y(n63845) );
  INVx1_ASAP7_75t_SL U63881 ( .A(n58406), .Y(n58748) );
  INVx1_ASAP7_75t_SL U63882 ( .A(n68194), .Y(n68196) );
  NAND2xp5_ASAP7_75t_SL U63883 ( .A(n59607), .B(n57409), .Y(n66352) );
  NAND2xp5_ASAP7_75t_SL U63884 ( .A(n53221), .B(n66352), .Y(n66355) );
  INVx1_ASAP7_75t_SL U63885 ( .A(n64736), .Y(n64737) );
  INVx3_ASAP7_75t_SL U63886 ( .A(n67839), .Y(n67264) );
  AOI21xp5_ASAP7_75t_SL U63887 ( .A1(n76273), .A2(n77031), .B(n64864), .Y(
        n77867) );
  INVx1_ASAP7_75t_SL U63888 ( .A(n68695), .Y(n68700) );
  NAND2x1p5_ASAP7_75t_SL U63889 ( .A(n69143), .B(n69148), .Y(n68695) );
  OAI22xp5_ASAP7_75t_SL U63890 ( .A1(n57099), .A2(n66766), .B1(n66765), .B2(
        n57165), .Y(n66823) );
  AOI21xp5_ASAP7_75t_SL U63891 ( .A1(n67741), .A2(n57179), .B(n66674), .Y(
        n66765) );
  BUFx3_ASAP7_75t_SL U63892 ( .A(n1862), .Y(n59547) );
  NOR2x1_ASAP7_75t_SL U63893 ( .A(n66889), .B(n66888), .Y(n67027) );
  OAI21xp5_ASAP7_75t_SL U63894 ( .A1(n59617), .A2(n67467), .B(n67466), .Y(
        n67693) );
  OAI22xp5_ASAP7_75t_SL U63895 ( .A1(n68383), .A2(n68381), .B1(n67693), .B2(
        n58903), .Y(n68398) );
  OAI21xp5_ASAP7_75t_SL U63896 ( .A1(n63021), .A2(n63446), .B(n63444), .Y(
        n58817) );
  OAI21xp5_ASAP7_75t_SL U63897 ( .A1(n63649), .A2(n63648), .B(n63652), .Y(
        n63793) );
  NAND2xp5_ASAP7_75t_SL U63898 ( .A(n75930), .B(n59165), .Y(n59416) );
  INVx1_ASAP7_75t_SL U63899 ( .A(n67940), .Y(n67941) );
  OAI22xp5_ASAP7_75t_SL U63900 ( .A1(n59192), .A2(n57156), .B1(n65053), .B2(
        n67974), .Y(n68164) );
  O2A1O1Ixp5_ASAP7_75t_SL U63901 ( .A1(n68265), .A2(n68267), .B(n68129), .C(
        n68130), .Y(n59270) );
  NAND2xp5_ASAP7_75t_SL U63902 ( .A(n67738), .B(n57394), .Y(n59149) );
  INVx1_ASAP7_75t_SL U63903 ( .A(n67552), .Y(n67554) );
  NOR2x1_ASAP7_75t_SL U63904 ( .A(n59967), .B(n59966), .Y(n77367) );
  OAI21xp5_ASAP7_75t_SL U63905 ( .A1(n60424), .A2(n59963), .B(n59962), .Y(
        n59967) );
  NAND2xp5_ASAP7_75t_SL U63906 ( .A(n2757), .B(n60401), .Y(n60317) );
  NAND2xp5_ASAP7_75t_SL U63907 ( .A(n4130), .B(n78261), .Y(icqmem_adr_qmem[14]) );
  INVx1_ASAP7_75t_SL U63908 ( .A(n69082), .Y(n58826) );
  INVx1_ASAP7_75t_SL U63909 ( .A(n66906), .Y(n66816) );
  NAND2xp5_ASAP7_75t_SL U63910 ( .A(n70782), .B(n70781), .Y(n70794) );
  NAND2xp5_ASAP7_75t_SL U63911 ( .A(n64798), .B(n75607), .Y(n64799) );
  INVx1_ASAP7_75t_SL U63912 ( .A(n75738), .Y(n75342) );
  OAI21xp5_ASAP7_75t_SL U63913 ( .A1(n59442), .A2(n57186), .B(n75917), .Y(
        n75983) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U63914 ( .A1(n59442), .A2(n57186), .B(n75917), 
        .C(n75980), .Y(n75920) );
  OAI21xp5_ASAP7_75t_SL U63915 ( .A1(n59559), .A2(n59020), .B(n62635), .Y(
        n68006) );
  OAI22xp5_ASAP7_75t_SL U63916 ( .A1(n62820), .A2(n62819), .B1(n62818), .B2(
        n62817), .Y(n62930) );
  NOR2x1_ASAP7_75t_SL U63917 ( .A(n59654), .B(n62757), .Y(n64025) );
  INVx1_ASAP7_75t_SL U63918 ( .A(n68054), .Y(n59177) );
  NAND2xp5_ASAP7_75t_SL U63919 ( .A(n59128), .B(n59127), .Y(n59126) );
  NAND2xp5_ASAP7_75t_SL U63920 ( .A(n67621), .B(n67447), .Y(n58967) );
  OAI22xp5_ASAP7_75t_SL U63921 ( .A1(n70180), .A2(n70179), .B1(n70178), .B2(
        n70177), .Y(n70181) );
  NOR2x1p5_ASAP7_75t_SL U63922 ( .A(n58729), .B(n58728), .Y(n58902) );
  BUFx3_ASAP7_75t_SL U63923 ( .A(n1819), .Y(n59543) );
  INVx1_ASAP7_75t_SL U63924 ( .A(n67670), .Y(n67674) );
  OAI21xp5_ASAP7_75t_SL U63925 ( .A1(n59654), .A2(n64509), .B(n58494), .Y(
        n58978) );
  AOI22xp5_ASAP7_75t_SL U63926 ( .A1(n68086), .A2(n63224), .B1(n63113), .B2(
        n57157), .Y(n63231) );
  NOR2x1p5_ASAP7_75t_SL U63927 ( .A(n58764), .B(n58763), .Y(n62558) );
  NOR2x1_ASAP7_75t_SL U63928 ( .A(n59414), .B(n58766), .Y(n58763) );
  INVx1_ASAP7_75t_SL U63929 ( .A(n67242), .Y(n59269) );
  INVx1_ASAP7_75t_SL U63930 ( .A(n66800), .Y(n66806) );
  INVx1_ASAP7_75t_SL U63931 ( .A(n63673), .Y(n63129) );
  NAND2xp5_ASAP7_75t_SL U63932 ( .A(n78206), .B(n4108), .Y(icqmem_adr_qmem[25]) );
  INVx1_ASAP7_75t_SL U63933 ( .A(n62774), .Y(n62776) );
  NOR2x1_ASAP7_75t_SL U63934 ( .A(n66663), .B(n66845), .Y(n66692) );
  NAND2xp5_ASAP7_75t_SL U63935 ( .A(n66692), .B(n66672), .Y(n66843) );
  NAND2x1p5_ASAP7_75t_SL U63936 ( .A(n58897), .B(n58405), .Y(n59610) );
  INVx1_ASAP7_75t_SL U63937 ( .A(n64920), .Y(n67475) );
  NAND2xp5_ASAP7_75t_SL U63938 ( .A(n2169), .B(n59559), .Y(n76204) );
  NOR2x1_ASAP7_75t_SL U63939 ( .A(n59719), .B(n59718), .Y(n75777) );
  AOI21xp5_ASAP7_75t_SL U63940 ( .A1(n76323), .A2(n59492), .B(n74032), .Y(
        n74038) );
  INVx1_ASAP7_75t_SL U63941 ( .A(n58943), .Y(n58832) );
  NAND2xp5_ASAP7_75t_SL U63942 ( .A(n66051), .B(n65968), .Y(n66078) );
  NOR2x1_ASAP7_75t_SL U63943 ( .A(n66049), .B(n65753), .Y(n65968) );
  NAND2xp5_ASAP7_75t_SL U63944 ( .A(n65482), .B(n65481), .Y(n65674) );
  NAND2x1_ASAP7_75t_SL U63945 ( .A(n67726), .B(n67727), .Y(n68353) );
  OAI21xp5_ASAP7_75t_SL U63946 ( .A1(n67699), .A2(n67698), .B(n56842), .Y(
        n67724) );
  NAND2xp5_ASAP7_75t_SL U63947 ( .A(n59640), .B(n67610), .Y(n67342) );
  OAI21xp5_ASAP7_75t_SL U63948 ( .A1(n74181), .A2(n74180), .B(n74144), .Y(
        n74191) );
  NAND2xp5_ASAP7_75t_SL U63949 ( .A(n73857), .B(n74303), .Y(n74305) );
  NAND2xp5_ASAP7_75t_SL U63950 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_3_), 
        .B(n74305), .Y(n74304) );
  INVx1_ASAP7_75t_SL U63951 ( .A(n67649), .Y(n67650) );
  XNOR2x1_ASAP7_75t_SL U63952 ( .A(n67651), .B(n67650), .Y(n67768) );
  NAND2xp5_ASAP7_75t_SL U63953 ( .A(n57078), .B(n57104), .Y(n66348) );
  OAI21xp5_ASAP7_75t_SL U63954 ( .A1(n66512), .A2(n66511), .B(n66371), .Y(
        n66439) );
  NAND2xp5_ASAP7_75t_SL U63955 ( .A(n53481), .B(n68327), .Y(n59489) );
  NOR2x1_ASAP7_75t_SL U63956 ( .A(n64734), .B(n64733), .Y(n74994) );
  INVx1_ASAP7_75t_SL U63957 ( .A(n64565), .Y(n64494) );
  NAND2xp5_ASAP7_75t_SL U63958 ( .A(n58025), .B(n64487), .Y(n64488) );
  NOR2x1_ASAP7_75t_SL U63959 ( .A(n66602), .B(n69301), .Y(n75059) );
  INVx1_ASAP7_75t_SL U63960 ( .A(n66586), .Y(n66536) );
  AOI22x1_ASAP7_75t_SL U63961 ( .A1(n67967), .A2(n66545), .B1(n66535), .B2(
        n67446), .Y(n66586) );
  INVx3_ASAP7_75t_SL U63962 ( .A(n59440), .Y(n67446) );
  INVx1_ASAP7_75t_SL U63963 ( .A(n66771), .Y(n66685) );
  INVx2_ASAP7_75t_SL U63964 ( .A(n67532), .Y(n67712) );
  BUFx3_ASAP7_75t_SL U63965 ( .A(n59609), .Y(n58931) );
  BUFx3_ASAP7_75t_SL U63966 ( .A(n1857), .Y(n59546) );
  INVx1_ASAP7_75t_SL U63967 ( .A(n70021), .Y(n69476) );
  INVx1_ASAP7_75t_SL U63968 ( .A(n68055), .Y(n67793) );
  NAND2x1p5_ASAP7_75t_SL U63969 ( .A(n66266), .B(n58791), .Y(n75894) );
  NAND2xp5_ASAP7_75t_SL U63970 ( .A(n57504), .B(n78167), .Y(n58791) );
  BUFx3_ASAP7_75t_SL U63971 ( .A(n59634), .Y(n59100) );
  OAI21xp5_ASAP7_75t_SL U63972 ( .A1(n58884), .A2(n58473), .B(n63093), .Y(
        n63132) );
  AOI21xp5_ASAP7_75t_SL U63973 ( .A1(n64507), .A2(n57214), .B(n62681), .Y(
        n75923) );
  INVx1_ASAP7_75t_SL U63974 ( .A(n63132), .Y(n63135) );
  NAND2xp5_ASAP7_75t_SL U63975 ( .A(n64944), .B(n64943), .Y(n64995) );
  OAI21xp5_ASAP7_75t_SL U63976 ( .A1(n64997), .A2(n64996), .B(n64995), .Y(
        n64998) );
  INVx1_ASAP7_75t_SL U63977 ( .A(n59031), .Y(n68421) );
  INVx1_ASAP7_75t_SL U63978 ( .A(n63644), .Y(n63607) );
  NAND2x1_ASAP7_75t_SL U63979 ( .A(n57113), .B(n57656), .Y(n67017) );
  AOI22xp5_ASAP7_75t_SL U63980 ( .A1(n67833), .A2(n67718), .B1(n57414), .B2(
        n68415), .Y(n68386) );
  INVx1_ASAP7_75t_SL U63981 ( .A(n63849), .Y(n63641) );
  NAND2xp5_ASAP7_75t_SL U63982 ( .A(n63633), .B(n63632), .Y(n63833) );
  OAI21xp5_ASAP7_75t_SL U63983 ( .A1(n66421), .A2(n66420), .B(n66484), .Y(
        n66492) );
  NAND2xp5_ASAP7_75t_SL U63984 ( .A(n67216), .B(n67215), .Y(n68693) );
  AOI22xp5_ASAP7_75t_SL U63985 ( .A1(n57163), .A2(n66455), .B1(n58336), .B2(
        n66461), .Y(n66491) );
  NAND2xp5_ASAP7_75t_SL U63986 ( .A(n58712), .B(n68110), .Y(n58714) );
  NAND2xp5_ASAP7_75t_SL U63987 ( .A(n75832), .B(n66300), .Y(n66303) );
  INVx1_ASAP7_75t_SL U63988 ( .A(n66303), .Y(n66311) );
  NAND2xp5_ASAP7_75t_SL U63989 ( .A(n77684), .B(n77683), .Y(or1200_du_N76) );
  INVx1_ASAP7_75t_SL U63990 ( .A(n68665), .Y(n58829) );
  O2A1O1Ixp5_ASAP7_75t_SL U63991 ( .A1(n67955), .A2(n68380), .B(n67954), .C(
        n67953), .Y(n68213) );
  NOR2x1_ASAP7_75t_SL U63992 ( .A(n67636), .B(n64684), .Y(n67635) );
  INVx1_ASAP7_75t_SL U63993 ( .A(n63165), .Y(n63168) );
  INVx1_ASAP7_75t_SL U63994 ( .A(n63059), .Y(n63061) );
  AOI21xp5_ASAP7_75t_SL U63995 ( .A1(n67452), .A2(n67451), .B(n67450), .Y(
        n67520) );
  OAI22xp5_ASAP7_75t_SL U63996 ( .A1(n67540), .A2(n67539), .B1(n67655), .B2(
        n67547), .Y(n67524) );
  INVx1_ASAP7_75t_SL U63997 ( .A(n67523), .Y(n67547) );
  OAI21xp5_ASAP7_75t_SL U63998 ( .A1(n64449), .A2(n53233), .B(n64686), .Y(
        n64465) );
  OAI21xp5_ASAP7_75t_SL U63999 ( .A1(n53233), .A2(n64687), .B(n64686), .Y(
        n64690) );
  NOR2x1_ASAP7_75t_SL U64000 ( .A(n64751), .B(n65122), .Y(n65115) );
  INVx2_ASAP7_75t_SL U64001 ( .A(n57500), .Y(n62738) );
  INVx1_ASAP7_75t_SL U64002 ( .A(n67779), .Y(n67780) );
  OAI21xp5_ASAP7_75t_SL U64003 ( .A1(n67438), .A2(n59491), .B(n58965), .Y(
        n67620) );
  OAI21xp5_ASAP7_75t_SL U64004 ( .A1(n69023), .A2(n69022), .B(n69021), .Y(
        n69112) );
  AOI21xp5_ASAP7_75t_SL U64005 ( .A1(n75291), .A2(n69211), .B(n69207), .Y(
        n74572) );
  NAND2x1_ASAP7_75t_SL U64006 ( .A(n59565), .B(n56861), .Y(n62591) );
  NAND2xp5_ASAP7_75t_SL U64007 ( .A(n58482), .B(n58802), .Y(n58646) );
  OAI21xp5_ASAP7_75t_SL U64008 ( .A1(n77013), .A2(n59843), .B(n59726), .Y(
        n77293) );
  NAND2xp5_ASAP7_75t_SL U64009 ( .A(n2157), .B(n59545), .Y(n76199) );
  NAND2xp5_ASAP7_75t_SL U64010 ( .A(n77732), .B(n61969), .Y(n66298) );
  NAND2xp5_ASAP7_75t_SL U64011 ( .A(n66298), .B(n66297), .Y(n64917) );
  NAND2xp5_ASAP7_75t_SL U64012 ( .A(n74936), .B(n74935), .Y(n63710) );
  NOR2x1p5_ASAP7_75t_SL U64013 ( .A(n57090), .B(n78009), .Y(n77374) );
  INVx1_ASAP7_75t_SL U64014 ( .A(n73960), .Y(n76658) );
  XNOR2x1_ASAP7_75t_SL U64015 ( .A(n68325), .B(n68326), .Y(n58687) );
  NAND2xp5_ASAP7_75t_SL U64016 ( .A(n77730), .B(n67354), .Y(n64649) );
  INVx1_ASAP7_75t_SL U64017 ( .A(n59070), .Y(n62656) );
  NAND2xp5_ASAP7_75t_SL U64018 ( .A(n73964), .B(n77217), .Y(n74036) );
  FAx1_ASAP7_75t_SL U64019 ( .A(n75793), .B(n59753), .CI(n59752), .CON(), .SN(
        n59754) );
  AOI21xp5_ASAP7_75t_SL U64020 ( .A1(n75792), .A2(n59751), .B(n75188), .Y(
        n59752) );
  NAND2xp5_ASAP7_75t_SL U64021 ( .A(n67553), .B(n67554), .Y(n67672) );
  AOI21xp5_ASAP7_75t_SL U64022 ( .A1(n75900), .A2(n59601), .B(n67385), .Y(
        n67402) );
  INVx1_ASAP7_75t_SL U64023 ( .A(n63805), .Y(n63665) );
  NOR2x1_ASAP7_75t_SL U64024 ( .A(n68008), .B(n67607), .Y(n58929) );
  AOI22xp5_ASAP7_75t_SL U64025 ( .A1(n53197), .A2(n67226), .B1(n67829), .B2(
        n67225), .Y(n67346) );
  OAI22xp5_ASAP7_75t_SL U64026 ( .A1(n66933), .A2(n59440), .B1(n66789), .B2(
        n59446), .Y(n68461) );
  NOR2x1_ASAP7_75t_SL U64027 ( .A(n76814), .B(n76815), .Y(n76813) );
  INVx1_ASAP7_75t_SL U64028 ( .A(n68203), .Y(n59303) );
  NOR2x1_ASAP7_75t_SL U64029 ( .A(n64751), .B(n64730), .Y(n64741) );
  NOR2x1_ASAP7_75t_SL U64030 ( .A(n66656), .B(n66421), .Y(n67096) );
  NOR2x1_ASAP7_75t_SL U64031 ( .A(n59598), .B(n59502), .Y(n58659) );
  NOR2x1_ASAP7_75t_SL U64032 ( .A(n61963), .B(n59546), .Y(n64482) );
  AOI21xp5_ASAP7_75t_SL U64033 ( .A1(n57186), .A2(n64482), .B(n66451), .Y(
        n64924) );
  NAND2xp5_ASAP7_75t_SL U64034 ( .A(n59986), .B(n60031), .Y(n60029) );
  NAND2xp5_ASAP7_75t_SL U64035 ( .A(n57100), .B(n77382), .Y(n4095) );
  OAI21xp5_ASAP7_75t_SL U64036 ( .A1(n58884), .A2(n67270), .B(n67269), .Y(
        n67296) );
  NAND2xp5_ASAP7_75t_SL U64037 ( .A(n2095), .B(n59541), .Y(n59941) );
  INVx2_ASAP7_75t_SL U64038 ( .A(n59662), .Y(n59190) );
  OAI21xp5_ASAP7_75t_SL U64039 ( .A1(n68011), .A2(n59664), .B(n59190), .Y(
        n67233) );
  INVx1_ASAP7_75t_SL U64040 ( .A(n64999), .Y(n64978) );
  INVx1_ASAP7_75t_SL U64041 ( .A(n63882), .Y(n63884) );
  INVx1_ASAP7_75t_SL U64042 ( .A(n63105), .Y(n63107) );
  XNOR2x1_ASAP7_75t_SL U64043 ( .A(n59355), .B(n59354), .Y(n68568) );
  INVx1_ASAP7_75t_SL U64044 ( .A(n67816), .Y(n67818) );
  AOI31xp67_ASAP7_75t_SL U64045 ( .A1(n70804), .A2(n70803), .A3(n70802), .B(
        n70801), .Y(n70841) );
  NAND2xp5_ASAP7_75t_SL U64046 ( .A(n71309), .B(n71350), .Y(n71325) );
  AOI22xp5_ASAP7_75t_SL U64047 ( .A1(n70725), .A2(n70931), .B1(n70724), .B2(
        n70985), .Y(n70743) );
  INVx1_ASAP7_75t_SL U64048 ( .A(n58328), .Y(n70985) );
  NAND2x1p5_ASAP7_75t_SL U64049 ( .A(n69026), .B(n68698), .Y(n69116) );
  AOI21xp5_ASAP7_75t_SL U64050 ( .A1(n66973), .A2(n53496), .B(n66971), .Y(
        n66974) );
  NOR2x1_ASAP7_75t_SL U64051 ( .A(n68350), .B(n68349), .Y(n68805) );
  NOR2x2_ASAP7_75t_SL U64052 ( .A(n59199), .B(n59198), .Y(n67846) );
  INVx2_ASAP7_75t_SL U64053 ( .A(n62749), .Y(n59198) );
  NAND2xp5_ASAP7_75t_SL U64054 ( .A(n59197), .B(n59411), .Y(n59199) );
  OAI21xp5_ASAP7_75t_SL U64055 ( .A1(n62671), .A2(n57122), .B(n59553), .Y(
        n59411) );
  OAI22xp5_ASAP7_75t_SL U64056 ( .A1(n67742), .A2(n59454), .B1(n57099), .B2(
        n67568), .Y(n67689) );
  INVx1_ASAP7_75t_SL U64057 ( .A(n67671), .Y(n67675) );
  NAND2xp5_ASAP7_75t_SL U64058 ( .A(n59263), .B(n61931), .Y(n59262) );
  NOR2x1_ASAP7_75t_SL U64059 ( .A(n68298), .B(n68300), .Y(n68324) );
  INVx1_ASAP7_75t_SL U64060 ( .A(n68178), .Y(n58742) );
  AOI22xp5_ASAP7_75t_SL U64061 ( .A1(n67842), .A2(n67843), .B1(n57380), .B2(
        n67844), .Y(n68178) );
  O2A1O1Ixp5_ASAP7_75t_SL U64062 ( .A1(n75922), .A2(n67738), .B(n63664), .C(
        n67898), .Y(n63800) );
  NOR2x1_ASAP7_75t_SL U64063 ( .A(n57234), .B(n64033), .Y(n67560) );
  NAND2xp5_ASAP7_75t_SL U64064 ( .A(n59455), .B(n64032), .Y(n64033) );
  INVx1_ASAP7_75t_SL U64065 ( .A(n68382), .Y(n66793) );
  OAI21xp5_ASAP7_75t_SL U64066 ( .A1(n75899), .A2(n67431), .B(n66632), .Y(
        n66633) );
  NAND2xp5_ASAP7_75t_SL U64067 ( .A(n60936), .B(n60935), .Y(n61228) );
  INVx1_ASAP7_75t_SL U64068 ( .A(n68499), .Y(n68457) );
  INVx1_ASAP7_75t_SL U64069 ( .A(n68495), .Y(n68475) );
  NAND2xp5_ASAP7_75t_SL U64070 ( .A(n58650), .B(n58649), .Y(n64026) );
  OAI22xp5_ASAP7_75t_SL U64071 ( .A1(n67752), .A2(n58658), .B1(n59491), .B2(
        n67753), .Y(n68391) );
  INVx1_ASAP7_75t_SL U64072 ( .A(n58754), .Y(n68028) );
  NAND2xp5_ASAP7_75t_SL U64073 ( .A(n67699), .B(n67698), .Y(n68419) );
  OAI21xp5_ASAP7_75t_SL U64074 ( .A1(n59607), .A2(n59510), .B(n66917), .Y(
        n67413) );
  INVx1_ASAP7_75t_SL U64075 ( .A(n66991), .Y(n66894) );
  NOR2x1_ASAP7_75t_SL U64076 ( .A(n66890), .B(n67027), .Y(n66991) );
  INVx1_ASAP7_75t_SL U64077 ( .A(n53612), .Y(n67431) );
  OAI21xp5_ASAP7_75t_SL U64078 ( .A1(n67434), .A2(n67097), .B(n66881), .Y(
        n67023) );
  OAI21xp5_ASAP7_75t_SL U64079 ( .A1(n53275), .A2(n67431), .B(n66880), .Y(
        n66881) );
  INVx1_ASAP7_75t_SL U64080 ( .A(n58842), .Y(n75473) );
  NAND2xp5_ASAP7_75t_SL U64081 ( .A(n66328), .B(n66327), .Y(n66329) );
  INVx1_ASAP7_75t_SL U64082 ( .A(n66591), .Y(n66563) );
  NOR2x1_ASAP7_75t_SL U64083 ( .A(n65107), .B(n65108), .Y(n68338) );
  NAND2x1p5_ASAP7_75t_SL U64084 ( .A(n64869), .B(n59281), .Y(n68735) );
  INVx1_ASAP7_75t_SL U64085 ( .A(n67833), .Y(n66829) );
  NAND2xp5_ASAP7_75t_SL U64086 ( .A(n77735), .B(n66297), .Y(n65017) );
  NAND2xp5_ASAP7_75t_SL U64087 ( .A(n58733), .B(n68345), .Y(n58732) );
  AOI21xp5_ASAP7_75t_SL U64088 ( .A1(n75918), .A2(n75917), .B(n75984), .Y(
        n75919) );
  NOR2x1_ASAP7_75t_SL U64089 ( .A(n57077), .B(n57133), .Y(n76004) );
  NAND2xp5_ASAP7_75t_SL U64090 ( .A(n75934), .B(n75945), .Y(n76166) );
  NAND2xp5_ASAP7_75t_SL U64091 ( .A(n76124), .B(n75933), .Y(n75945) );
  NAND2xp5_ASAP7_75t_SL U64092 ( .A(n59513), .B(n75921), .Y(n75988) );
  NAND2xp5_ASAP7_75t_SL U64093 ( .A(n59594), .B(n57941), .Y(n67458) );
  INVx1_ASAP7_75t_SL U64094 ( .A(n67537), .Y(n67690) );
  AOI21xp5_ASAP7_75t_SL U64095 ( .A1(n69138), .A2(n53500), .B(n66989), .Y(
        n69137) );
  INVx1_ASAP7_75t_SL U64096 ( .A(n58952), .Y(n58951) );
  INVx2_ASAP7_75t_SL U64097 ( .A(n58753), .Y(n66758) );
  AOI21xp5_ASAP7_75t_SL U64098 ( .A1(n78067), .A2(n60297), .B(n60296), .Y(
        n60298) );
  NAND2xp5_ASAP7_75t_SL U64099 ( .A(n60325), .B(n60311), .Y(n60401) );
  AOI21xp5_ASAP7_75t_SL U64100 ( .A1(n75644), .A2(n57310), .B(n66697), .Y(
        n67059) );
  NAND2xp5_ASAP7_75t_SL U64101 ( .A(n66254), .B(n66263), .Y(n59487) );
  OAI22xp5_ASAP7_75t_SL U64102 ( .A1(n67284), .A2(n66698), .B1(n67059), .B2(
        n75032), .Y(n66875) );
  OAI21x1_ASAP7_75t_SL U64103 ( .A1(n58775), .A2(n57441), .B(n66299), .Y(
        n67713) );
  INVx1_ASAP7_75t_SL U64104 ( .A(n67881), .Y(n66299) );
  INVx1_ASAP7_75t_SL U64105 ( .A(n65808), .Y(n65828) );
  OAI21x1_ASAP7_75t_SL U64106 ( .A1(n74208), .A2(n76976), .B(n65669), .Y(
        n65808) );
  NAND2xp5_ASAP7_75t_SL U64107 ( .A(n74206), .B(n76976), .Y(n65669) );
  OAI22xp5_ASAP7_75t_SL U64108 ( .A1(n67414), .A2(n66295), .B1(n59446), .B2(
        n59417), .Y(n66390) );
  AOI22xp5_ASAP7_75t_SL U64109 ( .A1(n67363), .A2(n57358), .B1(n57273), .B2(
        n59047), .Y(n67379) );
  BUFx3_ASAP7_75t_SL U64110 ( .A(n1656), .Y(n59534) );
  OAI21x1_ASAP7_75t_SL U64111 ( .A1(n59578), .A2(n58409), .B(n66452), .Y(
        n67467) );
  INVx1_ASAP7_75t_SL U64112 ( .A(n67379), .Y(n67651) );
  NAND2xp5_ASAP7_75t_SL U64113 ( .A(n67846), .B(n59600), .Y(n67389) );
  NOR2x1_ASAP7_75t_SL U64114 ( .A(n66676), .B(n66675), .Y(n67077) );
  INVx1_ASAP7_75t_SL U64115 ( .A(n64506), .Y(n64950) );
  INVx1_ASAP7_75t_SL U64116 ( .A(n67179), .Y(n67191) );
  NAND2x1_ASAP7_75t_SL U64117 ( .A(n59573), .B(n59574), .Y(n61214) );
  NAND2xp5_ASAP7_75t_SL U64118 ( .A(n57016), .B(n58708), .Y(n58710) );
  BUFx3_ASAP7_75t_SL U64119 ( .A(n2862), .Y(n59574) );
  XNOR2x1_ASAP7_75t_SL U64120 ( .A(n67814), .B(n67813), .Y(n59311) );
  NAND2xp5_ASAP7_75t_SL U64121 ( .A(n71127), .B(n71122), .Y(n71123) );
  NAND2xp5_ASAP7_75t_SL U64122 ( .A(n71132), .B(n71114), .Y(n71122) );
  AOI22xp5_ASAP7_75t_SL U64123 ( .A1(n58314), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[23]), .B1(n70681), 
        .B2(n70680), .Y(n70682) );
  INVx1_ASAP7_75t_SL U64124 ( .A(n67422), .Y(n67423) );
  NAND2xp5_ASAP7_75t_SL U64125 ( .A(n68484), .B(n68483), .Y(n68532) );
  NAND2x1_ASAP7_75t_SL U64126 ( .A(n59424), .B(n61914), .Y(n76430) );
  NOR2x1_ASAP7_75t_SL U64127 ( .A(n59367), .B(n59366), .Y(n64711) );
  NAND2x1p5_ASAP7_75t_SL U64128 ( .A(n77242), .B(n57117), .Y(n76679) );
  INVx4_ASAP7_75t_SL U64129 ( .A(n59565), .Y(n77242) );
  NAND2xp5_ASAP7_75t_SL U64130 ( .A(n65814), .B(n65813), .Y(n66007) );
  NAND2xp5_ASAP7_75t_SL U64131 ( .A(n59657), .B(n67639), .Y(n67879) );
  INVx1_ASAP7_75t_SL U64132 ( .A(n59036), .Y(n68115) );
  NAND2xp5_ASAP7_75t_SL U64133 ( .A(n67880), .B(n58716), .Y(n59360) );
  NAND2xp5_ASAP7_75t_SL U64134 ( .A(n58630), .B(n58629), .Y(n58716) );
  NAND2xp5_ASAP7_75t_SL U64135 ( .A(n58750), .B(n58749), .Y(n67880) );
  NOR2x1_ASAP7_75t_SL U64136 ( .A(n59508), .B(n59466), .Y(n66618) );
  AOI21xp5_ASAP7_75t_SL U64137 ( .A1(n68065), .A2(n58963), .B(n67886), .Y(
        n67887) );
  NOR2x1p5_ASAP7_75t_SL U64138 ( .A(n66618), .B(n59619), .Y(n67829) );
  INVx1_ASAP7_75t_SL U64139 ( .A(n64601), .Y(n64542) );
  NOR2x1_ASAP7_75t_SL U64140 ( .A(n64597), .B(n59240), .Y(n64601) );
  OAI21xp5_ASAP7_75t_SL U64141 ( .A1(n64410), .A2(n57158), .B(n64536), .Y(
        n64599) );
  NAND2xp5_ASAP7_75t_SL U64142 ( .A(n58155), .B(n64409), .Y(n64536) );
  OAI21xp5_ASAP7_75t_SL U64143 ( .A1(n70604), .A2(n70603), .B(n70602), .Y(
        n70610) );
  NOR2x1_ASAP7_75t_SL U64144 ( .A(n74383), .B(n74384), .Y(n74390) );
  NAND2xp5_ASAP7_75t_SL U64145 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_13_), .B(
        n74346), .Y(n74384) );
  NOR2x1_ASAP7_75t_SL U64146 ( .A(n76947), .B(n76962), .Y(n76934) );
  NAND2xp5_ASAP7_75t_SL U64147 ( .A(n74850), .B(n74901), .Y(n74904) );
  AOI21xp5_ASAP7_75t_SL U64148 ( .A1(n75901), .A2(n59600), .B(n67305), .Y(
        n67439) );
  INVx1_ASAP7_75t_SL U64149 ( .A(n68541), .Y(n68540) );
  INVx1_ASAP7_75t_SL U64150 ( .A(n59169), .Y(n67841) );
  BUFx2_ASAP7_75t_SL U64151 ( .A(n64368), .Y(n59488) );
  OAI21xp5_ASAP7_75t_SL U64152 ( .A1(n68417), .A2(n57029), .B(n68416), .Y(
        n68469) );
  INVx1_ASAP7_75t_SL U64153 ( .A(n77855), .Y(n76989) );
  OAI21xp5_ASAP7_75t_SL U64154 ( .A1(or1200_cpu_or1200_mult_mac_n124), .A2(
        n61826), .B(n60804), .Y(n61229) );
  OAI21xp5_ASAP7_75t_SL U64155 ( .A1(n74036), .A2(n74038), .B(n74035), .Y(
        or1200_cpu_or1200_except_n1742) );
  NAND2x1p5_ASAP7_75t_SL U64156 ( .A(n68591), .B(n69037), .Y(n69026) );
  XNOR2x2_ASAP7_75t_SL U64157 ( .A(n66952), .B(n66951), .Y(n68500) );
  OAI21xp5_ASAP7_75t_SL U64158 ( .A1(n59014), .A2(n68551), .B(n59015), .Y(
        n69034) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64159 ( .A1(n69149), .A2(n53206), .B(n57369), 
        .C(n69146), .Y(n69150) );
  INVx1_ASAP7_75t_SL U64160 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[11]), .Y(
        n73171) );
  OAI21xp5_ASAP7_75t_SL U64161 ( .A1(n4092), .A2(n77801), .B(n77800), .Y(n9472) );
  INVx2_ASAP7_75t_SL U64162 ( .A(n67930), .Y(n67990) );
  NAND2xp5_ASAP7_75t_SL U64163 ( .A(n75312), .B(n75313), .Y(n75311) );
  NAND2x1_ASAP7_75t_SL U64164 ( .A(n2073), .B(n59570), .Y(n59945) );
  INVx1_ASAP7_75t_SL U64165 ( .A(n62594), .Y(n62637) );
  INVx1_ASAP7_75t_SL U64166 ( .A(n62947), .Y(n63364) );
  BUFx6f_ASAP7_75t_SL U64167 ( .A(n66450), .Y(n59588) );
  INVx3_ASAP7_75t_SL U64168 ( .A(n59593), .Y(n59595) );
  OAI22xp5_ASAP7_75t_SL U64169 ( .A1(n63344), .A2(n62951), .B1(n62950), .B2(
        n62949), .Y(n63365) );
  NAND2xp5_ASAP7_75t_SL U64170 ( .A(n59595), .B(n67638), .Y(n62843) );
  INVx1_ASAP7_75t_SL U64171 ( .A(n68244), .Y(n68248) );
  INVx1_ASAP7_75t_SL U64172 ( .A(n68136), .Y(n68138) );
  INVx2_ASAP7_75t_SL U64173 ( .A(n1571), .Y(n77735) );
  INVx2_ASAP7_75t_SL U64174 ( .A(n59670), .Y(n58962) );
  NAND2xp5_ASAP7_75t_SL U64175 ( .A(n70182), .B(n70181), .Y(n70187) );
  NAND2xp5_ASAP7_75t_SL U64176 ( .A(n2461), .B(n59557), .Y(n76200) );
  INVx1_ASAP7_75t_SL U64177 ( .A(n76820), .Y(n77385) );
  NOR2x1_ASAP7_75t_SL U64178 ( .A(n59703), .B(n77249), .Y(n76820) );
  AOI22xp5_ASAP7_75t_SL U64179 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[1]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[0]), .B2(n57194), 
        .Y(n66080) );
  NAND2xp5_ASAP7_75t_SL U64180 ( .A(n67618), .B(n67619), .Y(n58969) );
  INVx1_ASAP7_75t_SL U64181 ( .A(n66271), .Y(n66256) );
  INVx1_ASAP7_75t_SL U64182 ( .A(n63605), .Y(n63606) );
  NAND2xp5_ASAP7_75t_SL U64183 ( .A(n67486), .B(n67485), .Y(n58971) );
  NAND2x1p5_ASAP7_75t_SL U64184 ( .A(n59323), .B(n59324), .Y(n66260) );
  INVx2_ASAP7_75t_SL U64185 ( .A(n58431), .Y(n75925) );
  XNOR2x2_ASAP7_75t_SL U64186 ( .A(n67208), .B(n67207), .Y(n75274) );
  BUFx3_ASAP7_75t_SL U64187 ( .A(n1640), .Y(n59532) );
  AOI21xp5_ASAP7_75t_SL U64188 ( .A1(n67196), .A2(n67195), .B(n67194), .Y(
        n67164) );
  NOR2x1_ASAP7_75t_SL U64189 ( .A(n74781), .B(n66635), .Y(n66638) );
  INVx1_ASAP7_75t_SL U64190 ( .A(n66634), .Y(n66635) );
  NAND2xp5_ASAP7_75t_SL U64191 ( .A(n53619), .B(n67489), .Y(n67729) );
  NAND2xp5_ASAP7_75t_SL U64192 ( .A(n67251), .B(n64626), .Y(n64485) );
  NOR2x1_ASAP7_75t_SL U64193 ( .A(n62591), .B(n76690), .Y(n62594) );
  O2A1O1Ixp5_ASAP7_75t_SL U64194 ( .A1(n67679), .A2(n67678), .B(n67677), .C(
        n67676), .Y(n68396) );
  AOI21xp5_ASAP7_75t_SL U64195 ( .A1(n67674), .A2(n67675), .B(n67673), .Y(
        n67677) );
  INVx1_ASAP7_75t_SL U64196 ( .A(n68904), .Y(n58887) );
  NAND2xp5_ASAP7_75t_SL U64197 ( .A(n59554), .B(n59543), .Y(n60737) );
  INVx1_ASAP7_75t_SL U64198 ( .A(n67353), .Y(n58923) );
  OAI22xp5_ASAP7_75t_SL U64199 ( .A1(n58402), .A2(n67971), .B1(n58232), .B2(
        n67972), .Y(n67561) );
  NAND2xp5_ASAP7_75t_SL U64200 ( .A(n65107), .B(n65108), .Y(n64739) );
  NOR2x1_ASAP7_75t_SL U64201 ( .A(n58647), .B(n62748), .Y(n67308) );
  AOI22xp5_ASAP7_75t_SL U64202 ( .A1(n58672), .A2(n57180), .B1(n59670), .B2(
        n58439), .Y(n59109) );
  OAI21xp5_ASAP7_75t_SL U64203 ( .A1(n68233), .A2(n58369), .B(n68231), .Y(
        n68237) );
  INVx2_ASAP7_75t_SL U64204 ( .A(n67805), .Y(n67984) );
  NAND2xp5_ASAP7_75t_SL U64205 ( .A(n69916), .B(n69915), .Y(n69963) );
  OAI21xp5_ASAP7_75t_SL U64206 ( .A1(n69862), .A2(n69861), .B(n69860), .Y(
        n69914) );
  AOI21xp5_ASAP7_75t_SL U64207 ( .A1(n69835), .A2(n69834), .B(n69833), .Y(
        n69861) );
  INVx1_ASAP7_75t_SL U64208 ( .A(n59519), .Y(n68602) );
  BUFx3_ASAP7_75t_SL U64209 ( .A(n68408), .Y(n59519) );
  NAND2xp5_ASAP7_75t_SL U64210 ( .A(n60554), .B(n59971), .Y(n61248) );
  NAND2x1_ASAP7_75t_SL U64211 ( .A(n2056), .B(n59538), .Y(n77011) );
  NAND2xp5_ASAP7_75t_SL U64212 ( .A(n2039), .B(n59560), .Y(n59926) );
  AOI21xp5_ASAP7_75t_SL U64213 ( .A1(n77584), .A2(n77128), .B(n60699), .Y(
        n61021) );
  NAND2xp5_ASAP7_75t_SL U64214 ( .A(n62052), .B(n60716), .Y(n77173) );
  NOR2x1_ASAP7_75t_SL U64215 ( .A(n62355), .B(n75841), .Y(n62519) );
  NAND2x1p5_ASAP7_75t_SL U64216 ( .A(n59708), .B(n59558), .Y(n62355) );
  NAND2xp5_ASAP7_75t_SL U64217 ( .A(n73557), .B(n73556), .Y(n73574) );
  NAND2xp5_ASAP7_75t_SL U64218 ( .A(n73537), .B(n73536), .Y(n73544) );
  NAND2xp5_ASAP7_75t_SL U64219 ( .A(n73593), .B(n73583), .Y(n73582) );
  NAND2xp5_ASAP7_75t_SL U64220 ( .A(n3331), .B(n73708), .Y(n73528) );
  NAND2xp5_ASAP7_75t_SL U64221 ( .A(n1900), .B(n59535), .Y(n75299) );
  OAI21xp5_ASAP7_75t_SL U64222 ( .A1(n63652), .A2(n63651), .B(n63650), .Y(
        n63794) );
  NAND2xp5_ASAP7_75t_SL U64223 ( .A(n63234), .B(n63233), .Y(n63645) );
  OAI21xp5_ASAP7_75t_SL U64224 ( .A1(n63122), .A2(n67315), .B(n63121), .Y(
        n63233) );
  INVx2_ASAP7_75t_SL U64225 ( .A(n57182), .Y(n59468) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64226 ( .A1(n59578), .A2(n75734), .B(n75338), 
        .C(n59561), .Y(n64309) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64227 ( .A1(n59532), .A2(n75734), .B(n75338), 
        .C(n59531), .Y(n74613) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64228 ( .A1(n59582), .A2(n75734), .B(n75338), 
        .C(n59579), .Y(n61892) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64229 ( .A1(n57312), .A2(n75734), .B(n75338), 
        .C(n59486), .Y(n62516) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64230 ( .A1(n59563), .A2(n75595), .B(n75593), 
        .C(n75872), .Y(n75597) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64231 ( .A1(n59536), .A2(n75734), .B(n75338), 
        .C(n59535), .Y(n75339) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64232 ( .A1(n59552), .A2(n75734), .B(n62340), 
        .C(n59560), .Y(n60867) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64233 ( .A1(n59569), .A2(n75734), .B(n64830), 
        .C(n59554), .Y(n62337) );
  NAND2xp5_ASAP7_75t_SL U64234 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_24_), .B(
        n74298), .Y(n74332) );
  OAI21xp5_ASAP7_75t_SL U64235 ( .A1(n74295), .A2(n74297), .B(n72560), .Y(
        n74298) );
  INVx1_ASAP7_75t_SL U64236 ( .A(n64368), .Y(n64358) );
  INVx1_ASAP7_75t_SL U64237 ( .A(n68542), .Y(n68545) );
  NAND2xp5_ASAP7_75t_SL U64238 ( .A(n59357), .B(n59608), .Y(n67908) );
  OAI21xp5_ASAP7_75t_SL U64239 ( .A1(n76279), .A2(n62295), .B(n60771), .Y(
        n62309) );
  NAND2xp5_ASAP7_75t_SL U64240 ( .A(n59545), .B(n60768), .Y(n62295) );
  INVx1_ASAP7_75t_SL U64241 ( .A(n65003), .Y(n64977) );
  INVx1_ASAP7_75t_SL U64242 ( .A(n67962), .Y(n76077) );
  NOR2x1p5_ASAP7_75t_SL U64243 ( .A(n58882), .B(n64025), .Y(n65034) );
  OAI21xp5_ASAP7_75t_SL U64244 ( .A1(n68688), .A2(n59449), .B(n74111), .Y(
        n68689) );
  INVx1_ASAP7_75t_SL U64245 ( .A(n58903), .Y(n66794) );
  NAND2x1p5_ASAP7_75t_SL U64246 ( .A(n67356), .B(n64649), .Y(n75897) );
  INVx1_ASAP7_75t_SL U64247 ( .A(n67843), .Y(n68123) );
  XOR2x2_ASAP7_75t_SL U64248 ( .A(n68190), .B(n68189), .Y(n58452) );
  NAND2xp5_ASAP7_75t_SL U64249 ( .A(n68707), .B(n68714), .Y(n58772) );
  INVx1_ASAP7_75t_SL U64250 ( .A(n68534), .Y(n66976) );
  NAND2xp5_ASAP7_75t_SL U64251 ( .A(n65342), .B(n65337), .Y(n65344) );
  NOR2x1_ASAP7_75t_SL U64252 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_18_), .B(n65375), .Y(
        n65337) );
  INVx1_ASAP7_75t_SL U64253 ( .A(n64983), .Y(n59281) );
  AOI21xp5_ASAP7_75t_SL U64254 ( .A1(n59087), .A2(n64589), .B(n58994), .Y(
        n58993) );
  NAND2xp5_ASAP7_75t_SL U64255 ( .A(n68235), .B(n68234), .Y(n68029) );
  INVx4_ASAP7_75t_SL U64256 ( .A(n59605), .Y(n59604) );
  INVx1_ASAP7_75t_SL U64257 ( .A(n64948), .Y(n64949) );
  OAI21xp5_ASAP7_75t_SL U64258 ( .A1(n64951), .A2(n64648), .B(n64948), .Y(
        n59050) );
  INVx1_ASAP7_75t_SL U64259 ( .A(n68316), .Y(n68317) );
  NAND2x1_ASAP7_75t_SL U64260 ( .A(n67646), .B(n67647), .Y(n67802) );
  INVx1_ASAP7_75t_SL U64261 ( .A(n64658), .Y(n64660) );
  AOI21xp5_ASAP7_75t_SL U64262 ( .A1(n67663), .A2(n68054), .B(n67662), .Y(
        n67664) );
  INVx2_ASAP7_75t_SL U64263 ( .A(n59548), .Y(n74781) );
  BUFx3_ASAP7_75t_SL U64264 ( .A(n1865), .Y(n59548) );
  INVx2_ASAP7_75t_SL U64265 ( .A(n67657), .Y(n67655) );
  NOR2x1_ASAP7_75t_SL U64266 ( .A(n59377), .B(n59375), .Y(n67657) );
  AOI21xp5_ASAP7_75t_SL U64267 ( .A1(n73478), .A2(n73252), .B(n73251), .Y(
        n73469) );
  OAI22xp5_ASAP7_75t_SL U64268 ( .A1(n73472), .A2(n73473), .B1(n73250), .B2(
        n73249), .Y(n73251) );
  OAI21xp5_ASAP7_75t_SL U64269 ( .A1(n59631), .A2(n73227), .B(n73226), .Y(
        n73235) );
  INVx1_ASAP7_75t_SL U64270 ( .A(n68585), .Y(n74556) );
  INVx1_ASAP7_75t_SL U64271 ( .A(n75096), .Y(n75097) );
  BUFx6f_ASAP7_75t_SL U64272 ( .A(n2949), .Y(n59578) );
  INVx1_ASAP7_75t_SL U64273 ( .A(n63608), .Y(n63611) );
  OAI21xp5_ASAP7_75t_SL U64274 ( .A1(n67944), .A2(n59230), .B(n63213), .Y(
        n63630) );
  NAND2xp5_ASAP7_75t_SL U64275 ( .A(n75930), .B(n59230), .Y(n63213) );
  INVx2_ASAP7_75t_SL U64276 ( .A(n59464), .Y(n60623) );
  INVx4_ASAP7_75t_SL U64277 ( .A(n59602), .Y(n59230) );
  INVx1_ASAP7_75t_SL U64278 ( .A(n68392), .Y(n59000) );
  INVx1_ASAP7_75t_SL U64279 ( .A(n68510), .Y(n68511) );
  OAI22xp5_ASAP7_75t_SL U64280 ( .A1(n59468), .A2(n67467), .B1(n67963), .B2(
        n67383), .Y(n67515) );
  NAND2xp5_ASAP7_75t_SL U64281 ( .A(n62903), .B(n62902), .Y(n63310) );
  INVx3_ASAP7_75t_SL U64282 ( .A(n59442), .Y(n59443) );
  XNOR2x2_ASAP7_75t_SL U64283 ( .A(n58441), .B(n68207), .Y(n68300) );
  OAI21xp5_ASAP7_75t_SL U64284 ( .A1(n59466), .A2(n68087), .B(n64938), .Y(
        n67843) );
  INVx1_ASAP7_75t_SL U64285 ( .A(n64712), .Y(n64722) );
  NAND2xp5_ASAP7_75t_SL U64286 ( .A(n53219), .B(n64030), .Y(n63862) );
  INVx1_ASAP7_75t_SL U64287 ( .A(n68222), .Y(n65008) );
  NAND2xp5_ASAP7_75t_SL U64288 ( .A(n64929), .B(n67322), .Y(n65005) );
  BUFx6f_ASAP7_75t_SL U64289 ( .A(n58143), .Y(n58863) );
  INVx1_ASAP7_75t_SL U64290 ( .A(n66910), .Y(n58722) );
  NAND2xp5_ASAP7_75t_SL U64291 ( .A(n71386), .B(n58312), .Y(n71372) );
  NAND2x1p5_ASAP7_75t_SL U64292 ( .A(n59508), .B(n59467), .Y(n67826) );
  XNOR2x1_ASAP7_75t_SL U64293 ( .A(n58435), .B(n59120), .Y(n68516) );
  XNOR2x2_ASAP7_75t_SL U64294 ( .A(n59456), .B(n75947), .Y(n66930) );
  NAND2xp5_ASAP7_75t_SL U64295 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_16_), 
        .B(n74394), .Y(n74405) );
  NOR2x1_ASAP7_75t_SL U64296 ( .A(n74386), .B(n74387), .Y(n74394) );
  NAND2xp5_ASAP7_75t_SL U64297 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_7_), 
        .B(n74373), .Y(n74372) );
  INVx2_ASAP7_75t_SL U64298 ( .A(n59502), .Y(n59283) );
  BUFx3_ASAP7_75t_SL U64299 ( .A(n68410), .Y(n59502) );
  NAND2xp5_ASAP7_75t_SL U64300 ( .A(n63793), .B(n63794), .Y(n63796) );
  NOR2x1_ASAP7_75t_SL U64301 ( .A(n67217), .B(n67218), .Y(n68711) );
  OAI22xp5_ASAP7_75t_SL U64302 ( .A1(n67442), .A2(n67018), .B1(n58903), .B2(
        n66853), .Y(n67005) );
  INVx2_ASAP7_75t_SL U64303 ( .A(n59446), .Y(n59447) );
  INVx2_ASAP7_75t_SL U64304 ( .A(n67902), .Y(n67866) );
  NAND2xp5_ASAP7_75t_SL U64305 ( .A(n64732), .B(n64736), .Y(n64735) );
  BUFx6f_ASAP7_75t_SL U64306 ( .A(n59350), .Y(n59352) );
  AOI21xp5_ASAP7_75t_SL U64307 ( .A1(n75102), .A2(n75103), .B(n75101), .Y(
        n75115) );
  OAI21xp5_ASAP7_75t_SL U64308 ( .A1(n57414), .A2(n58476), .B(n66423), .Y(
        n66484) );
  OAI21xp5_ASAP7_75t_SL U64309 ( .A1(n67937), .A2(n67796), .B(n67936), .Y(
        n67648) );
  BUFx3_ASAP7_75t_SL U64310 ( .A(n1584), .Y(n59529) );
  INVx1_ASAP7_75t_SL U64311 ( .A(n68346), .Y(n58733) );
  INVx1_ASAP7_75t_SL U64312 ( .A(n68101), .Y(n65043) );
  INVx1_ASAP7_75t_SL U64313 ( .A(n63881), .Y(n63886) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64314 ( .A1(n59503), .A2(n59514), .B(n67460), 
        .C(n62784), .Y(n62786) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64315 ( .A1(n68008), .A2(n56827), .B(n57104), 
        .C(n68007), .Y(n68009) );
  INVx1_ASAP7_75t_SL U64316 ( .A(n67460), .Y(n63068) );
  NAND2xp5_ASAP7_75t_SL U64317 ( .A(n57272), .B(n59595), .Y(n67460) );
  INVx2_ASAP7_75t_SL U64318 ( .A(n56827), .Y(n59593) );
  NAND2xp5_ASAP7_75t_SL U64319 ( .A(n75289), .B(n75288), .Y(n78171) );
  NOR2x1_ASAP7_75t_SL U64320 ( .A(n58895), .B(n69100), .Y(n69118) );
  INVx1_ASAP7_75t_SL U64321 ( .A(n66984), .Y(n66904) );
  NAND2xp5_ASAP7_75t_SL U64322 ( .A(n59321), .B(n62555), .Y(n59323) );
  INVx1_ASAP7_75t_SL U64323 ( .A(n67163), .Y(n67161) );
  NAND2xp5_ASAP7_75t_SL U64324 ( .A(n59604), .B(n67360), .Y(n59048) );
  INVx1_ASAP7_75t_SL U64325 ( .A(n62711), .Y(n62999) );
  NAND2xp5_ASAP7_75t_SL U64326 ( .A(n59557), .B(n59465), .Y(n62640) );
  NAND2x1_ASAP7_75t_SL U64327 ( .A(n67230), .B(n58929), .Y(n67457) );
  NAND2xp5_ASAP7_75t_SL U64328 ( .A(n68397), .B(n59090), .Y(n59022) );
  OAI21xp5_ASAP7_75t_SL U64329 ( .A1(n70754), .A2(n70755), .B(n70741), .Y(
        n70751) );
  NAND2xp5_ASAP7_75t_SL U64330 ( .A(n71026), .B(n58326), .Y(n70982) );
  NAND2xp5_ASAP7_75t_SL U64331 ( .A(n70590), .B(n70601), .Y(n70586) );
  NAND2xp5_ASAP7_75t_SL U64332 ( .A(n70577), .B(n70608), .Y(n70590) );
  NAND2xp5_ASAP7_75t_SL U64333 ( .A(n70578), .B(n70600), .Y(n70601) );
  NOR2x1_ASAP7_75t_SL U64334 ( .A(n74399), .B(n74400), .Y(n74409) );
  NAND2xp5_ASAP7_75t_SL U64335 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_19_), .B(
        n74413), .Y(n74423) );
  NOR2x1_ASAP7_75t_SL U64336 ( .A(n74307), .B(n74408), .Y(n74413) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64337 ( .A1(n67227), .A2(n67451), .B(n68101), 
        .C(n62876), .Y(n62875) );
  INVx1_ASAP7_75t_SL U64338 ( .A(n68630), .Y(n68631) );
  AOI22xp5_ASAP7_75t_SL U64339 ( .A1(n66601), .A2(n66600), .B1(n66599), .B2(
        n66598), .Y(n68630) );
  NOR2x1_ASAP7_75t_SL U64340 ( .A(n63876), .B(n63875), .Y(n64699) );
  BUFx6f_ASAP7_75t_SL U64341 ( .A(n1813), .Y(n59542) );
  NAND2x1p5_ASAP7_75t_SL U64342 ( .A(n57302), .B(n64896), .Y(n67868) );
  AOI21xp5_ASAP7_75t_SL U64343 ( .A1(n59353), .A2(n58469), .B(n64515), .Y(
        n67030) );
  OAI21xp5_ASAP7_75t_SL U64344 ( .A1(n71089), .A2(n71281), .B(n71088), .Y(
        n71210) );
  NAND2xp5_ASAP7_75t_SL U64345 ( .A(n71352), .B(n71351), .Y(n71407) );
  INVx1_ASAP7_75t_SL U64346 ( .A(n63238), .Y(n63150) );
  NAND2xp5_ASAP7_75t_SL U64347 ( .A(n63133), .B(n63132), .Y(n63238) );
  OAI21xp5_ASAP7_75t_SL U64348 ( .A1(n63477), .A2(n63476), .B(n63448), .Y(
        n58814) );
  NAND2xp5_ASAP7_75t_SL U64349 ( .A(n60199), .B(n61999), .Y(n60197) );
  NAND2xp5_ASAP7_75t_SL U64350 ( .A(n60193), .B(n77996), .Y(n61287) );
  AOI21xp5_ASAP7_75t_SL U64351 ( .A1(n53440), .A2(n77369), .B(n76844), .Y(
        n65211) );
  INVx4_ASAP7_75t_SL U64352 ( .A(n59456), .Y(n67963) );
  INVx2_ASAP7_75t_SL U64353 ( .A(n68053), .Y(n59354) );
  BUFx3_ASAP7_75t_SL U64354 ( .A(n1836), .Y(n59544) );
  BUFx6f_ASAP7_75t_SL U64355 ( .A(n2789), .Y(n59567) );
  INVx1_ASAP7_75t_SL U64356 ( .A(n68555), .Y(n68558) );
  INVx3_ASAP7_75t_SL U64357 ( .A(n59659), .Y(n58851) );
  AND2x6_ASAP7_75t_SL U64358 ( .A(n58978), .B(n58977), .Y(n59659) );
  NAND2x1_ASAP7_75t_SL U64359 ( .A(n68587), .B(n68588), .Y(n69028) );
  INVx1_ASAP7_75t_SL U64360 ( .A(n68268), .Y(n65065) );
  INVx1_ASAP7_75t_SL U64361 ( .A(n68019), .Y(n67741) );
  NAND2xp5_ASAP7_75t_SL U64362 ( .A(n64924), .B(n64923), .Y(n68019) );
  INVx1_ASAP7_75t_SL U64363 ( .A(n68955), .Y(n69005) );
  OAI21xp5_ASAP7_75t_SL U64364 ( .A1(n75912), .A2(n59599), .B(n67289), .Y(
        n67387) );
  INVx2_ASAP7_75t_SL U64365 ( .A(n59551), .Y(n77705) );
  INVx1_ASAP7_75t_SL U64366 ( .A(n68579), .Y(n58998) );
  OAI21xp5_ASAP7_75t_SL U64367 ( .A1(n67844), .A2(n57158), .B(n59040), .Y(
        n67895) );
  INVx2_ASAP7_75t_SL U64368 ( .A(n76078), .Y(n59041) );
  AOI21xp5_ASAP7_75t_SL U64369 ( .A1(n71033), .A2(n71032), .B(n71031), .Y(
        n71053) );
  NAND2xp5_ASAP7_75t_SL U64370 ( .A(n69083), .B(n69298), .Y(n58852) );
  INVx1_ASAP7_75t_SL U64371 ( .A(n67111), .Y(n66509) );
  NAND2xp5_ASAP7_75t_SL U64372 ( .A(n66524), .B(n66523), .Y(n74111) );
  AOI21xp5_ASAP7_75t_SL U64373 ( .A1(n66505), .A2(n66504), .B(n66503), .Y(
        n66516) );
  INVx1_ASAP7_75t_SL U64374 ( .A(n63233), .Y(n63647) );
  OAI21xp5_ASAP7_75t_SL U64375 ( .A1(n64746), .A2(n64745), .B(n65102), .Y(
        n64748) );
  OAI21xp5_ASAP7_75t_SL U64376 ( .A1(n76880), .A2(n68807), .B(n76881), .Y(
        n59346) );
  INVx1_ASAP7_75t_SL U64377 ( .A(n64657), .Y(n64662) );
  INVx1_ASAP7_75t_SL U64378 ( .A(n64523), .Y(n64378) );
  NAND2xp5_ASAP7_75t_SL U64379 ( .A(n63876), .B(n63875), .Y(n64728) );
  INVx2_ASAP7_75t_SL U64380 ( .A(n59610), .Y(n59608) );
  NAND2x1_ASAP7_75t_SL U64381 ( .A(n68955), .B(n59382), .Y(n68975) );
  INVx1_ASAP7_75t_SL U64382 ( .A(n68068), .Y(n68072) );
  NAND2xp5_ASAP7_75t_SL U64383 ( .A(or1200_cpu_rf_rdb), .B(n77407), .Y(n77363)
         );
  AOI31xp67_ASAP7_75t_SL U64384 ( .A1(n60213), .A2(n60214), .A3(n60212), .B(
        n60211), .Y(n76538) );
  NAND2xp5_ASAP7_75t_SL U64385 ( .A(n59883), .B(n59882), .Y(n60212) );
  INVx1_ASAP7_75t_SL U64386 ( .A(n62948), .Y(n63344) );
  NAND2xp5_ASAP7_75t_SL U64387 ( .A(n62869), .B(n62850), .Y(n62855) );
  OAI21xp5_ASAP7_75t_SL U64388 ( .A1(n66695), .A2(n66694), .B(n66693), .Y(
        n66707) );
  INVx2_ASAP7_75t_SL U64389 ( .A(n59663), .Y(n59666) );
  OAI21xp5_ASAP7_75t_SL U64390 ( .A1(n77214), .A2(n1739), .B(n60262), .Y(
        or1200_cpu_to_sr[2]) );
  NAND2xp5_ASAP7_75t_SL U64391 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_20_), 
        .B(n74416), .Y(n74426) );
  INVx1_ASAP7_75t_SL U64392 ( .A(n63003), .Y(n62969) );
  INVx3_ASAP7_75t_SL U64393 ( .A(n75901), .Y(n75903) );
  NOR2x1p5_ASAP7_75t_SL U64394 ( .A(n62583), .B(n67625), .Y(n75901) );
  NOR2x1_ASAP7_75t_SL U64395 ( .A(n66204), .B(n76950), .Y(n76949) );
  NOR2x1_ASAP7_75t_SL U64396 ( .A(n74058), .B(n74201), .Y(n74179) );
  XNOR2x1_ASAP7_75t_SL U64397 ( .A(n59091), .B(n59027), .Y(n68428) );
  INVx1_ASAP7_75t_SL U64398 ( .A(n68437), .Y(n59091) );
  NAND2xp5_ASAP7_75t_SL U64399 ( .A(n62599), .B(n57186), .Y(n62600) );
  INVx1_ASAP7_75t_SL U64400 ( .A(n68255), .Y(n65068) );
  NAND2x1p5_ASAP7_75t_SL U64401 ( .A(n64609), .B(n53291), .Y(n67951) );
  NAND2xp5_ASAP7_75t_SL U64402 ( .A(n60053), .B(n60054), .Y(n60079) );
  NAND2xp5_ASAP7_75t_SL U64403 ( .A(n59987), .B(n60016), .Y(n60014) );
  INVx1_ASAP7_75t_SL U64404 ( .A(n68565), .Y(n68252) );
  INVx1_ASAP7_75t_SL U64405 ( .A(n66494), .Y(n66406) );
  INVx3_ASAP7_75t_SL U64406 ( .A(n59553), .Y(n59387) );
  BUFx3_ASAP7_75t_SL U64407 ( .A(n1941), .Y(n59553) );
  NOR2x1_ASAP7_75t_SL U64408 ( .A(n74347), .B(n74348), .Y(n74385) );
  NOR2x1_ASAP7_75t_SL U64409 ( .A(n74222), .B(n74223), .Y(n74450) );
  NOR2x1_ASAP7_75t_SL U64410 ( .A(n74432), .B(n74433), .Y(n74431) );
  NOR2x1_ASAP7_75t_SL U64411 ( .A(n74342), .B(n74343), .Y(n74371) );
  AOI21xp5_ASAP7_75t_SL U64412 ( .A1(n75464), .A2(n75096), .B(n75086), .Y(
        n75087) );
  NOR2x1_ASAP7_75t_SL U64413 ( .A(n58852), .B(n58826), .Y(n68662) );
  NAND2xp5_ASAP7_75t_SL U64414 ( .A(n66742), .B(n66741), .Y(n66968) );
  NAND2xp5_ASAP7_75t_SL U64415 ( .A(n59112), .B(n59111), .Y(n66741) );
  INVx1_ASAP7_75t_SL U64416 ( .A(n75440), .Y(n59767) );
  BUFx6f_ASAP7_75t_SL U64417 ( .A(n1842), .Y(n59545) );
  OAI22xp5_ASAP7_75t_SL U64418 ( .A1(n68015), .A2(n67315), .B1(n68383), .B2(
        n67314), .Y(n67893) );
  INVx1_ASAP7_75t_SL U64419 ( .A(n59394), .Y(n63124) );
  NAND2x1_ASAP7_75t_SL U64420 ( .A(n68517), .B(n68516), .Y(n69012) );
  BUFx6f_ASAP7_75t_SL U64421 ( .A(n3115), .Y(n59580) );
  NAND2xp5_ASAP7_75t_SL U64422 ( .A(n68736), .B(n58854), .Y(n68806) );
  OAI21xp5_ASAP7_75t_SL U64423 ( .A1(n75089), .A2(n75088), .B(n75087), .Y(
        n75090) );
  NOR2x1_ASAP7_75t_SL U64424 ( .A(n75107), .B(n75088), .Y(n75470) );
  NAND2xp5_ASAP7_75t_SL U64425 ( .A(n75103), .B(n75138), .Y(n75080) );
  NAND2xp5_ASAP7_75t_SL U64426 ( .A(n75062), .B(n75061), .Y(n75103) );
  INVx1_ASAP7_75t_SL U64427 ( .A(n68066), .Y(n68067) );
  AOI21xp5_ASAP7_75t_SL U64428 ( .A1(n68919), .A2(n68920), .B(n68663), .Y(
        n68664) );
  INVx1_ASAP7_75t_SL U64429 ( .A(n58723), .Y(n68527) );
  NAND2xp5_ASAP7_75t_SL U64430 ( .A(n69006), .B(n69029), .Y(n69011) );
  NAND2xp5_ASAP7_75t_SL U64431 ( .A(n68539), .B(n68540), .Y(n69006) );
  OAI21xp5_ASAP7_75t_SL U64432 ( .A1(n57179), .A2(n67432), .B(n66787), .Y(
        n66928) );
  NAND2xp5_ASAP7_75t_SL U64433 ( .A(n73944), .B(n73937), .Y(n75814) );
  NAND2xp5_ASAP7_75t_SL U64434 ( .A(n75223), .B(n75222), .Y(n75751) );
  INVx3_ASAP7_75t_SL U64435 ( .A(n59579), .Y(n76486) );
  BUFx6f_ASAP7_75t_SL U64436 ( .A(n2956), .Y(n59579) );
  OAI21xp5_ASAP7_75t_SL U64437 ( .A1(n58471), .A2(n75095), .B(n59422), .Y(
        n59421) );
  BUFx3_ASAP7_75t_SL U64438 ( .A(n75983), .Y(n59514) );
  INVx3_ASAP7_75t_SL U64439 ( .A(n59586), .Y(n59585) );
  INVx1_ASAP7_75t_SL U64440 ( .A(n64233), .Y(n59586) );
  AOI21xp5_ASAP7_75t_SL U64441 ( .A1(n67617), .A2(n67616), .B(n67615), .Y(
        n59114) );
  INVx2_ASAP7_75t_SL U64442 ( .A(n59569), .Y(n76653) );
  BUFx6f_ASAP7_75t_SL U64443 ( .A(n2830), .Y(n59569) );
  NAND2x1p5_ASAP7_75t_SL U64444 ( .A(n76881), .B(n68904), .Y(n68920) );
  NAND2xp5_ASAP7_75t_SL U64445 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_15_), .B(
        n74390), .Y(n74400) );
  NAND2xp5_ASAP7_75t_SL U64446 ( .A(n70617), .B(n70616), .Y(n70618) );
  NAND2xp5_ASAP7_75t_SL U64447 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[7]), .B(
        n70607), .Y(n70617) );
  NAND2xp5_ASAP7_75t_SL U64448 ( .A(n70613), .B(n70612), .Y(n70616) );
  AOI21xp5_ASAP7_75t_SL U64449 ( .A1(n71305), .A2(n71299), .B(n71292), .Y(
        n71276) );
  AOI21xp5_ASAP7_75t_SL U64450 ( .A1(n70839), .A2(n70838), .B(n70837), .Y(
        n70878) );
  AOI21xp5_ASAP7_75t_SL U64451 ( .A1(n71157), .A2(n71156), .B(n71155), .Y(
        n71299) );
  XNOR2x1_ASAP7_75t_SL U64452 ( .A(n75643), .B(n58406), .Y(n75044) );
  INVx1_ASAP7_75t_SL U64453 ( .A(n67347), .Y(n67348) );
  BUFx6f_ASAP7_75t_SL U64454 ( .A(n2939), .Y(n59577) );
  NAND2xp5_ASAP7_75t_SL U64455 ( .A(n68265), .B(n68267), .Y(n58891) );
  XOR2x2_ASAP7_75t_SL U64456 ( .A(n57169), .B(n58402), .Y(n58492) );
  XNOR2x2_ASAP7_75t_SL U64457 ( .A(n57169), .B(n59594), .Y(n62654) );
  XNOR2x2_ASAP7_75t_SL U64458 ( .A(n57169), .B(n59603), .Y(n63823) );
  NAND2xp5_ASAP7_75t_SL U64459 ( .A(n67188), .B(n58327), .Y(n67187) );
  NAND2xp5_ASAP7_75t_SL U64460 ( .A(n68563), .B(n68567), .Y(n68254) );
  OAI21xp5_ASAP7_75t_SL U64461 ( .A1(n58402), .A2(n59510), .B(n64960), .Y(
        n67849) );
  BUFx6f_ASAP7_75t_SL U64462 ( .A(n76632), .Y(n59505) );
  BUFx6f_ASAP7_75t_SL U64463 ( .A(n1995), .Y(n59559) );
  OAI21xp5_ASAP7_75t_SL U64464 ( .A1(n67434), .A2(n67718), .B(n67277), .Y(
        n67471) );
  INVx1_ASAP7_75t_SL U64465 ( .A(n67724), .Y(n68425) );
  NAND2xp5_ASAP7_75t_SL U64466 ( .A(n59403), .B(n58902), .Y(n59404) );
  INVx1_ASAP7_75t_SL U64467 ( .A(n65027), .Y(n64653) );
  INVx1_ASAP7_75t_SL U64468 ( .A(n68296), .Y(n68341) );
  INVx3_ASAP7_75t_SL U64469 ( .A(n59649), .Y(n59648) );
  INVx1_ASAP7_75t_SL U64470 ( .A(n64729), .Y(n65104) );
  INVx1_ASAP7_75t_SL U64471 ( .A(n58735), .Y(n64076) );
  AND2x4_ASAP7_75t_SL U64472 ( .A(n59476), .B(n62649), .Y(n58440) );
  OAI21xp5_ASAP7_75t_SL U64473 ( .A1(n68661), .A2(n68662), .B(n68660), .Y(
        n52010) );
  AOI21xp5_ASAP7_75t_SL U64474 ( .A1(n68662), .A2(n68659), .B(n68658), .Y(
        n68660) );
  NAND2xp5_ASAP7_75t_SL U64475 ( .A(n71344), .B(n71325), .Y(n71326) );
  INVx2_ASAP7_75t_SL U64476 ( .A(n71284), .Y(n71315) );
  NAND2x1_ASAP7_75t_SL U64477 ( .A(n58790), .B(n67445), .Y(n67923) );
  O2A1O1Ixp33_ASAP7_75t_SRAM U64478 ( .A1(n76049), .A2(n59615), .B(n63202), 
        .C(n68079), .Y(n63203) );
  INVx1_ASAP7_75t_SL U64479 ( .A(n68549), .Y(n68551) );
  OAI21xp5_ASAP7_75t_SL U64480 ( .A1(n58919), .A2(n75438), .B(n66725), .Y(
        n67752) );
  NAND2xp5_ASAP7_75t_SL U64481 ( .A(n58384), .B(n58919), .Y(n66725) );
  INVx6_ASAP7_75t_SL U64482 ( .A(n59660), .Y(n58919) );
  OR2x6_ASAP7_75t_SL U64483 ( .A(n59181), .B(n59180), .Y(n59660) );
  NAND2xp5_ASAP7_75t_SL U64484 ( .A(n58847), .B(n58846), .Y(n67760) );
  INVx3_ASAP7_75t_SL U64485 ( .A(n68100), .Y(n67736) );
  INVx1_ASAP7_75t_SL U64486 ( .A(n68061), .Y(n68060) );
  INVx1_ASAP7_75t_SL U64487 ( .A(n67373), .Y(n67613) );
  INVx1_ASAP7_75t_SL U64488 ( .A(n68493), .Y(n58988) );
  OAI21xp5_ASAP7_75t_SL U64489 ( .A1(n59024), .A2(n59023), .B(n59022), .Y(
        n59021) );
  BUFx6f_ASAP7_75t_SL U64490 ( .A(n2841), .Y(n59571) );
  BUFx6f_ASAP7_75t_SL U64491 ( .A(n1566), .Y(n59528) );
  INVx1_ASAP7_75t_SL U64492 ( .A(n75464), .Y(n75088) );
  INVx3_ASAP7_75t_SL U64493 ( .A(n67709), .Y(n59446) );
  NAND2xp5_ASAP7_75t_SL U64494 ( .A(n75042), .B(n75041), .Y(n75106) );
  NAND2xp5_ASAP7_75t_SL U64495 ( .A(n68640), .B(n68639), .Y(n75042) );
  AOI21xp5_ASAP7_75t_SL U64496 ( .A1(n67804), .A2(n67801), .B(n58896), .Y(
        n67939) );
  NAND2xp5_ASAP7_75t_SL U64497 ( .A(n68593), .B(n68592), .Y(n69025) );
  INVx1_ASAP7_75t_SL U64498 ( .A(n69300), .Y(n68666) );
  NOR2x1_ASAP7_75t_SL U64499 ( .A(n59654), .B(n62682), .Y(n67860) );
  XNOR2x2_ASAP7_75t_SL U64500 ( .A(n67941), .B(n59428), .Y(n68050) );
  OAI21xp5_ASAP7_75t_SL U64501 ( .A1(n58334), .A2(n58737), .B(n57557), .Y(
        n68049) );
  OAI21xp5_ASAP7_75t_SL U64502 ( .A1(n73397), .A2(n73396), .B(n73395), .Y(
        n73403) );
  OAI21xp5_ASAP7_75t_SL U64503 ( .A1(n59630), .A2(n73229), .B(n73228), .Y(
        n73234) );
  NAND2xp5_ASAP7_75t_SL U64504 ( .A(n59343), .B(n59345), .Y(n59342) );
  INVx1_ASAP7_75t_SL U64505 ( .A(n59094), .Y(n58689) );
  BUFx3_ASAP7_75t_SL U64506 ( .A(n68006), .Y(n59437) );
  INVx3_ASAP7_75t_SL U64507 ( .A(n59568), .Y(n76690) );
  BUFx6f_ASAP7_75t_SL U64508 ( .A(n2802), .Y(n59568) );
  NAND2xp5_ASAP7_75t_SL U64509 ( .A(n68972), .B(n69005), .Y(n59385) );
  NAND2xp5_ASAP7_75t_SL U64510 ( .A(n67221), .B(n59390), .Y(n75112) );
  INVx2_ASAP7_75t_SL U64511 ( .A(n67846), .Y(n76057) );
  NAND2xp5_ASAP7_75t_SL U64512 ( .A(n64735), .B(n74994), .Y(n65110) );
  NOR2x1_ASAP7_75t_SL U64513 ( .A(n64741), .B(n64740), .Y(n68902) );
  NAND2xp5_ASAP7_75t_SL U64514 ( .A(n64738), .B(n64737), .Y(n74991) );
  OAI22xp5_ASAP7_75t_SL U64515 ( .A1(n59698), .A2(n71375), .B1(n57211), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_45_), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n238) );
  INVx1_ASAP7_75t_SL U64516 ( .A(n69304), .Y(n59196) );
  NOR2x1_ASAP7_75t_SL U64517 ( .A(n68632), .B(n68631), .Y(n69304) );
  OAI21xp5_ASAP7_75t_SL U64518 ( .A1(n59273), .A2(n59274), .B(n59272), .Y(
        n75085) );
  AND2x4_ASAP7_75t_SL U64519 ( .A(n75915), .B(n66244), .Y(n58433) );
  OAI21x1_ASAP7_75t_SL U64520 ( .A1(n59142), .A2(n58516), .B(n58633), .Y(
        n66557) );
  INVx1_ASAP7_75t_SL U64521 ( .A(n59449), .Y(n74113) );
  BUFx2_ASAP7_75t_SL U64522 ( .A(n69238), .Y(n59449) );
  AOI21xp5_ASAP7_75t_SL U64523 ( .A1(n74559), .A2(n68586), .B(n68585), .Y(
        n68674) );
  OAI21xp5_ASAP7_75t_SL U64524 ( .A1(n57158), .A2(n66469), .B(n58859), .Y(
        n67144) );
  OAI21xp5_ASAP7_75t_SL U64525 ( .A1(n67434), .A2(n67020), .B(n58525), .Y(
        n58858) );
  INVx1_ASAP7_75t_SL U64526 ( .A(n68717), .Y(n68914) );
  AOI21xp5_ASAP7_75t_SL U64527 ( .A1(n66778), .A2(n66779), .B(n66780), .Y(
        n66820) );
  INVx1_ASAP7_75t_SL U64528 ( .A(n75287), .Y(n68714) );
  INVx1_ASAP7_75t_SL U64529 ( .A(n69095), .Y(n58895) );
  INVx1_ASAP7_75t_SL U64530 ( .A(n66989), .Y(n66983) );
  NAND2xp5_ASAP7_75t_SL U64531 ( .A(n53505), .B(n68909), .Y(n68869) );
  NAND2xp5_ASAP7_75t_SL U64532 ( .A(n68906), .B(n68578), .Y(n68909) );
  NOR2x1_ASAP7_75t_SL U64533 ( .A(n68538), .B(n68537), .Y(n69008) );
  BUFx5_ASAP7_75t_SL U64534 ( .A(n67806), .Y(n59506) );
  OAI21xp5_ASAP7_75t_SL U64535 ( .A1(n71306), .A2(n71305), .B(n71304), .Y(
        n71307) );
  AOI21xp5_ASAP7_75t_SL U64536 ( .A1(n68750), .A2(n68804), .B(n57269), .Y(
        n68738) );
  INVx1_ASAP7_75t_SL U64537 ( .A(n68806), .Y(n68750) );
  INVx1_ASAP7_75t_SL U64538 ( .A(n63025), .Y(n63026) );
  NOR2x1_ASAP7_75t_SL U64539 ( .A(n74309), .B(n74401), .Y(n74308) );
  NAND2xp5_ASAP7_75t_SL U64540 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_37_), .B(
        n74402), .Y(n74401) );
  NAND2xp5_ASAP7_75t_SL U64541 ( .A(n71110), .B(n71109), .Y(n71114) );
  OAI21xp5_ASAP7_75t_SL U64542 ( .A1(n71100), .A2(n71099), .B(n71098), .Y(
        n71109) );
  NOR2x1_ASAP7_75t_SL U64543 ( .A(n68975), .B(n68958), .Y(n68976) );
  NAND2xp5_ASAP7_75t_SL U64544 ( .A(n68837), .B(n68836), .Y(n68908) );
  NOR2x1_ASAP7_75t_SL U64545 ( .A(n57130), .B(n58831), .Y(n59457) );
  INVx1_ASAP7_75t_SL U64546 ( .A(n68351), .Y(n68352) );
  OAI21xp5_ASAP7_75t_SL U64547 ( .A1(n66442), .A2(n66443), .B(n66441), .Y(
        n66530) );
  NAND2xp5_ASAP7_75t_SL U64548 ( .A(n66443), .B(n66442), .Y(n66441) );
  OAI21xp5_ASAP7_75t_SL U64549 ( .A1(n66427), .A2(n66426), .B(n66428), .Y(
        n66446) );
  NAND2xp5_ASAP7_75t_SL U64550 ( .A(n66426), .B(n66427), .Y(n66428) );
  INVx2_ASAP7_75t_SL U64551 ( .A(n59166), .Y(n74788) );
  NOR2x1_ASAP7_75t_SL U64552 ( .A(n68560), .B(n68726), .Y(n58688) );
  INVx1_ASAP7_75t_SL U64553 ( .A(n68554), .Y(n66979) );
  INVx2_ASAP7_75t_SL U64554 ( .A(n69114), .Y(n69102) );
  OAI21xp5_ASAP7_75t_SL U64555 ( .A1(n62081), .A2(n64273), .B(n62080), .Y(
        n62501) );
  NOR2x1_ASAP7_75t_SL U64556 ( .A(n76320), .B(n76319), .Y(n76324) );
  OAI21xp5_ASAP7_75t_SL U64557 ( .A1(n59557), .A2(n60759), .B(n61399), .Y(
        n61560) );
  AOI22xp5_ASAP7_75t_SL U64558 ( .A1(n64694), .A2(n64551), .B1(n64550), .B2(
        n64693), .Y(n64984) );
  OAI22xp5_ASAP7_75t_SL U64559 ( .A1(n64502), .A2(n58884), .B1(n59012), .B2(
        n65061), .Y(n64639) );
  INVx1_ASAP7_75t_SL U64560 ( .A(n68975), .Y(n68967) );
  INVx2_ASAP7_75t_SL U64561 ( .A(n68102), .Y(n67609) );
  INVx1_ASAP7_75t_SL U64562 ( .A(n67067), .Y(n67069) );
  AOI21xp5_ASAP7_75t_SL U64563 ( .A1(n67169), .A2(n67178), .B(n67186), .Y(
        n67193) );
  BUFx6f_ASAP7_75t_SL U64564 ( .A(n1981), .Y(n59558) );
  OAI21xp5_ASAP7_75t_SL U64565 ( .A1(n63292), .A2(n63310), .B(n62912), .Y(
        n63366) );
  AOI21xp5_ASAP7_75t_SL U64566 ( .A1(n63311), .A2(n62911), .B(n63345), .Y(
        n62912) );
  NAND2x1_ASAP7_75t_SL U64567 ( .A(n63280), .B(n63281), .Y(n63298) );
  NOR2x1_ASAP7_75t_SL U64568 ( .A(n62893), .B(n62892), .Y(n63281) );
  AOI21xp5_ASAP7_75t_SL U64569 ( .A1(n69160), .A2(n69157), .B(n69156), .Y(
        n69158) );
  XNOR2x2_ASAP7_75t_SL U64570 ( .A(n59603), .B(n59510), .Y(n64379) );
  INVx1_ASAP7_75t_SL U64571 ( .A(n69117), .Y(n69083) );
  NOR2x1_ASAP7_75t_SL U64572 ( .A(n58313), .B(n59404), .Y(n68900) );
  XNOR2x1_ASAP7_75t_SL U64573 ( .A(n68330), .B(n59329), .Y(n68327) );
  OAI21xp5_ASAP7_75t_SL U64574 ( .A1(n67944), .A2(n67740), .B(n59416), .Y(
        n65042) );
  INVx3_ASAP7_75t_SL U64575 ( .A(n67444), .Y(n67944) );
  INVx4_ASAP7_75t_SL U64576 ( .A(n58408), .Y(n75930) );
  INVx4_ASAP7_75t_SL U64577 ( .A(n59605), .Y(n59603) );
  INVx1_ASAP7_75t_SL U64578 ( .A(n68567), .Y(n68835) );
  NAND2xp5_ASAP7_75t_SL U64579 ( .A(n68565), .B(n68566), .Y(n68567) );
  BUFx6f_ASAP7_75t_SL U64580 ( .A(n1602), .Y(n59530) );
  NAND2xp5_ASAP7_75t_SL U64581 ( .A(n75094), .B(n75093), .Y(n78168) );
  INVx2_ASAP7_75t_SL U64582 ( .A(n59636), .Y(n59635) );
  OAI21xp5_ASAP7_75t_SL U64583 ( .A1(n59207), .A2(n59342), .B(n58522), .Y(
        n59208) );
  NAND2x1_ASAP7_75t_SL U64584 ( .A(n68808), .B(n57063), .Y(n59345) );
  NAND2xp5_ASAP7_75t_SL U64585 ( .A(n68871), .B(n68870), .Y(n51995) );
  NAND2xp5_ASAP7_75t_SL U64586 ( .A(n59594), .B(n59459), .Y(n64606) );
  INVx2_ASAP7_75t_SL U64587 ( .A(n67276), .Y(n59459) );
  NAND2xp5_ASAP7_75t_SL U64588 ( .A(n59389), .B(n59391), .Y(n69241) );
  INVx1_ASAP7_75t_SL U64589 ( .A(n69241), .Y(n68686) );
  NAND2xp5_ASAP7_75t_SL U64590 ( .A(n68735), .B(n64870), .Y(n68761) );
  NAND2x1_ASAP7_75t_SL U64591 ( .A(n74111), .B(n68684), .Y(n69235) );
  OAI21xp5_ASAP7_75t_SL U64592 ( .A1(n68646), .A2(n68647), .B(n59420), .Y(
        n51987) );
  NAND2xp5_ASAP7_75t_SL U64593 ( .A(n58445), .B(n68673), .Y(n75107) );
  INVx1_ASAP7_75t_SL U64594 ( .A(n64996), .Y(n64946) );
  BUFx6f_ASAP7_75t_SL U64595 ( .A(n1956), .Y(n59555) );
  INVx1_ASAP7_75t_SL U64596 ( .A(n68920), .Y(n68721) );
  INVx5_ASAP7_75t_SL U64597 ( .A(n59665), .Y(n59664) );
  NAND2xp5_ASAP7_75t_SL U64598 ( .A(n59196), .B(n68667), .Y(n59195) );
  AOI22xp5_ASAP7_75t_SL U64599 ( .A1(n66597), .A2(n66596), .B1(n66595), .B2(
        n66594), .Y(n66604) );
  OAI21xp5_ASAP7_75t_SL U64600 ( .A1(n57032), .A2(n66809), .B(n58438), .Y(
        n66910) );
  NAND2xp5_ASAP7_75t_SL U64601 ( .A(n66816), .B(n66907), .Y(n67041) );
  NOR2x1_ASAP7_75t_SL U64602 ( .A(n68697), .B(n68696), .Y(n74562) );
  NAND2xp5_ASAP7_75t_SL U64603 ( .A(n67044), .B(n66905), .Y(n67210) );
  BUFx6f_ASAP7_75t_SL U64604 ( .A(n1971), .Y(n59557) );
  INVx1_ASAP7_75t_SL U64605 ( .A(n59025), .Y(n68492) );
  INVx2_ASAP7_75t_SL U64606 ( .A(n1989), .Y(n59441) );
  INVx1_ASAP7_75t_SL U64607 ( .A(n65049), .Y(n64903) );
  XOR2x2_ASAP7_75t_SL U64608 ( .A(n69138), .B(n66867), .Y(n66982) );
  INVx1_ASAP7_75t_SL U64609 ( .A(n69139), .Y(n66867) );
  INVx3_ASAP7_75t_SL U64610 ( .A(n59670), .Y(n58672) );
  AO21x2_ASAP7_75t_SL U64611 ( .A1(n58474), .A2(n58909), .B(n58908), .Y(n58404) );
  INVx8_ASAP7_75t_SL U64612 ( .A(n59597), .Y(n59598) );
  INVxp33_ASAP7_75t_SRAM U64613 ( .A(n78165), .Y(n77995) );
  INVxp33_ASAP7_75t_SRAM U64614 ( .A(n4139), .Y(n78175) );
  INVxp33_ASAP7_75t_SRAM U64615 ( .A(n1192), .Y(dwb_adr_o[30]) );
  OAI21xp33_ASAP7_75t_SRAM U64616 ( .A1(n77748), .A2(n4240), .B(n77747), .Y(
        dwb_dat_o[31]) );
  INVxp33_ASAP7_75t_SRAM U64617 ( .A(n1341), .Y(dwb_cyc_o) );
  INVxp33_ASAP7_75t_SRAM U64618 ( .A(n1187), .Y(dwb_adr_o[31]) );
  INVxp33_ASAP7_75t_SRAM U64619 ( .A(n1046), .Y(iwb_adr_o[5]) );
  INVxp33_ASAP7_75t_SRAM U64620 ( .A(n1035), .Y(iwb_adr_o[4]) );
  INVxp33_ASAP7_75t_SRAM U64621 ( .A(n1057), .Y(iwb_adr_o[6]) );
  INVxp33_ASAP7_75t_SRAM U64622 ( .A(n1068), .Y(iwb_adr_o[7]) );
  INVxp33_ASAP7_75t_SRAM U64623 ( .A(n2773), .Y(iwb_stb_o) );
  INVxp33_ASAP7_75t_SRAM U64624 ( .A(n1349), .Y(dwb_we_o) );
  INVxp33_ASAP7_75t_SRAM U64625 ( .A(n833), .Y(iwb_adr_o[2]) );
  INVxp33_ASAP7_75t_SRAM U64626 ( .A(n1079), .Y(iwb_adr_o[8]) );
  INVxp33_ASAP7_75t_SRAM U64627 ( .A(n1090), .Y(iwb_adr_o[9]) );
  INVxp33_ASAP7_75t_SRAM U64628 ( .A(n1101), .Y(iwb_adr_o[10]) );
  INVxp33_ASAP7_75t_SRAM U64629 ( .A(n2769), .Y(iwb_adr_o[11]) );
  INVxp33_ASAP7_75t_SRAM U64630 ( .A(n849), .Y(iwb_adr_o[12]) );
  OAI21xp33_ASAP7_75t_SRAM U64631 ( .A1(n77748), .A2(n4302), .B(n77698), .Y(
        dwb_dat_o[10]) );
  INVxp33_ASAP7_75t_SRAM U64632 ( .A(n2536), .Y(dbg_is_o[0]) );
  INVxp33_ASAP7_75t_SRAM U64633 ( .A(n1508), .Y(dbg_bp_o) );
  INVxp33_ASAP7_75t_SRAM U64634 ( .A(n1181), .Y(sig_tick) );
  INVxp33_ASAP7_75t_SRAM U64635 ( .A(n1222), .Y(dwb_adr_o[24]) );
  INVxp33_ASAP7_75t_SRAM U64636 ( .A(n1252), .Y(dwb_adr_o[18]) );
  INVxp33_ASAP7_75t_SRAM U64637 ( .A(n1262), .Y(dwb_adr_o[16]) );
  INVxp33_ASAP7_75t_SRAM U64638 ( .A(n1277), .Y(dwb_adr_o[13]) );
  INVxp33_ASAP7_75t_SRAM U64639 ( .A(n1297), .Y(dwb_adr_o[11]) );
  INVxp33_ASAP7_75t_SRAM U64640 ( .A(n1302), .Y(dwb_adr_o[10]) );
  INVxp33_ASAP7_75t_SRAM U64641 ( .A(n1307), .Y(dwb_adr_o[9]) );
  INVxp33_ASAP7_75t_SRAM U64642 ( .A(n1312), .Y(dwb_adr_o[8]) );
  INVxp33_ASAP7_75t_SRAM U64643 ( .A(n1317), .Y(dwb_adr_o[7]) );
  INVxp33_ASAP7_75t_SRAM U64644 ( .A(n1322), .Y(dwb_adr_o[6]) );
  INVxp33_ASAP7_75t_SRAM U64645 ( .A(n1327), .Y(dwb_adr_o[5]) );
  INVxp33_ASAP7_75t_SRAM U64646 ( .A(n1332), .Y(dwb_adr_o[4]) );
  INVxp33_ASAP7_75t_SRAM U64647 ( .A(n1337), .Y(dwb_adr_o[3]) );
  OAI21xp33_ASAP7_75t_SRAM U64648 ( .A1(n77748), .A2(n4265), .B(n77720), .Y(
        dwb_dat_o[22]) );
  INVxp33_ASAP7_75t_SRAM U64649 ( .A(n77723), .Y(n77721) );
  INVxp33_ASAP7_75t_SRAM U64650 ( .A(n1287), .Y(dwb_adr_o[1]) );
  OAI21xp33_ASAP7_75t_SRAM U64651 ( .A1(n77748), .A2(n4256), .B(n77731), .Y(
        dwb_dat_o[24]) );
  OAI21xp33_ASAP7_75t_SRAM U64652 ( .A1(n77748), .A2(n4254), .B(n77733), .Y(
        dwb_dat_o[25]) );
  INVxp33_ASAP7_75t_SRAM U64653 ( .A(n1292), .Y(dwb_adr_o[0]) );
  OAI21xp33_ASAP7_75t_SRAM U64654 ( .A1(n77748), .A2(n4242), .B(n77743), .Y(
        dwb_dat_o[30]) );
  OAI21xp33_ASAP7_75t_SRAM U64655 ( .A1(n77748), .A2(n4252), .B(n77736), .Y(
        dwb_dat_o[26]) );
  INVxp33_ASAP7_75t_SRAM U64656 ( .A(n77742), .Y(n77744) );
  INVxp33_ASAP7_75t_SRAM U64657 ( .A(n77741), .Y(n77746) );
  OAI21xp33_ASAP7_75t_SRAM U64658 ( .A1(n77748), .A2(n4250), .B(n77737), .Y(
        dwb_dat_o[27]) );
  INVxp33_ASAP7_75t_SRAM U64659 ( .A(n3100), .Y(dwb_stb_o) );
  OAI21xp33_ASAP7_75t_SRAM U64660 ( .A1(n77748), .A2(n4248), .B(n77739), .Y(
        dwb_dat_o[28]) );
  OAI21xp33_ASAP7_75t_SRAM U64661 ( .A1(n77748), .A2(n4246), .B(n77740), .Y(
        dwb_dat_o[29]) );
  INVxp33_ASAP7_75t_SRAM U64662 ( .A(n77728), .Y(n77727) );
  INVxp33_ASAP7_75t_SRAM U64663 ( .A(n1022), .Y(iwb_adr_o[31]) );
  INVxp33_ASAP7_75t_SRAM U64664 ( .A(n887), .Y(iwb_adr_o[16]) );
  INVxp33_ASAP7_75t_SRAM U64665 ( .A(n1013), .Y(iwb_adr_o[30]) );
  INVxp33_ASAP7_75t_SRAM U64666 ( .A(n977), .Y(iwb_adr_o[26]) );
  INVxp33_ASAP7_75t_SRAM U64667 ( .A(n959), .Y(iwb_adr_o[24]) );
  INVxp33_ASAP7_75t_SRAM U64668 ( .A(n950), .Y(iwb_adr_o[23]) );
  INVxp33_ASAP7_75t_SRAM U64669 ( .A(n941), .Y(iwb_adr_o[22]) );
  INVxp33_ASAP7_75t_SRAM U64670 ( .A(n932), .Y(iwb_adr_o[21]) );
  INVxp33_ASAP7_75t_SRAM U64671 ( .A(n2767), .Y(iwb_cyc_o) );
  INVxp33_ASAP7_75t_SRAM U64672 ( .A(n923), .Y(iwb_adr_o[20]) );
  INVxp33_ASAP7_75t_SRAM U64673 ( .A(n905), .Y(iwb_adr_o[18]) );
  INVxp33_ASAP7_75t_SRAM U64674 ( .A(n914), .Y(iwb_adr_o[19]) );
  INVxp33_ASAP7_75t_SRAM U64675 ( .A(n878), .Y(iwb_adr_o[15]) );
  INVxp33_ASAP7_75t_SRAM U64676 ( .A(n860), .Y(iwb_adr_o[13]) );
  INVxp33_ASAP7_75t_SRAM U64677 ( .A(n896), .Y(iwb_adr_o[17]) );
  INVxp33_ASAP7_75t_SRAM U64678 ( .A(n869), .Y(iwb_adr_o[14]) );
  OAI21xp33_ASAP7_75t_SRAM U64679 ( .A1(n2410), .A2(n74780), .B(n74779), .Y(
        n1497) );
  NOR2xp33_ASAP7_75t_SL U64680 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_start_i), .B(n70650), .Y(
        n70648) );
  INVx1_ASAP7_75t_SL U64681 ( .A(n70530), .Y(n70526) );
  AOI22xp33_ASAP7_75t_SRAM U64682 ( .A1(n57217), .A2(n3310), .B1(n73667), .B2(
        n57205), .Y(n73643) );
  NAND2xp33_ASAP7_75t_SRAM U64683 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_5_), .Y(n62038) );
  NOR2xp33_ASAP7_75t_SL U64684 ( .A(n62047), .B(n62049), .Y(n62059) );
  OAI22xp33_ASAP7_75t_SRAM U64685 ( .A1(n70327), .A2(n70440), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_), .B2(
        n70540), .Y(n70308) );
  OAI22xp33_ASAP7_75t_SRAM U64686 ( .A1(n74664), .A2(n70440), .B1(n74654), 
        .B2(n70540), .Y(n70338) );
  OAI22xp33_ASAP7_75t_SRAM U64687 ( .A1(n74662), .A2(n70440), .B1(n70297), 
        .B2(n70540), .Y(n70300) );
  AOI22xp33_ASAP7_75t_SRAM U64688 ( .A1(n74680), .A2(n74644), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .B2(
        n74686), .Y(n70306) );
  AOI21xp33_ASAP7_75t_SRAM U64689 ( .A1(n74680), .A2(n70311), .B(n74706), .Y(
        n70274) );
  OAI22xp33_ASAP7_75t_SRAM U64690 ( .A1(n74659), .A2(n70440), .B1(n70439), 
        .B2(n70540), .Y(n70425) );
  OAI22xp33_ASAP7_75t_SRAM U64691 ( .A1(n70486), .A2(n70440), .B1(n74659), 
        .B2(n70540), .Y(n70441) );
  AOI22xp33_ASAP7_75t_SRAM U64692 ( .A1(n74680), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_16_), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_), .B2(
        n70543), .Y(n70325) );
  AOI22xp33_ASAP7_75t_SRAM U64693 ( .A1(n74680), .A2(n74660), .B1(n74655), 
        .B2(n70543), .Y(n70395) );
  NOR2xp33_ASAP7_75t_SL U64694 ( .A(n70251), .B(n70252), .Y(n70485) );
  NOR2xp33_ASAP7_75t_SL U64695 ( .A(n70440), .B(n70487), .Y(n70272) );
  INVx1_ASAP7_75t_SL U64696 ( .A(n74680), .Y(n70440) );
  NOR2xp33_ASAP7_75t_SL U64697 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_), .B(
        n74682), .Y(n70542) );
  OAI21xp33_ASAP7_75t_SRAM U64698 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[14]), .A2(n3309), .B(
        n73817), .Y(n73804) );
  OAI21xp33_ASAP7_75t_SRAM U64699 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[15]), .A2(n3309), .B(
        n73817), .Y(n73801) );
  NAND2xp33_ASAP7_75t_SRAM U64700 ( .A(n72093), .B(n72065), .Y(n72066) );
  OAI21xp33_ASAP7_75t_SRAM U64701 ( .A1(n72281), .A2(n72282), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .Y(
        n72075) );
  OAI21xp33_ASAP7_75t_SRAM U64702 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .A2(
        n72238), .B(n72242), .Y(n72000) );
  OAI22xp33_ASAP7_75t_SRAM U64703 ( .A1(n72059), .A2(n72147), .B1(n72355), 
        .B2(n72068), .Y(n71990) );
  OAI21xp33_ASAP7_75t_SRAM U64704 ( .A1(n72441), .A2(n72440), .B(n57192), .Y(
        n72442) );
  OAI22xp33_ASAP7_75t_SRAM U64705 ( .A1(n72435), .A2(n72434), .B1(n59623), 
        .B2(n72432), .Y(n72439) );
  OAI21xp33_ASAP7_75t_SRAM U64706 ( .A1(n72027), .A2(n72050), .B(n58599), .Y(
        n71981) );
  AOI22xp33_ASAP7_75t_SRAM U64707 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_), 
        .A2(n57216), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_), 
        .B2(n57207), .Y(n71763) );
  AOI22xp33_ASAP7_75t_SRAM U64708 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), 
        .A2(n71888), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .B2(n58611), .Y(n71764) );
  AOI22xp33_ASAP7_75t_SRAM U64709 ( .A1(n72062), .A2(n72039), .B1(n72286), 
        .B2(n72038), .Y(n72043) );
  AOI22xp33_ASAP7_75t_SRAM U64710 ( .A1(n72093), .A2(n72091), .B1(n72105), 
        .B2(n72094), .Y(n72011) );
  AOI22xp33_ASAP7_75t_SRAM U64711 ( .A1(n72095), .A2(n72009), .B1(n72126), 
        .B2(n72092), .Y(n72012) );
  OAI21xp33_ASAP7_75t_SRAM U64712 ( .A1(n72367), .A2(n72309), .B(n57123), .Y(
        n72297) );
  AOI22xp33_ASAP7_75t_SRAM U64713 ( .A1(n72062), .A2(n72109), .B1(n72286), 
        .B2(n72125), .Y(n72018) );
  OAI21xp33_ASAP7_75t_SRAM U64714 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_), 
        .A2(n58422), .B(n71759), .Y(n71760) );
  OAI22xp33_ASAP7_75t_SRAM U64715 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_37_), 
        .A2(n57208), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_35_), 
        .B2(n71890), .Y(n71761) );
  AOI22xp33_ASAP7_75t_SRAM U64716 ( .A1(n72286), .A2(n72065), .B1(n72116), 
        .B2(n71924), .Y(n71925) );
  AOI22xp33_ASAP7_75t_SRAM U64717 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .A2(n57216), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), 
        .B2(n57207), .Y(n71854) );
  AOI22xp33_ASAP7_75t_SRAM U64718 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_), 
        .A2(n71888), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_), 
        .B2(n58611), .Y(n71855) );
  OAI22xp33_ASAP7_75t_SRAM U64719 ( .A1(n71984), .A2(n58608), .B1(n71952), 
        .B2(n58422), .Y(n71892) );
  AOI22xp33_ASAP7_75t_SRAM U64720 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .A2(n57216), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .B2(n57207), .Y(n71826) );
  AOI22xp33_ASAP7_75t_SRAM U64721 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_), 
        .A2(n71888), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_), 
        .B2(n58611), .Y(n71827) );
  OAI21xp33_ASAP7_75t_SRAM U64722 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_), 
        .A2(n71890), .B(n71857), .Y(n71858) );
  NOR2xp33_ASAP7_75t_SL U64723 ( .A(n72331), .B(n71906), .Y(n72020) );
  AOI22xp33_ASAP7_75t_SRAM U64724 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .A2(
        n72054), .B1(n71995), .B2(n71894), .Y(n71895) );
  NOR2xp33_ASAP7_75t_SL U64725 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        n72355), .Y(n72095) );
  AOI21xp33_ASAP7_75t_SRAM U64726 ( .A1(n72401), .A2(n72400), .B(n72399), .Y(
        n72408) );
  AOI22xp33_ASAP7_75t_SRAM U64727 ( .A1(n72286), .A2(n72092), .B1(n72110), 
        .B2(n71942), .Y(n71945) );
  O2A1O1Ixp5_ASAP7_75t_SL U64728 ( .A1(n72312), .A2(n72516), .B(n72247), .C(
        n72246), .Y(n72463) );
  AOI22xp33_ASAP7_75t_SRAM U64729 ( .A1(n72286), .A2(n72103), .B1(n72110), 
        .B2(n72125), .Y(n71889) );
  AOI21xp33_ASAP7_75t_SRAM U64730 ( .A1(n71943), .A2(n72286), .B(n71834), .Y(
        n71840) );
  OAI22xp33_ASAP7_75t_SRAM U64731 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_), 
        .A2(n57125), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_), 
        .B2(n57203), .Y(n72188) );
  AOI22xp33_ASAP7_75t_SRAM U64732 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_22_), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_), .B2(n71899), .Y(n71849) );
  AOI22xp33_ASAP7_75t_SRAM U64733 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_), 
        .A2(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_), 
        .B2(n71894), .Y(n71898) );
  AOI22xp33_ASAP7_75t_SRAM U64734 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), .B2(n72517), .Y(n71918) );
  OAI22xp33_ASAP7_75t_SRAM U64735 ( .A1(n72162), .A2(n57127), .B1(n57203), 
        .B2(n72132), .Y(n72134) );
  OAI22xp33_ASAP7_75t_SRAM U64736 ( .A1(n72147), .A2(n72087), .B1(n72355), 
        .B2(n72086), .Y(n72088) );
  NOR2xp33_ASAP7_75t_SL U64737 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .B(
        n72242), .Y(n72381) );
  OAI21xp33_ASAP7_75t_SRAM U64738 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .A2(
        n72341), .B(n71770), .Y(n71877) );
  OAI21xp33_ASAP7_75t_SRAM U64739 ( .A1(n72309), .A2(n58422), .B(n71753), .Y(
        n71754) );
  OAI22xp33_ASAP7_75t_SRAM U64740 ( .A1(n72307), .A2(n57208), .B1(n71890), 
        .B2(n72316), .Y(n71755) );
  NOR2xp33_ASAP7_75t_SL U64741 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .Y(
        n72286) );
  NOR2xp33_ASAP7_75t_SL U64742 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        n57192), .Y(n72393) );
  OAI21xp33_ASAP7_75t_SRAM U64743 ( .A1(n72367), .A2(n71952), .B(n57203), .Y(
        n71935) );
  INVxp33_ASAP7_75t_SRAM U64744 ( .A(n71702), .Y(n71699) );
  NOR2xp33_ASAP7_75t_SL U64745 ( .A(n59705), .B(n73689), .Y(n73786) );
  NOR2xp33_ASAP7_75t_SL U64746 ( .A(n73618), .B(n73817), .Y(n73793) );
  XNOR2xp5_ASAP7_75t_SL U64747 ( .A(n70213), .B(n70212), .Y(n70597) );
  NOR2xp33_ASAP7_75t_SL U64748 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[7]), .B(
        n70599), .Y(n70598) );
  NOR2xp33_ASAP7_75t_SL U64749 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[3]), .B(
        n70238), .Y(n70237) );
  NOR2xp33_ASAP7_75t_SL U64750 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[1]), .B(
        n70569), .Y(n70568) );
  NOR2xp33_ASAP7_75t_SL U64751 ( .A(n72242), .B(n72412), .Y(n72426) );
  NOR2xp33_ASAP7_75t_SL U64752 ( .A(n72175), .B(n57192), .Y(n72412) );
  NOR2xp33_ASAP7_75t_SL U64753 ( .A(n71983), .B(n57192), .Y(n72242) );
  NOR2xp33_ASAP7_75t_SL U64754 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .B(
        n57192), .Y(n72104) );
  NOR2xp33_ASAP7_75t_SL U64755 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        n72147), .Y(n72105) );
  NOR2xp33_ASAP7_75t_SL U64756 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .B(
        n57127), .Y(n71768) );
  NOR2xp33_ASAP7_75t_SL U64757 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .B(
        n72437), .Y(n72502) );
  OAI22xp33_ASAP7_75t_SRAM U64758 ( .A1(n72197), .A2(n57127), .B1(n57203), 
        .B2(n72162), .Y(n72166) );
  NOR2xp33_ASAP7_75t_SL U64759 ( .A(n71868), .B(n71867), .Y(n72322) );
  O2A1O1Ixp5_ASAP7_75t_SL U64760 ( .A1(n66128), .A2(n65625), .B(n65589), .C(
        n66090), .Y(n65607) );
  OAI21xp33_ASAP7_75t_SRAM U64761 ( .A1(n65653), .A2(n65578), .B(n65516), .Y(
        n66103) );
  AOI22xp33_ASAP7_75t_SRAM U64762 ( .A1(n66146), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[27]), .B1(n65593), 
        .B2(n66145), .Y(n65511) );
  OAI21xp33_ASAP7_75t_SRAM U64763 ( .A1(n65653), .A2(n65583), .B(n65509), .Y(
        n66102) );
  AOI22xp33_ASAP7_75t_SRAM U64764 ( .A1(n66146), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[31]), .B1(n65600), 
        .B2(n66145), .Y(n65504) );
  INVxp33_ASAP7_75t_SRAM U64765 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[15]), .Y(n65644) );
  O2A1O1Ixp5_ASAP7_75t_SL U64766 ( .A1(n59562), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[34]), .B(n66181), 
        .C(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[36]), .Y(n66163)
         );
  NOR2xp33_ASAP7_75t_SL U64767 ( .A(n65534), .B(n66111), .Y(n66137) );
  NOR2xp33_ASAP7_75t_SL U64768 ( .A(n74142), .B(n66135), .Y(n66166) );
  NAND3xp33_ASAP7_75t_SL U64769 ( .A(n65515), .B(n65642), .C(n65514), .Y(
        n66160) );
  NOR2xp33_ASAP7_75t_SL U64770 ( .A(n66150), .B(n65595), .Y(n66162) );
  AOI22xp33_ASAP7_75t_SRAM U64771 ( .A1(n66146), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[36]), .B1(n65611), 
        .B2(n66145), .Y(n65572) );
  OAI21xp33_ASAP7_75t_SRAM U64772 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]), .A2(n65805), .B(
        n65563), .Y(n66096) );
  NOR2xp33_ASAP7_75t_SL U64773 ( .A(n66095), .B(n65515), .Y(n66113) );
  NOR2xp33_ASAP7_75t_SL U64774 ( .A(n66091), .B(n66090), .Y(n66155) );
  AO21x1_ASAP7_75t_SL U64775 ( .A1(n71698), .A2(n71697), .B(n71712), .Y(n71710) );
  NOR2xp33_ASAP7_75t_SL U64776 ( .A(n72588), .B(n74232), .Y(n74245) );
  NOR2xp33_ASAP7_75t_SL U64777 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_3_), .B(
        n72582), .Y(n74235) );
  NOR2xp33_ASAP7_75t_SL U64778 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_0_), .B(
        n72564), .Y(n74098) );
  OAI21xp33_ASAP7_75t_SRAM U64779 ( .A1(n3088), .A2(n77480), .B(n61298), .Y(
        n9382) );
  OAI22xp33_ASAP7_75t_SRAM U64780 ( .A1(n65462), .A2(n65461), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[47]), .B2(n65460), 
        .Y(n65463) );
  AO21x1_ASAP7_75t_SL U64781 ( .A1(n77483), .A2(n3088), .B(n77482), .Y(n58421)
         );
  AOI211xp5_ASAP7_75t_SL U64782 ( .A1(n70033), .A2(n69907), .B(n69906), .C(
        n69905), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[16]) );
  O2A1O1Ixp5_ASAP7_75t_SL U64783 ( .A1(n66193), .A2(n65541), .B(n65540), .C(
        n65539), .Y(n65556) );
  XNOR2xp5_ASAP7_75t_SL U64784 ( .A(n72640), .B(n72639), .Y(n27982) );
  NOR2xp33_ASAP7_75t_SL U64785 ( .A(n69769), .B(n69768), .Y(n70067) );
  O2A1O1Ixp5_ASAP7_75t_SL U64786 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[6]), .A2(n65784), 
        .B(n65823), .C(n65431), .Y(n65432) );
  XNOR2xp5_ASAP7_75t_SL U64787 ( .A(n70131), .B(n70130), .Y(n3262) );
  NOR2xp33_ASAP7_75t_SL U64788 ( .A(n65404), .B(n65478), .Y(n65416) );
  NOR2xp33_ASAP7_75t_SL U64789 ( .A(n65452), .B(n65450), .Y(n65543) );
  O2A1O1Ixp5_ASAP7_75t_SL U64790 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]), .A2(n65761), 
        .B(n65831), .C(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), 
        .Y(n65412) );
  NOR2xp33_ASAP7_75t_SL U64791 ( .A(n65380), .B(n65660), .Y(n65423) );
  NOR2xp33_ASAP7_75t_SL U64792 ( .A(n65379), .B(n65456), .Y(n65409) );
  NOR2xp33_ASAP7_75t_SL U64793 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[46]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[45]), .Y(n65457) );
  NOR2xp33_ASAP7_75t_SL U64794 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[44]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .Y(n65421) );
  NOR3xp33_ASAP7_75t_SL U64795 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[47]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .Y(n65377) );
  NOR2xp33_ASAP7_75t_SL U64796 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[36]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[38]), .Y(n65544) );
  NOR2xp33_ASAP7_75t_SL U64797 ( .A(n78329), .B(n69560), .Y(n69900) );
  AOI21xp33_ASAP7_75t_SRAM U64798 ( .A1(n66052), .A2(n66070), .B(n65900), .Y(
        n65906) );
  XNOR2xp5_ASAP7_75t_SL U64799 ( .A(n72626), .B(n72632), .Y(n27981) );
  XNOR2xp5_ASAP7_75t_SL U64800 ( .A(n72616), .B(n72631), .Y(n72626) );
  NOR2xp33_ASAP7_75t_SL U64801 ( .A(n69897), .B(n69902), .Y(n70083) );
  NOR2xp33_ASAP7_75t_SL U64802 ( .A(n69458), .B(n69457), .Y(n69512) );
  AOI21xp33_ASAP7_75t_SRAM U64803 ( .A1(n66052), .A2(n65987), .B(n65811), .Y(
        n65812) );
  NOR2xp33_ASAP7_75t_SL U64804 ( .A(n69741), .B(n69740), .Y(n70043) );
  AOI21xp33_ASAP7_75t_SRAM U64805 ( .A1(n66052), .A2(n65991), .B(n65875), .Y(
        n65876) );
  OAI21xp33_ASAP7_75t_SRAM U64806 ( .A1(n65974), .A2(n65872), .B(n65968), .Y(
        n65873) );
  NOR2xp33_ASAP7_75t_SL U64807 ( .A(n66053), .B(n66052), .Y(n66057) );
  NOR2xp33_ASAP7_75t_SL U64808 ( .A(n66060), .B(n66051), .Y(n66053) );
  NOR2xp33_ASAP7_75t_SL U64809 ( .A(n69441), .B(n69440), .Y(n69943) );
  NAND2xp33_ASAP7_75t_SRAM U64810 ( .A(n65881), .B(n66052), .Y(n65884) );
  AOI22xp33_ASAP7_75t_SRAM U64811 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[13]), .A2(
        n69874), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]), .B2(
        n70038), .Y(n69875) );
  NOR2xp33_ASAP7_75t_SL U64812 ( .A(n69450), .B(n69449), .Y(n69811) );
  NOR2xp33_ASAP7_75t_SL U64813 ( .A(n69433), .B(n69432), .Y(n69809) );
  OAI22xp33_ASAP7_75t_SRAM U64814 ( .A1(n78345), .A2(n69564), .B1(n78343), 
        .B2(n69496), .Y(n69432) );
  NOR2xp33_ASAP7_75t_SL U64815 ( .A(n78341), .B(n69497), .Y(n69433) );
  NOR2xp33_ASAP7_75t_SL U64816 ( .A(n69424), .B(n69423), .Y(n69942) );
  OAI21xp33_ASAP7_75t_SRAM U64817 ( .A1(n66027), .A2(n65973), .B(n65968), .Y(
        n65923) );
  NOR2xp33_ASAP7_75t_SL U64818 ( .A(n66040), .B(n65980), .Y(n65950) );
  OAI21xp33_ASAP7_75t_SRAM U64819 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_), 
        .A2(n71993), .B(n71953), .Y(n71606) );
  AOI21xp33_ASAP7_75t_SRAM U64820 ( .A1(n72263), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_), 
        .Y(n71603) );
  NOR2xp33_ASAP7_75t_SL U64821 ( .A(n65797), .B(n65796), .Y(n65987) );
  NOR2xp33_ASAP7_75t_SL U64822 ( .A(n65795), .B(n65794), .Y(n65929) );
  NOR2xp33_ASAP7_75t_SL U64823 ( .A(n65895), .B(n65894), .Y(n66070) );
  NOR2xp33_ASAP7_75t_SL U64824 ( .A(n65790), .B(n65789), .Y(n65953) );
  NOR2xp33_ASAP7_75t_SL U64825 ( .A(n66060), .B(n66052), .Y(n66086) );
  NOR2xp33_ASAP7_75t_SL U64826 ( .A(n65749), .B(n66001), .Y(n65750) );
  OAI22xp33_ASAP7_75t_SRAM U64827 ( .A1(n65980), .A2(n65848), .B1(n65847), 
        .B2(n66052), .Y(n65869) );
  O2A1O1Ixp5_ASAP7_75t_SL U64828 ( .A1(n70021), .A2(n78333), .B(n69569), .C(
        n69568), .Y(n69883) );
  NOR2xp33_ASAP7_75t_SL U64829 ( .A(n71531), .B(n71532), .Y(n71537) );
  NOR2xp33_ASAP7_75t_SL U64830 ( .A(n71534), .B(n71535), .Y(n71533) );
  NOR2xp33_ASAP7_75t_SL U64831 ( .A(n71524), .B(n71523), .Y(n71527) );
  O2A1O1Ixp5_ASAP7_75t_SL U64832 ( .A1(n70079), .A2(n70118), .B(n69485), .C(
        n69484), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[45]) );
  O2A1O1Ixp5_ASAP7_75t_SL U64833 ( .A1(n69941), .A2(n69823), .B(n69483), .C(
        n69824), .Y(n69484) );
  NOR2xp33_ASAP7_75t_SL U64834 ( .A(n70114), .B(n69421), .Y(n70019) );
  NOR2xp33_ASAP7_75t_SL U64835 ( .A(n65764), .B(n65763), .Y(n66020) );
  NOR2xp33_ASAP7_75t_SL U64836 ( .A(n65748), .B(n65747), .Y(n65909) );
  NAND3xp33_ASAP7_75t_SL U64837 ( .A(n65756), .B(n65755), .C(n65754), .Y(
        n66047) );
  XNOR2xp5_ASAP7_75t_SL U64838 ( .A(n72633), .B(n72660), .Y(n27980) );
  XNOR2xp5_ASAP7_75t_SL U64839 ( .A(n72661), .B(n72662), .Y(n72633) );
  O2A1O1Ixp5_ASAP7_75t_SL U64840 ( .A1(n77642), .A2(n77641), .B(n77675), .C(
        n77640), .Y(n1704) );
  O2A1O1Ixp5_ASAP7_75t_SL U64841 ( .A1(n76472), .A2(n76473), .B(n74813), .C(
        n74784), .Y(n74785) );
  AOI21xp33_ASAP7_75t_SRAM U64842 ( .A1(n65723), .A2(n66052), .B(n65722), .Y(
        n65724) );
  AOI22xp33_ASAP7_75t_SRAM U64843 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .B2(n57194), .Y(n65717) );
  INVx1_ASAP7_75t_SL U64844 ( .A(n66060), .Y(n66049) );
  AOI22xp33_ASAP7_75t_SRAM U64845 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[45]), .A2(n57187), 
        .B1(n57188), .B2(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[44]), .Y(n65709) );
  AOI22xp33_ASAP7_75t_SRAM U64846 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[47]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[46]), .B2(n57194), .Y(n65710) );
  NOR2xp33_ASAP7_75t_SL U64847 ( .A(n58573), .B(n65696), .Y(n66075) );
  AO22x1_ASAP7_75t_SL U64848 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[3]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[2]), .B2(n57194), 
        .Y(n58573) );
  NOR2xp33_ASAP7_75t_SL U64849 ( .A(n65485), .B(n65484), .Y(n65691) );
  NOR2xp33_ASAP7_75t_SL U64850 ( .A(n58578), .B(n65679), .Y(n65966) );
  XNOR2xp5_ASAP7_75t_SL U64851 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[3]), .B(n65482), .Y(
        n65676) );
  OR2x2_ASAP7_75t_SL U64852 ( .A(n65828), .B(n65841), .Y(n58571) );
  OR2x2_ASAP7_75t_SL U64853 ( .A(n65808), .B(n65841), .Y(n58418) );
  OR2x2_ASAP7_75t_SL U64854 ( .A(n65828), .B(n65830), .Y(n58419) );
  OR2x2_ASAP7_75t_SL U64855 ( .A(n65808), .B(n65830), .Y(n58582) );
  NOR2xp33_ASAP7_75t_SL U64856 ( .A(n65496), .B(n65486), .Y(n65500) );
  NOR2xp33_ASAP7_75t_SL U64857 ( .A(n65665), .B(n65664), .Y(n66063) );
  NOR2xp33_ASAP7_75t_SL U64858 ( .A(n74894), .B(n65663), .Y(n65664) );
  AOI21xp33_ASAP7_75t_SRAM U64859 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_1_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_0_), .B(n78435), .Y(
        n65366) );
  INVxp33_ASAP7_75t_SRAM U64860 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_18_), .Y(n65367) );
  NOR2xp33_ASAP7_75t_SL U64861 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_0_), .B(
        n78437), .Y(n74817) );
  NOR2xp33_ASAP7_75t_SL U64862 ( .A(n74754), .B(n74808), .Y(n74920) );
  O2A1O1Ixp5_ASAP7_75t_SL U64863 ( .A1(n74807), .A2(n74806), .B(n74805), .C(
        n74804), .Y(n74826) );
  NAND2xp33_ASAP7_75t_SRAM U64864 ( .A(n59629), .B(n73006), .Y(n3339) );
  AOI22xp33_ASAP7_75t_SRAM U64865 ( .A1(n72993), .A2(n72992), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), 
        .B2(n72991), .Y(n72998) );
  NOR2xp33_ASAP7_75t_SL U64866 ( .A(n72853), .B(n73020), .Y(n72720) );
  AOI22xp33_ASAP7_75t_SRAM U64867 ( .A1(n73030), .A2(n72923), .B1(n73024), 
        .B2(n72921), .Y(n72871) );
  AOI22xp33_ASAP7_75t_SRAM U64868 ( .A1(n73030), .A2(n72912), .B1(n73028), 
        .B2(n72891), .Y(n72767) );
  O2A1O1Ixp5_ASAP7_75t_SL U64869 ( .A1(n77475), .A2(n77474), .B(n77473), .C(
        n77472), .Y(n77477) );
  INVxp33_ASAP7_75t_SRAM U64870 ( .A(n3086), .Y(n77471) );
  O2A1O1Ixp5_ASAP7_75t_SL U64871 ( .A1(n57189), .A2(n4092), .B(n7192), .C(
        n59700), .Y(n77804) );
  NOR2xp33_ASAP7_75t_SL U64872 ( .A(n833), .B(n77793), .Y(n77803) );
  XOR2xp5_ASAP7_75t_SL U64873 ( .A(n63313), .B(n63312), .Y(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N6) );
  NOR2xp33_ASAP7_75t_SL U64874 ( .A(n1125), .B(n75029), .Y(n75647) );
  NOR2xp33_ASAP7_75t_SL U64875 ( .A(n1129), .B(n66238), .Y(n75027) );
  NOR2xp33_ASAP7_75t_SL U64876 ( .A(n1133), .B(n66231), .Y(n66233) );
  NOR2xp33_ASAP7_75t_SL U64877 ( .A(n1137), .B(n66225), .Y(n66226) );
  NOR2xp33_ASAP7_75t_SL U64878 ( .A(n1143), .B(n1141), .Y(n75395) );
  NOR2xp33_ASAP7_75t_SL U64879 ( .A(n71698), .B(n71678), .Y(n71679) );
  NOR2xp33_ASAP7_75t_SL U64880 ( .A(n71653), .B(n71688), .Y(n71680) );
  NOR2xp33_ASAP7_75t_SL U64881 ( .A(n71787), .B(n71786), .Y(n71793) );
  AO21x1_ASAP7_75t_SL U64882 ( .A1(n71712), .A2(n71674), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_9_), .Y(
        n71799) );
  NOR2xp33_ASAP7_75t_SL U64883 ( .A(n71643), .B(n71636), .Y(n71662) );
  NOR2xp33_ASAP7_75t_SL U64884 ( .A(n71656), .B(n71645), .Y(n71670) );
  XNOR2xp5_ASAP7_75t_SL U64885 ( .A(n70180), .B(n70179), .Y(n3259) );
  NAND2xp33_ASAP7_75t_SRAM U64886 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .B(
        n72788), .Y(n72790) );
  O2A1O1Ixp5_ASAP7_75t_SL U64887 ( .A1(n72993), .A2(n72907), .B(n72753), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .Y(
        n72754) );
  NOR2xp33_ASAP7_75t_SL U64888 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_), 
        .B(n71547), .Y(n71599) );
  NOR2xp33_ASAP7_75t_SL U64889 ( .A(n71459), .B(n71635), .Y(n71616) );
  NOR2xp33_ASAP7_75t_SL U64890 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_22_), 
        .B(n71541), .Y(n71587) );
  NOR2xp33_ASAP7_75t_SL U64891 ( .A(n71632), .B(n71580), .Y(n71574) );
  NAND4xp25_ASAP7_75t_SL U64892 ( .A(n71542), .B(n71583), .C(n72005), .D(
        n72054), .Y(n71565) );
  NOR3xp33_ASAP7_75t_SL U64893 ( .A(n71551), .B(n71550), .C(n71549), .Y(n71542) );
  NOR2xp33_ASAP7_75t_SL U64894 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_), 
        .Y(n71561) );
  NOR2xp33_ASAP7_75t_SL U64895 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_), 
        .B(n71487), .Y(n71491) );
  NOR2xp33_ASAP7_75t_SL U64896 ( .A(n71471), .B(n71496), .Y(n71452) );
  NOR2xp33_ASAP7_75t_SL U64897 ( .A(n71437), .B(n71494), .Y(n71485) );
  NOR2xp33_ASAP7_75t_SL U64898 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .B(n71481), .Y(n71470) );
  NOR2xp33_ASAP7_75t_SL U64899 ( .A(n71418), .B(n71419), .Y(n71424) );
  NOR2xp33_ASAP7_75t_SL U64900 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_), 
        .B(n71480), .Y(n71428) );
  NOR2xp33_ASAP7_75t_SL U64901 ( .A(n71459), .B(n71462), .Y(n71505) );
  NOR2xp33_ASAP7_75t_SL U64902 ( .A(n71417), .B(n71474), .Y(n71469) );
  NAND3xp33_ASAP7_75t_SL U64903 ( .A(n71438), .B(n71548), .C(n72263), .Y(
        n71474) );
  NOR2xp33_ASAP7_75t_SL U64904 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_), 
        .Y(n71548) );
  NOR2xp33_ASAP7_75t_SL U64905 ( .A(n71601), .B(n71468), .Y(n71438) );
  NOR2xp33_ASAP7_75t_SL U64906 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_1_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_0_), 
        .Y(n71478) );
  NOR2xp33_ASAP7_75t_SL U64907 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_2_), 
        .Y(n71501) );
  NOR2xp33_ASAP7_75t_SL U64908 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_10_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_), 
        .Y(n71576) );
  NAND2xp33_ASAP7_75t_SRAM U64909 ( .A(n57081), .B(n70531), .Y(n70529) );
  NOR2xp33_ASAP7_75t_SL U64910 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .Y(
        n72876) );
  O2A1O1Ixp5_ASAP7_75t_SL U64911 ( .A1(n69773), .A2(n69772), .B(n69771), .C(
        n69774), .Y(n69782) );
  OAI21xp33_ASAP7_75t_SRAM U64912 ( .A1(n57081), .A2(n69937), .B(n69936), .Y(
        n69938) );
  NOR2xp33_ASAP7_75t_SL U64913 ( .A(n61305), .B(n61304), .Y(n77484) );
  O2A1O1Ixp5_ASAP7_75t_SL U64914 ( .A1(n62032), .A2(n62031), .B(n57073), .C(
        n62030), .Y(n62033) );
  O2A1O1Ixp5_ASAP7_75t_SL U64915 ( .A1(or1200_cpu_or1200_mult_mac_ex_freeze_r), 
        .A2(n75220), .B(n62029), .C(n62028), .Y(n62030) );
  INVxp33_ASAP7_75t_SRAM U64916 ( .A(n1494), .Y(n62027) );
  XNOR2xp5_ASAP7_75t_SL U64917 ( .A(n70751), .B(n70747), .Y(n70748) );
  O2A1O1Ixp5_ASAP7_75t_SL U64918 ( .A1(n65394), .A2(n65392), .B(n65355), .C(
        n65354), .Y(n65356) );
  O2A1O1Ixp5_ASAP7_75t_SL U64919 ( .A1(n70376), .A2(n70455), .B(n78234), .C(
        n70477), .Y(n70367) );
  O2A1O1Ixp5_ASAP7_75t_SL U64920 ( .A1(n70376), .A2(n70409), .B(n70334), .C(
        n70477), .Y(n70335) );
  O2A1O1Ixp5_ASAP7_75t_SL U64921 ( .A1(n70376), .A2(n70438), .B(n78235), .C(
        n70477), .Y(n70353) );
  O2A1O1Ixp5_ASAP7_75t_SL U64922 ( .A1(n70376), .A2(n70394), .B(n78236), .C(
        n70477), .Y(n70324) );
  O2A1O1Ixp5_ASAP7_75t_SL U64923 ( .A1(n70376), .A2(n70481), .B(n78233), .C(
        n70477), .Y(n70377) );
  O2A1O1Ixp5_ASAP7_75t_SL U64924 ( .A1(n70478), .A2(n70438), .B(n70436), .C(
        n70477), .Y(n70437) );
  O2A1O1Ixp5_ASAP7_75t_SL U64925 ( .A1(n70478), .A2(n70409), .B(n78231), .C(
        n70477), .Y(n70408) );
  O2A1O1Ixp5_ASAP7_75t_SL U64926 ( .A1(n70478), .A2(n70455), .B(n78230), .C(
        n70477), .Y(n70454) );
  O2A1O1Ixp5_ASAP7_75t_SL U64927 ( .A1(n70478), .A2(n70394), .B(n78232), .C(
        n70477), .Y(n70393) );
  O2A1O1Ixp5_ASAP7_75t_SL U64928 ( .A1(n70478), .A2(n70481), .B(n78229), .C(
        n70477), .Y(n70479) );
  O2A1O1Ixp5_ASAP7_75t_SL U64929 ( .A1(n70303), .A2(n70419), .B(n78240), .C(
        n70477), .Y(n70271) );
  O2A1O1Ixp5_ASAP7_75t_SL U64930 ( .A1(n70303), .A2(n70438), .B(n78239), .C(
        n70477), .Y(n70282) );
  O2A1O1Ixp5_ASAP7_75t_SL U64931 ( .A1(n70303), .A2(n70394), .B(n78241), .C(
        n70477), .Y(n70256) );
  O2A1O1Ixp5_ASAP7_75t_SL U64932 ( .A1(n70303), .A2(n70455), .B(n78238), .C(
        n70477), .Y(n70290) );
  O2A1O1Ixp5_ASAP7_75t_SL U64933 ( .A1(n70303), .A2(n70409), .B(n70262), .C(
        n70477), .Y(n70263) );
  O2A1O1Ixp5_ASAP7_75t_SL U64934 ( .A1(n70303), .A2(n70481), .B(n78237), .C(
        n70477), .Y(n70304) );
  OAI21xp33_ASAP7_75t_SRAM U64935 ( .A1(n57081), .A2(n69990), .B(n69989), .Y(
        n69991) );
  O2A1O1Ixp5_ASAP7_75t_SL U64936 ( .A1(n63507), .A2(n63510), .B(n63492), .C(
        n76897), .Y(n63493) );
  NAND2xp33_ASAP7_75t_SRAM U64937 ( .A(n59629), .B(n72985), .Y(n1546) );
  NOR2xp33_ASAP7_75t_SL U64938 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .B(
        n72727), .Y(n72744) );
  NOR2xp33_ASAP7_75t_SL U64939 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), .B(
        n72999), .Y(n73028) );
  NOR2xp33_ASAP7_75t_SL U64940 ( .A(n72862), .B(n72861), .Y(n72974) );
  NOR2xp33_ASAP7_75t_SL U64941 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .B(
        n72993), .Y(n73030) );
  NOR2xp33_ASAP7_75t_SL U64942 ( .A(n72990), .B(n72976), .Y(n73037) );
  AOI22xp33_ASAP7_75t_SRAM U64943 ( .A1(n72961), .A2(n73040), .B1(n73042), 
        .B2(n72956), .Y(n72957) );
  NOR2xp33_ASAP7_75t_SL U64944 ( .A(n72954), .B(n72953), .Y(n72961) );
  NAND2xp33_ASAP7_75t_SRAM U64945 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .B(
        n72955), .Y(n72950) );
  NOR2xp33_ASAP7_75t_SL U64946 ( .A(n72949), .B(n72948), .Y(n72952) );
  NOR2xp33_ASAP7_75t_SL U64947 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), .Y(
        n73024) );
  NOR2xp33_ASAP7_75t_SL U64948 ( .A(n72932), .B(n72931), .Y(n72943) );
  AOI21xp33_ASAP7_75t_SRAM U64949 ( .A1(n72927), .A2(n73008), .B(n72921), .Y(
        n72922) );
  NOR2xp33_ASAP7_75t_SL U64950 ( .A(n72923), .B(n72920), .Y(n72947) );
  NAND2xp33_ASAP7_75t_SRAM U64951 ( .A(n72915), .B(n72935), .Y(n72895) );
  NOR2xp33_ASAP7_75t_SL U64952 ( .A(n72772), .B(n72771), .Y(n72915) );
  NOR2xp33_ASAP7_75t_SL U64953 ( .A(n78341), .B(n57190), .Y(n72772) );
  NOR2xp33_ASAP7_75t_SL U64954 ( .A(n78432), .B(n57190), .Y(n72722) );
  NOR2xp33_ASAP7_75t_SL U64955 ( .A(n78352), .B(n57190), .Y(n72740) );
  NOR2xp33_ASAP7_75t_SL U64956 ( .A(n72698), .B(n72697), .Y(n72898) );
  NOR2xp33_ASAP7_75t_SL U64957 ( .A(n78357), .B(n57190), .Y(n72698) );
  NOR2xp33_ASAP7_75t_SL U64958 ( .A(n72684), .B(n72683), .Y(n72886) );
  NOR2xp33_ASAP7_75t_SL U64959 ( .A(n78369), .B(n57190), .Y(n72684) );
  NOR2xp33_ASAP7_75t_SL U64960 ( .A(n72686), .B(n72685), .Y(n72888) );
  NOR2xp33_ASAP7_75t_SL U64961 ( .A(n78365), .B(n57190), .Y(n72686) );
  NOR2xp33_ASAP7_75t_SL U64962 ( .A(n72858), .B(n72857), .Y(n73029) );
  NOR2xp33_ASAP7_75t_SL U64963 ( .A(n78434), .B(n59626), .Y(n72858) );
  INVx1_ASAP7_75t_SL U64964 ( .A(n59629), .Y(n59628) );
  O2A1O1Ixp5_ASAP7_75t_SL U64965 ( .A1(n68799), .A2(n68815), .B(n76884), .C(
        n76906), .Y(n68800) );
  O2A1O1Ixp5_ASAP7_75t_SL U64966 ( .A1(n68820), .A2(n74999), .B(n68785), .C(
        n68784), .Y(n68786) );
  XNOR2xp5_ASAP7_75t_SL U64967 ( .A(or1200_cpu_or1200_mult_mac_n315), .B(
        n63485), .Y(n63507) );
  O2A1O1Ixp5_ASAP7_75t_SL U64968 ( .A1(n63786), .A2(n63785), .B(n63784), .C(
        n76906), .Y(n63787) );
  O2A1O1Ixp5_ASAP7_75t_SL U64969 ( .A1(n63773), .A2(n63772), .B(n63771), .C(
        n76897), .Y(n63788) );
  O2A1O1Ixp5_ASAP7_75t_SL U64970 ( .A1(n65156), .A2(n76906), .B(n65155), .C(
        n65154), .Y(n65157) );
  O2A1O1Ixp5_ASAP7_75t_SL U64971 ( .A1(n75019), .A2(n76906), .B(n75003), .C(
        n75002), .Y(n75004) );
  O2A1O1Ixp5_ASAP7_75t_SL U64972 ( .A1(n63356), .A2(n63355), .B(n63354), .C(
        n76897), .Y(n63357) );
  O2A1O1Ixp5_ASAP7_75t_SL U64973 ( .A1(n63330), .A2(n63336), .B(n63329), .C(
        n76906), .Y(n63331) );
  O2A1O1Ixp5_ASAP7_75t_SL U64974 ( .A1(n63328), .A2(n63318), .B(n63317), .C(
        n76897), .Y(n63332) );
  XOR2xp5_ASAP7_75t_SL U64975 ( .A(n63305), .B(n63287), .Y(n63288) );
  XOR2xp5_ASAP7_75t_SL U64976 ( .A(n63389), .B(n63284), .Y(n63290) );
  XOR2xp5_ASAP7_75t_SL U64977 ( .A(n63426), .B(n63415), .Y(n63407) );
  NAND2xp5_ASAP7_75t_SL U64978 ( .A(n59493), .B(n63266), .Y(n68787) );
  NOR2xp33_ASAP7_75t_SL U64979 ( .A(n72625), .B(n72624), .Y(n72636) );
  INVx1_ASAP7_75t_SL U64980 ( .A(n59629), .Y(n59627) );
  NOR2xp33_ASAP7_75t_SL U64981 ( .A(n72629), .B(n72657), .Y(n72662) );
  NOR2xp33_ASAP7_75t_SL U64982 ( .A(n72645), .B(n1558), .Y(n72657) );
  NOR2xp33_ASAP7_75t_SL U64983 ( .A(n72628), .B(n72667), .Y(n72629) );
  INVx1_ASAP7_75t_SL U64984 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_29_), 
        .Y(n78363) );
  NOR2xp33_ASAP7_75t_SL U64985 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_), .B(n78381), .Y(
        n72600) );
  NOR2xp33_ASAP7_75t_SL U64986 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_), .B(n78371), .Y(n72602)
         );
  AOI22xp33_ASAP7_75t_SRAM U64987 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_), .A2(n78376), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_), .B2(n78379), .Y(
        n72598) );
  NOR2xp33_ASAP7_75t_SL U64988 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_30_), .B(n78382), .Y(n72609)
         );
  NOR2xp33_ASAP7_75t_SL U64989 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_), .Y(n72654) );
  NOR2xp33_ASAP7_75t_SL U64990 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_29_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_), .Y(n72643) );
  NOR2xp33_ASAP7_75t_SL U64991 ( .A(n72665), .B(n72664), .Y(n72663) );
  NOR2xp33_ASAP7_75t_SL U64992 ( .A(n72614), .B(n72619), .Y(n72642) );
  NOR2xp33_ASAP7_75t_SL U64993 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_), .Y(n72621) );
  NOR2xp33_ASAP7_75t_SL U64994 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .Y(n72620) );
  OR2x2_ASAP7_75t_SL U64995 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_27_), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_), .Y(n72665) );
  NOR2xp33_ASAP7_75t_SL U64996 ( .A(n72964), .B(n58572), .Y(n72645) );
  XNOR2xp5_ASAP7_75t_SL U64997 ( .A(n70196), .B(n53435), .Y(n3257) );
  NOR2xp33_ASAP7_75t_SL U64998 ( .A(n63348), .B(n63347), .Y(n63369) );
  XOR2xp5_ASAP7_75t_SL U64999 ( .A(n63344), .B(n63343), .Y(n63348) );
  XNOR2xp5_ASAP7_75t_SL U65000 ( .A(n69181), .B(n75291), .Y(n69186) );
  O2A1O1Ixp5_ASAP7_75t_SL U65001 ( .A1(n57074), .A2(n2093), .B(n77553), .C(
        n77552), .Y(n9223) );
  O2A1O1Ixp5_ASAP7_75t_SL U65002 ( .A1(n59689), .A2(n2165), .B(n77534), .C(
        n77552), .Y(n9229) );
  AOI22xp33_ASAP7_75t_SRAM U65003 ( .A1(n65357), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_5_), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_r_a), .B2(n65401), .Y(
        n65350) );
  NOR2xp33_ASAP7_75t_SL U65004 ( .A(n1776), .B(n59689), .Y(n61123) );
  NOR2xp33_ASAP7_75t_SL U65005 ( .A(or1200_cpu_or1200_except_n687), .B(n76669), 
        .Y(n76676) );
  NOR2xp33_ASAP7_75t_SL U65006 ( .A(n69131), .B(n69133), .Y(n69132) );
  O2A1O1Ixp5_ASAP7_75t_SL U65007 ( .A1(n1145), .A2(n75390), .B(n74977), .C(
        n75645), .Y(n74978) );
  NOR2xp33_ASAP7_75t_SL U65008 ( .A(n1149), .B(n74975), .Y(n62551) );
  NOR2xp33_ASAP7_75t_SL U65009 ( .A(n76805), .B(n76806), .Y(n77282) );
  OAI21xp33_ASAP7_75t_SRAM U65010 ( .A1(n74716), .A2(n74715), .B(n74714), .Y(
        n74717) );
  NOR2xp33_ASAP7_75t_SL U65011 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_), .Y(
        n74680) );
  AOI21xp33_ASAP7_75t_SRAM U65012 ( .A1(n74679), .A2(n74682), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_5_), .Y(
        n74675) );
  OAI21xp33_ASAP7_75t_SRAM U65013 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .A2(
        n2345), .B(n74646), .Y(n74647) );
  OAI21xp33_ASAP7_75t_SRAM U65014 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_), .A2(
        n74645), .B(n2335), .Y(n74649) );
  XNOR2xp5_ASAP7_75t_SL U65015 ( .A(n63450), .B(n63449), .Y(n52048) );
  INVx1_ASAP7_75t_SL U65016 ( .A(n77233), .Y(n59680) );
  NOR4xp25_ASAP7_75t_SL U65017 ( .A(n77206), .B(n77200), .C(n77161), .D(n76540), .Y(n77683) );
  NOR2xp33_ASAP7_75t_SL U65018 ( .A(n76539), .B(n76609), .Y(n77160) );
  NOR2xp33_ASAP7_75t_SL U65019 ( .A(n1753), .B(n1961), .Y(n76609) );
  NOR2xp33_ASAP7_75t_SL U65020 ( .A(n62210), .B(n62209), .Y(n75649) );
  NOR2xp33_ASAP7_75t_SL U65021 ( .A(n63915), .B(n63914), .Y(n75386) );
  NAND4xp25_ASAP7_75t_SL U65022 ( .A(n63913), .B(n63912), .C(n63911), .D(
        n63910), .Y(n63914) );
  NOR2xp33_ASAP7_75t_SL U65023 ( .A(n1175), .B(n1149), .Y(n63910) );
  NOR2xp33_ASAP7_75t_SL U65024 ( .A(n1151), .B(n1169), .Y(n63911) );
  NOR4xp25_ASAP7_75t_SL U65025 ( .A(n1155), .B(n1159), .C(n1173), .D(n1167), 
        .Y(n63907) );
  NOR4xp25_ASAP7_75t_SL U65026 ( .A(n1153), .B(n1183), .C(n1157), .D(n1171), 
        .Y(n63908) );
  NOR2xp33_ASAP7_75t_SL U65027 ( .A(n75648), .B(n62549), .Y(n74975) );
  NOR2xp33_ASAP7_75t_SL U65028 ( .A(n1151), .B(n62496), .Y(n62549) );
  NOR2xp33_ASAP7_75t_SL U65029 ( .A(n1155), .B(n62488), .Y(n62491) );
  NOR2xp33_ASAP7_75t_SL U65030 ( .A(n1183), .B(n62407), .Y(n62483) );
  NOR2xp33_ASAP7_75t_SL U65031 ( .A(n1169), .B(n62233), .Y(n62303) );
  NOR2xp33_ASAP7_75t_SL U65032 ( .A(n62219), .B(n62218), .Y(n62228) );
  NOR2xp33_ASAP7_75t_SL U65033 ( .A(n1179), .B(n1177), .Y(n63912) );
  NOR2xp33_ASAP7_75t_SL U65034 ( .A(n1428), .B(n62201), .Y(n62203) );
  NOR2xp33_ASAP7_75t_SL U65035 ( .A(n74974), .B(n75645), .Y(n74976) );
  NAND4xp25_ASAP7_75t_SL U65036 ( .A(n62191), .B(n62190), .C(n62189), .D(
        n62188), .Y(n62192) );
  XNOR2xp5_ASAP7_75t_SL U65037 ( .A(n1179), .B(n1486), .Y(n62188) );
  XNOR2xp5_ASAP7_75t_SL U65038 ( .A(n1147), .B(n1452), .Y(n62189) );
  XNOR2xp5_ASAP7_75t_SL U65039 ( .A(n1171), .B(n1478), .Y(n62190) );
  XNOR2xp5_ASAP7_75t_SL U65040 ( .A(n1135), .B(n1440), .Y(n62191) );
  NAND4xp25_ASAP7_75t_SL U65041 ( .A(n62187), .B(n62186), .C(n62185), .D(
        n62184), .Y(n62193) );
  XNOR2xp5_ASAP7_75t_SL U65042 ( .A(n1149), .B(n1454), .Y(n62184) );
  XNOR2xp5_ASAP7_75t_SL U65043 ( .A(n1173), .B(n1480), .Y(n62185) );
  XNOR2xp5_ASAP7_75t_SL U65044 ( .A(n1161), .B(n1468), .Y(n62186) );
  XNOR2xp5_ASAP7_75t_SL U65045 ( .A(n1169), .B(n1476), .Y(n62187) );
  NAND4xp25_ASAP7_75t_SL U65046 ( .A(n62183), .B(n62182), .C(n62181), .D(
        n62180), .Y(n62194) );
  XNOR2xp5_ASAP7_75t_SL U65047 ( .A(n1157), .B(n1462), .Y(n62180) );
  XNOR2xp5_ASAP7_75t_SL U65048 ( .A(n1139), .B(n1444), .Y(n62181) );
  XNOR2xp5_ASAP7_75t_SL U65049 ( .A(n1151), .B(n1456), .Y(n62182) );
  XNOR2xp5_ASAP7_75t_SL U65050 ( .A(n1159), .B(n1466), .Y(n62183) );
  XNOR2xp5_ASAP7_75t_SL U65051 ( .A(n1141), .B(n1446), .Y(n62174) );
  XNOR2xp5_ASAP7_75t_SL U65052 ( .A(n1137), .B(n1442), .Y(n62175) );
  XNOR2xp5_ASAP7_75t_SL U65053 ( .A(n1133), .B(n1438), .Y(n62176) );
  XNOR2xp5_ASAP7_75t_SL U65054 ( .A(n1145), .B(n1450), .Y(n62177) );
  XNOR2xp5_ASAP7_75t_SL U65055 ( .A(n1163), .B(n1470), .Y(n62170) );
  XNOR2xp5_ASAP7_75t_SL U65056 ( .A(n1131), .B(n1436), .Y(n62171) );
  XNOR2xp5_ASAP7_75t_SL U65057 ( .A(n1155), .B(n1460), .Y(n62172) );
  XNOR2xp5_ASAP7_75t_SL U65058 ( .A(n1129), .B(n1434), .Y(n62173) );
  NOR2xp33_ASAP7_75t_SL U65059 ( .A(n62169), .B(n62168), .Y(n62197) );
  NAND4xp25_ASAP7_75t_SL U65060 ( .A(n62167), .B(n62166), .C(n62165), .D(
        n62164), .Y(n62168) );
  XNOR2xp5_ASAP7_75t_SL U65061 ( .A(n1177), .B(n1484), .Y(n62164) );
  XNOR2xp5_ASAP7_75t_SL U65062 ( .A(n1143), .B(n1448), .Y(n62165) );
  XNOR2xp5_ASAP7_75t_SL U65063 ( .A(n1167), .B(n1474), .Y(n62166) );
  XNOR2xp5_ASAP7_75t_SL U65064 ( .A(n1127), .B(n1432), .Y(n62167) );
  NAND4xp25_ASAP7_75t_SL U65065 ( .A(n62163), .B(n62162), .C(n62161), .D(
        n62160), .Y(n62169) );
  XNOR2xp5_ASAP7_75t_SL U65066 ( .A(n1153), .B(n1458), .Y(n62160) );
  XNOR2xp5_ASAP7_75t_SL U65067 ( .A(n1183), .B(n1464), .Y(n62161) );
  XNOR2xp5_ASAP7_75t_SL U65068 ( .A(n1165), .B(n1472), .Y(n62162) );
  XNOR2xp5_ASAP7_75t_SL U65069 ( .A(n1175), .B(n1482), .Y(n62163) );
  O2A1O1Ixp5_ASAP7_75t_SL U65070 ( .A1(n76958), .A2(n76957), .B(n76956), .C(
        n76955), .Y(n76960) );
  INVxp33_ASAP7_75t_SRAM U65071 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_22_), .Y(n76938)
         );
  INVxp33_ASAP7_75t_SRAM U65072 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_20_), .Y(n76966)
         );
  XNOR2xp5_ASAP7_75t_SL U65073 ( .A(or1200_cpu_or1200_mult_mac_n255), .B(
        or1200_cpu_or1200_mult_mac_n401), .Y(n69314) );
  NOR2xp33_ASAP7_75t_SL U65074 ( .A(n68945), .B(n68944), .Y(n68993) );
  NOR2xp33_ASAP7_75t_SL U65075 ( .A(n68844), .B(n68843), .Y(n68878) );
  NOR2xp33_ASAP7_75t_SL U65076 ( .A(n3092), .B(n77486), .Y(n61998) );
  O2A1O1Ixp5_ASAP7_75t_SL U65077 ( .A1(n69331), .A2(n2755), .B(n69330), .C(
        n77454), .Y(n9392) );
  NOR2xp33_ASAP7_75t_SL U65078 ( .A(n65499), .B(n65498), .Y(n76977) );
  NOR2xp33_ASAP7_75t_SL U65079 ( .A(n66197), .B(n65533), .Y(n65498) );
  NOR2xp33_ASAP7_75t_SL U65080 ( .A(n65525), .B(n65492), .Y(n65499) );
  O2A1O1Ixp5_ASAP7_75t_SL U65081 ( .A1(n74941), .A2(n58559), .B(n74940), .C(
        n74939), .Y(n77446) );
  AOI211xp5_ASAP7_75t_SL U65082 ( .A1(n77125), .A2(n61374), .B(n61373), .C(
        n77122), .Y(n61375) );
  XNOR2xp5_ASAP7_75t_SL U65083 ( .A(or1200_cpu_or1200_except_n506), .B(n62333), 
        .Y(n61364) );
  O2A1O1Ixp5_ASAP7_75t_SL U65084 ( .A1(n59543), .A2(n75227), .B(n61346), .C(
        n59542), .Y(n61352) );
  NOR2xp33_ASAP7_75t_SL U65085 ( .A(n61345), .B(n62250), .Y(n77612) );
  INVxp33_ASAP7_75t_SRAM U65086 ( .A(n1392), .Y(n61328) );
  OAI21xp33_ASAP7_75t_SRAM U65087 ( .A1(n1390), .A2(n76716), .B(n61325), .Y(
        n61332) );
  AOI22xp33_ASAP7_75t_SRAM U65088 ( .A1(n1468), .A2(n76712), .B1(n76711), .B2(
        n1161), .Y(n61324) );
  O2A1O1Ixp5_ASAP7_75t_SL U65089 ( .A1(n61753), .A2(n61609), .B(n61608), .C(
        n61607), .Y(n61611) );
  OAI22xp33_ASAP7_75t_SRAM U65090 ( .A1(or1200_cpu_or1200_mult_mac_n151), .A2(
        n64275), .B1(or1200_cpu_or1200_mult_mac_n215), .B2(n77633), .Y(n61604)
         );
  INVxp33_ASAP7_75t_SRAM U65091 ( .A(or1200_cpu_or1200_mult_mac_n112), .Y(
        n62365) );
  O2A1O1Ixp5_ASAP7_75t_SL U65092 ( .A1(n62351), .A2(n62350), .B(n76750), .C(
        n62349), .Y(n62352) );
  AOI22xp33_ASAP7_75t_SRAM U65093 ( .A1(n76713), .A2(n62316), .B1(n76634), 
        .B2(n63253), .Y(n62323) );
  INVxp33_ASAP7_75t_SRAM U65094 ( .A(n3141), .Y(n62326) );
  NOR2xp33_ASAP7_75t_SL U65095 ( .A(n62298), .B(n62297), .Y(n76628) );
  NOR2xp33_ASAP7_75t_SL U65096 ( .A(n62251), .B(n62250), .Y(n77602) );
  AOI21xp33_ASAP7_75t_SRAM U65097 ( .A1(n76735), .A2(n62244), .B(n62243), .Y(
        n62245) );
  OAI22xp33_ASAP7_75t_SRAM U65098 ( .A1(or1200_cpu_or1200_mult_mac_n217), .A2(
        n77633), .B1(n1404), .B2(n77035), .Y(n62238) );
  AOI22xp33_ASAP7_75t_SRAM U65099 ( .A1(n1474), .A2(n76712), .B1(n76711), .B2(
        n1167), .Y(n62235) );
  INVxp33_ASAP7_75t_SRAM U65100 ( .A(n1536), .Y(n62244) );
  NOR2xp33_ASAP7_75t_SL U65101 ( .A(n63498), .B(n63497), .Y(n63499) );
  O2A1O1Ixp5_ASAP7_75t_SL U65102 ( .A1(n59558), .A2(n75227), .B(n61524), .C(
        n59557), .Y(n61537) );
  XNOR2xp5_ASAP7_75t_SL U65103 ( .A(n61487), .B(n62288), .Y(n61517) );
  INVxp33_ASAP7_75t_SRAM U65104 ( .A(n1416), .Y(n61474) );
  INVxp33_ASAP7_75t_SRAM U65105 ( .A(n1480), .Y(n61470) );
  INVxp33_ASAP7_75t_SRAM U65106 ( .A(n3418), .Y(n61464) );
  AOI211xp5_ASAP7_75t_SL U65107 ( .A1(n76735), .A2(n61390), .B(n61389), .C(
        n61388), .Y(n61392) );
  OAI22xp33_ASAP7_75t_SRAM U65108 ( .A1(or1200_cpu_or1200_mult_mac_n149), .A2(
        n64275), .B1(n1412), .B2(n77035), .Y(n61383) );
  OAI21xp33_ASAP7_75t_SRAM U65109 ( .A1(n1410), .A2(n76716), .B(n61380), .Y(
        n61385) );
  AOI22xp33_ASAP7_75t_SRAM U65110 ( .A1(n1478), .A2(n76712), .B1(n76711), .B2(
        n1171), .Y(n61379) );
  O2A1O1Ixp5_ASAP7_75t_SL U65111 ( .A1(n76790), .A2(n76789), .B(n57126), .C(
        n76788), .Y(n76800) );
  O2A1O1Ixp5_ASAP7_75t_SL U65112 ( .A1(n76758), .A2(n76757), .B(n76756), .C(
        n76755), .Y(n76790) );
  NOR2xp33_ASAP7_75t_SL U65113 ( .A(n61263), .B(n61262), .Y(n61267) );
  INVxp33_ASAP7_75t_SRAM U65114 ( .A(n1420), .Y(n61250) );
  OAI21xp33_ASAP7_75t_SRAM U65115 ( .A1(n1418), .A2(n76716), .B(n61247), .Y(
        n61254) );
  AOI22xp33_ASAP7_75t_SRAM U65116 ( .A1(n1482), .A2(n76712), .B1(n76711), .B2(
        n1175), .Y(n61246) );
  O2A1O1Ixp5_ASAP7_75t_SL U65117 ( .A1(n59568), .A2(n75227), .B(n76775), .C(
        n59708), .Y(n61217) );
  AOI211xp5_ASAP7_75t_SL U65118 ( .A1(n77128), .A2(n77665), .B(n64854), .C(
        n58286), .Y(n64861) );
  O2A1O1Ixp5_ASAP7_75t_SL U65119 ( .A1(n57212), .A2(n75735), .B(n64830), .C(
        n1571), .Y(n64831) );
  AOI21xp33_ASAP7_75t_SRAM U65120 ( .A1(n64829), .A2(n57126), .B(n64828), .Y(
        n64833) );
  O2A1O1Ixp5_ASAP7_75t_SL U65121 ( .A1(n75701), .A2(n74607), .B(n77078), .C(
        n75699), .Y(n60852) );
  INVxp33_ASAP7_75t_SRAM U65122 ( .A(n1374), .Y(n60820) );
  O2A1O1Ixp5_ASAP7_75t_SL U65123 ( .A1(n73969), .A2(n73992), .B(n75852), .C(
        n60793), .Y(n60794) );
  O2A1O1Ixp5_ASAP7_75t_SL U65124 ( .A1(n59573), .A2(n75227), .B(n76775), .C(
        n59548), .Y(n73939) );
  INVxp33_ASAP7_75t_SRAM U65125 ( .A(or1200_cpu_or1200_mult_mac_n195), .Y(
        n73920) );
  O2A1O1Ixp5_ASAP7_75t_SL U65126 ( .A1(n3132), .A2(n77133), .B(n57073), .C(
        n77132), .Y(n77135) );
  INVxp33_ASAP7_75t_SRAM U65127 ( .A(n3392), .Y(n69346) );
  AOI21xp33_ASAP7_75t_SRAM U65128 ( .A1(n76735), .A2(n61688), .B(n61687), .Y(
        n61689) );
  OAI22xp33_ASAP7_75t_SRAM U65129 ( .A1(or1200_cpu_or1200_mult_mac_n163), .A2(
        n64275), .B1(n1384), .B2(n77035), .Y(n61682) );
  OAI21xp33_ASAP7_75t_SRAM U65130 ( .A1(n1115), .A2(n76716), .B(n61679), .Y(
        n61684) );
  AOI22xp33_ASAP7_75t_SRAM U65131 ( .A1(n1464), .A2(n76712), .B1(n76711), .B2(
        n1183), .Y(n61678) );
  INVxp33_ASAP7_75t_SRAM U65132 ( .A(n1112), .Y(n61688) );
  O2A1O1Ixp5_ASAP7_75t_SL U65133 ( .A1(n63586), .A2(n75735), .B(n75338), .C(
        n59533), .Y(n63587) );
  INVxp33_ASAP7_75t_SRAM U65134 ( .A(n1358), .Y(n63552) );
  OAI21xp33_ASAP7_75t_SRAM U65135 ( .A1(n76232), .A2(n62515), .B(n77082), .Y(
        n62541) );
  NOR2xp33_ASAP7_75t_SL U65136 ( .A(n62513), .B(n62512), .Y(n77649) );
  OAI22xp33_ASAP7_75t_SRAM U65137 ( .A1(n1366), .A2(n77035), .B1(n1364), .B2(
        n75364), .Y(n62504) );
  INVx3_ASAP7_75t_SL U65138 ( .A(n59695), .Y(n59688) );
  NOR2xp33_ASAP7_75t_SL U65139 ( .A(n62468), .B(n62467), .Y(n77902) );
  AOI21xp33_ASAP7_75t_SRAM U65140 ( .A1(n73921), .A2(n63452), .B(n62428), .Y(
        n62429) );
  OAI22xp33_ASAP7_75t_SRAM U65141 ( .A1(or1200_cpu_or1200_mult_mac_n229), .A2(
        n74587), .B1(n1380), .B2(n75364), .Y(n62410) );
  OAI22xp33_ASAP7_75t_SRAM U65142 ( .A1(or1200_cpu_or1200_mult_mac_n165), .A2(
        n64275), .B1(n1382), .B2(n77035), .Y(n62411) );
  XNOR2xp5_ASAP7_75t_SL U65143 ( .A(n61830), .B(n61763), .Y(n61794) );
  NOR2xp33_ASAP7_75t_SL U65144 ( .A(n61181), .B(n61180), .Y(n64853) );
  NOR2xp33_ASAP7_75t_SL U65145 ( .A(n61344), .B(n61618), .Y(n62250) );
  INVxp33_ASAP7_75t_SRAM U65146 ( .A(or1200_cpu_or1200_mult_mac_n161), .Y(
        n61777) );
  INVxp33_ASAP7_75t_SRAM U65147 ( .A(n1388), .Y(n61748) );
  INVxp33_ASAP7_75t_SRAM U65148 ( .A(n1466), .Y(n61744) );
  AOI211xp5_ASAP7_75t_SL U65149 ( .A1(n77128), .A2(n77653), .B(n64143), .C(
        n64216), .Y(n64144) );
  INVxp33_ASAP7_75t_SRAM U65150 ( .A(or1200_cpu_or1200_mult_mac_n88), .Y(
        n64124) );
  NAND3xp33_ASAP7_75t_SL U65151 ( .A(n61310), .B(n58613), .C(n61147), .Y(
        n76557) );
  NAND2xp33_ASAP7_75t_SRAM U65152 ( .A(n62382), .B(n61084), .Y(n61093) );
  NOR2xp33_ASAP7_75t_SL U65153 ( .A(n60882), .B(n77122), .Y(n62459) );
  NOR2xp33_ASAP7_75t_SL U65154 ( .A(n2607), .B(n76787), .Y(n77122) );
  O2A1O1Ixp5_ASAP7_75t_SL U65155 ( .A1(n73916), .A2(n62447), .B(n77065), .C(
        n75872), .Y(n60882) );
  OAI22xp33_ASAP7_75t_SRAM U65156 ( .A1(n76729), .A2(n77638), .B1(
        or1200_cpu_or1200_mult_mac_n167), .B2(n64275), .Y(n61066) );
  OAI21xp33_ASAP7_75t_SRAM U65157 ( .A1(or1200_cpu_or1200_mult_mac_n231), .A2(
        n74587), .B(n77632), .Y(n61063) );
  O2A1O1Ixp5_ASAP7_75t_SL U65158 ( .A1(n64246), .A2(n64245), .B(n57126), .C(
        n64244), .Y(n64247) );
  AOI31xp33_ASAP7_75t_SL U65159 ( .A1(n64215), .A2(n64214), .A3(n64213), .B(
        n64212), .Y(n77664) );
  O2A1O1Ixp5_ASAP7_75t_SL U65160 ( .A1(n75334), .A2(n75333), .B(n75332), .C(
        n75331), .Y(n75344) );
  INVx1_ASAP7_75t_SL U65161 ( .A(n74582), .Y(n77035) );
  XNOR2xp5_ASAP7_75t_SL U65162 ( .A(n75361), .B(n75360), .Y(n75374) );
  O2A1O1Ixp5_ASAP7_75t_SL U65163 ( .A1(n59563), .A2(n59547), .B(n75852), .C(
        n75589), .Y(n75595) );
  NOR2xp33_ASAP7_75t_SL U65164 ( .A(n75886), .B(n75885), .Y(n77187) );
  AOI211xp5_ASAP7_75t_SL U65165 ( .A1(or1200_cpu_or1200_except_n544), .A2(
        n75884), .B(n76791), .C(n75883), .Y(n75885) );
  AOI22xp33_ASAP7_75t_SRAM U65166 ( .A1(n75854), .A2(n75853), .B1(n76345), 
        .B2(n75852), .Y(n75857) );
  NOR2xp33_ASAP7_75t_SL U65167 ( .A(n75830), .B(n75829), .Y(n77667) );
  OAI22xp33_ASAP7_75t_SRAM U65168 ( .A1(n1125), .A2(n75818), .B1(n1181), .B2(
        n75817), .Y(n75821) );
  O2A1O1Ixp5_ASAP7_75t_SL U65169 ( .A1(n59567), .A2(n64773), .B(n64772), .C(
        n75863), .Y(n64794) );
  AOI31xp33_ASAP7_75t_SL U65170 ( .A1(n62535), .A2(n62534), .A3(n62533), .B(
        n62532), .Y(n75833) );
  O2A1O1Ixp5_ASAP7_75t_SL U65171 ( .A1(n76627), .A2(n59712), .B(n59443), .C(
        n62356), .Y(n62358) );
  NOR2xp33_ASAP7_75t_SL U65172 ( .A(n70202), .B(n70204), .Y(n70203) );
  NOR2xp33_ASAP7_75t_SL U65173 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[7]), .Y(
        n70205) );
  NOR2xp33_ASAP7_75t_SL U65174 ( .A(n70144), .B(n70143), .Y(n70164) );
  XNOR2xp5_ASAP7_75t_SL U65175 ( .A(n70116), .B(n70126), .Y(n70130) );
  NOR2xp33_ASAP7_75t_SL U65176 ( .A(n70115), .B(n70123), .Y(n70126) );
  NOR2xp33_ASAP7_75t_SL U65177 ( .A(n70112), .B(n70111), .Y(n70115) );
  NOR2xp33_ASAP7_75t_SL U65178 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_21_), .B(n69420), .Y(
        n69421) );
  OAI21xp33_ASAP7_75t_SRAM U65179 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_8_), .A2(n69414), .B(
        n78345), .Y(n69415) );
  NOR4xp25_ASAP7_75t_SL U65180 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_9_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_7_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_3_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_5_), .Y(n69412) );
  NOR2xp33_ASAP7_75t_SL U65181 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_), .B(n78429), .Y(
        n69413) );
  XNOR2xp5_ASAP7_75t_SL U65182 ( .A(n70162), .B(n70163), .Y(n70144) );
  XNOR2xp5_ASAP7_75t_SL U65183 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[1]), .B(
        n70110), .Y(n70113) );
  NOR2xp33_ASAP7_75t_SL U65184 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_22_), .B(n69582), .Y(
        n69410) );
  NOR2xp33_ASAP7_75t_SL U65185 ( .A(n69404), .B(n69403), .Y(n69446) );
  NAND2xp33_ASAP7_75t_SRAM U65186 ( .A(n69392), .B(n69391), .Y(n69398) );
  INVxp33_ASAP7_75t_SRAM U65187 ( .A(n69390), .Y(n69391) );
  INVxp33_ASAP7_75t_SRAM U65188 ( .A(n69393), .Y(n69387) );
  INVxp33_ASAP7_75t_SRAM U65189 ( .A(n69394), .Y(n69389) );
  NOR2xp33_ASAP7_75t_SL U65190 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[5]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[3]), .Y(n69549)
         );
  NOR2xp33_ASAP7_75t_SL U65191 ( .A(n70119), .B(n70118), .Y(n70139) );
  NOR2xp33_ASAP7_75t_SL U65192 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_21_), .B(n69443), .Y(
        n69574) );
  NOR2xp33_ASAP7_75t_SL U65193 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[10]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[11]), .Y(n69536) );
  OAI21xp33_ASAP7_75t_SRAM U65194 ( .A1(n69535), .A2(n69534), .B(n69533), .Y(
        n69539) );
  XOR2xp5_ASAP7_75t_SL U65195 ( .A(n70147), .B(n70149), .Y(n70162) );
  XNOR2xp5_ASAP7_75t_SL U65196 ( .A(n70175), .B(n70176), .Y(n70180) );
  NOR2xp33_ASAP7_75t_SL U65197 ( .A(n70161), .B(n70173), .Y(n70176) );
  XNOR2xp5_ASAP7_75t_SL U65198 ( .A(n70145), .B(n70146), .Y(n70147) );
  NOR3xp33_ASAP7_75t_SL U65199 ( .A(n69439), .B(n69438), .C(n69437), .Y(n69445) );
  NOR2xp33_ASAP7_75t_SL U65200 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_20_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_22_), .Y(n69425) );
  XNOR2xp5_ASAP7_75t_SL U65201 ( .A(n70137), .B(n70153), .Y(n70146) );
  XNOR2xp5_ASAP7_75t_SL U65202 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[3]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[3]), .Y(
        n70137) );
  NOR2xp33_ASAP7_75t_SL U65203 ( .A(n69927), .B(n70080), .Y(n70135) );
  NOR2xp33_ASAP7_75t_SL U65204 ( .A(n69977), .B(n69903), .Y(n70080) );
  NOR2xp33_ASAP7_75t_SL U65205 ( .A(n69525), .B(n69977), .Y(n69927) );
  XNOR2xp5_ASAP7_75t_SL U65206 ( .A(n70186), .B(n70188), .Y(n70182) );
  NOR2xp33_ASAP7_75t_SL U65207 ( .A(n70165), .B(n70169), .Y(n70171) );
  NOR2xp33_ASAP7_75t_SL U65208 ( .A(n70174), .B(n70173), .Y(n70188) );
  NOR2xp33_ASAP7_75t_SL U65209 ( .A(n70160), .B(n70159), .Y(n70173) );
  XNOR2xp5_ASAP7_75t_SL U65210 ( .A(n70155), .B(n70166), .Y(n70160) );
  NOR2xp33_ASAP7_75t_SL U65211 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_29_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_28_), .Y(n69406) );
  NOR2xp33_ASAP7_75t_SL U65212 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_27_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_24_), .Y(n69407) );
  INVx1_ASAP7_75t_SL U65213 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_30_), .Y(n78382) );
  NOR2xp33_ASAP7_75t_SL U65214 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_), .Y(n69405) );
  XNOR2xp5_ASAP7_75t_SL U65215 ( .A(n70197), .B(n70194), .Y(n70196) );
  NAND3xp33_ASAP7_75t_SL U65216 ( .A(n78383), .B(n78370), .C(n69519), .Y(
        n69520) );
  NOR2xp33_ASAP7_75t_SL U65217 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_), .Y(n69519) );
  INVx1_ASAP7_75t_SL U65218 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_), 
        .Y(n78370) );
  NAND3xp33_ASAP7_75t_SL U65219 ( .A(n69518), .B(n78381), .C(n78372), .Y(
        n69521) );
  INVx1_ASAP7_75t_SL U65220 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_), 
        .Y(n78372) );
  INVx1_ASAP7_75t_SL U65221 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_27_), 
        .Y(n78381) );
  NOR2xp33_ASAP7_75t_SL U65222 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_29_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_), .Y(n69518) );
  NOR2xp33_ASAP7_75t_SL U65223 ( .A(n70190), .B(n70206), .Y(n70191) );
  INVxp33_ASAP7_75t_SRAM U65224 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_r_a), .Y(n65284) );
  XNOR2xp5_ASAP7_75t_SL U65225 ( .A(n71158), .B(n71276), .Y(n71159) );
  XNOR2xp5_ASAP7_75t_SL U65226 ( .A(n71170), .B(n71169), .Y(n71158) );
  NOR2xp33_ASAP7_75t_SL U65227 ( .A(n75181), .B(n77389), .Y(n75182) );
  NOR2xp33_ASAP7_75t_SL U65228 ( .A(n77390), .B(n77389), .Y(n77391) );
  XOR2xp5_ASAP7_75t_SL U65229 ( .A(n2037), .B(or1200_cpu_or1200_except_n667), 
        .Y(n77387) );
  NOR2xp33_ASAP7_75t_SL U65230 ( .A(n2071), .B(or1200_cpu_or1200_except_n652), 
        .Y(n65228) );
  NOR2xp33_ASAP7_75t_SL U65231 ( .A(n65227), .B(n65226), .Y(n65229) );
  XNOR2xp5_ASAP7_75t_SL U65232 ( .A(n2071), .B(or1200_cpu_or1200_except_n652), 
        .Y(n65226) );
  NOR2xp33_ASAP7_75t_SL U65233 ( .A(id_insn_22_), .B(n65218), .Y(n65227) );
  NOR2xp33_ASAP7_75t_SL U65234 ( .A(n2671), .B(or1200_cpu_or1200_except_n637), 
        .Y(n75415) );
  NOR2xp33_ASAP7_75t_SL U65235 ( .A(n2685), .B(or1200_cpu_or1200_except_n643), 
        .Y(n75541) );
  AOI211xp5_ASAP7_75t_SL U65236 ( .A1(n63963), .A2(n63980), .B(n63966), .C(
        n63965), .Y(n63976) );
  XNOR2xp5_ASAP7_75t_SL U65237 ( .A(n2623), .B(or1200_cpu_or1200_except_n616), 
        .Y(n63965) );
  NOR2xp33_ASAP7_75t_SL U65238 ( .A(or1200_cpu_or1200_except_n613), .B(n2098), 
        .Y(n63966) );
  NOR2xp33_ASAP7_75t_SL U65239 ( .A(n2110), .B(or1200_cpu_or1200_except_n610), 
        .Y(n63963) );
  AND2x2_ASAP7_75t_SL U65240 ( .A(or1200_cpu_or1200_except_n616), .B(n2623), 
        .Y(n63977) );
  NOR2xp33_ASAP7_75t_SL U65241 ( .A(n63761), .B(n63762), .Y(n63756) );
  NOR3xp33_ASAP7_75t_SL U65242 ( .A(n63762), .B(n76519), .C(n63760), .Y(n63757) );
  NOR2xp33_ASAP7_75t_SL U65243 ( .A(n2148), .B(or1200_cpu_or1200_except_n601), 
        .Y(n63760) );
  XNOR2xp5_ASAP7_75t_SL U65244 ( .A(n2134), .B(or1200_cpu_or1200_except_n604), 
        .Y(n76519) );
  XNOR2xp5_ASAP7_75t_SL U65245 ( .A(n2122), .B(or1200_cpu_or1200_except_n607), 
        .Y(n63762) );
  NOR2xp33_ASAP7_75t_SL U65246 ( .A(n76579), .B(n76578), .Y(n76577) );
  NOR2xp33_ASAP7_75t_SL U65247 ( .A(n3390), .B(or1200_cpu_or1200_except_n583), 
        .Y(n76579) );
  XNOR2xp5_ASAP7_75t_SL U65248 ( .A(n2172), .B(or1200_cpu_or1200_except_n595), 
        .Y(n76601) );
  AND2x2_ASAP7_75t_SL U65249 ( .A(or1200_cpu_or1200_except_n595), .B(n2172), 
        .Y(n58558) );
  XNOR2xp5_ASAP7_75t_SL U65250 ( .A(n2160), .B(or1200_cpu_or1200_except_n598), 
        .Y(n76814) );
  XOR2xp5_ASAP7_75t_SL U65251 ( .A(or1200_cpu_or1200_except_n601), .B(n2148), 
        .Y(n76841) );
  XNOR2xp5_ASAP7_75t_SL U65252 ( .A(n2110), .B(or1200_cpu_or1200_except_n610), 
        .Y(n76529) );
  AND2x2_ASAP7_75t_SL U65253 ( .A(n2630), .B(or1200_cpu_or1200_except_n619), 
        .Y(n63994) );
  XNOR2xp5_ASAP7_75t_SL U65254 ( .A(n2644), .B(or1200_cpu_or1200_except_n625), 
        .Y(n64003) );
  AND2x2_ASAP7_75t_SL U65255 ( .A(or1200_cpu_or1200_except_n625), .B(n2644), 
        .Y(n58592) );
  XNOR2xp5_ASAP7_75t_SL U65256 ( .A(n3392), .B(or1200_cpu_or1200_except_n628), 
        .Y(n64009) );
  AND2x2_ASAP7_75t_SL U65257 ( .A(n3392), .B(or1200_cpu_or1200_except_n628), 
        .Y(n58601) );
  XNOR2xp5_ASAP7_75t_SL U65258 ( .A(n2657), .B(or1200_cpu_or1200_except_n631), 
        .Y(n74967) );
  AND2x2_ASAP7_75t_SL U65259 ( .A(or1200_cpu_or1200_except_n631), .B(n2657), 
        .Y(n58604) );
  XOR2xp5_ASAP7_75t_SL U65260 ( .A(or1200_cpu_or1200_except_n634), .B(n2664), 
        .Y(n64163) );
  NOR2xp33_ASAP7_75t_SL U65261 ( .A(n65202), .B(n75543), .Y(n65204) );
  XNOR2xp5_ASAP7_75t_SL U65262 ( .A(n3117), .B(or1200_cpu_or1200_except_n646), 
        .Y(n75543) );
  XNOR2xp5_ASAP7_75t_SL U65263 ( .A(n2671), .B(or1200_cpu_or1200_except_n637), 
        .Y(n64265) );
  XNOR2xp5_ASAP7_75t_SL U65264 ( .A(n2054), .B(or1200_cpu_or1200_except_n655), 
        .Y(n75157) );
  O2A1O1Ixp5_ASAP7_75t_SL U65265 ( .A1(n65278), .A2(n65274), .B(n65273), .C(
        n65331), .Y(n2484) );
  NOR4xp25_ASAP7_75t_SL U65266 ( .A(n75504), .B(n75503), .C(n75502), .D(n75501), .Y(n75505) );
  NAND4xp25_ASAP7_75t_SL U65267 ( .A(or1200_cpu_or1200_mult_mac_n315), .B(
        or1200_cpu_or1200_mult_mac_n307), .C(or1200_cpu_or1200_mult_mac_n301), 
        .D(or1200_cpu_or1200_mult_mac_n333), .Y(n75501) );
  NAND4xp25_ASAP7_75t_SL U65268 ( .A(or1200_cpu_or1200_mult_mac_n309), .B(
        or1200_cpu_or1200_mult_mac_n289), .C(or1200_cpu_or1200_mult_mac_n291), 
        .D(or1200_cpu_or1200_mult_mac_n293), .Y(n75503) );
  NAND4xp25_ASAP7_75t_SL U65269 ( .A(or1200_cpu_or1200_mult_mac_n343), .B(
        or1200_cpu_or1200_mult_mac_n303), .C(or1200_cpu_or1200_mult_mac_n337), 
        .D(or1200_cpu_or1200_mult_mac_n341), .Y(n75504) );
  NOR4xp25_ASAP7_75t_SL U65270 ( .A(n75500), .B(n75499), .C(n75498), .D(n75497), .Y(n75506) );
  NAND4xp25_ASAP7_75t_SL U65271 ( .A(or1200_cpu_or1200_mult_mac_n317), .B(
        or1200_cpu_or1200_mult_mac_n321), .C(or1200_cpu_or1200_mult_mac_n347), 
        .D(or1200_cpu_or1200_mult_mac_n297), .Y(n75497) );
  NAND4xp25_ASAP7_75t_SL U65272 ( .A(or1200_cpu_or1200_mult_mac_n311), .B(
        or1200_cpu_or1200_mult_mac_n313), .C(or1200_cpu_or1200_mult_mac_n299), 
        .D(or1200_cpu_or1200_mult_mac_n305), .Y(n75498) );
  NAND4xp25_ASAP7_75t_SL U65273 ( .A(or1200_cpu_or1200_mult_mac_n323), .B(
        or1200_cpu_or1200_mult_mac_n319), .C(or1200_cpu_or1200_mult_mac_n325), 
        .D(or1200_cpu_or1200_mult_mac_n329), .Y(n75499) );
  NAND4xp25_ASAP7_75t_SL U65274 ( .A(or1200_cpu_or1200_mult_mac_n327), .B(
        or1200_cpu_or1200_mult_mac_n331), .C(or1200_cpu_or1200_mult_mac_n335), 
        .D(or1200_cpu_or1200_mult_mac_n339), .Y(n75500) );
  NOR4xp25_ASAP7_75t_SL U65275 ( .A(n75496), .B(n75495), .C(n75494), .D(n75493), .Y(n75513) );
  NAND4xp25_ASAP7_75t_SL U65276 ( .A(or1200_cpu_or1200_mult_mac_n353), .B(
        or1200_cpu_or1200_mult_mac_n351), .C(or1200_cpu_or1200_mult_mac_n357), 
        .D(or1200_cpu_or1200_mult_mac_n355), .Y(n75493) );
  NAND4xp25_ASAP7_75t_SL U65277 ( .A(or1200_cpu_or1200_mult_mac_n363), .B(
        or1200_cpu_or1200_mult_mac_n359), .C(or1200_cpu_or1200_mult_mac_n361), 
        .D(or1200_cpu_or1200_mult_mac_n365), .Y(n75494) );
  NAND4xp25_ASAP7_75t_SL U65278 ( .A(or1200_cpu_or1200_mult_mac_n371), .B(
        or1200_cpu_or1200_mult_mac_n367), .C(or1200_cpu_or1200_mult_mac_n369), 
        .D(or1200_cpu_or1200_mult_mac_n373), .Y(n75495) );
  NAND4xp25_ASAP7_75t_SL U65279 ( .A(or1200_cpu_or1200_mult_mac_n375), .B(
        or1200_cpu_or1200_mult_mac_n377), .C(or1200_cpu_or1200_mult_mac_n379), 
        .D(or1200_cpu_or1200_mult_mac_n385), .Y(n75496) );
  NOR4xp25_ASAP7_75t_SL U65280 ( .A(n75492), .B(n75491), .C(n75490), .D(n75489), .Y(n75514) );
  NAND4xp25_ASAP7_75t_SL U65281 ( .A(or1200_cpu_or1200_mult_mac_n395), .B(
        or1200_cpu_or1200_mult_mac_n409), .C(or1200_cpu_or1200_mult_mac_n411), 
        .D(or1200_cpu_or1200_mult_mac_n413), .Y(n75489) );
  NAND4xp25_ASAP7_75t_SL U65282 ( .A(or1200_cpu_or1200_mult_mac_n397), .B(
        or1200_cpu_or1200_mult_mac_n383), .C(or1200_cpu_or1200_mult_mac_n387), 
        .D(or1200_cpu_or1200_mult_mac_n391), .Y(n75490) );
  NAND4xp25_ASAP7_75t_SL U65283 ( .A(or1200_cpu_or1200_mult_mac_n407), .B(
        or1200_cpu_or1200_mult_mac_n381), .C(or1200_cpu_or1200_mult_mac_n393), 
        .D(or1200_cpu_or1200_mult_mac_n389), .Y(n75491) );
  NAND4xp25_ASAP7_75t_SL U65284 ( .A(or1200_cpu_or1200_mult_mac_n405), .B(
        or1200_cpu_or1200_mult_mac_n403), .C(or1200_cpu_or1200_mult_mac_n401), 
        .D(or1200_cpu_or1200_mult_mac_n399), .Y(n75492) );
  AND2x2_ASAP7_75t_SL U65285 ( .A(or1200_cpu_or1200_mult_mac_n265), .B(
        or1200_cpu_or1200_mult_mac_n411), .Y(n76900) );
  NOR2xp33_ASAP7_75t_SL U65286 ( .A(or1200_cpu_or1200_mult_mac_n265), .B(
        or1200_cpu_or1200_mult_mac_n411), .Y(n76896) );
  XOR2xp5_ASAP7_75t_SL U65287 ( .A(or1200_cpu_or1200_mult_mac_n413), .B(
        or1200_cpu_or1200_mult_mac_n267), .Y(n76911) );
  AOI211xp5_ASAP7_75t_SL U65288 ( .A1(or1200_cpu_rf_datab[21]), .A2(n57091), 
        .B(n77184), .C(n62140), .Y(n62141) );
  AOI211xp5_ASAP7_75t_SL U65289 ( .A1(n77128), .A2(n58557), .B(n62136), .C(
        n74626), .Y(n62137) );
  NOR2xp33_ASAP7_75t_SL U65290 ( .A(n75872), .B(n73915), .Y(n62135) );
  AOI211xp5_ASAP7_75t_SL U65291 ( .A1(n75727), .A2(n62116), .B(n62115), .C(
        n62114), .Y(n62117) );
  AOI22xp33_ASAP7_75t_SRAM U65292 ( .A1(or1200_cpu_or1200_fpu_result_arith[21]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[21]), .Y(
        n62113) );
  INVxp33_ASAP7_75t_SRAM U65293 ( .A(or1200_cpu_or1200_mult_mac_n86), .Y(
        n62116) );
  OAI21xp33_ASAP7_75t_SRAM U65294 ( .A1(n75433), .A2(n62104), .B(n77082), .Y(
        n62132) );
  INVxp33_ASAP7_75t_SRAM U65295 ( .A(n64107), .Y(n62104) );
  OAI22xp33_ASAP7_75t_SRAM U65296 ( .A1(n1139), .A2(n77033), .B1(n1444), .B2(
        n77034), .Y(n62097) );
  NOR2xp33_ASAP7_75t_SL U65297 ( .A(n64097), .B(n74595), .Y(n64321) );
  NOR2xp33_ASAP7_75t_SL U65298 ( .A(n63563), .B(n63562), .Y(n74596) );
  HB1xp67_ASAP7_75t_SL U65299 ( .A(n76903), .Y(n59673) );
  AND2x2_ASAP7_75t_SL U65300 ( .A(or1200_cpu_or1200_mult_mac_n263), .B(
        or1200_cpu_or1200_mult_mac_n409), .Y(n75663) );
  NOR2xp33_ASAP7_75t_SL U65301 ( .A(or1200_cpu_or1200_mult_mac_n263), .B(
        or1200_cpu_or1200_mult_mac_n409), .Y(n75659) );
  NOR2xp33_ASAP7_75t_SL U65302 ( .A(or1200_cpu_or1200_mult_mac_n261), .B(
        or1200_cpu_or1200_mult_mac_n407), .Y(n75660) );
  AND2x2_ASAP7_75t_SL U65303 ( .A(or1200_cpu_or1200_mult_mac_n257), .B(
        or1200_cpu_or1200_mult_mac_n403), .Y(n75121) );
  NOR2xp33_ASAP7_75t_SL U65304 ( .A(or1200_cpu_or1200_mult_mac_n253), .B(
        or1200_cpu_or1200_mult_mac_n399), .Y(n69311) );
  AO21x1_ASAP7_75t_SL U65305 ( .A1(n69292), .A2(n69291), .B(n69290), .Y(n69313) );
  NOR2xp33_ASAP7_75t_SL U65306 ( .A(or1200_cpu_or1200_mult_mac_n251), .B(
        or1200_cpu_or1200_mult_mac_n397), .Y(n69290) );
  NOR2xp33_ASAP7_75t_SL U65307 ( .A(n69243), .B(n69242), .Y(n69258) );
  NOR2xp33_ASAP7_75t_SL U65308 ( .A(or1200_cpu_or1200_mult_mac_n245), .B(
        or1200_cpu_or1200_mult_mac_n391), .Y(n69242) );
  NOR2xp33_ASAP7_75t_SL U65309 ( .A(or1200_cpu_or1200_mult_mac_n241), .B(
        or1200_cpu_or1200_mult_mac_n387), .Y(n74570) );
  NOR2xp33_ASAP7_75t_SL U65310 ( .A(n75293), .B(n69187), .Y(n69207) );
  NOR2xp33_ASAP7_75t_SL U65311 ( .A(n75292), .B(n75294), .Y(n69187) );
  NOR2xp33_ASAP7_75t_SL U65312 ( .A(or1200_cpu_or1200_mult_mac_n239), .B(
        or1200_cpu_or1200_mult_mac_n385), .Y(n75294) );
  NOR2xp33_ASAP7_75t_SL U65313 ( .A(or1200_cpu_or1200_mult_mac_n237), .B(
        or1200_cpu_or1200_mult_mac_n383), .Y(n75292) );
  NOR2xp33_ASAP7_75t_SL U65314 ( .A(or1200_cpu_or1200_mult_mac_n233), .B(
        or1200_cpu_or1200_mult_mac_n379), .Y(n69277) );
  NOR2xp33_ASAP7_75t_SL U65315 ( .A(or1200_cpu_or1200_mult_mac_n235), .B(
        or1200_cpu_or1200_mult_mac_n381), .Y(n69278) );
  AND2x2_ASAP7_75t_SL U65316 ( .A(or1200_cpu_or1200_mult_mac_n227), .B(
        or1200_cpu_or1200_mult_mac_n373), .Y(n69106) );
  NOR2xp33_ASAP7_75t_SL U65317 ( .A(or1200_cpu_or1200_mult_mac_n225), .B(
        or1200_cpu_or1200_mult_mac_n371), .Y(n69089) );
  NOR2xp33_ASAP7_75t_SL U65318 ( .A(or1200_cpu_or1200_mult_mac_n227), .B(
        or1200_cpu_or1200_mult_mac_n373), .Y(n69090) );
  NOR2xp33_ASAP7_75t_SL U65319 ( .A(or1200_cpu_or1200_mult_mac_n223), .B(
        or1200_cpu_or1200_mult_mac_n369), .Y(n69088) );
  AND2x2_ASAP7_75t_SL U65320 ( .A(or1200_cpu_or1200_mult_mac_n219), .B(
        or1200_cpu_or1200_mult_mac_n365), .Y(n68997) );
  NOR2xp33_ASAP7_75t_SL U65321 ( .A(or1200_cpu_or1200_mult_mac_n217), .B(
        or1200_cpu_or1200_mult_mac_n363), .Y(n68995) );
  NOR2xp33_ASAP7_75t_SL U65322 ( .A(or1200_cpu_or1200_mult_mac_n219), .B(
        or1200_cpu_or1200_mult_mac_n365), .Y(n68996) );
  NOR2xp33_ASAP7_75t_SL U65323 ( .A(or1200_cpu_or1200_mult_mac_n215), .B(
        or1200_cpu_or1200_mult_mac_n361), .Y(n68994) );
  AND2x2_ASAP7_75t_SL U65324 ( .A(or1200_cpu_or1200_mult_mac_n209), .B(
        or1200_cpu_or1200_mult_mac_n355), .Y(n68882) );
  NOR2xp33_ASAP7_75t_SL U65325 ( .A(or1200_cpu_or1200_mult_mac_n205), .B(
        or1200_cpu_or1200_mult_mac_n351), .Y(n68845) );
  NOR2xp33_ASAP7_75t_SL U65326 ( .A(n76885), .B(n68880), .Y(n68890) );
  AND2x2_ASAP7_75t_SL U65327 ( .A(or1200_cpu_or1200_mult_mac_n203), .B(
        or1200_cpu_or1200_mult_mac_n349), .Y(n76885) );
  NOR2xp33_ASAP7_75t_SL U65328 ( .A(or1200_cpu_or1200_mult_mac_n343), .B(
        or1200_cpu_or1200_mult_mac_n197), .Y(n75009) );
  NOR2xp33_ASAP7_75t_SL U65329 ( .A(or1200_cpu_or1200_mult_mac_n345), .B(
        or1200_cpu_or1200_mult_mac_n199), .Y(n75006) );
  NOR2xp33_ASAP7_75t_SL U65330 ( .A(n68780), .B(n68779), .Y(n68781) );
  XNOR2xp5_ASAP7_75t_SL U65331 ( .A(or1200_cpu_or1200_mult_mac_n341), .B(
        or1200_cpu_or1200_mult_mac_n195), .Y(n68779) );
  AND2x2_ASAP7_75t_SL U65332 ( .A(or1200_cpu_or1200_mult_mac_n193), .B(
        or1200_cpu_or1200_mult_mac_n339), .Y(n68780) );
  AOI211xp5_ASAP7_75t_SL U65333 ( .A1(n65174), .A2(n65173), .B(n65172), .C(
        n65171), .Y(n65178) );
  NOR2xp33_ASAP7_75t_SL U65334 ( .A(or1200_cpu_or1200_mult_mac_n335), .B(
        or1200_cpu_or1200_mult_mac_n189), .Y(n65171) );
  NOR2xp33_ASAP7_75t_SL U65335 ( .A(or1200_cpu_or1200_mult_mac_n333), .B(
        or1200_cpu_or1200_mult_mac_n187), .Y(n65172) );
  NOR2xp33_ASAP7_75t_SL U65336 ( .A(or1200_cpu_or1200_mult_mac_n327), .B(
        or1200_cpu_or1200_mult_mac_n181), .Y(n65128) );
  NOR2xp33_ASAP7_75t_SL U65337 ( .A(or1200_cpu_or1200_mult_mac_n329), .B(
        or1200_cpu_or1200_mult_mac_n183), .Y(n65129) );
  AOI31xp33_ASAP7_75t_SL U65338 ( .A1(n65089), .A2(n65088), .A3(n65087), .B(
        n65086), .Y(n65179) );
  NOR2xp33_ASAP7_75t_SL U65339 ( .A(or1200_cpu_or1200_mult_mac_n319), .B(
        or1200_cpu_or1200_mult_mac_n173), .Y(n63888) );
  NOR2xp33_ASAP7_75t_SL U65340 ( .A(n63487), .B(n63486), .Y(n63533) );
  NOR2xp33_ASAP7_75t_SL U65341 ( .A(or1200_cpu_or1200_mult_mac_n311), .B(
        or1200_cpu_or1200_mult_mac_n165), .Y(n63486) );
  NOR2xp33_ASAP7_75t_SL U65342 ( .A(or1200_cpu_or1200_mult_mac_n309), .B(
        or1200_cpu_or1200_mult_mac_n163), .Y(n63487) );
  NOR2xp33_ASAP7_75t_SL U65343 ( .A(n63432), .B(n63431), .Y(n63460) );
  NOR2xp33_ASAP7_75t_SL U65344 ( .A(or1200_cpu_or1200_mult_mac_n303), .B(
        or1200_cpu_or1200_mult_mac_n157), .Y(n63431) );
  NOR2xp33_ASAP7_75t_SL U65345 ( .A(or1200_cpu_or1200_mult_mac_n301), .B(
        or1200_cpu_or1200_mult_mac_n155), .Y(n63432) );
  NOR2xp33_ASAP7_75t_SL U65346 ( .A(n63372), .B(n63371), .Y(n63378) );
  NOR2xp33_ASAP7_75t_SL U65347 ( .A(or1200_cpu_or1200_mult_mac_n299), .B(
        or1200_cpu_or1200_mult_mac_n153), .Y(n63371) );
  NOR2xp33_ASAP7_75t_SL U65348 ( .A(or1200_cpu_or1200_mult_mac_n297), .B(
        or1200_cpu_or1200_mult_mac_n151), .Y(n63372) );
  NOR2xp33_ASAP7_75t_SL U65349 ( .A(n63338), .B(n63337), .Y(n63373) );
  NOR2xp33_ASAP7_75t_SL U65350 ( .A(or1200_cpu_or1200_mult_mac_n293), .B(
        or1200_cpu_or1200_mult_mac_n147), .Y(n63337) );
  NOR2xp33_ASAP7_75t_SL U65351 ( .A(or1200_cpu_or1200_mult_mac_n295), .B(
        or1200_cpu_or1200_mult_mac_n149), .Y(n63338) );
  NOR2xp33_ASAP7_75t_SL U65352 ( .A(or1200_cpu_or1200_mult_mac_n287), .B(
        or1200_cpu_or1200_mult_mac_n141), .Y(n63275) );
  AOI211xp5_ASAP7_75t_SL U65353 ( .A1(n63459), .A2(n63458), .B(n63457), .C(
        n63522), .Y(n65088) );
  AND2x2_ASAP7_75t_SL U65354 ( .A(or1200_cpu_or1200_mult_mac_n307), .B(
        or1200_cpu_or1200_mult_mac_n161), .Y(n63457) );
  NOR2xp33_ASAP7_75t_SL U65355 ( .A(n63456), .B(n63455), .Y(n63459) );
  NOR2xp33_ASAP7_75t_SL U65356 ( .A(or1200_cpu_or1200_mult_mac_n305), .B(
        or1200_cpu_or1200_mult_mac_n159), .Y(n63455) );
  NOR2xp33_ASAP7_75t_SL U65357 ( .A(or1200_cpu_or1200_mult_mac_n307), .B(
        or1200_cpu_or1200_mult_mac_n161), .Y(n63456) );
  NOR2xp33_ASAP7_75t_SL U65358 ( .A(or1200_cpu_or1200_mult_mac_n315), .B(
        or1200_cpu_or1200_mult_mac_n169), .Y(n63511) );
  NOR2xp33_ASAP7_75t_SL U65359 ( .A(or1200_cpu_or1200_mult_mac_n313), .B(
        or1200_cpu_or1200_mult_mac_n167), .Y(n63512) );
  NOR2xp33_ASAP7_75t_SL U65360 ( .A(n65076), .B(n65075), .Y(n65083) );
  NOR2xp33_ASAP7_75t_SL U65361 ( .A(or1200_cpu_or1200_mult_mac_n325), .B(
        or1200_cpu_or1200_mult_mac_n179), .Y(n65075) );
  NOR2xp33_ASAP7_75t_SL U65362 ( .A(or1200_cpu_or1200_mult_mac_n323), .B(
        or1200_cpu_or1200_mult_mac_n177), .Y(n65076) );
  NOR2xp33_ASAP7_75t_SL U65363 ( .A(or1200_cpu_or1200_mult_mac_n321), .B(
        or1200_cpu_or1200_mult_mac_n175), .Y(n63887) );
  NOR2xp33_ASAP7_75t_SL U65364 ( .A(n65132), .B(n65131), .Y(n65147) );
  NOR2xp33_ASAP7_75t_SL U65365 ( .A(or1200_cpu_or1200_mult_mac_n331), .B(
        or1200_cpu_or1200_mult_mac_n185), .Y(n65132) );
  XNOR2xp5_ASAP7_75t_SL U65366 ( .A(or1200_cpu_or1200_mult_mac_n343), .B(
        or1200_cpu_or1200_mult_mac_n197), .Y(n68820) );
  AND2x2_ASAP7_75t_SL U65367 ( .A(or1200_cpu_or1200_mult_mac_n233), .B(
        or1200_cpu_or1200_mult_mac_n379), .Y(n69282) );
  NOR2xp33_ASAP7_75t_SL U65368 ( .A(n58612), .B(n69244), .Y(n69284) );
  AND2x2_ASAP7_75t_SL U65369 ( .A(or1200_cpu_or1200_mult_mac_n245), .B(
        or1200_cpu_or1200_mult_mac_n391), .Y(n69244) );
  AND2x2_ASAP7_75t_SL U65370 ( .A(or1200_cpu_or1200_mult_mac_n247), .B(
        or1200_cpu_or1200_mult_mac_n393), .Y(n58612) );
  NAND4xp25_ASAP7_75t_SL U65371 ( .A(n69211), .B(n74571), .C(n69210), .D(
        n69209), .Y(n69279) );
  NOR2xp33_ASAP7_75t_SL U65372 ( .A(n75293), .B(n75290), .Y(n69211) );
  AND2x2_ASAP7_75t_SL U65373 ( .A(or1200_cpu_or1200_mult_mac_n237), .B(
        or1200_cpu_or1200_mult_mac_n383), .Y(n75290) );
  AND2x2_ASAP7_75t_SL U65374 ( .A(or1200_cpu_or1200_mult_mac_n239), .B(
        or1200_cpu_or1200_mult_mac_n385), .Y(n75293) );
  NOR2xp33_ASAP7_75t_SL U65375 ( .A(n69274), .B(n69273), .Y(n69292) );
  AND2x2_ASAP7_75t_SL U65376 ( .A(or1200_cpu_or1200_mult_mac_n249), .B(
        or1200_cpu_or1200_mult_mac_n395), .Y(n69273) );
  AND2x2_ASAP7_75t_SL U65377 ( .A(or1200_cpu_or1200_mult_mac_n251), .B(
        or1200_cpu_or1200_mult_mac_n397), .Y(n69274) );
  AND2x2_ASAP7_75t_SL U65378 ( .A(or1200_cpu_or1200_mult_mac_n255), .B(
        or1200_cpu_or1200_mult_mac_n401), .Y(n58617) );
  NOR2xp33_ASAP7_75t_SL U65379 ( .A(or1200_cpu_or1200_mult_mac_n259), .B(
        or1200_cpu_or1200_mult_mac_n405), .Y(n75662) );
  NOR2xp33_ASAP7_75t_SL U65380 ( .A(or1200_cpu_or1200_mult_mac_n253), .B(
        n69309), .Y(n69323) );
  NOR2xp33_ASAP7_75t_SL U65381 ( .A(n69246), .B(n69245), .Y(n69251) );
  NOR2xp33_ASAP7_75t_SL U65382 ( .A(or1200_cpu_or1200_mult_mac_n391), .B(
        n74114), .Y(n69245) );
  NOR2xp33_ASAP7_75t_SL U65383 ( .A(or1200_cpu_or1200_mult_mac_n389), .B(
        n74573), .Y(n69246) );
  NOR2xp33_ASAP7_75t_SL U65384 ( .A(n69171), .B(n69170), .Y(n69177) );
  NOR2xp33_ASAP7_75t_SL U65385 ( .A(n69172), .B(n69164), .Y(n69176) );
  NOR2xp33_ASAP7_75t_SL U65386 ( .A(or1200_cpu_or1200_mult_mac_n377), .B(
        n69126), .Y(n69164) );
  NOR2xp33_ASAP7_75t_SL U65387 ( .A(or1200_cpu_or1200_mult_mac_n381), .B(
        n77042), .Y(n69172) );
  NAND4xp25_ASAP7_75t_SL U65388 ( .A(n69068), .B(n69067), .C(n69066), .D(
        n69065), .Y(n69069) );
  AOI31xp33_ASAP7_75t_SL U65389 ( .A1(n68795), .A2(n68794), .A3(n68793), .B(
        n68792), .Y(n74998) );
  NOR2xp33_ASAP7_75t_SL U65390 ( .A(or1200_cpu_or1200_mult_mac_n327), .B(
        n65079), .Y(n65094) );
  NOR2xp33_ASAP7_75t_SL U65391 ( .A(n64170), .B(n64169), .Y(n65098) );
  NOR2xp33_ASAP7_75t_SL U65392 ( .A(or1200_cpu_or1200_mult_mac_n325), .B(
        n74584), .Y(n64169) );
  NOR2xp33_ASAP7_75t_SL U65393 ( .A(or1200_cpu_or1200_mult_mac_n323), .B(
        n63892), .Y(n64170) );
  NOR2xp33_ASAP7_75t_SL U65394 ( .A(or1200_cpu_or1200_mult_mac_n305), .B(
        n63410), .Y(n63425) );
  NOR2xp33_ASAP7_75t_SL U65395 ( .A(or1200_cpu_or1200_mult_mac_n317), .B(
        n77038), .Y(n63523) );
  XNOR2xp5_ASAP7_75t_SL U65396 ( .A(or1200_cpu_or1200_mult_mac_n309), .B(
        or1200_cpu_or1200_mult_mac_n163), .Y(n63522) );
  NOR2xp33_ASAP7_75t_SL U65397 ( .A(n63518), .B(n63517), .Y(n63527) );
  NOR2xp33_ASAP7_75t_SL U65398 ( .A(or1200_cpu_or1200_mult_mac_n301), .B(
        n76722), .Y(n63400) );
  AOI211xp5_ASAP7_75t_SL U65399 ( .A1(n63397), .A2(n63396), .B(n63395), .C(
        n63394), .Y(n63402) );
  NOR2xp33_ASAP7_75t_SL U65400 ( .A(or1200_cpu_or1200_mult_mac_n155), .B(
        n76754), .Y(n63395) );
  XNOR2xp5_ASAP7_75t_SL U65401 ( .A(or1200_cpu_or1200_mult_mac_n289), .B(
        or1200_cpu_or1200_mult_mac_n143), .Y(n63273) );
  NOR2xp33_ASAP7_75t_SL U65402 ( .A(n63305), .B(n63388), .Y(n63387) );
  NOR2xp33_ASAP7_75t_SL U65403 ( .A(n63304), .B(n63303), .Y(n63388) );
  XNOR2xp5_ASAP7_75t_SL U65404 ( .A(or1200_cpu_or1200_mult_mac_n291), .B(
        or1200_cpu_or1200_mult_mac_n145), .Y(n63303) );
  XOR2xp5_ASAP7_75t_SL U65405 ( .A(or1200_cpu_or1200_mult_mac_n293), .B(
        or1200_cpu_or1200_mult_mac_n147), .Y(n63305) );
  NOR2xp33_ASAP7_75t_SL U65406 ( .A(n63385), .B(n63384), .Y(n63398) );
  NOR2xp33_ASAP7_75t_SL U65407 ( .A(n63322), .B(n63321), .Y(n63323) );
  NOR2xp33_ASAP7_75t_SL U65408 ( .A(or1200_cpu_or1200_mult_mac_n297), .B(
        n63314), .Y(n63321) );
  NOR2xp33_ASAP7_75t_SL U65409 ( .A(or1200_cpu_or1200_mult_mac_n295), .B(
        n63325), .Y(n63322) );
  NOR2xp33_ASAP7_75t_SL U65410 ( .A(n63424), .B(n63423), .Y(n63427) );
  NOR2xp33_ASAP7_75t_SL U65411 ( .A(or1200_cpu_or1200_mult_mac_n157), .B(
        n63411), .Y(n63424) );
  AOI211xp5_ASAP7_75t_SL U65412 ( .A1(n69059), .A2(n69058), .B(n69057), .C(
        n69056), .Y(n69067) );
  NOR2xp33_ASAP7_75t_SL U65413 ( .A(or1200_cpu_or1200_mult_mac_n221), .B(
        n68985), .Y(n69056) );
  NOR2xp33_ASAP7_75t_SL U65414 ( .A(or1200_cpu_or1200_mult_mac_n223), .B(
        n69022), .Y(n69057) );
  NOR2xp33_ASAP7_75t_SL U65415 ( .A(n68988), .B(n68987), .Y(n68991) );
  NOR2xp33_ASAP7_75t_SL U65416 ( .A(or1200_cpu_or1200_mult_mac_n217), .B(
        n68938), .Y(n68988) );
  NOR2xp33_ASAP7_75t_SL U65417 ( .A(n68873), .B(n68872), .Y(n68875) );
  NOR2xp33_ASAP7_75t_SL U65418 ( .A(or1200_cpu_or1200_mult_mac_n205), .B(
        n68830), .Y(n68841) );
  NOR2xp33_ASAP7_75t_SL U65419 ( .A(or1200_cpu_or1200_mult_mac_n207), .B(
        n68847), .Y(n68842) );
  NOR2xp33_ASAP7_75t_SL U65420 ( .A(n69052), .B(n68941), .Y(n68943) );
  NOR2xp33_ASAP7_75t_SL U65421 ( .A(or1200_cpu_or1200_mult_mac_n359), .B(
        n68892), .Y(n68941) );
  NOR2xp33_ASAP7_75t_SL U65422 ( .A(or1200_cpu_or1200_mult_mac_n355), .B(
        n68849), .Y(n68877) );
  NOR2xp33_ASAP7_75t_SL U65423 ( .A(or1200_cpu_or1200_mult_mac_n361), .B(
        n68932), .Y(n69052) );
  NOR2xp33_ASAP7_75t_SL U65424 ( .A(or1200_cpu_or1200_mult_mac_n357), .B(
        n68864), .Y(n68874) );
  NOR2xp33_ASAP7_75t_SL U65425 ( .A(or1200_cpu_or1200_mult_mac_n373), .B(
        n69084), .Y(n69086) );
  NOR2xp33_ASAP7_75t_SL U65426 ( .A(n69200), .B(n69199), .Y(n69204) );
  NOR2xp33_ASAP7_75t_SL U65427 ( .A(or1200_cpu_or1200_mult_mac_n385), .B(
        n75363), .Y(n69199) );
  NOR2xp33_ASAP7_75t_SL U65428 ( .A(or1200_cpu_or1200_mult_mac_n395), .B(
        n69256), .Y(n69255) );
  NOR2xp33_ASAP7_75t_SL U65429 ( .A(or1200_cpu_or1200_mult_mac_n251), .B(
        n69270), .Y(n69272) );
  NOR2xp33_ASAP7_75t_SL U65430 ( .A(or1200_cpu_or1200_mult_mac_n401), .B(
        n69324), .Y(n75127) );
  XNOR2xp5_ASAP7_75t_SL U65431 ( .A(or1200_cpu_or1200_mult_mac_n261), .B(
        or1200_cpu_or1200_mult_mac_n407), .Y(n75652) );
  INVx1_ASAP7_75t_SL U65432 ( .A(n65398), .Y(n65402) );
  O2A1O1Ixp5_ASAP7_75t_SL U65433 ( .A1(n75866), .A2(n75575), .B(n61891), .C(
        n73925), .Y(n61893) );
  INVxp33_ASAP7_75t_SRAM U65434 ( .A(or1200_cpu_or1200_mult_mac_n66), .Y(
        n61865) );
  AOI31xp33_ASAP7_75t_SL U65435 ( .A1(n61851), .A2(n61850), .A3(n61849), .B(
        n61848), .Y(n77676) );
  O2A1O1Ixp5_ASAP7_75t_SL U65436 ( .A1(n74270), .A2(n74269), .B(n74268), .C(
        n74267), .Y(n2876) );
  O2A1O1Ixp5_ASAP7_75t_SL U65437 ( .A1(n70099), .A2(n70501), .B(n70101), .C(
        n58553), .Y(n70100) );
  INVx3_ASAP7_75t_SL U65438 ( .A(n59695), .Y(n59689) );
  AND2x2_ASAP7_75t_SL U65439 ( .A(n73589), .B(n3275), .Y(n73616) );
  NOR2xp33_ASAP7_75t_SL U65440 ( .A(n73572), .B(n73559), .Y(n73585) );
  NOR2xp33_ASAP7_75t_SL U65441 ( .A(n73558), .B(n73658), .Y(n73559) );
  NOR2xp33_ASAP7_75t_SL U65442 ( .A(n73659), .B(n73656), .Y(n73573) );
  NOR2xp33_ASAP7_75t_SL U65443 ( .A(n73549), .B(n73548), .Y(n73583) );
  AO21x1_ASAP7_75t_SL U65444 ( .A1(n73542), .A2(n73569), .B(n73541), .Y(n73577) );
  NOR2xp33_ASAP7_75t_SL U65445 ( .A(n73551), .B(n73550), .Y(n73548) );
  NOR2xp33_ASAP7_75t_SL U65446 ( .A(n73535), .B(n73593), .Y(n73537) );
  NOR2xp33_ASAP7_75t_SL U65447 ( .A(n73595), .B(n73594), .Y(n73593) );
  NOR2xp33_ASAP7_75t_SL U65448 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[2]), .B(n73534), 
        .Y(n73535) );
  INVxp33_ASAP7_75t_SRAM U65449 ( .A(n73521), .Y(n73527) );
  NOR2xp33_ASAP7_75t_SL U65450 ( .A(n73541), .B(n73540), .Y(n73570) );
  NOR2xp33_ASAP7_75t_SL U65451 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[0]), .B(n73606), 
        .Y(n73540) );
  NOR2xp33_ASAP7_75t_SL U65452 ( .A(n73536), .B(n73505), .Y(n73569) );
  NOR2xp33_ASAP7_75t_SL U65453 ( .A(n73601), .B(n73504), .Y(n73536) );
  NOR2xp33_ASAP7_75t_SL U65454 ( .A(n73613), .B(n73591), .Y(n73555) );
  NOR2xp33_ASAP7_75t_SL U65455 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[5]), .B(n73554), 
        .Y(n73571) );
  NOR2xp33_ASAP7_75t_SL U65456 ( .A(n70943), .B(n70948), .Y(n70944) );
  NOR2xp33_ASAP7_75t_SL U65457 ( .A(n75266), .B(n75270), .Y(n77860) );
  O2A1O1Ixp5_ASAP7_75t_SL U65458 ( .A1(n76755), .A2(n75256), .B(n75255), .C(
        n75872), .Y(n75257) );
  NOR4xp25_ASAP7_75t_SL U65459 ( .A(n62108), .B(n62107), .C(n62106), .D(n62105), .Y(n75350) );
  O2A1O1Ixp5_ASAP7_75t_SL U65460 ( .A1(n75866), .A2(n75244), .B(n75243), .C(
        n75863), .Y(n75253) );
  NOR4xp25_ASAP7_75t_SL U65461 ( .A(n61105), .B(n61496), .C(n61104), .D(n61510), .Y(n75330) );
  NOR4xp25_ASAP7_75t_SL U65462 ( .A(n61098), .B(n61509), .C(n61097), .D(n61506), .Y(n75324) );
  NOR4xp25_ASAP7_75t_SL U65463 ( .A(n61505), .B(n61096), .C(n61095), .D(n61094), .Y(n75327) );
  O2A1O1Ixp5_ASAP7_75t_SL U65464 ( .A1(n75236), .A2(n75235), .B(n75591), .C(
        n75234), .Y(n75237) );
  O2A1O1Ixp5_ASAP7_75t_SL U65465 ( .A1(n59575), .A2(n75227), .B(n76775), .C(
        n59549), .Y(n75228) );
  O2A1O1Ixp5_ASAP7_75t_SL U65466 ( .A1(n75223), .A2(n75222), .B(n75751), .C(
        n75221), .Y(n75256) );
  INVxp33_ASAP7_75t_SRAM U65467 ( .A(n63444), .Y(n63450) );
  NOR2xp33_ASAP7_75t_SL U65468 ( .A(n61058), .B(n61056), .Y(n60729) );
  NOR2xp33_ASAP7_75t_SL U65469 ( .A(n61012), .B(n61011), .Y(n61013) );
  NOR2xp33_ASAP7_75t_SL U65470 ( .A(n60718), .B(n60505), .Y(n61315) );
  NOR2xp33_ASAP7_75t_SL U65471 ( .A(n62020), .B(n60504), .Y(n61310) );
  NOR3xp33_ASAP7_75t_SL U65472 ( .A(n61009), .B(n61012), .C(n61010), .Y(n77185) );
  NOR3xp33_ASAP7_75t_SL U65473 ( .A(n61008), .B(n61007), .C(n61006), .Y(n61010) );
  XOR2xp5_ASAP7_75t_SL U65474 ( .A(n2623), .B(n2572), .Y(n61006) );
  XOR2xp5_ASAP7_75t_SL U65475 ( .A(n3392), .B(n2023), .Y(n61007) );
  NAND4xp25_ASAP7_75t_SL U65476 ( .A(n61005), .B(n61004), .C(n61003), .D(
        n61002), .Y(n61008) );
  NOR2xp33_ASAP7_75t_SL U65477 ( .A(n2188), .B(n61125), .Y(n61002) );
  XNOR2xp5_ASAP7_75t_SL U65478 ( .A(n2644), .B(n2042), .Y(n61003) );
  XNOR2xp5_ASAP7_75t_SL U65479 ( .A(n2630), .B(n2076), .Y(n61004) );
  XNOR2xp5_ASAP7_75t_SL U65480 ( .A(n2637), .B(n2059), .Y(n61005) );
  NOR2xp33_ASAP7_75t_SL U65481 ( .A(or1200_cpu_or1200_mult_mac_n112), .B(
        n61826), .Y(n62350) );
  NOR2xp33_ASAP7_75t_SL U65482 ( .A(or1200_cpu_or1200_mult_mac_n114), .B(
        n61826), .Y(n62347) );
  NOR2xp33_ASAP7_75t_SL U65483 ( .A(n60809), .B(n60808), .Y(n62289) );
  NOR3xp33_ASAP7_75t_SL U65484 ( .A(n61825), .B(n64316), .C(n75361), .Y(n61836) );
  O2A1O1Ixp5_ASAP7_75t_SL U65485 ( .A1(n75742), .A2(n75741), .B(n75740), .C(
        n75739), .Y(n75743) );
  O2A1O1Ixp5_ASAP7_75t_SL U65486 ( .A1(n75733), .A2(n75732), .B(n75731), .C(
        n75730), .Y(n75744) );
  NOR2xp33_ASAP7_75t_SL U65487 ( .A(n63267), .B(n61858), .Y(n75847) );
  INVxp33_ASAP7_75t_SRAM U65488 ( .A(or1200_cpu_or1200_mult_mac_n68), .Y(
        n75726) );
  NOR2xp33_ASAP7_75t_SL U65489 ( .A(n75707), .B(n60858), .Y(n75729) );
  O2A1O1Ixp5_ASAP7_75t_SL U65490 ( .A1(n59528), .A2(n59645), .B(n75703), .C(
        n75702), .Y(n75704) );
  AOI31xp33_ASAP7_75t_SL U65491 ( .A1(n60863), .A2(n58589), .A3(n61191), .B(
        n60862), .Y(n75705) );
  NOR2xp33_ASAP7_75t_SL U65492 ( .A(n77726), .B(n62134), .Y(n75214) );
  NAND4xp25_ASAP7_75t_SL U65493 ( .A(n60881), .B(n60880), .C(n60879), .D(
        n60878), .Y(n77124) );
  NOR2xp33_ASAP7_75t_SL U65494 ( .A(n2607), .B(n61852), .Y(n61853) );
  NOR2xp33_ASAP7_75t_SL U65495 ( .A(n77060), .B(n62133), .Y(n73915) );
  NOR2xp33_ASAP7_75t_SL U65496 ( .A(n60825), .B(n60824), .Y(n61156) );
  NAND4xp25_ASAP7_75t_SL U65497 ( .A(n2542), .B(ex_insn[16]), .C(n2614), .D(
        n2819), .Y(n60824) );
  NAND3xp33_ASAP7_75t_SL U65498 ( .A(ex_insn[28]), .B(ex_insn[26]), .C(n2594), 
        .Y(n60825) );
  NAND3xp33_ASAP7_75t_SL U65499 ( .A(n77080), .B(n77021), .C(n77153), .Y(
        n77081) );
  NOR2xp33_ASAP7_75t_SL U65500 ( .A(or1200_cpu_or1200_except_n502), .B(n76792), 
        .Y(n76795) );
  NOR2xp33_ASAP7_75t_SL U65501 ( .A(or1200_cpu_or1200_except_n498), .B(n61651), 
        .Y(n62263) );
  NOR2xp33_ASAP7_75t_SL U65502 ( .A(or1200_cpu_or1200_except_n526), .B(
        or1200_cpu_or1200_except_n528), .Y(n61838) );
  NOR2xp33_ASAP7_75t_SL U65503 ( .A(n60841), .B(n58607), .Y(n77082) );
  OR2x2_ASAP7_75t_SL U65504 ( .A(n61001), .B(n61009), .Y(n77137) );
  INVx2_ASAP7_75t_SL U65505 ( .A(n59695), .Y(n59692) );
  NOR2xp33_ASAP7_75t_SL U65506 ( .A(n61000), .B(n60999), .Y(n61012) );
  NAND4xp25_ASAP7_75t_SL U65507 ( .A(n60998), .B(n60997), .C(n60996), .D(
        n60995), .Y(n60999) );
  XNOR2xp5_ASAP7_75t_SL U65508 ( .A(n2644), .B(n2045), .Y(n60996) );
  XNOR2xp5_ASAP7_75t_SL U65509 ( .A(n2637), .B(n2062), .Y(n60997) );
  XNOR2xp5_ASAP7_75t_SL U65510 ( .A(n2623), .B(n2575), .Y(n60998) );
  XNOR2xp5_ASAP7_75t_SL U65511 ( .A(n2630), .B(n2079), .Y(n60993) );
  XNOR2xp5_ASAP7_75t_SL U65512 ( .A(n3392), .B(n2026), .Y(n60994) );
  O2A1O1Ixp5_ASAP7_75t_SL U65513 ( .A1(n60288), .A2(n60287), .B(n60286), .C(
        n77352), .Y(n60289) );
  NOR2xp33_ASAP7_75t_SL U65514 ( .A(n60501), .B(n60500), .Y(n62020) );
  O2A1O1Ixp5_ASAP7_75t_SL U65515 ( .A1(or1200_cpu_or1200_if_insn_saved[16]), 
        .A2(n59682), .B(n60507), .C(n77357), .Y(n2700) );
  NOR2xp33_ASAP7_75t_SL U65516 ( .A(n70949), .B(n70948), .Y(n70963) );
  XNOR2xp5_ASAP7_75t_SL U65517 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[6]), .B(
        n70600), .Y(n70596) );
  NOR2xp33_ASAP7_75t_SL U65518 ( .A(n70074), .B(n70075), .Y(n70089) );
  NOR2xp33_ASAP7_75t_SL U65519 ( .A(n70071), .B(n70070), .Y(n70075) );
  NOR2xp33_ASAP7_75t_SL U65520 ( .A(n70050), .B(n70051), .Y(n70070) );
  NOR2xp33_ASAP7_75t_SL U65521 ( .A(n70047), .B(n70046), .Y(n70051) );
  AOI31xp33_ASAP7_75t_SL U65522 ( .A1(n70010), .A2(n70009), .A3(n70008), .B(
        n70007), .Y(n70046) );
  NOR2xp33_ASAP7_75t_SL U65523 ( .A(n70002), .B(n70047), .Y(n70004) );
  NOR2xp33_ASAP7_75t_SL U65524 ( .A(n69985), .B(n70006), .Y(n70005) );
  AO21x1_ASAP7_75t_SL U65525 ( .A1(n69964), .A2(n69963), .B(n69962), .Y(n70010) );
  NOR2xp33_ASAP7_75t_SL U65526 ( .A(n69933), .B(n69961), .Y(n69960) );
  NOR2xp33_ASAP7_75t_SL U65527 ( .A(n69891), .B(n69890), .Y(n69909) );
  NOR2xp33_ASAP7_75t_SL U65528 ( .A(n69884), .B(n69911), .Y(n69910) );
  NOR2xp33_ASAP7_75t_SL U65529 ( .A(n69829), .B(n69849), .Y(n69830) );
  NOR2xp33_ASAP7_75t_SL U65530 ( .A(n69816), .B(n69832), .Y(n69831) );
  NOR2xp33_ASAP7_75t_SL U65531 ( .A(n69773), .B(n69770), .Y(n69756) );
  NOR2xp33_ASAP7_75t_SL U65532 ( .A(n69748), .B(n69758), .Y(n69757) );
  NOR2xp33_ASAP7_75t_SL U65533 ( .A(n69799), .B(n69817), .Y(n69804) );
  NOR2xp33_ASAP7_75t_SL U65534 ( .A(n69908), .B(n69958), .Y(n69916) );
  OR2x2_ASAP7_75t_SL U65535 ( .A(n70502), .B(n70372), .Y(n58553) );
  O2A1O1Ixp5_ASAP7_75t_SL U65536 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[25]), .A2(n69714), .B(
        n59520), .C(n70098), .Y(n69715) );
  NOR2xp33_ASAP7_75t_SL U65537 ( .A(n69702), .B(n69701), .Y(n70002) );
  NOR2xp33_ASAP7_75t_SL U65538 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_20_), .B(n70011), 
        .Y(n70047) );
  NOR2xp33_ASAP7_75t_SL U65539 ( .A(n69696), .B(n69695), .Y(n70011) );
  NOR2xp33_ASAP7_75t_SL U65540 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_19_), .B(n69988), 
        .Y(n70006) );
  NOR2xp33_ASAP7_75t_SL U65541 ( .A(n69692), .B(n69691), .Y(n69988) );
  NOR2xp33_ASAP7_75t_SL U65542 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_18_), .B(n69965), 
        .Y(n70003) );
  NOR2xp33_ASAP7_75t_SL U65543 ( .A(n69681), .B(n69684), .Y(n69965) );
  NOR2xp33_ASAP7_75t_SL U65544 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_17_), .B(n69935), 
        .Y(n69961) );
  NOR2xp33_ASAP7_75t_SL U65545 ( .A(n69679), .B(n69678), .Y(n69935) );
  NOR2xp33_ASAP7_75t_SL U65546 ( .A(n69678), .B(n69674), .Y(n69933) );
  NOR2xp33_ASAP7_75t_SL U65547 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_16_), .B(n69917), 
        .Y(n69958) );
  NOR2xp33_ASAP7_75t_SL U65548 ( .A(n69671), .B(n69670), .Y(n69908) );
  NOR2xp33_ASAP7_75t_SL U65549 ( .A(n69669), .B(n69668), .Y(n69917) );
  NOR2xp33_ASAP7_75t_SL U65550 ( .A(n69665), .B(n69664), .Y(n69891) );
  NOR2xp33_ASAP7_75t_SL U65551 ( .A(n69663), .B(n69662), .Y(n69884) );
  NOR2xp33_ASAP7_75t_SL U65552 ( .A(n69911), .B(n69656), .Y(n69913) );
  NOR2xp33_ASAP7_75t_SL U65553 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_14_), .B(n69887), 
        .Y(n69911) );
  NOR2xp33_ASAP7_75t_SL U65554 ( .A(n69653), .B(n69652), .Y(n69887) );
  NOR2xp33_ASAP7_75t_SL U65555 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_15_), .B(n69893), 
        .Y(n69890) );
  NOR2xp33_ASAP7_75t_SL U65556 ( .A(n69649), .B(n69648), .Y(n69893) );
  NOR2xp33_ASAP7_75t_SL U65557 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_11_), .B(n69838), 
        .Y(n69849) );
  NOR2xp33_ASAP7_75t_SL U65558 ( .A(n69643), .B(n69642), .Y(n69838) );
  INVxp33_ASAP7_75t_SRAM U65559 ( .A(n69829), .Y(n69634) );
  NOR2xp33_ASAP7_75t_SL U65560 ( .A(n69643), .B(n69633), .Y(n69829) );
  NOR2xp33_ASAP7_75t_SL U65561 ( .A(n69821), .B(n70103), .Y(n69643) );
  INVxp33_ASAP7_75t_SRAM U65562 ( .A(n69816), .Y(n69635) );
  NOR2xp33_ASAP7_75t_SL U65563 ( .A(n69630), .B(n69629), .Y(n69816) );
  INVxp33_ASAP7_75t_SRAM U65564 ( .A(n69834), .Y(n69636) );
  NOR2xp33_ASAP7_75t_SL U65565 ( .A(n69832), .B(n69817), .Y(n69834) );
  NOR2xp33_ASAP7_75t_SL U65566 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_9_), .B(n69805), .Y(
        n69817) );
  NOR2xp33_ASAP7_75t_SL U65567 ( .A(n69626), .B(n69625), .Y(n69805) );
  NOR2xp33_ASAP7_75t_SL U65568 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_10_), .B(n69819), 
        .Y(n69832) );
  NOR2xp33_ASAP7_75t_SL U65569 ( .A(n69627), .B(n69630), .Y(n69819) );
  NOR2xp33_ASAP7_75t_SL U65570 ( .A(n69626), .B(n69623), .Y(n69799) );
  NOR2xp33_ASAP7_75t_SL U65571 ( .A(n69620), .B(n70103), .Y(n69626) );
  NOR2xp33_ASAP7_75t_SL U65572 ( .A(n69788), .B(n70515), .Y(n69802) );
  INVxp33_ASAP7_75t_SRAM U65573 ( .A(n69800), .Y(n69617) );
  NOR2xp33_ASAP7_75t_SL U65574 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_5_), .B(n69753), .Y(
        n69770) );
  NOR2xp33_ASAP7_75t_SL U65575 ( .A(n69615), .B(n69614), .Y(n69753) );
  NOR2xp33_ASAP7_75t_SL U65576 ( .A(n69608), .B(n69607), .Y(n69748) );
  NOR2xp33_ASAP7_75t_SL U65577 ( .A(n69615), .B(n69604), .Y(n69773) );
  NOR2xp33_ASAP7_75t_SL U65578 ( .A(n69602), .B(n59521), .Y(n69614) );
  NOR2xp33_ASAP7_75t_SL U65579 ( .A(n69752), .B(n70103), .Y(n69615) );
  NOR2xp33_ASAP7_75t_SL U65580 ( .A(n69600), .B(n69599), .Y(n69785) );
  NOR2xp33_ASAP7_75t_SL U65581 ( .A(n69608), .B(n69605), .Y(n69751) );
  NOR2xp33_ASAP7_75t_SL U65582 ( .A(n69598), .B(n59520), .Y(n69605) );
  NOR2xp33_ASAP7_75t_SL U65583 ( .A(n69597), .B(n70103), .Y(n69608) );
  NOR2xp33_ASAP7_75t_SL U65584 ( .A(n69755), .B(n69596), .Y(n69750) );
  AOI31xp33_ASAP7_75t_SL U65585 ( .A1(n69728), .A2(n69595), .A3(n69726), .B(
        n69727), .Y(n69735) );
  NOR2xp33_ASAP7_75t_SL U65586 ( .A(n69594), .B(n69730), .Y(n69727) );
  NOR2xp33_ASAP7_75t_SL U65587 ( .A(n69589), .B(n69755), .Y(n69734) );
  NOR2xp33_ASAP7_75t_SL U65588 ( .A(n69588), .B(n69587), .Y(n69589) );
  NOR2xp33_ASAP7_75t_SL U65589 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_3_), .B(n69736), .Y(
        n69755) );
  NOR2xp33_ASAP7_75t_SL U65590 ( .A(n69586), .B(n69585), .Y(n69736) );
  NOR2xp33_ASAP7_75t_SL U65591 ( .A(n69731), .B(n70103), .Y(n69586) );
  INVxp33_ASAP7_75t_SRAM U65592 ( .A(n63878), .Y(n63256) );
  INVxp33_ASAP7_75t_SRAM U65593 ( .A(n63883), .Y(n63244) );
  NOR2xp33_ASAP7_75t_SL U65594 ( .A(n65112), .B(n65111), .Y(n65121) );
  O2A1O1Ixp5_ASAP7_75t_SL U65595 ( .A1(n60497), .A2(n60496), .B(n77566), .C(
        n60495), .Y(n60498) );
  NOR2xp33_ASAP7_75t_SL U65596 ( .A(n65261), .B(n65267), .Y(n65271) );
  O2A1O1Ixp5_ASAP7_75t_SL U65597 ( .A1(n77427), .A2(n61149), .B(n61155), .C(
        n61148), .Y(n61150) );
  INVxp33_ASAP7_75t_SRAM U65598 ( .A(n1753), .Y(n62009) );
  NAND2xp33_ASAP7_75t_SRAM U65599 ( .A(n62016), .B(n61139), .Y(n61143) );
  NAND2xp33_ASAP7_75t_SRAM U65600 ( .A(n3390), .B(n2517), .Y(n62014) );
  AOI211xp5_ASAP7_75t_SL U65601 ( .A1(n76926), .A2(n76565), .B(n76564), .C(
        n76563), .Y(n76567) );
  INVxp33_ASAP7_75t_SRAM U65602 ( .A(or1200_ic_top_from_icram[24]), .Y(n60485)
         );
  INVxp33_ASAP7_75t_SRAM U65603 ( .A(or1200_ic_top_from_icram[2]), .Y(n60350)
         );
  INVxp33_ASAP7_75t_SRAM U65604 ( .A(or1200_ic_top_from_icram[5]), .Y(n61594)
         );
  INVxp33_ASAP7_75t_SRAM U65605 ( .A(or1200_ic_top_from_icram[10]), .Y(n77380)
         );
  INVxp33_ASAP7_75t_SRAM U65606 ( .A(or1200_ic_top_from_icram[3]), .Y(n60357)
         );
  INVxp33_ASAP7_75t_SRAM U65607 ( .A(or1200_ic_top_from_icram[1]), .Y(n60378)
         );
  INVxp33_ASAP7_75t_SRAM U65608 ( .A(or1200_ic_top_from_icram[4]), .Y(n60896)
         );
  INVxp33_ASAP7_75t_SRAM U65609 ( .A(or1200_ic_top_from_icram[8]), .Y(n60394)
         );
  INVxp33_ASAP7_75t_SRAM U65610 ( .A(or1200_ic_top_from_icram[9]), .Y(n60400)
         );
  INVxp33_ASAP7_75t_SRAM U65611 ( .A(or1200_ic_top_from_icram[25]), .Y(n60476)
         );
  INVxp33_ASAP7_75t_SRAM U65612 ( .A(or1200_ic_top_from_icram[23]), .Y(n60415)
         );
  INVxp33_ASAP7_75t_SRAM U65613 ( .A(or1200_ic_top_from_icram[0]), .Y(n60368)
         );
  INVxp33_ASAP7_75t_SRAM U65614 ( .A(or1200_ic_top_from_icram[6]), .Y(n61027)
         );
  INVxp33_ASAP7_75t_SRAM U65615 ( .A(or1200_ic_top_from_icram[7]), .Y(n60388)
         );
  NAND3xp33_ASAP7_75t_SL U65616 ( .A(n78250), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_2_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r2_0_), .Y(n65398) );
  NOR2xp33_ASAP7_75t_SL U65617 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_16_), .B(n65298), .Y(
        n65289) );
  NOR2xp33_ASAP7_75t_SL U65618 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_0_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_1_), .Y(n65396) );
  AOI31xp33_ASAP7_75t_SL U65619 ( .A1(n62001), .A2(n77425), .A3(n61028), .B(
        n60719), .Y(n77461) );
  NOR3xp33_ASAP7_75t_SL U65620 ( .A(n57093), .B(n60723), .C(n60718), .Y(n60719) );
  NOR2xp33_ASAP7_75t_SL U65621 ( .A(n62024), .B(n57072), .Y(n62001) );
  XNOR2xp5_ASAP7_75t_SL U65622 ( .A(n77173), .B(n77172), .Y(n77458) );
  NOR2xp33_ASAP7_75t_SL U65623 ( .A(n69339), .B(n69340), .Y(n77172) );
  NOR2xp33_ASAP7_75t_SL U65624 ( .A(n2517), .B(n69338), .Y(n69340) );
  NOR2xp33_ASAP7_75t_SL U65625 ( .A(n69337), .B(n69336), .Y(n69339) );
  O2A1O1Ixp5_ASAP7_75t_SL U65626 ( .A1(n59442), .A2(n75227), .B(n61524), .C(
        n59564), .Y(n60969) );
  OAI21xp33_ASAP7_75t_SRAM U65627 ( .A1(or1200_cpu_or1200_mult_mac_n289), .A2(
        n77073), .B(n60966), .Y(n60967) );
  NOR4xp25_ASAP7_75t_SL U65628 ( .A(n75224), .B(n61870), .C(n75236), .D(n60956), .Y(n75346) );
  NOR2xp33_ASAP7_75t_SL U65629 ( .A(n61873), .B(n60942), .Y(n75233) );
  NOR2xp33_ASAP7_75t_SL U65630 ( .A(n61878), .B(n60937), .Y(n62123) );
  NOR2xp33_ASAP7_75t_SL U65631 ( .A(n60792), .B(n61854), .Y(n77060) );
  XOR2xp5_ASAP7_75t_SL U65632 ( .A(n60936), .B(n60935), .Y(n60951) );
  O2A1O1Ixp5_ASAP7_75t_SL U65633 ( .A1(n62604), .A2(n60934), .B(n62644), .C(
        n60933), .Y(n60953) );
  NOR2xp33_ASAP7_75t_SL U65634 ( .A(n60912), .B(n60911), .Y(n64248) );
  INVx1_ASAP7_75t_SL U65635 ( .A(n77128), .Y(n76744) );
  OAI22xp33_ASAP7_75t_SRAM U65636 ( .A1(n1983), .A2(n61226), .B1(n1985), .B2(
        n76717), .Y(n60977) );
  AOI211xp5_ASAP7_75t_SL U65637 ( .A1(n61595), .A2(n60900), .B(n60899), .C(
        n60898), .Y(n60902) );
  OAI22xp33_ASAP7_75t_SRAM U65638 ( .A1(n1177), .A2(n61597), .B1(n1422), .B2(
        n60897), .Y(n60898) );
  INVxp33_ASAP7_75t_SRAM U65639 ( .A(n1484), .Y(n60900) );
  NOR2xp33_ASAP7_75t_SL U65640 ( .A(n2814), .B(n60338), .Y(n60720) );
  NOR2xp33_ASAP7_75t_SL U65641 ( .A(n2616), .B(n2609), .Y(n61030) );
  NAND4xp25_ASAP7_75t_SL U65642 ( .A(n60713), .B(n60712), .C(n60711), .D(
        n60710), .Y(n61056) );
  XNOR2xp5_ASAP7_75t_SL U65643 ( .A(n2685), .B(n2023), .Y(n60710) );
  XNOR2xp5_ASAP7_75t_SL U65644 ( .A(n2657), .B(n2572), .Y(n60711) );
  NOR2xp33_ASAP7_75t_SL U65645 ( .A(n2188), .B(n60709), .Y(n60712) );
  NOR2xp33_ASAP7_75t_SL U65646 ( .A(n60708), .B(n60707), .Y(n60713) );
  NAND3xp33_ASAP7_75t_SL U65647 ( .A(n60841), .B(n2807), .C(n2567), .Y(n60690)
         );
  NOR2xp33_ASAP7_75t_SL U65648 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_3_), .B(
        n78436), .Y(n74802) );
  NOR2xp33_ASAP7_75t_SL U65649 ( .A(n60688), .B(n60687), .Y(n75876) );
  NOR2xp33_ASAP7_75t_SL U65650 ( .A(n77763), .B(n77726), .Y(n60687) );
  NOR2xp33_ASAP7_75t_SL U65651 ( .A(n77751), .B(n77756), .Y(n77726) );
  NOR2xp33_ASAP7_75t_SL U65652 ( .A(n60671), .B(n60672), .Y(n76775) );
  O2A1O1Ixp5_ASAP7_75t_SL U65653 ( .A1(n60666), .A2(n63668), .B(n60946), .C(
        n60665), .Y(n60675) );
  NOR4xp25_ASAP7_75t_SL U65654 ( .A(n64304), .B(n60664), .C(n64836), .D(n64110), .Y(n64113) );
  AOI31xp33_ASAP7_75t_SL U65655 ( .A1(n60863), .A2(n60661), .A3(n60660), .B(
        n60659), .Y(n62366) );
  O2A1O1Ixp5_ASAP7_75t_SL U65656 ( .A1(n59565), .A2(n59183), .B(n59568), .C(
        n59079), .Y(n60655) );
  NOR2xp33_ASAP7_75t_SL U65657 ( .A(n2587), .B(n61858), .Y(n75853) );
  O2A1O1Ixp5_ASAP7_75t_SL U65658 ( .A1(n60641), .A2(n75740), .B(n61411), .C(
        n60640), .Y(n60649) );
  O2A1O1Ixp5_ASAP7_75t_SL U65659 ( .A1(n59528), .A2(n75832), .B(n59574), .C(
        n57215), .Y(n60641) );
  NOR4xp25_ASAP7_75t_SL U65660 ( .A(n75706), .B(n60637), .C(n75482), .D(n60636), .Y(n64132) );
  INVxp33_ASAP7_75t_SRAM U65661 ( .A(n64858), .Y(n76749) );
  NOR2xp33_ASAP7_75t_SL U65662 ( .A(n60621), .B(n60672), .Y(n61697) );
  INVxp33_ASAP7_75t_SRAM U65663 ( .A(n3123), .Y(n61336) );
  NOR2xp33_ASAP7_75t_SL U65664 ( .A(n60619), .B(n61649), .Y(n61215) );
  NOR2xp33_ASAP7_75t_SL U65665 ( .A(n60616), .B(n61408), .Y(n61429) );
  NOR2xp33_ASAP7_75t_SL U65666 ( .A(n60614), .B(n60854), .Y(n60872) );
  O2A1O1Ixp5_ASAP7_75t_SL U65667 ( .A1(n59559), .A2(n59079), .B(n59568), .C(
        n59183), .Y(n60606) );
  NOR2xp33_ASAP7_75t_SL U65668 ( .A(n60591), .B(n61852), .Y(n77125) );
  NOR2xp33_ASAP7_75t_SL U65669 ( .A(n3423), .B(n77708), .Y(n77751) );
  NOR2xp33_ASAP7_75t_SL U65670 ( .A(n77729), .B(n61852), .Y(n62292) );
  OR2x2_ASAP7_75t_SL U65671 ( .A(n77763), .B(n60688), .Y(n61852) );
  NAND3xp33_ASAP7_75t_SL U65672 ( .A(n60590), .B(n2581), .C(n2567), .Y(n60688)
         );
  INVx1_ASAP7_75t_SL U65673 ( .A(n3076), .Y(n77763) );
  NOR2xp33_ASAP7_75t_SL U65674 ( .A(n2569), .B(n60589), .Y(n77756) );
  NOR2xp33_ASAP7_75t_SL U65675 ( .A(n60588), .B(n60587), .Y(n64796) );
  NOR2xp33_ASAP7_75t_SL U65676 ( .A(n2843), .B(n77770), .Y(n77752) );
  NOR2xp33_ASAP7_75t_SL U65677 ( .A(n62254), .B(n61546), .Y(n61544) );
  NOR2xp33_ASAP7_75t_SL U65678 ( .A(n3419), .B(n2843), .Y(n60875) );
  INVxp33_ASAP7_75t_SRAM U65679 ( .A(or1200_cpu_or1200_mult_mac_n205), .Y(
        n60563) );
  AOI21xp33_ASAP7_75t_SRAM U65680 ( .A1(n77039), .A2(n63270), .B(n60562), .Y(
        n60565) );
  O2A1O1Ixp5_ASAP7_75t_SL U65681 ( .A1(n1486), .A2(n62418), .B(n60561), .C(
        n61746), .Y(n60562) );
  INVxp33_ASAP7_75t_SRAM U65682 ( .A(n1179), .Y(n60560) );
  NOR2xp33_ASAP7_75t_SL U65683 ( .A(n60555), .B(n60899), .Y(n60566) );
  INVxp33_ASAP7_75t_SRAM U65684 ( .A(n76735), .Y(n60570) );
  NOR2xp33_ASAP7_75t_SL U65685 ( .A(n60706), .B(n60705), .Y(n61058) );
  NAND4xp25_ASAP7_75t_SL U65686 ( .A(n60704), .B(n60703), .C(n60702), .D(
        n60995), .Y(n60705) );
  XNOR2xp5_ASAP7_75t_SL U65687 ( .A(n2657), .B(n2575), .Y(n60702) );
  XNOR2xp5_ASAP7_75t_SL U65688 ( .A(n2671), .B(n2062), .Y(n60703) );
  XNOR2xp5_ASAP7_75t_SL U65689 ( .A(n2678), .B(n2045), .Y(n60704) );
  XNOR2xp5_ASAP7_75t_SL U65690 ( .A(n2664), .B(n2079), .Y(n60700) );
  XNOR2xp5_ASAP7_75t_SL U65691 ( .A(n2685), .B(n2026), .Y(n60701) );
  NOR2xp33_ASAP7_75t_SL U65692 ( .A(n73426), .B(n73427), .Y(n73425) );
  NOR2xp33_ASAP7_75t_SL U65693 ( .A(n73423), .B(n73432), .Y(n73427) );
  INVxp33_ASAP7_75t_SRAM U65694 ( .A(n51956), .Y(n73836) );
  NOR2xp33_ASAP7_75t_SL U65695 ( .A(n73462), .B(n73463), .Y(n73461) );
  NOR2xp33_ASAP7_75t_SL U65696 ( .A(n73455), .B(n73468), .Y(n73463) );
  INVxp33_ASAP7_75t_SRAM U65697 ( .A(n78219), .Y(n73846) );
  NOR2xp33_ASAP7_75t_SL U65698 ( .A(n73354), .B(n73396), .Y(n73398) );
  NOR2xp33_ASAP7_75t_SL U65699 ( .A(n73390), .B(n73389), .Y(n73399) );
  AOI31xp33_ASAP7_75t_SL U65700 ( .A1(n73357), .A2(n73408), .A3(n73358), .B(
        n73353), .Y(n73396) );
  AOI31xp33_ASAP7_75t_SL U65701 ( .A1(n73348), .A2(n73347), .A3(n73346), .B(
        n73345), .Y(n73358) );
  NOR2xp33_ASAP7_75t_SL U65702 ( .A(n73336), .B(n73339), .Y(n73348) );
  NOR2xp33_ASAP7_75t_SL U65703 ( .A(n73340), .B(n59630), .Y(n73339) );
  AOI31xp33_ASAP7_75t_SL U65704 ( .A1(n73352), .A2(n73351), .A3(n73350), .B(
        n73335), .Y(n73408) );
  NOR2xp33_ASAP7_75t_SL U65705 ( .A(n73316), .B(n73315), .Y(n73363) );
  NOR2xp33_ASAP7_75t_SL U65706 ( .A(n73310), .B(n73309), .Y(n73316) );
  AOI31xp33_ASAP7_75t_SL U65707 ( .A1(n73320), .A2(n73319), .A3(n73318), .B(
        n73306), .Y(n73366) );
  AOI31xp33_ASAP7_75t_SL U65708 ( .A1(n73453), .A2(n73454), .A3(n73452), .B(
        n73270), .Y(n73420) );
  AOI211xp5_ASAP7_75t_SL U65709 ( .A1(n73470), .A2(n73263), .B(n73262), .C(
        n73261), .Y(n73454) );
  XNOR2xp5_ASAP7_75t_SL U65710 ( .A(n73256), .B(n73255), .Y(n73470) );
  NOR2xp33_ASAP7_75t_SL U65711 ( .A(n73473), .B(n73471), .Y(n73252) );
  NOR2xp33_ASAP7_75t_SL U65712 ( .A(n73475), .B(n73476), .Y(n73263) );
  XNOR2xp5_ASAP7_75t_SL U65713 ( .A(n73225), .B(n73224), .Y(n73476) );
  NOR2xp33_ASAP7_75t_SL U65714 ( .A(n73222), .B(n59631), .Y(n73259) );
  NOR2xp33_ASAP7_75t_SL U65715 ( .A(n73253), .B(n73254), .Y(n73475) );
  NOR2xp33_ASAP7_75t_SL U65716 ( .A(n73216), .B(n73215), .Y(n73253) );
  NOR2xp33_ASAP7_75t_SL U65717 ( .A(n73217), .B(n59630), .Y(n73215) );
  XNOR2xp5_ASAP7_75t_SL U65718 ( .A(n73206), .B(n73205), .Y(n73462) );
  NOR2xp33_ASAP7_75t_SL U65719 ( .A(n73456), .B(n73465), .Y(n73269) );
  NOR2xp33_ASAP7_75t_SL U65720 ( .A(n73196), .B(n73195), .Y(n73201) );
  NOR2xp33_ASAP7_75t_SL U65721 ( .A(n73211), .B(n59631), .Y(n73195) );
  NOR2xp33_ASAP7_75t_SL U65722 ( .A(n73203), .B(n73204), .Y(n73456) );
  NOR2xp33_ASAP7_75t_SL U65723 ( .A(n73190), .B(n73189), .Y(n73203) );
  AOI31xp33_ASAP7_75t_SL U65724 ( .A1(n73278), .A2(n73277), .A3(n73276), .B(
        n73187), .Y(n73416) );
  AOI22xp33_ASAP7_75t_SRAM U65725 ( .A1(n73379), .A2(n73185), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[13]), .B2(
        n73382), .Y(n73278) );
  AOI31xp33_ASAP7_75t_SL U65726 ( .A1(n73274), .A2(n73273), .A3(n73272), .B(
        n73182), .Y(n73417) );
  O2A1O1Ixp5_ASAP7_75t_SL U65727 ( .A1(n73180), .A2(n57185), .B(n73179), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[12]), .Y(
        n73181) );
  NOR2xp33_ASAP7_75t_SL U65728 ( .A(n73167), .B(n73170), .Y(n73178) );
  NOR2xp33_ASAP7_75t_SL U65729 ( .A(n73169), .B(n59630), .Y(n73167) );
  NOR2xp33_ASAP7_75t_SL U65730 ( .A(n73415), .B(n73440), .Y(n73289) );
  NOR2xp33_ASAP7_75t_SL U65731 ( .A(n73144), .B(n59630), .Y(n73151) );
  NOR2xp33_ASAP7_75t_SL U65732 ( .A(n73435), .B(n73445), .Y(n73301) );
  AOI31xp33_ASAP7_75t_SL U65733 ( .A1(n73299), .A2(n73298), .A3(n73297), .B(
        n73137), .Y(n73295) );
  AOI31xp33_ASAP7_75t_SL U65734 ( .A1(n73324), .A2(n73323), .A3(n73322), .B(
        n73125), .Y(n73359) );
  O2A1O1Ixp5_ASAP7_75t_SL U65735 ( .A1(n73123), .A2(n57185), .B(n73122), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[20]), .Y(
        n73124) );
  AOI31xp33_ASAP7_75t_SL U65736 ( .A1(n73327), .A2(n73326), .A3(n73325), .B(
        n73121), .Y(n73367) );
  NOR2xp33_ASAP7_75t_SL U65737 ( .A(n73113), .B(n73112), .Y(n73390) );
  AOI31xp33_ASAP7_75t_SL U65738 ( .A1(n73393), .A2(n73392), .A3(n73391), .B(
        n73387), .Y(n73400) );
  XNOR2xp5_ASAP7_75t_SL U65739 ( .A(n27420), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n254), .Y(n59525) );
  XOR2xp5_ASAP7_75t_SL U65740 ( .A(n74502), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[26]), .Y(
        n73375) );
  XNOR2xp5_ASAP7_75t_SL U65741 ( .A(n3128), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1[0]), .Y(n76983) );
  OAI22xp33_ASAP7_75t_SRAM U65742 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[15]), .A2(
        n73144), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[16]), .B2(
        n73128), .Y(n73087) );
  NOR2xp33_ASAP7_75t_SL U65743 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[22]), .B(
        n73340), .Y(n73086) );
  AOI22xp33_ASAP7_75t_SRAM U65744 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[18]), .A2(
        n73308), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[17]), .B2(
        n73076), .Y(n73077) );
  NOR2xp33_ASAP7_75t_SL U65745 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[17]), .B(
        n73076), .Y(n73134) );
  NAND2xp33_ASAP7_75t_SRAM U65746 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[16]), .B(
        n73128), .Y(n73078) );
  AOI211xp5_ASAP7_75t_SL U65747 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[14]), .A2(
        n73140), .B(n73083), .C(n73147), .Y(n73081) );
  NOR2xp33_ASAP7_75t_SL U65748 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[15]), .B(
        n73150), .Y(n73147) );
  NOR2xp33_ASAP7_75t_SL U65749 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[21]), .B(
        n73119), .Y(n73083) );
  OAI22xp33_ASAP7_75t_SRAM U65750 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[10]), .A2(
        n73163), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[9]), .B2(
        n73156), .Y(n73074) );
  NAND2xp33_ASAP7_75t_SRAM U65751 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[10]), .B(
        n73163), .Y(n73066) );
  NAND2xp33_ASAP7_75t_SRAM U65752 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[11]), .B(
        n73171), .Y(n73067) );
  NOR2xp33_ASAP7_75t_SL U65753 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[8]), .B(
        n73211), .Y(n73208) );
  NOR2xp33_ASAP7_75t_SL U65754 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[7]), .B(
        n73191), .Y(n73052) );
  NOR2xp33_ASAP7_75t_SL U65755 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[6]), .B(
        n73265), .Y(n73054) );
  NOR2xp33_ASAP7_75t_SL U65756 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[5]), .B(
        n73221), .Y(n73257) );
  OAI22xp33_ASAP7_75t_SRAM U65757 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[4]), .A2(
        n73219), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[3]), .B2(
        n73238), .Y(n73051) );
  OAI22xp33_ASAP7_75t_SRAM U65758 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[3]), .A2(
        n73239), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[2]), .B2(
        n73244), .Y(n73061) );
  OAI22xp33_ASAP7_75t_SRAM U65759 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[2]), .A2(
        n73241), .B1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[1]), .B2(
        n73229), .Y(n73048) );
  NOR2xp33_ASAP7_75t_SL U65760 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[0]), .B(
        n73231), .Y(n73483) );
  NOR3xp33_ASAP7_75t_SL U65761 ( .A(n69438), .B(n69437), .C(n65236), .Y(n70154) );
  NOR2xp33_ASAP7_75t_SL U65762 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_21_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_20_), .Y(n69385) );
  NOR2xp33_ASAP7_75t_SL U65763 ( .A(n69404), .B(n69395), .Y(n69435) );
  OR2x2_ASAP7_75t_SL U65764 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_17_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_16_), .Y(n69395) );
  NOR2xp33_ASAP7_75t_SL U65765 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_15_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_14_), .Y(n69400) );
  NOR2xp33_ASAP7_75t_SL U65766 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_13_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_12_), .Y(n69386) );
  NOR2xp33_ASAP7_75t_SL U65767 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_9_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_8_), .Y(n69388) );
  NOR2xp33_ASAP7_75t_SL U65768 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_11_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_10_), .Y(n69393) );
  NOR2xp33_ASAP7_75t_SL U65769 ( .A(n69428), .B(n69426), .Y(n69439) );
  NOR2xp33_ASAP7_75t_SL U65770 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_7_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_6_), .Y(n69394) );
  NOR2xp33_ASAP7_75t_SL U65771 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_3_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_), .Y(n69392) );
  NOR2xp33_ASAP7_75t_SL U65772 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_0_), .Y(n69390) );
  NOR2xp33_ASAP7_75t_SL U65773 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[17]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[16]), .Y(n69541) );
  NOR2xp33_ASAP7_75t_SL U65774 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[18]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[19]), .Y(n69547) );
  NOR2xp33_ASAP7_75t_SL U65775 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[20]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[21]), .Y(n69545) );
  INVx1_ASAP7_75t_SL U65776 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[22]), .Y(n78364) );
  NOR2xp33_ASAP7_75t_SL U65777 ( .A(n69529), .B(n69527), .Y(n74499) );
  NOR2xp33_ASAP7_75t_SL U65778 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[14]), .Y(n69540) );
  NOR2xp33_ASAP7_75t_SL U65779 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[12]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[13]), .Y(n69543) );
  NAND3xp33_ASAP7_75t_SL U65780 ( .A(n69523), .B(n78344), .C(n78348), .Y(
        n69529) );
  NOR2xp33_ASAP7_75t_SL U65781 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[8]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[11]), .Y(n69523) );
  NOR2xp33_ASAP7_75t_SL U65782 ( .A(n69526), .B(n69530), .Y(n74500) );
  NOR2xp33_ASAP7_75t_SL U65783 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[1]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[0]), .Y(n69535)
         );
  NOR2xp33_ASAP7_75t_SL U65784 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[3]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[2]), .Y(n69532)
         );
  NOR2xp33_ASAP7_75t_SL U65785 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[6]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[7]), .Y(n69538)
         );
  NOR2xp33_ASAP7_75t_SL U65786 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[5]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[4]), .Y(n69533)
         );
  INVxp33_ASAP7_75t_SRAM U65787 ( .A(n74497), .Y(n74501) );
  XNOR2xp5_ASAP7_75t_SL U65788 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_31_), .B(n74518), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n254) );
  INVx1_ASAP7_75t_SL U65789 ( .A(n3128), .Y(n74518) );
  INVx1_ASAP7_75t_SL U65790 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r1[0]), .Y(n27420) );
  AOI211xp5_ASAP7_75t_SL U65791 ( .A1(n77373), .A2(n60510), .B(n60509), .C(
        n60508), .Y(n9589) );
  INVxp33_ASAP7_75t_SRAM U65792 ( .A(n74257), .Y(n74259) );
  NOR2xp33_ASAP7_75t_SL U65793 ( .A(n57269), .B(n68748), .Y(n68752) );
  AND2x2_ASAP7_75t_SL U65794 ( .A(n2616), .B(n2609), .Y(n62142) );
  NOR2xp33_ASAP7_75t_SL U65795 ( .A(n2589), .B(n61145), .Y(n61312) );
  NOR2xp33_ASAP7_75t_SL U65796 ( .A(n74994), .B(n75788), .Y(n74995) );
  NOR2xp33_ASAP7_75t_SL U65797 ( .A(n75789), .B(n75790), .Y(n75788) );
  NAND2xp33_ASAP7_75t_SRAM U65798 ( .A(n74992), .B(n74991), .Y(n74996) );
  OAI22xp33_ASAP7_75t_SRAM U65799 ( .A1(or1200_cpu_or1200_except_n170), .A2(
        n57070), .B1(n76828), .B2(n77294), .Y(n76640) );
  OAI22xp33_ASAP7_75t_SRAM U65800 ( .A1(or1200_cpu_or1200_except_n178), .A2(
        n57070), .B1(n77594), .B2(n77294), .Y(n76998) );
  OAI22xp33_ASAP7_75t_SRAM U65801 ( .A1(or1200_cpu_or1200_except_n172), .A2(
        n57070), .B1(n77603), .B2(n77294), .Y(n76697) );
  XNOR2xp5_ASAP7_75t_SL U65802 ( .A(n76696), .B(n76695), .Y(n77982) );
  OAI22xp33_ASAP7_75t_SRAM U65803 ( .A1(or1200_cpu_or1200_except_n166), .A2(
        n57070), .B1(n75781), .B2(n77294), .Y(n75782) );
  OAI22xp33_ASAP7_75t_SRAM U65804 ( .A1(or1200_cpu_or1200_except_n174), .A2(
        n57070), .B1(n77600), .B2(n77294), .Y(n76618) );
  INVxp33_ASAP7_75t_SRAM U65805 ( .A(n74240), .Y(n74241) );
  NAND2xp5_ASAP7_75t_SL U65806 ( .A(n60335), .B(n76538), .Y(n60337) );
  OAI22xp33_ASAP7_75t_SRAM U65807 ( .A1(or1200_cpu_or1200_except_n164), .A2(
        n57070), .B1(n77615), .B2(n77294), .Y(n76552) );
  NOR2xp33_ASAP7_75t_SL U65808 ( .A(n76245), .B(n76244), .Y(n77990) );
  OAI22xp33_ASAP7_75t_SRAM U65809 ( .A1(or1200_cpu_or1200_except_n130), .A2(
        n57070), .B1(n77177), .B2(n77294), .Y(n77178) );
  OAI22xp33_ASAP7_75t_SRAM U65810 ( .A1(or1200_cpu_or1200_except_n182), .A2(
        n57070), .B1(n76688), .B2(n77294), .Y(n76684) );
  OAI22xp33_ASAP7_75t_SRAM U65811 ( .A1(or1200_cpu_or1200_except_n132), .A2(
        n57070), .B1(n75796), .B2(n77294), .Y(n75797) );
  O2A1O1Ixp5_ASAP7_75t_SL U65812 ( .A1(n76836), .A2(n76835), .B(n76834), .C(
        n77269), .Y(n77262) );
  OAI22xp33_ASAP7_75t_SRAM U65813 ( .A1(or1200_cpu_or1200_except_n142), .A2(
        n57070), .B1(n75447), .B2(n77294), .Y(n75448) );
  OAI22xp33_ASAP7_75t_SRAM U65814 ( .A1(or1200_cpu_or1200_except_n128), .A2(
        n57070), .B1(n75198), .B2(n77294), .Y(n75199) );
  OAI22xp33_ASAP7_75t_SRAM U65815 ( .A1(or1200_cpu_or1200_except_n156), .A2(
        n57070), .B1(n77646), .B2(n77294), .Y(n77152) );
  OAI22xp33_ASAP7_75t_SRAM U65816 ( .A1(or1200_cpu_or1200_except_n126), .A2(
        n57070), .B1(n75675), .B2(n77294), .Y(n75676) );
  OAI22xp33_ASAP7_75t_SRAM U65817 ( .A1(or1200_cpu_or1200_except_n124), .A2(
        n57070), .B1(n77673), .B2(n77294), .Y(n76919) );
  OAI22xp33_ASAP7_75t_SRAM U65818 ( .A1(or1200_cpu_or1200_except_n154), .A2(
        n57070), .B1(n76235), .B2(n77294), .Y(n76231) );
  OAI22xp33_ASAP7_75t_SRAM U65819 ( .A1(or1200_cpu_or1200_except_n158), .A2(
        n57070), .B1(n77019), .B2(n77294), .Y(n77020) );
  OAI22xp33_ASAP7_75t_SRAM U65820 ( .A1(or1200_cpu_or1200_except_n180), .A2(
        n57070), .B1(n77591), .B2(n77294), .Y(n76863) );
  OAI22xp33_ASAP7_75t_SRAM U65821 ( .A1(or1200_cpu_or1200_except_n162), .A2(
        n57070), .B1(n77295), .B2(n77294), .Y(n77297) );
  OAI22xp33_ASAP7_75t_SRAM U65822 ( .A1(or1200_cpu_or1200_except_n160), .A2(
        n57070), .B1(n77637), .B2(n77294), .Y(n77226) );
  NOR2xp33_ASAP7_75t_SL U65823 ( .A(n78154), .B(n78155), .Y(n77225) );
  NOR2xp33_ASAP7_75t_SL U65824 ( .A(n60817), .B(n77165), .Y(n77048) );
  NOR2xp33_ASAP7_75t_SL U65825 ( .A(or1200_cpu_or1200_except_n266), .B(n76507), 
        .Y(n76510) );
  NOR2xp33_ASAP7_75t_SL U65826 ( .A(n76663), .B(n76731), .Y(n62155) );
  OAI21xp33_ASAP7_75t_SRAM U65827 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_1_), 
        .A2(n76489), .B(n78436), .Y(n76488) );
  NOR2xp33_ASAP7_75t_SL U65828 ( .A(n76476), .B(n76475), .Y(n76493) );
  NOR2xp33_ASAP7_75t_SL U65829 ( .A(n76399), .B(n74007), .Y(n76464) );
  NOR2xp33_ASAP7_75t_SL U65830 ( .A(n74011), .B(n74012), .Y(n76448) );
  NOR2xp33_ASAP7_75t_SL U65831 ( .A(n76436), .B(n76435), .Y(n76774) );
  NOR2xp33_ASAP7_75t_SL U65832 ( .A(n76358), .B(n76360), .Y(n76439) );
  NOR2xp33_ASAP7_75t_SL U65833 ( .A(n61099), .B(n73990), .Y(n76432) );
  AOI22xp33_ASAP7_75t_SRAM U65834 ( .A1(n76472), .A2(n76428), .B1(n76424), 
        .B2(n76423), .Y(n76481) );
  AOI31xp33_ASAP7_75t_SL U65835 ( .A1(n76420), .A2(n76419), .A3(n76422), .B(
        n76418), .Y(n76484) );
  AOI211xp5_ASAP7_75t_SL U65836 ( .A1(n76416), .A2(n76415), .B(n76482), .C(
        n76414), .Y(n76417) );
  INVxp33_ASAP7_75t_SRAM U65837 ( .A(n76410), .Y(n76412) );
  OAI21xp33_ASAP7_75t_SRAM U65838 ( .A1(n59168), .A2(n59167), .B(n76409), .Y(
        n76482) );
  NOR2xp33_ASAP7_75t_SL U65839 ( .A(n74783), .B(n74782), .Y(n74798) );
  AOI21xp33_ASAP7_75t_SRAM U65840 ( .A1(n76386), .A2(n76385), .B(n76384), .Y(
        n76390) );
  NAND2xp33_ASAP7_75t_SRAM U65841 ( .A(n76465), .B(n76365), .Y(n76387) );
  NOR2xp33_ASAP7_75t_SL U65842 ( .A(n74778), .B(n74777), .Y(n76404) );
  NOR2xp33_ASAP7_75t_SL U65843 ( .A(n76326), .B(n76499), .Y(n76495) );
  NOR2xp33_ASAP7_75t_SL U65844 ( .A(n3123), .B(n77142), .Y(n76499) );
  NOR2xp33_ASAP7_75t_SL U65845 ( .A(n75475), .B(n73960), .Y(n77142) );
  NAND2xp33_ASAP7_75t_SRAM U65846 ( .A(n1868), .B(n75890), .Y(n75851) );
  O2A1O1Ixp5_ASAP7_75t_SL U65847 ( .A1(n59533), .A2(n75318), .B(n77713), .C(
        n74006), .Y(n74009) );
  INVxp33_ASAP7_75t_SRAM U65848 ( .A(n73998), .Y(n76452) );
  NOR2xp33_ASAP7_75t_SL U65849 ( .A(n77064), .B(n73992), .Y(n76465) );
  NAND2xp33_ASAP7_75t_SRAM U65850 ( .A(n73991), .B(n76381), .Y(n76364) );
  NAND2xp33_ASAP7_75t_SRAM U65851 ( .A(n76451), .B(n73986), .Y(n76384) );
  NAND2xp33_ASAP7_75t_SRAM U65852 ( .A(n76445), .B(n73985), .Y(n76368) );
  NAND2xp33_ASAP7_75t_SRAM U65853 ( .A(n73981), .B(n73980), .Y(n76367) );
  NOR2xp33_ASAP7_75t_SL U65854 ( .A(n73974), .B(n73976), .Y(n76354) );
  AOI21xp33_ASAP7_75t_SRAM U65855 ( .A1(n73970), .A2(n76366), .B(n76436), .Y(
        n76374) );
  NAND2xp33_ASAP7_75t_SRAM U65856 ( .A(n76377), .B(n76466), .Y(n73987) );
  NOR2xp33_ASAP7_75t_SL U65857 ( .A(n77063), .B(n73969), .Y(n76466) );
  NAND2xp33_ASAP7_75t_SRAM U65858 ( .A(n76442), .B(n73989), .Y(n76389) );
  NAND2xp33_ASAP7_75t_SRAM U65859 ( .A(n1588), .B(n64241), .Y(n73965) );
  AOI22xp33_ASAP7_75t_SRAM U65860 ( .A1(n59549), .A2(n57215), .B1(n59550), 
        .B2(n75740), .Y(n76343) );
  NOR2xp33_ASAP7_75t_SL U65861 ( .A(n1868), .B(n75890), .Y(n75849) );
  NOR2xp33_ASAP7_75t_SL U65862 ( .A(n64151), .B(n64150), .Y(n76315) );
  NOR2xp33_ASAP7_75t_SL U65863 ( .A(n64149), .B(n64148), .Y(n64151) );
  NAND4xp25_ASAP7_75t_SL U65864 ( .A(n76296), .B(n76295), .C(n76294), .D(
        n76293), .Y(n76297) );
  NOR4xp25_ASAP7_75t_SL U65865 ( .A(n76292), .B(n76291), .C(n76290), .D(n76289), .Y(n76294) );
  XNOR2xp5_ASAP7_75t_SL U65866 ( .A(n76431), .B(n60752), .Y(n76289) );
  XNOR2xp5_ASAP7_75t_SL U65867 ( .A(n61560), .B(n61559), .Y(n76292) );
  XNOR2xp5_ASAP7_75t_SL U65868 ( .A(n62296), .B(n76278), .Y(n76296) );
  O2A1O1Ixp5_ASAP7_75t_SL U65869 ( .A1(n76279), .A2(n62312), .B(n62311), .C(
        n62310), .Y(n62314) );
  O2A1O1Ixp5_ASAP7_75t_SL U65870 ( .A1(n76288), .A2(n76287), .B(n76286), .C(
        n76285), .Y(n76804) );
  NOR2xp33_ASAP7_75t_SL U65871 ( .A(n61675), .B(n61674), .Y(n61799) );
  XNOR2xp5_ASAP7_75t_SL U65872 ( .A(n58206), .B(n61798), .Y(n61800) );
  XNOR2xp5_ASAP7_75t_SL U65873 ( .A(n61954), .B(n61120), .Y(n76304) );
  NOR2xp33_ASAP7_75t_SL U65874 ( .A(n76276), .B(n76275), .Y(n76309) );
  NOR2xp33_ASAP7_75t_SL U65875 ( .A(n63548), .B(n75307), .Y(n63549) );
  AOI31xp33_ASAP7_75t_SL U65876 ( .A1(n75813), .A2(n75812), .A3(n75811), .B(
        n75810), .Y(n76314) );
  AOI31xp33_ASAP7_75t_SL U65877 ( .A1(n64201), .A2(n64200), .A3(n64199), .B(
        n64198), .Y(n76271) );
  NOR2xp33_ASAP7_75t_SL U65878 ( .A(n73949), .B(n75808), .Y(n73952) );
  NOR2xp33_ASAP7_75t_SL U65879 ( .A(n64810), .B(n64809), .Y(n75808) );
  O2A1O1Ixp5_ASAP7_75t_SL U65880 ( .A1(n76263), .A2(n76262), .B(n76261), .C(
        n76260), .Y(n77030) );
  NOR2xp33_ASAP7_75t_SL U65881 ( .A(n64190), .B(n64756), .Y(n76269) );
  NOR2xp33_ASAP7_75t_SL U65882 ( .A(n75679), .B(n75680), .Y(n75683) );
  NOR2xp33_ASAP7_75t_SL U65883 ( .A(n75811), .B(n75812), .Y(n75806) );
  XNOR2xp5_ASAP7_75t_SL U65884 ( .A(n75890), .B(n61983), .Y(n75812) );
  NOR2xp33_ASAP7_75t_SL U65885 ( .A(n73949), .B(n73950), .Y(n61981) );
  NOR2xp33_ASAP7_75t_SL U65886 ( .A(n57212), .B(n61978), .Y(n73949) );
  AO21x1_ASAP7_75t_SL U65887 ( .A1(n61977), .A2(n65017), .B(n61976), .Y(n61978) );
  NOR2xp33_ASAP7_75t_SL U65888 ( .A(n62081), .B(n61960), .Y(n64269) );
  NOR2xp33_ASAP7_75t_SL U65889 ( .A(n64188), .B(n64185), .Y(n64196) );
  NAND2xp33_ASAP7_75t_SRAM U65890 ( .A(n78170), .B(n61906), .Y(n61907) );
  OAI21xp33_ASAP7_75t_SRAM U65891 ( .A1(n59550), .A2(n57120), .B(n61905), .Y(
        n61906) );
  NOR2xp33_ASAP7_75t_SL U65892 ( .A(n75517), .B(n74029), .Y(n61987) );
  NOR2xp33_ASAP7_75t_SL U65893 ( .A(n76486), .B(n61904), .Y(n74029) );
  NAND2xp33_ASAP7_75t_SRAM U65894 ( .A(n57120), .B(n78170), .Y(n61903) );
  NOR2xp33_ASAP7_75t_SL U65895 ( .A(n64146), .B(n64147), .Y(n64150) );
  NOR2xp33_ASAP7_75t_SL U65896 ( .A(n61934), .B(n63546), .Y(n61935) );
  AOI211xp5_ASAP7_75t_SL U65897 ( .A1(n61950), .A2(n76258), .B(n62499), .C(
        n62500), .Y(n62080) );
  NOR2xp33_ASAP7_75t_SL U65898 ( .A(n59572), .B(n76259), .Y(n62499) );
  XNOR2xp5_ASAP7_75t_SL U65899 ( .A(n76627), .B(n60770), .Y(n76279) );
  NOR2xp33_ASAP7_75t_SL U65900 ( .A(n78005), .B(n57120), .Y(n60761) );
  NOR2xp33_ASAP7_75t_SL U65901 ( .A(n60754), .B(n60753), .Y(n60756) );
  NOR2xp33_ASAP7_75t_SL U65902 ( .A(n76431), .B(n60752), .Y(n60753) );
  NOR2xp33_ASAP7_75t_SL U65903 ( .A(n60844), .B(n73971), .Y(n76431) );
  NOR2xp33_ASAP7_75t_SL U65904 ( .A(n59710), .B(n77242), .Y(n73971) );
  OAI21xp33_ASAP7_75t_SRAM U65905 ( .A1(n59708), .A2(n59646), .B(n57120), .Y(
        n60750) );
  NOR2xp33_ASAP7_75t_SL U65906 ( .A(n76653), .B(n60736), .Y(n61321) );
  NOR2xp33_ASAP7_75t_SL U65907 ( .A(n61954), .B(n61917), .Y(n62076) );
  AOI31xp33_ASAP7_75t_SL U65908 ( .A1(n57128), .A2(n60783), .A3(n60782), .B(
        n60781), .Y(n62466) );
  NOR2xp33_ASAP7_75t_SL U65909 ( .A(n57128), .B(n60780), .Y(n60781) );
  NAND2xp33_ASAP7_75t_SRAM U65910 ( .A(n59542), .B(n60775), .Y(n61673) );
  NOR2xp33_ASAP7_75t_SL U65911 ( .A(n60743), .B(n60744), .Y(n60745) );
  NAND2xp33_ASAP7_75t_SRAM U65912 ( .A(n59540), .B(n60742), .Y(n60743) );
  NOR2xp33_ASAP7_75t_SL U65913 ( .A(n61937), .B(n76263), .Y(n61950) );
  NOR2xp33_ASAP7_75t_SL U65914 ( .A(n57210), .B(n61938), .Y(n61937) );
  O2A1O1Ixp5_ASAP7_75t_SL U65915 ( .A1(n53455), .A2(n62757), .B(n60733), .C(
        n57116), .Y(n61936) );
  XNOR2xp5_ASAP7_75t_SL U65916 ( .A(n57641), .B(n60735), .Y(n61954) );
  INVxp33_ASAP7_75t_SRAM U65917 ( .A(n75477), .Y(n60731) );
  OAI22xp33_ASAP7_75t_SRAM U65918 ( .A1(or1200_cpu_or1200_except_n136), .A2(
        n57070), .B1(n74079), .B2(n77294), .Y(n74080) );
  NOR2xp33_ASAP7_75t_SL U65919 ( .A(n74417), .B(n74505), .Y(n74427) );
  OAI22xp33_ASAP7_75t_SRAM U65920 ( .A1(or1200_cpu_or1200_except_n146), .A2(
        n57070), .B1(n74127), .B2(n77294), .Y(n74128) );
  OAI22xp33_ASAP7_75t_SRAM U65921 ( .A1(or1200_cpu_or1200_except_n134), .A2(
        n57070), .B1(n69371), .B2(n77294), .Y(n69372) );
  OAI22xp33_ASAP7_75t_SRAM U65922 ( .A1(or1200_cpu_or1200_except_n138), .A2(
        n57070), .B1(n74045), .B2(n77294), .Y(n74046) );
  NOR2xp33_ASAP7_75t_SL U65923 ( .A(n58621), .B(n77235), .Y(n77289) );
  NOR2xp33_ASAP7_75t_SL U65924 ( .A(n73907), .B(n60550), .Y(n77852) );
  NOR2xp33_ASAP7_75t_SL U65925 ( .A(n58574), .B(n60547), .Y(n61481) );
  XNOR2xp5_ASAP7_75t_SL U65926 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_6_), 
        .B(n74345), .Y(n74375) );
  AOI31xp33_ASAP7_75t_SL U65927 ( .A1(n74227), .A2(n73861), .A3(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_26_), 
        .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_27_), 
        .Y(n73862) );
  NAND3xp33_ASAP7_75t_SL U65928 ( .A(n74358), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_10_), 
        .C(or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_9_), .Y(n74322) );
  NOR2xp33_ASAP7_75t_SL U65929 ( .A(n73858), .B(n74345), .Y(n74373) );
  XNOR2xp5_ASAP7_75t_SL U65930 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1[0]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_sign_o), .Y(n73855) );
  NOR2xp33_ASAP7_75t_SL U65931 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_0_), 
        .B(n73854), .Y(n74302) );
  NOR2xp33_ASAP7_75t_SL U65932 ( .A(n3310), .B(n3337), .Y(n73854) );
  NOR2xp33_ASAP7_75t_SL U65933 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_2_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_1_), .Y(n74731) );
  NOR2xp33_ASAP7_75t_SL U65934 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[26]), .B(n73486), .Y(
        n73491) );
  AOI31xp33_ASAP7_75t_SL U65935 ( .A1(n73502), .A2(n73743), .A3(n73753), .B(
        n73501), .Y(n73873) );
  NOR2xp33_ASAP7_75t_SL U65936 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[19]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[20]), .Y(n73497) );
  NOR2xp33_ASAP7_75t_SL U65937 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[15]), .B(n73642), .Y(
        n73499) );
  NOR2xp33_ASAP7_75t_SL U65938 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[14]), .Y(n73493) );
  OAI21xp33_ASAP7_75t_SRAM U65939 ( .A1(n73522), .A2(n73523), .B(n73492), .Y(
        n73494) );
  NOR2xp33_ASAP7_75t_SL U65940 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[11]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[12]), .Y(n73492) );
  NOR2xp33_ASAP7_75t_SL U65941 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[7]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[8]), .Y(n73522) );
  OAI21xp33_ASAP7_75t_SRAM U65942 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[1]), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[2]), .B(n73521), .Y(
        n73495) );
  NOR2xp33_ASAP7_75t_SL U65943 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[3]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[4]), .Y(n73521) );
  NOR2xp33_ASAP7_75t_SL U65944 ( .A(n73528), .B(n73523), .Y(n73496) );
  NOR2xp33_ASAP7_75t_SL U65945 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[22]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[20]), .Y(n73515) );
  AOI21xp33_ASAP7_75t_SRAM U65946 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[15]), .A2(n3321), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[17]), .Y(n73511) );
  NOR2xp33_ASAP7_75t_SL U65947 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[14]), .B(n73642), .Y(
        n73508) );
  INVxp33_ASAP7_75t_SRAM U65948 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[12]), .Y(n73509) );
  AOI21xp33_ASAP7_75t_SRAM U65949 ( .A1(n73828), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[2]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[4]), .Y(n73507) );
  NOR4xp25_ASAP7_75t_SL U65950 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[11]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[9]), .C(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]), .D(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[7]), .Y(n73514) );
  OR2x2_ASAP7_75t_SL U65951 ( .A(n61162), .B(n77454), .Y(n77362) );
  NOR2xp33_ASAP7_75t_SL U65952 ( .A(n71196), .B(n71195), .Y(n71197) );
  NOR2xp33_ASAP7_75t_SL U65953 ( .A(n71200), .B(n71185), .Y(n71195) );
  NOR2xp33_ASAP7_75t_SL U65954 ( .A(n62479), .B(n62478), .Y(n77295) );
  NOR2xp33_ASAP7_75t_SL U65955 ( .A(n71238), .B(n71239), .Y(n71215) );
  NOR2xp33_ASAP7_75t_SL U65956 ( .A(n71206), .B(n71205), .Y(n71239) );
  NOR2xp33_ASAP7_75t_SL U65957 ( .A(n63738), .B(n63737), .Y(n4138) );
  O2A1O1Ixp5_ASAP7_75t_SL U65958 ( .A1(n76825), .A2(n77260), .B(
        or1200_cpu_or1200_genpc_pcreg_default[7]), .C(n63734), .Y(n63735) );
  AND2x2_ASAP7_75t_SL U65959 ( .A(n4058), .B(n4057), .Y(n77603) );
  NOR2xp33_ASAP7_75t_SL U65960 ( .A(n76605), .B(n76604), .Y(n4089) );
  O2A1O1Ixp5_ASAP7_75t_SL U65961 ( .A1(n61171), .A2(n77260), .B(n61170), .C(
        n76825), .Y(n61172) );
  AND2x2_ASAP7_75t_SL U65962 ( .A(n4062), .B(n4061), .Y(n77600) );
  NOR2xp33_ASAP7_75t_SL U65963 ( .A(n61574), .B(n61573), .Y(n4091) );
  AND2x2_ASAP7_75t_SL U65964 ( .A(n4071), .B(n4070), .Y(n77594) );
  NOR2xp33_ASAP7_75t_SL U65965 ( .A(n76532), .B(n76531), .Y(n4134) );
  NOR2xp33_ASAP7_75t_SL U65966 ( .A(n74960), .B(n74959), .Y(n76530) );
  O2A1O1Ixp5_ASAP7_75t_SL U65967 ( .A1(n1106), .A2(n77260), .B(n74958), .C(
        n74957), .Y(n74959) );
  NOR2xp33_ASAP7_75t_SL U65968 ( .A(or1200_cpu_or1200_except_n116), .B(
        or1200_cpu_or1200_except_n286), .Y(n74950) );
  NOR2xp33_ASAP7_75t_SL U65969 ( .A(n63697), .B(n63696), .Y(n4135) );
  AND2x2_ASAP7_75t_SL U65970 ( .A(n4046), .B(n4045), .Y(n75781) );
  NOR2xp33_ASAP7_75t_SL U65971 ( .A(n58567), .B(n61277), .Y(n4136) );
  AND2x2_ASAP7_75t_SL U65972 ( .A(n4050), .B(n4049), .Y(n76508) );
  XNOR2xp5_ASAP7_75t_SL U65973 ( .A(n61268), .B(n76822), .Y(n61269) );
  NOR2xp33_ASAP7_75t_SL U65974 ( .A(n77274), .B(n77273), .Y(n4090) );
  AND2x2_ASAP7_75t_SL U65975 ( .A(n4067), .B(n4066), .Y(n77597) );
  NOR2xp33_ASAP7_75t_SL U65976 ( .A(n71389), .B(n71404), .Y(n71406) );
  XNOR2xp5_ASAP7_75t_SL U65977 ( .A(n75984), .B(n59514), .Y(n75985) );
  XOR2xp5_ASAP7_75t_SL U65978 ( .A(n76177), .B(n76176), .Y(n76178) );
  NOR2xp33_ASAP7_75t_SL U65979 ( .A(n76843), .B(n58560), .Y(n78059) );
  AND2x2_ASAP7_75t_SL U65980 ( .A(n4054), .B(n4053), .Y(n76828) );
  OR2x2_ASAP7_75t_SL U65981 ( .A(n61168), .B(n61577), .Y(n77251) );
  NAND2xp33_ASAP7_75t_SRAM U65982 ( .A(n60459), .B(n77456), .Y(n61036) );
  NOR2xp33_ASAP7_75t_SL U65983 ( .A(n70611), .B(n70610), .Y(n70612) );
  XNOR2xp5_ASAP7_75t_SL U65984 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_output_o_31_), .Y(
        n70565) );
  NOR2xp33_ASAP7_75t_SL U65985 ( .A(n70564), .B(n70563), .Y(n74285) );
  NAND4xp25_ASAP7_75t_SL U65986 ( .A(n70562), .B(n70561), .C(n70560), .D(
        n70559), .Y(n70563) );
  NOR4xp25_ASAP7_75t_SL U65987 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_23_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_16_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_15_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_13_), .Y(
        n70559) );
  NOR4xp25_ASAP7_75t_SL U65988 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_1_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_0_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_24_), .Y(
        n70560) );
  NOR4xp25_ASAP7_75t_SL U65989 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_6_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_5_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_4_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_3_), .Y(
        n70561) );
  NOR4xp25_ASAP7_75t_SL U65990 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_14_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_9_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_8_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_7_), .Y(
        n70562) );
  NAND4xp25_ASAP7_75t_SL U65991 ( .A(n70558), .B(n70557), .C(n70556), .D(
        n70555), .Y(n70564) );
  NOR3xp33_ASAP7_75t_SL U65992 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_10_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_0_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_1_), .Y(
        n70555) );
  NOR2xp33_ASAP7_75t_SL U65993 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_12_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_11_), .Y(
        n70556) );
  NOR4xp25_ASAP7_75t_SL U65994 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_20_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_19_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_18_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_17_), .Y(
        n70557) );
  NOR4xp25_ASAP7_75t_SL U65995 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_26_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_25_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_22_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_rmndr_i_21_), .Y(
        n70558) );
  NOR2xp33_ASAP7_75t_SL U65996 ( .A(n71342), .B(n71345), .Y(n71392) );
  NOR2xp33_ASAP7_75t_SL U65997 ( .A(n71367), .B(n71368), .Y(n71345) );
  NOR2xp33_ASAP7_75t_SL U65998 ( .A(n71297), .B(n71296), .Y(n71298) );
  NOR2xp33_ASAP7_75t_SL U65999 ( .A(n78226), .B(n71145), .Y(n71155) );
  NOR2xp33_ASAP7_75t_SL U66000 ( .A(n78225), .B(n71184), .Y(n71200) );
  NOR2xp33_ASAP7_75t_SL U66001 ( .A(n71083), .B(n71082), .Y(n71153) );
  NOR2xp33_ASAP7_75t_SL U66002 ( .A(n71048), .B(n71047), .Y(n71061) );
  NOR2xp33_ASAP7_75t_SL U66003 ( .A(n71071), .B(n71072), .Y(n71083) );
  NOR2xp33_ASAP7_75t_SL U66004 ( .A(n78400), .B(n71413), .Y(n71071) );
  NOR2xp33_ASAP7_75t_SL U66005 ( .A(n71095), .B(n71094), .Y(n71113) );
  NOR2xp33_ASAP7_75t_SL U66006 ( .A(n78399), .B(n71413), .Y(n71095) );
  NOR2xp33_ASAP7_75t_SL U66007 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_27_), .B(n71084), 
        .Y(n71136) );
  NOR2xp33_ASAP7_75t_SL U66008 ( .A(n78411), .B(n71413), .Y(n70855) );
  NOR2xp33_ASAP7_75t_SL U66009 ( .A(n70797), .B(n70796), .Y(n70798) );
  NOR2xp33_ASAP7_75t_SL U66010 ( .A(n70757), .B(n70756), .Y(n70800) );
  NOR2xp33_ASAP7_75t_SL U66011 ( .A(n78419), .B(n71413), .Y(n70754) );
  NOR2xp33_ASAP7_75t_SL U66012 ( .A(n70698), .B(n70699), .Y(n70712) );
  NOR2xp33_ASAP7_75t_SL U66013 ( .A(n70697), .B(n70696), .Y(n70700) );
  XNOR2xp5_ASAP7_75t_SL U66014 ( .A(n70701), .B(n70702), .Y(n70703) );
  O2A1O1Ixp5_ASAP7_75t_SL U66015 ( .A1(n70737), .A2(n70705), .B(n70692), .C(
        n57115), .Y(n70693) );
  NOR2xp33_ASAP7_75t_SL U66016 ( .A(n70750), .B(n70749), .Y(n70804) );
  NOR2xp33_ASAP7_75t_SL U66017 ( .A(n70728), .B(n70727), .Y(n70750) );
  NOR2xp33_ASAP7_75t_SL U66018 ( .A(n78422), .B(n71413), .Y(n70726) );
  NOR2xp33_ASAP7_75t_SL U66019 ( .A(n70782), .B(n70781), .Y(n70816) );
  NOR2xp33_ASAP7_75t_SL U66020 ( .A(n70792), .B(n70793), .Y(n70817) );
  NOR2xp33_ASAP7_75t_SL U66021 ( .A(n78415), .B(n71413), .Y(n70792) );
  NOR2xp33_ASAP7_75t_SL U66022 ( .A(n78416), .B(n71413), .Y(n70782) );
  NOR2xp33_ASAP7_75t_SL U66023 ( .A(n70770), .B(n70769), .Y(n70773) );
  NOR2xp33_ASAP7_75t_SL U66024 ( .A(n53473), .B(n70896), .Y(n70777) );
  NOR2xp33_ASAP7_75t_SL U66025 ( .A(n78414), .B(n71413), .Y(n70815) );
  NOR2xp33_ASAP7_75t_SL U66026 ( .A(n70858), .B(n70857), .Y(n70875) );
  NOR2xp33_ASAP7_75t_SL U66027 ( .A(n70832), .B(n70831), .Y(n70857) );
  NOR2xp33_ASAP7_75t_SL U66028 ( .A(n78413), .B(n71413), .Y(n70829) );
  NOR2xp33_ASAP7_75t_SL U66029 ( .A(n78412), .B(n71413), .Y(n70847) );
  NAND4xp25_ASAP7_75t_SL U66030 ( .A(n70975), .B(n70968), .C(n70967), .D(
        n70966), .Y(n71032) );
  NOR2xp33_ASAP7_75t_SL U66031 ( .A(n70965), .B(n70971), .Y(n70968) );
  NOR2xp33_ASAP7_75t_SL U66032 ( .A(n70959), .B(n70958), .Y(n70971) );
  NOR2xp33_ASAP7_75t_SL U66033 ( .A(n70918), .B(n70919), .Y(n70937) );
  NOR2xp33_ASAP7_75t_SL U66034 ( .A(n78407), .B(n71413), .Y(n70918) );
  NOR2xp33_ASAP7_75t_SL U66035 ( .A(n70905), .B(n70904), .Y(n70969) );
  NOR2xp33_ASAP7_75t_SL U66036 ( .A(n78406), .B(n71413), .Y(n70935) );
  NOR2xp33_ASAP7_75t_SL U66037 ( .A(n70887), .B(n70886), .Y(n70888) );
  NOR2xp33_ASAP7_75t_SL U66038 ( .A(n78405), .B(n71413), .Y(n70959) );
  NOR2xp33_ASAP7_75t_SL U66039 ( .A(n78403), .B(n71413), .Y(n71005) );
  AOI211xp5_ASAP7_75t_SL U66040 ( .A1(n71263), .A2(n71376), .B(n71233), .C(
        n71232), .Y(n71234) );
  NOR2xp33_ASAP7_75t_SL U66041 ( .A(n71335), .B(n71230), .Y(n71233) );
  NOR2xp33_ASAP7_75t_SL U66042 ( .A(n71413), .B(n71178), .Y(n71271) );
  NOR2xp33_ASAP7_75t_SL U66043 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_33_), .B(n71166), 
        .Y(n71178) );
  NOR2xp33_ASAP7_75t_SL U66044 ( .A(n71413), .B(n71204), .Y(n71272) );
  NOR2xp33_ASAP7_75t_SL U66045 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_34_), .B(n71183), 
        .Y(n71204) );
  NOR2xp33_ASAP7_75t_SL U66046 ( .A(n70705), .B(n57115), .Y(n70707) );
  NOR2xp33_ASAP7_75t_SL U66047 ( .A(n71293), .B(n71292), .Y(n71295) );
  NOR2xp33_ASAP7_75t_SL U66048 ( .A(n71144), .B(n71143), .Y(n71145) );
  NOR2xp33_ASAP7_75t_SL U66049 ( .A(n53473), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .Y(n59522) );
  NOR2xp33_ASAP7_75t_SL U66050 ( .A(n53473), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .Y(n70996) );
  NOR2xp33_ASAP7_75t_SL U66051 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_4_), .B(n71015), .Y(
        n71087) );
  NOR2xp33_ASAP7_75t_SL U66052 ( .A(n71251), .B(n71252), .Y(n71293) );
  NOR2xp33_ASAP7_75t_SL U66053 ( .A(n71324), .B(n71343), .Y(n71309) );
  NOR2xp33_ASAP7_75t_SL U66054 ( .A(n71291), .B(n71290), .Y(n71343) );
  NOR2xp33_ASAP7_75t_SL U66055 ( .A(n71289), .B(n71288), .Y(n71324) );
  NOR2xp33_ASAP7_75t_SL U66056 ( .A(n71287), .B(n71286), .Y(n71290) );
  NOR2xp33_ASAP7_75t_SL U66057 ( .A(n70843), .B(n57115), .Y(n70825) );
  NOR2xp33_ASAP7_75t_SL U66058 ( .A(n71340), .B(n71346), .Y(n71327) );
  NOR2xp33_ASAP7_75t_SL U66059 ( .A(n71321), .B(n71320), .Y(n71340) );
  NOR2xp33_ASAP7_75t_SL U66060 ( .A(n70823), .B(n57115), .Y(n70811) );
  NOR2xp33_ASAP7_75t_SL U66061 ( .A(n71413), .B(n71384), .Y(n71390) );
  NOR2xp33_ASAP7_75t_SL U66062 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_45_), .B(n71366), 
        .Y(n71384) );
  OR2x2_ASAP7_75t_SL U66063 ( .A(n59526), .B(n58315), .Y(n71149) );
  NAND4xp25_ASAP7_75t_SL U66064 ( .A(n70679), .B(n71245), .C(n70678), .D(
        n70677), .Y(n70680) );
  NAND3xp33_ASAP7_75t_SL U66065 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_count_0_), .B(n59526), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[19]), .Y(n70678) );
  NOR2xp33_ASAP7_75t_SL U66066 ( .A(n53473), .B(n71314), .Y(n70665) );
  NOR2xp33_ASAP7_75t_SL U66067 ( .A(n58315), .B(n53473), .Y(n70666) );
  NOR2xp33_ASAP7_75t_SL U66068 ( .A(n71314), .B(n71015), .Y(n70667) );
  NOR2xp33_ASAP7_75t_SL U66069 ( .A(n58315), .B(n71015), .Y(n70668) );
  HB1xp67_ASAP7_75t_SL U66070 ( .A(n3351), .Y(n59701) );
  NOR2xp33_ASAP7_75t_SL U66071 ( .A(n57090), .B(n60458), .Y(n77395) );
  NOR2xp33_ASAP7_75t_SL U66072 ( .A(n77841), .B(n60462), .Y(n61040) );
  NOR2xp33_ASAP7_75t_SL U66073 ( .A(n61045), .B(n61044), .Y(n77397) );
  NOR2xp33_ASAP7_75t_SL U66074 ( .A(n77448), .B(n60301), .Y(n60302) );
  INVx1_ASAP7_75t_SL U66075 ( .A(or1200_cpu_or1200_except_n116), .Y(n77448) );
  INVxp33_ASAP7_75t_SRAM U66076 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_4_), .Y(
        n72538) );
  XNOR2xp5_ASAP7_75t_SL U66077 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .B(
        n72547), .Y(n72543) );
  AND2x2_ASAP7_75t_SL U66078 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .Y(
        n72534) );
  NOR2xp33_ASAP7_75t_SL U66079 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .B(
        n72528), .Y(n72535) );
  NOR2xp33_ASAP7_75t_SL U66080 ( .A(n72524), .B(n57203), .Y(n72528) );
  NAND2xp33_ASAP7_75t_SRAM U66081 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_), .Y(
        n72524) );
  INVxp33_ASAP7_75t_SRAM U66082 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_2_), .Y(
        n72527) );
  OAI21xp33_ASAP7_75t_SRAM U66083 ( .A1(n72517), .A2(n74265), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .Y(
        n72518) );
  INVxp33_ASAP7_75t_SRAM U66084 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_1_), .Y(
        n72521) );
  NOR2xp33_ASAP7_75t_SL U66085 ( .A(n61580), .B(n61579), .Y(n77591) );
  NAND2xp33_ASAP7_75t_SRAM U66086 ( .A(n68754), .B(n68753), .Y(n68763) );
  NOR2xp33_ASAP7_75t_SL U66087 ( .A(n68757), .B(n65071), .Y(n68765) );
  INVxp33_ASAP7_75t_SRAM U66088 ( .A(n68758), .Y(n64988) );
  NOR2xp33_ASAP7_75t_SL U66089 ( .A(n68337), .B(n64985), .Y(n68755) );
  INVxp33_ASAP7_75t_SRAM U66090 ( .A(n68345), .Y(n64985) );
  NAND2xp33_ASAP7_75t_SRAM U66091 ( .A(n68756), .B(n58733), .Y(n68757) );
  XNOR2xp5_ASAP7_75t_SL U66092 ( .A(n75998), .B(n75997), .Y(n75999) );
  OAI21xp33_ASAP7_75t_SRAM U66093 ( .A1(n2779), .A2(n77339), .B(n2777), .Y(
        n77506) );
  INVxp33_ASAP7_75t_SRAM U66094 ( .A(n77353), .Y(n77339) );
  O2A1O1Ixp5_ASAP7_75t_SL U66095 ( .A1(n77503), .A2(n77502), .B(n77501), .C(
        n22057), .Y(n77504) );
  INVx1_ASAP7_75t_SL U66096 ( .A(n62153), .Y(n77451) );
  NOR2xp33_ASAP7_75t_SL U66097 ( .A(n60177), .B(n60176), .Y(n74079) );
  NOR2xp33_ASAP7_75t_SL U66098 ( .A(n62477), .B(n1588), .Y(n60176) );
  NOR2xp33_ASAP7_75t_SL U66099 ( .A(n60159), .B(n60158), .Y(n77019) );
  NOR2xp33_ASAP7_75t_SL U66100 ( .A(n60155), .B(n64096), .Y(n78258) );
  NOR2xp33_ASAP7_75t_SL U66101 ( .A(n60136), .B(n60135), .Y(n74984) );
  NOR2xp33_ASAP7_75t_SL U66102 ( .A(n60127), .B(n60126), .Y(n74639) );
  O2A1O1Ixp5_ASAP7_75t_SL U66103 ( .A1(n807), .A2(n59703), .B(n60114), .C(
        n76821), .Y(n60109) );
  O2A1O1Ixp5_ASAP7_75t_SL U66104 ( .A1(n77346), .A2(n60105), .B(n60104), .C(
        n60103), .Y(n60106) );
  OAI21xp33_ASAP7_75t_SRAM U66105 ( .A1(n77429), .A2(
        or1200_cpu_or1200_except_n116), .B(n3426), .Y(n60103) );
  NOR2xp33_ASAP7_75t_SL U66106 ( .A(n60092), .B(n60091), .Y(n77646) );
  INVx1_ASAP7_75t_SL U66107 ( .A(n60317), .Y(n61162) );
  NOR2xp33_ASAP7_75t_SL U66108 ( .A(n60073), .B(n60072), .Y(n75620) );
  NOR2xp33_ASAP7_75t_SL U66109 ( .A(n60062), .B(n60061), .Y(n75431) );
  NOR2xp33_ASAP7_75t_SL U66110 ( .A(n60045), .B(n60044), .Y(n77637) );
  NOR2xp33_ASAP7_75t_SL U66111 ( .A(n823), .B(n63939), .Y(n60156) );
  NOR2xp33_ASAP7_75t_SL U66112 ( .A(n1106), .B(n74954), .Y(n74957) );
  XNOR2xp5_ASAP7_75t_SL U66113 ( .A(n65213), .B(n60171), .Y(n60040) );
  XNOR2xp5_ASAP7_75t_SL U66114 ( .A(n765), .B(icqmem_adr_qmem[28]), .Y(n60189)
         );
  XNOR2xp5_ASAP7_75t_SL U66115 ( .A(n761), .B(icqmem_adr_qmem[29]), .Y(n60190)
         );
  OR2x2_ASAP7_75t_SL U66116 ( .A(n59703), .B(n76821), .Y(n77260) );
  XOR2xp5_ASAP7_75t_SL U66117 ( .A(icqmem_adr_qmem[31]), .B(n753), .Y(n60269)
         );
  NOR2xp33_ASAP7_75t_SL U66118 ( .A(n791), .B(n60147), .Y(n60054) );
  NAND3xp33_ASAP7_75t_SL U66119 ( .A(n59980), .B(n59979), .C(n58544), .Y(
        n60041) );
  AND2x2_ASAP7_75t_SL U66120 ( .A(or1200_cpu_or1200_genpc_pcreg_default[5]), 
        .B(or1200_cpu_or1200_genpc_pcreg_default[2]), .Y(n58544) );
  NOR2xp33_ASAP7_75t_SL U66121 ( .A(n1073), .B(n61167), .Y(n59980) );
  NAND4xp25_ASAP7_75t_SL U66122 ( .A(n59978), .B(n59977), .C(n59976), .D(
        n59975), .Y(n59981) );
  NOR2xp33_ASAP7_75t_SL U66123 ( .A(n819), .B(n59703), .Y(n59975) );
  NOR2xp33_ASAP7_75t_SL U66124 ( .A(n1095), .B(n1084), .Y(n59976) );
  NOR2xp33_ASAP7_75t_SL U66125 ( .A(n823), .B(n815), .Y(n59977) );
  NOR2xp33_ASAP7_75t_SL U66126 ( .A(n847), .B(n1106), .Y(n59978) );
  NOR2xp33_ASAP7_75t_SL U66127 ( .A(n779), .B(n775), .Y(n59985) );
  NOR2xp33_ASAP7_75t_SL U66128 ( .A(n77309), .B(n60287), .Y(n60283) );
  AND2x2_ASAP7_75t_SL U66129 ( .A(n1851), .B(n1849), .Y(n77309) );
  NOR2xp33_ASAP7_75t_SL U66130 ( .A(n76062), .B(n76126), .Y(n76088) );
  NOR2xp33_ASAP7_75t_SL U66131 ( .A(n76061), .B(n76060), .Y(n76126) );
  NOR2xp33_ASAP7_75t_SL U66132 ( .A(n76026), .B(n76025), .Y(n76060) );
  NOR2xp33_ASAP7_75t_SL U66133 ( .A(n58297), .B(n76013), .Y(n76025) );
  AOI211xp5_ASAP7_75t_SL U66134 ( .A1(n76191), .A2(n58962), .B(n75972), .C(
        n75971), .Y(n75975) );
  NOR2xp33_ASAP7_75t_SL U66135 ( .A(n58569), .B(n76185), .Y(n75971) );
  OAI21xp33_ASAP7_75t_SRAM U66136 ( .A1(n59662), .A2(n58569), .B(n76194), .Y(
        n75972) );
  OAI21xp33_ASAP7_75t_SRAM U66137 ( .A1(n75965), .A2(n75964), .B(n59662), .Y(
        n75966) );
  NOR2xp33_ASAP7_75t_SL U66138 ( .A(n76098), .B(n76100), .Y(n75936) );
  NOR2xp33_ASAP7_75t_SL U66139 ( .A(or1200_cpu_or1200_mult_mac_n32), .B(n57310), .Y(n76100) );
  NOR2xp33_ASAP7_75t_SL U66140 ( .A(or1200_cpu_or1200_mult_mac_n30), .B(n59660), .Y(n76098) );
  NAND2xp33_ASAP7_75t_SRAM U66141 ( .A(n75935), .B(n57315), .Y(n76090) );
  NOR2xp33_ASAP7_75t_SL U66142 ( .A(or1200_cpu_or1200_mult_mac_n28), .B(n59653), .Y(n76114) );
  NOR3xp33_ASAP7_75t_SL U66143 ( .A(n76128), .B(n76132), .C(n76122), .Y(n76138) );
  NOR2xp33_ASAP7_75t_SL U66144 ( .A(or1200_cpu_or1200_mult_mac_n26), .B(n59459), .Y(n76122) );
  NOR2xp33_ASAP7_75t_SL U66145 ( .A(n76061), .B(n76089), .Y(n75932) );
  NOR2xp33_ASAP7_75t_SL U66146 ( .A(n76027), .B(n76031), .Y(n76040) );
  NOR2xp33_ASAP7_75t_SL U66147 ( .A(or1200_cpu_or1200_mult_mac_n48), .B(n76028), .Y(n76031) );
  NOR2xp33_ASAP7_75t_SL U66148 ( .A(or1200_cpu_or1200_mult_mac_n50), .B(n75930), .Y(n76027) );
  NOR2xp33_ASAP7_75t_SL U66149 ( .A(n76019), .B(n76021), .Y(n75929) );
  XNOR2xp5_ASAP7_75t_SL U66150 ( .A(or1200_cpu_or1200_mult_mac_n50), .B(n75930), .Y(n76021) );
  NOR2xp33_ASAP7_75t_SL U66151 ( .A(n75928), .B(n75927), .Y(n76019) );
  NOR2xp33_ASAP7_75t_SL U66152 ( .A(n75926), .B(n76003), .Y(n76011) );
  XNOR2xp5_ASAP7_75t_SL U66153 ( .A(or1200_cpu_or1200_mult_mac_n52), .B(n75927), .Y(n76008) );
  AOI211xp5_ASAP7_75t_SL U66154 ( .A1(n76125), .A2(n76062), .B(n76087), .C(
        n75914), .Y(n76124) );
  NOR2xp33_ASAP7_75t_SL U66155 ( .A(n76085), .B(n75912), .Y(n76097) );
  AOI21xp33_ASAP7_75t_SRAM U66156 ( .A1(n59041), .A2(
        or1200_cpu_or1200_mult_mac_n34), .B(n76081), .Y(n75910) );
  NOR2xp33_ASAP7_75t_SL U66157 ( .A(n76069), .B(n75907), .Y(n76075) );
  NOR2xp33_ASAP7_75t_SL U66158 ( .A(n76058), .B(n76057), .Y(n76069) );
  AO21x1_ASAP7_75t_SL U66159 ( .A1(n76041), .A2(n75931), .B(n75905), .Y(n76062) );
  OAI21xp33_ASAP7_75t_SRAM U66160 ( .A1(n76045), .A2(n59510), .B(n76048), .Y(
        n75905) );
  NAND2xp33_ASAP7_75t_SRAM U66161 ( .A(or1200_cpu_or1200_mult_mac_n44), .B(
        n75904), .Y(n76048) );
  NOR2xp33_ASAP7_75t_SL U66162 ( .A(n76047), .B(n76042), .Y(n75931) );
  NOR2xp33_ASAP7_75t_SL U66163 ( .A(or1200_cpu_or1200_mult_mac_n44), .B(n75904), .Y(n76047) );
  NOR2xp33_ASAP7_75t_SL U66164 ( .A(n75902), .B(n75901), .Y(n76034) );
  NOR2xp33_ASAP7_75t_SL U66165 ( .A(n76023), .B(n57169), .Y(n76033) );
  AOI21xp33_ASAP7_75t_SRAM U66166 ( .A1(or1200_cpu_or1200_mult_mac_n16), .A2(
        n59651), .B(n76159), .Y(n75898) );
  AND2x2_ASAP7_75t_SL U66167 ( .A(or1200_cpu_or1200_mult_mac_n18), .B(n59648), 
        .Y(n76159) );
  NOR2xp33_ASAP7_75t_SL U66168 ( .A(or1200_cpu_or1200_mult_mac_n20), .B(n58753), .Y(n76151) );
  NOR2xp33_ASAP7_75t_SL U66169 ( .A(or1200_cpu_or1200_mult_mac_n18), .B(n59647), .Y(n76149) );
  NAND2xp33_ASAP7_75t_SRAM U66170 ( .A(or1200_cpu_or1200_mult_mac_n20), .B(
        n58753), .Y(n76147) );
  XNOR2xp5_ASAP7_75t_SL U66171 ( .A(or1200_cpu_or1200_mult_mac_n22), .B(n57394), .Y(n76132) );
  NOR2xp33_ASAP7_75t_SL U66172 ( .A(n76129), .B(n57311), .Y(n75896) );
  NOR2xp33_ASAP7_75t_SL U66173 ( .A(or1200_cpu_or1200_mult_mac_n16), .B(n57325), .Y(n75941) );
  NOR2xp33_ASAP7_75t_SL U66174 ( .A(n75957), .B(n53310), .Y(n75948) );
  XNOR2xp5_ASAP7_75t_SL U66175 ( .A(n75924), .B(n59504), .Y(n75998) );
  NOR2xp33_ASAP7_75t_SL U66176 ( .A(or1200_cpu_or1200_mult_mac_n58), .B(n58701), .Y(n75994) );
  NOR2xp33_ASAP7_75t_SL U66177 ( .A(n76005), .B(n58431), .Y(n76009) );
  NOR2xp33_ASAP7_75t_SL U66178 ( .A(n63245), .B(n75760), .Y(n63247) );
  NAND2xp33_ASAP7_75t_SRAM U66179 ( .A(n59550), .B(n66249), .Y(n78170) );
  NOR2xp33_ASAP7_75t_SL U66180 ( .A(or1200_cpu_or1200_mult_mac_div_cntr_4_), 
        .B(n61812), .Y(n75759) );
  NOR2xp33_ASAP7_75t_SL U66181 ( .A(or1200_cpu_or1200_mult_mac_div_cntr_1_), 
        .B(or1200_cpu_or1200_mult_mac_div_cntr_0_), .Y(n61811) );
  NAND2xp33_ASAP7_75t_SRAM U66182 ( .A(n68836), .B(n68852), .Y(n68829) );
  NOR2xp33_ASAP7_75t_SL U66183 ( .A(n77956), .B(n77955), .Y(n77961) );
  OAI22xp33_ASAP7_75t_SRAM U66184 ( .A1(or1200_ic_top_from_icram[16]), .A2(
        n77954), .B1(or1200_cpu_or1200_if_insn_saved[16]), .B2(n78009), .Y(
        n77955) );
  NOR2xp33_ASAP7_75t_SL U66185 ( .A(n60515), .B(n60514), .Y(n77947) );
  NOR2xp33_ASAP7_75t_SL U66186 ( .A(n60522), .B(n60521), .Y(n77938) );
  AND2x2_ASAP7_75t_SL U66187 ( .A(n77842), .B(n59686), .Y(n77952) );
  NOR2xp33_ASAP7_75t_SL U66188 ( .A(n77424), .B(n78006), .Y(n60451) );
  XNOR2xp5_ASAP7_75t_SL U66189 ( .A(n60293), .B(n60292), .Y(n78067) );
  INVx1_ASAP7_75t_SL U66190 ( .A(n22057), .Y(n77833) );
  NOR2xp33_ASAP7_75t_SL U66191 ( .A(n77432), .B(n77436), .Y(n62153) );
  INVx1_ASAP7_75t_SL U66192 ( .A(or1200_cpu_or1200_except_n288), .Y(n77432) );
  NOR4xp25_ASAP7_75t_SL U66193 ( .A(n63767), .B(n76227), .C(pic_ints_i[1]), 
        .D(pic_ints_i[0]), .Y(n60256) );
  NOR2xp33_ASAP7_75t_SL U66194 ( .A(n60255), .B(n1366), .Y(n76227) );
  AND2x2_ASAP7_75t_SL U66195 ( .A(pic_ints_i[19]), .B(or1200_pic_picmr_19_), 
        .Y(n63767) );
  NOR4xp25_ASAP7_75t_SL U66196 ( .A(n77010), .B(n74973), .C(n76610), .D(n76635), .Y(n60257) );
  NOR2xp33_ASAP7_75t_SL U66197 ( .A(n60254), .B(n1396), .Y(n76635) );
  NOR2xp33_ASAP7_75t_SL U66198 ( .A(n60253), .B(n1404), .Y(n76610) );
  NOR2xp33_ASAP7_75t_SL U66199 ( .A(n60252), .B(n1358), .Y(n74973) );
  NOR2xp33_ASAP7_75t_SL U66200 ( .A(n60251), .B(n1374), .Y(n77010) );
  NOR4xp25_ASAP7_75t_SL U66201 ( .A(n77207), .B(n77286), .C(n75773), .D(n76993), .Y(n60258) );
  NOR2xp33_ASAP7_75t_SL U66202 ( .A(n60250), .B(n1412), .Y(n76993) );
  NOR2xp33_ASAP7_75t_SL U66203 ( .A(n60249), .B(n1388), .Y(n75773) );
  NOR2xp33_ASAP7_75t_SL U66204 ( .A(n60248), .B(n1382), .Y(n77286) );
  NOR2xp33_ASAP7_75t_SL U66205 ( .A(n60247), .B(n1378), .Y(n77207) );
  NOR4xp25_ASAP7_75t_SL U66206 ( .A(n76545), .B(n76243), .C(n63255), .D(n76694), .Y(n60245) );
  NOR2xp33_ASAP7_75t_SL U66207 ( .A(n60244), .B(n1400), .Y(n76694) );
  NOR2xp33_ASAP7_75t_SL U66208 ( .A(n60243), .B(n1362), .Y(n63255) );
  NOR2xp33_ASAP7_75t_SL U66209 ( .A(n60242), .B(n1392), .Y(n76243) );
  NOR2xp33_ASAP7_75t_SL U66210 ( .A(n60241), .B(n1384), .Y(n76545) );
  NOR4xp25_ASAP7_75t_SL U66211 ( .A(n76856), .B(n77141), .C(n76687), .D(n76197), .Y(n60246) );
  NOR2xp33_ASAP7_75t_SL U66212 ( .A(n60240), .B(n1408), .Y(n76197) );
  NOR2xp33_ASAP7_75t_SL U66213 ( .A(n60239), .B(n1420), .Y(n76687) );
  NOR2xp33_ASAP7_75t_SL U66214 ( .A(n60238), .B(n1370), .Y(n77141) );
  NOR2xp33_ASAP7_75t_SL U66215 ( .A(n60237), .B(n1416), .Y(n76856) );
  AOI31xp33_ASAP7_75t_SL U66216 ( .A1(n60235), .A2(n58588), .A3(n60236), .B(
        n1717), .Y(n76544) );
  AND2x2_ASAP7_75t_SL U66217 ( .A(n3141), .B(n1536), .Y(n58588) );
  NOR2xp33_ASAP7_75t_SL U66218 ( .A(n61381), .B(n75767), .Y(n74937) );
  NOR2xp33_ASAP7_75t_SL U66219 ( .A(n60818), .B(n64207), .Y(n60227) );
  NOR2xp33_ASAP7_75t_SL U66220 ( .A(n60224), .B(n60223), .Y(n61064) );
  AO21x1_ASAP7_75t_SL U66221 ( .A1(n76492), .A2(n76327), .B(n62002), .Y(n76498) );
  NOR2xp33_ASAP7_75t_SL U66222 ( .A(n75518), .B(n76751), .Y(n75522) );
  NOR2xp33_ASAP7_75t_SL U66223 ( .A(n60222), .B(n76538), .Y(n62149) );
  NOR2xp33_ASAP7_75t_SL U66224 ( .A(n61133), .B(n59970), .Y(n59971) );
  NOR2xp33_ASAP7_75t_SL U66225 ( .A(n59969), .B(n75687), .Y(n59970) );
  NOR2xp33_ASAP7_75t_SL U66226 ( .A(n77623), .B(n64208), .Y(n59969) );
  INVx1_ASAP7_75t_SL U66227 ( .A(n77994), .Y(n61133) );
  NOR2xp33_ASAP7_75t_SL U66228 ( .A(n69368), .B(n60218), .Y(n74926) );
  NOR2xp33_ASAP7_75t_SL U66229 ( .A(n1753), .B(n62237), .Y(n69368) );
  NOR2xp33_ASAP7_75t_SL U66230 ( .A(n60208), .B(n3100), .Y(n77418) );
  XNOR2xp5_ASAP7_75t_SL U66231 ( .A(n3375), .B(n3095), .Y(n60209) );
  INVx1_ASAP7_75t_SL U66232 ( .A(or1200_cpu_or1200_except_n567), .Y(n77208) );
  NAND2xp33_ASAP7_75t_SRAM U66233 ( .A(n59822), .B(n59922), .Y(n59826) );
  INVxp33_ASAP7_75t_SRAM U66234 ( .A(or1200_dc_top_tag_3_), .Y(n59822) );
  NOR2xp33_ASAP7_75t_SL U66235 ( .A(or1200_dc_top_tag_11_), .B(n74041), .Y(
        n59807) );
  XNOR2xp5_ASAP7_75t_SL U66236 ( .A(or1200_dc_top_tag_13_), .B(n78094), .Y(
        n59800) );
  XNOR2xp5_ASAP7_75t_SL U66237 ( .A(or1200_dc_top_tag_7_), .B(n74574), .Y(
        n59795) );
  NOR2xp33_ASAP7_75t_SL U66238 ( .A(n59794), .B(n59855), .Y(n74574) );
  NOR2xp33_ASAP7_75t_SL U66239 ( .A(n77148), .B(n77150), .Y(n77017) );
  NOR3xp33_ASAP7_75t_SL U66240 ( .A(n59778), .B(n59777), .C(
        or1200_dc_top_tag_19_), .Y(n59776) );
  NOR2xp33_ASAP7_75t_SL U66241 ( .A(or1200_dc_top_tag_18_), .B(n60291), .Y(
        n59778) );
  XOR2xp5_ASAP7_75t_SL U66242 ( .A(n59574), .B(n1879), .Y(n59774) );
  NOR2xp33_ASAP7_75t_SL U66243 ( .A(or1200_dc_top_tag_15_), .B(n75190), .Y(
        n59773) );
  XOR2xp5_ASAP7_75t_SL U66244 ( .A(n59528), .B(n1882), .Y(n59763) );
  NOR2xp33_ASAP7_75t_SL U66245 ( .A(n75188), .B(n69366), .Y(n69365) );
  NOR2xp33_ASAP7_75t_SL U66246 ( .A(n75189), .B(n75190), .Y(n75793) );
  AO21x1_ASAP7_75t_SL U66247 ( .A1(n59748), .A2(n59870), .B(n59871), .Y(n59750) );
  NOR2xp33_ASAP7_75t_SL U66248 ( .A(n59787), .B(n75424), .Y(n74125) );
  XOR2xp5_ASAP7_75t_SL U66249 ( .A(n57377), .B(n1891), .Y(n59758) );
  NOR2xp33_ASAP7_75t_SL U66250 ( .A(or1200_dc_top_tag_7_), .B(n59855), .Y(
        n59747) );
  XNOR2xp5_ASAP7_75t_SL U66251 ( .A(or1200_dc_top_tag_17_), .B(n75192), .Y(
        n59738) );
  NOR2xp33_ASAP7_75t_SL U66252 ( .A(n74121), .B(n74981), .Y(n75300) );
  NOR2xp33_ASAP7_75t_SL U66253 ( .A(n76546), .B(n59845), .Y(n59725) );
  NOR2xp33_ASAP7_75t_SL U66254 ( .A(n78166), .B(n59885), .Y(n60582) );
  NOR2xp33_ASAP7_75t_SL U66255 ( .A(n78166), .B(n59891), .Y(n78001) );
  NOR2xp33_ASAP7_75t_SL U66256 ( .A(n3086), .B(n77481), .Y(n61285) );
  INVx1_ASAP7_75t_SL U66257 ( .A(n3090), .Y(n77481) );
  XNOR2xp5_ASAP7_75t_SL U66258 ( .A(n3097), .B(n3376), .Y(n59876) );
  NOR2xp33_ASAP7_75t_SL U66259 ( .A(n59953), .B(n59952), .Y(n77304) );
  XOR2xp5_ASAP7_75t_SL U66260 ( .A(n2763), .B(n2765), .Y(n59952) );
  AOI31xp33_ASAP7_75t_SL U66261 ( .A1(n77758), .A2(n3076), .A3(n2607), .B(
        n77460), .Y(n60191) );
  AND2x2_ASAP7_75t_SL U66262 ( .A(n3423), .B(n2569), .Y(n77758) );
  NOR2xp33_ASAP7_75t_SL U66263 ( .A(n59871), .B(n75195), .Y(n59873) );
  NOR2xp33_ASAP7_75t_SL U66264 ( .A(n1918), .B(n59575), .Y(n59871) );
  NOR2xp33_ASAP7_75t_SL U66265 ( .A(n69356), .B(n74041), .Y(n75618) );
  AOI211xp5_ASAP7_75t_SL U66266 ( .A1(n74041), .A2(n74043), .B(n59864), .C(
        n69361), .Y(n78090) );
  NAND2xp33_ASAP7_75t_SRAM U66267 ( .A(n1912), .B(n59529), .Y(n59799) );
  NOR2xp33_ASAP7_75t_SL U66268 ( .A(n69357), .B(n59864), .Y(n74043) );
  AOI211xp5_ASAP7_75t_SL U66269 ( .A1(n59861), .A2(n75426), .B(n75439), .C(
        n75440), .Y(n59862) );
  NOR2xp33_ASAP7_75t_SL U66270 ( .A(n59858), .B(n74124), .Y(n59859) );
  AOI31xp33_ASAP7_75t_SL U66271 ( .A1(n59857), .A2(n74122), .A3(n59856), .B(
        n59855), .Y(n74124) );
  NOR2xp33_ASAP7_75t_SL U66272 ( .A(n1900), .B(n59535), .Y(n74121) );
  NAND2xp33_ASAP7_75t_SRAM U66273 ( .A(n74118), .B(n59851), .Y(n59853) );
  AOI21xp33_ASAP7_75t_SRAM U66274 ( .A1(n59922), .A2(n77148), .B(n59850), .Y(
        n74119) );
  NOR2xp33_ASAP7_75t_SL U66275 ( .A(n59715), .B(n76206), .Y(n76615) );
  INVxp33_ASAP7_75t_SRAM U66276 ( .A(n76199), .Y(n59715) );
  NOR2xp33_ASAP7_75t_SL U66277 ( .A(n76205), .B(n76611), .Y(n76860) );
  NOR2xp33_ASAP7_75t_SL U66278 ( .A(n76682), .B(n76683), .Y(n76861) );
  NOR2xp33_ASAP7_75t_SL U66279 ( .A(n59714), .B(n76613), .Y(n59719) );
  NOR2xp33_ASAP7_75t_SL U66280 ( .A(n59934), .B(n76638), .Y(n59716) );
  NOR2xp33_ASAP7_75t_SL U66281 ( .A(n59724), .B(n59723), .Y(n59845) );
  NOR2xp33_ASAP7_75t_SL U66282 ( .A(n75779), .B(n76548), .Y(n59724) );
  NOR2xp33_ASAP7_75t_SL U66283 ( .A(n76550), .B(n59721), .Y(n59722) );
  NOR2xp33_ASAP7_75t_SL U66284 ( .A(n59860), .B(n74120), .Y(n75425) );
  NOR2xp33_ASAP7_75t_SL U66285 ( .A(n59842), .B(n59844), .Y(n74120) );
  NOR2xp33_ASAP7_75t_SL U66286 ( .A(n77015), .B(n59841), .Y(n59844) );
  NAND2xp33_ASAP7_75t_SRAM U66287 ( .A(n59922), .B(n59926), .Y(n59841) );
  NAND2xp33_ASAP7_75t_SRAM U66288 ( .A(n77011), .B(n59945), .Y(n59840) );
  NAND4xp25_ASAP7_75t_SL U66289 ( .A(n76229), .B(n59854), .C(n59851), .D(
        n75299), .Y(n59860) );
  NOR2xp33_ASAP7_75t_SL U66290 ( .A(n74118), .B(n59821), .Y(n76229) );
  NOR2xp33_ASAP7_75t_SL U66291 ( .A(n59839), .B(n75424), .Y(n59861) );
  NOR2xp33_ASAP7_75t_SL U66292 ( .A(n1936), .B(n1117), .Y(n75763) );
  NOR2xp33_ASAP7_75t_SL U66293 ( .A(n60307), .B(n69334), .Y(n60422) );
  AO21x1_ASAP7_75t_SL U66294 ( .A1(n60306), .A2(n60305), .B(n77678), .Y(n69334) );
  NAND3xp33_ASAP7_75t_SL U66295 ( .A(n59993), .B(n59961), .C(n2598), .Y(n76657) );
  NOR2xp33_ASAP7_75t_SL U66296 ( .A(n77370), .B(n76844), .Y(n60305) );
  AND2x2_ASAP7_75t_SL U66297 ( .A(n64209), .B(n59965), .Y(n76844) );
  NOR2xp33_ASAP7_75t_SL U66298 ( .A(n62476), .B(n60826), .Y(n59965) );
  NAND3xp33_ASAP7_75t_SL U66299 ( .A(n77853), .B(n77931), .C(n60546), .Y(
        n60557) );
  NOR2xp33_ASAP7_75t_SL U66300 ( .A(n77937), .B(n77851), .Y(n60546) );
  NOR2xp33_ASAP7_75t_SL U66301 ( .A(n59943), .B(n59942), .Y(n77851) );
  NOR2xp33_ASAP7_75t_SL U66302 ( .A(n59940), .B(n59939), .Y(n77937) );
  NOR2xp33_ASAP7_75t_SL U66303 ( .A(n59938), .B(n59937), .Y(n77931) );
  NOR2xp33_ASAP7_75t_SL U66304 ( .A(n60545), .B(n59936), .Y(n77853) );
  NOR2xp33_ASAP7_75t_SL U66305 ( .A(n59924), .B(n59923), .Y(n64282) );
  NOR2xp33_ASAP7_75t_SL U66306 ( .A(n59993), .B(n75475), .Y(n59991) );
  INVx1_ASAP7_75t_SL U66307 ( .A(n77210), .Y(n75475) );
  OAI31xp33_ASAP7_75t_SL U66308 ( .A1(n2598), .A2(n3123), .A3(n2691), .B(
        n59957), .Y(n59990) );
  AOI31xp33_ASAP7_75t_SL U66309 ( .A1(or1200_cpu_or1200_except_n292), .A2(
        or1200_cpu_or1200_except_n286), .A3(or1200_cpu_except_type_1_), .B(
        or1200_cpu_or1200_except_n116), .Y(n59955) );
  NOR2xp33_ASAP7_75t_SL U66310 ( .A(n2970), .B(n2598), .Y(n59956) );
  AOI31xp33_ASAP7_75t_SL U66311 ( .A1(n77425), .A2(n77427), .A3(n59960), .B(
        n77677), .Y(n60306) );
  NOR2xp33_ASAP7_75t_SL U66312 ( .A(n76672), .B(n59959), .Y(n77677) );
  NOR2xp33_ASAP7_75t_SL U66313 ( .A(n2657), .B(n62024), .Y(n59960) );
  NOR2xp33_ASAP7_75t_SL U66314 ( .A(n2609), .B(n59958), .Y(n77425) );
  NOR3xp33_ASAP7_75t_SL U66315 ( .A(n60304), .B(n2693), .C(n2972), .Y(n60307)
         );
  NOR2xp33_ASAP7_75t_SL U66316 ( .A(n59951), .B(n60105), .Y(n60311) );
  NOR2xp33_ASAP7_75t_SL U66317 ( .A(n59950), .B(n77348), .Y(n60105) );
  NAND3xp33_ASAP7_75t_SL U66318 ( .A(n59919), .B(n59918), .C(n59917), .Y(
        n77348) );
  NOR4xp25_ASAP7_75t_SL U66319 ( .A(n59916), .B(n59915), .C(n59914), .D(n59913), .Y(n59917) );
  XNOR2xp5_ASAP7_75t_SL U66320 ( .A(or1200_ic_top_tag[19]), .B(n1025), .Y(
        n59913) );
  XNOR2xp5_ASAP7_75t_SL U66321 ( .A(or1200_ic_top_tag[9]), .B(n935), .Y(n59914) );
  XNOR2xp5_ASAP7_75t_SL U66322 ( .A(or1200_ic_top_tag[6]), .B(n908), .Y(n59915) );
  XNOR2xp5_ASAP7_75t_SL U66323 ( .A(or1200_ic_top_tag[7]), .B(n917), .Y(n59916) );
  NOR4xp25_ASAP7_75t_SL U66324 ( .A(n59912), .B(n59911), .C(n59910), .D(n59909), .Y(n59918) );
  XNOR2xp5_ASAP7_75t_SL U66325 ( .A(or1200_ic_top_tag[8]), .B(n926), .Y(n59909) );
  XNOR2xp5_ASAP7_75t_SL U66326 ( .A(or1200_ic_top_tag[15]), .B(n989), .Y(
        n59910) );
  XNOR2xp5_ASAP7_75t_SL U66327 ( .A(or1200_ic_top_tag[14]), .B(n980), .Y(
        n59911) );
  XNOR2xp5_ASAP7_75t_SL U66328 ( .A(or1200_ic_top_tag[2]), .B(n872), .Y(n59912) );
  NOR3xp33_ASAP7_75t_SL U66329 ( .A(n59908), .B(n59907), .C(n59906), .Y(n59919) );
  NAND4xp25_ASAP7_75t_SL U66330 ( .A(n59905), .B(n59904), .C(n59903), .D(
        n59902), .Y(n59906) );
  XOR2xp5_ASAP7_75t_SL U66331 ( .A(n1016), .B(or1200_ic_top_tag[18]), .Y(
        n59902) );
  XOR2xp5_ASAP7_75t_SL U66332 ( .A(n971), .B(or1200_ic_top_tag[13]), .Y(n59903) );
  XOR2xp5_ASAP7_75t_SL U66333 ( .A(n962), .B(or1200_ic_top_tag[12]), .Y(n59904) );
  XOR2xp5_ASAP7_75t_SL U66334 ( .A(n953), .B(or1200_ic_top_tag[11]), .Y(n59905) );
  NAND4xp25_ASAP7_75t_SL U66335 ( .A(n59901), .B(n59900), .C(n59899), .D(
        n59898), .Y(n59907) );
  XOR2xp5_ASAP7_75t_SL U66336 ( .A(n890), .B(or1200_ic_top_tag[4]), .Y(n59898)
         );
  XOR2xp5_ASAP7_75t_SL U66337 ( .A(n998), .B(or1200_ic_top_tag[16]), .Y(n59899) );
  XOR2xp5_ASAP7_75t_SL U66338 ( .A(n944), .B(or1200_ic_top_tag[10]), .Y(n59900) );
  XOR2xp5_ASAP7_75t_SL U66339 ( .A(n899), .B(or1200_ic_top_tag[5]), .Y(n59901)
         );
  NAND4xp25_ASAP7_75t_SL U66340 ( .A(n59897), .B(n59896), .C(n59895), .D(
        or1200_ic_top_tag_v), .Y(n59908) );
  XOR2xp5_ASAP7_75t_SL U66341 ( .A(n863), .B(or1200_ic_top_tag[1]), .Y(n59895)
         );
  XOR2xp5_ASAP7_75t_SL U66342 ( .A(n852), .B(or1200_ic_top_tag[0]), .Y(n59896)
         );
  NOR2xp33_ASAP7_75t_SL U66343 ( .A(n59894), .B(n59893), .Y(n59897) );
  XNOR2xp5_ASAP7_75t_SL U66344 ( .A(or1200_ic_top_tag[3]), .B(n881), .Y(n59893) );
  XNOR2xp5_ASAP7_75t_SL U66345 ( .A(or1200_ic_top_tag[17]), .B(n1007), .Y(
        n59894) );
  NOR2xp33_ASAP7_75t_SL U66346 ( .A(n77349), .B(n77401), .Y(n77345) );
  INVx1_ASAP7_75t_SL U66347 ( .A(n2781), .Y(n77338) );
  NOR2xp33_ASAP7_75t_SL U66348 ( .A(n60102), .B(n22057), .Y(n59951) );
  NOR2xp33_ASAP7_75t_SL U66349 ( .A(n77337), .B(n77401), .Y(n60102) );
  INVx1_ASAP7_75t_SL U66350 ( .A(n2757), .Y(n60421) );
  NOR2xp33_ASAP7_75t_SL U66351 ( .A(n77403), .B(n2773), .Y(n60273) );
  NOR2xp33_ASAP7_75t_SL U66352 ( .A(n58546), .B(n74113), .Y(n58838) );
  NAND2xp33_ASAP7_75t_SRAM U66353 ( .A(n68917), .B(n68916), .Y(n68924) );
  NOR2xp33_ASAP7_75t_SL U66354 ( .A(n74852), .B(n74872), .Y(n74858) );
  NOR2xp33_ASAP7_75t_SL U66355 ( .A(n74216), .B(n74872), .Y(n74867) );
  NOR2xp33_ASAP7_75t_SL U66356 ( .A(n74843), .B(n74872), .Y(n74845) );
  NOR2xp33_ASAP7_75t_SL U66357 ( .A(n74908), .B(n74907), .Y(n74909) );
  NOR2xp33_ASAP7_75t_SL U66358 ( .A(n77171), .B(n74906), .Y(n78189) );
  NAND2xp33_ASAP7_75t_SRAM U66359 ( .A(n52489), .B(n52498), .Y(n74908) );
  NAND2xp33_ASAP7_75t_SRAM U66360 ( .A(n1520), .B(n74889), .Y(n74893) );
  NOR2xp33_ASAP7_75t_SL U66361 ( .A(n74859), .B(n74872), .Y(n74860) );
  XNOR2xp5_ASAP7_75t_SL U66362 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_1_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_0_), .Y(n74053) );
  XNOR2xp5_ASAP7_75t_SL U66363 ( .A(n74181), .B(n74180), .Y(n74183) );
  XOR2xp5_ASAP7_75t_SL U66364 ( .A(n74090), .B(n74089), .Y(n74091) );
  NOR2xp33_ASAP7_75t_SL U66365 ( .A(n66220), .B(n74190), .Y(n74187) );
  NOR2xp33_ASAP7_75t_SL U66366 ( .A(n74158), .B(n66212), .Y(n66213) );
  AND2x2_ASAP7_75t_SL U66367 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_20_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_19_), .Y(n76965)
         );
  AOI31xp33_ASAP7_75t_SL U66368 ( .A1(n66202), .A2(n76976), .A3(n74749), .B(
        n66201), .Y(n74838) );
  NOR2xp33_ASAP7_75t_SL U66369 ( .A(n65538), .B(n65541), .Y(n66199) );
  NOR2xp33_ASAP7_75t_SL U66370 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[10]), .B(n65446), 
        .Y(n65537) );
  NAND4xp25_ASAP7_75t_SL U66371 ( .A(n66193), .B(n66192), .C(n66191), .D(
        n66190), .Y(n66194) );
  NOR2xp33_ASAP7_75t_SL U66372 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[4]), .Y(n66190) );
  NOR3xp33_ASAP7_75t_SL U66373 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[0]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[3]), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .Y(n66191) );
  NOR2xp33_ASAP7_75t_SL U66374 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[1]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[2]), .Y(n66192) );
  NOR2xp33_ASAP7_75t_SL U66375 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[6]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[8]), .Y(n66193) );
  NOR2xp33_ASAP7_75t_SL U66376 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[14]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[13]), .Y(n65447) );
  NOR2xp33_ASAP7_75t_SL U66377 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[15]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[16]), .Y(n65449) );
  NOR2xp33_ASAP7_75t_SL U66378 ( .A(n65425), .B(n65468), .Y(n65469) );
  NOR2xp33_ASAP7_75t_SL U66379 ( .A(n74158), .B(n66216), .Y(n74163) );
  NOR2xp33_ASAP7_75t_SL U66380 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_24_), .B(n66208), .Y(n74745) );
  NOR4xp25_ASAP7_75t_SL U66381 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_12_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_13_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_14_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_15_), .Y(n66173) );
  NOR4xp25_ASAP7_75t_SL U66382 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_8_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_9_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_10_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_11_), .Y(n66174) );
  NOR4xp25_ASAP7_75t_SL U66383 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_4_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_5_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_6_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_7_), .Y(n66171)
         );
  NOR4xp25_ASAP7_75t_SL U66384 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_0_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_1_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_2_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_3_), .Y(n66172)
         );
  NOR4xp25_ASAP7_75t_SL U66385 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_20_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_21_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_22_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_23_), .Y(n66169) );
  NOR4xp25_ASAP7_75t_SL U66386 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_16_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_17_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_18_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_19_), .Y(n66170) );
  NAND3xp33_ASAP7_75t_SL U66387 ( .A(n74884), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_13_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_14_), .Y(n74887)
         );
  AND2x2_ASAP7_75t_SL U66388 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_9_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_8_), .Y(n76942)
         );
  NOR2xp33_ASAP7_75t_SL U66389 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]), .B(n74749), .Y(
        n74213) );
  NOR2xp33_ASAP7_75t_SL U66390 ( .A(n74173), .B(n74174), .Y(n74747) );
  NOR2xp33_ASAP7_75t_SL U66391 ( .A(n66207), .B(n74189), .Y(n74166) );
  NAND2xp33_ASAP7_75t_SRAM U66392 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]), .B(n74152), .Y(
        n74155) );
  NOR2xp33_ASAP7_75t_SL U66393 ( .A(n74150), .B(n74149), .Y(n74151) );
  XNOR2xp5_ASAP7_75t_SL U66394 ( .A(n74150), .B(n74148), .Y(n74192) );
  XNOR2xp5_ASAP7_75t_SL U66395 ( .A(n74147), .B(n74146), .Y(n74148) );
  NOR2xp33_ASAP7_75t_SL U66396 ( .A(n66189), .B(n66188), .Y(n74139) );
  NOR2xp33_ASAP7_75t_SL U66397 ( .A(n74137), .B(n66183), .Y(n66187) );
  NOR2xp33_ASAP7_75t_SL U66398 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[2]), .B(n66182), .Y(
        n66183) );
  NOR2xp33_ASAP7_75t_SL U66399 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_2_), .B(n66178), .Y(
        n66186) );
  NOR2xp33_ASAP7_75t_SL U66400 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_1_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_N398), .Y(n66184) );
  NOR2xp33_ASAP7_75t_SL U66401 ( .A(n74135), .B(n74145), .Y(n74141) );
  OAI21xp33_ASAP7_75t_SRAM U66402 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .A2(n74137), .B(
        n74133), .Y(n74135) );
  INVx1_ASAP7_75t_SL U66403 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_0_), .Y(n65487) );
  NOR2xp33_ASAP7_75t_SL U66404 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[2]), .B(n65653), .Y(
        n65529) );
  OR2x2_ASAP7_75t_SL U66405 ( .A(n59562), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]), .Y(n65653) );
  AND4x1_ASAP7_75t_SL U66406 ( .A(n65488), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[0]), .Y(n65525) );
  AOI31xp33_ASAP7_75t_SL U66407 ( .A1(n65493), .A2(n65491), .A3(n65490), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]), .Y(n65526) );
  NOR2xp33_ASAP7_75t_SL U66408 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_inf_d), .B(n65497), .Y(n65533)
         );
  NOR2xp33_ASAP7_75t_SL U66409 ( .A(n76978), .B(n74152), .Y(n65497) );
  NOR2xp33_ASAP7_75t_SL U66410 ( .A(n65496), .B(n74134), .Y(n74152) );
  NOR2xp33_ASAP7_75t_SL U66411 ( .A(n65489), .B(n65506), .Y(n65493) );
  AND2x2_ASAP7_75t_SL U66412 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[3]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .Y(n65495) );
  NOR2xp33_ASAP7_75t_SL U66413 ( .A(n69235), .B(n69231), .Y(n69229) );
  INVxp33_ASAP7_75t_SRAM U66414 ( .A(n68735), .Y(n58855) );
  NOR2xp33_ASAP7_75t_SL U66415 ( .A(n68748), .B(n68734), .Y(n68804) );
  NAND2xp33_ASAP7_75t_SRAM U66416 ( .A(n59063), .B(n59451), .Y(n59062) );
  NAND2xp33_ASAP7_75t_SRAM U66417 ( .A(n69299), .B(n59196), .Y(n69303) );
  NOR2xp33_ASAP7_75t_SL U66418 ( .A(n58485), .B(n69296), .Y(n59214) );
  NOR2xp33_ASAP7_75t_SL U66419 ( .A(n69119), .B(n69118), .Y(n69151) );
  INVxp33_ASAP7_75t_SRAM U66420 ( .A(n59392), .Y(n69155) );
  NOR2xp33_ASAP7_75t_SL U66421 ( .A(n69304), .B(n69301), .Y(n68654) );
  NAND2xp33_ASAP7_75t_SRAM U66422 ( .A(n69012), .B(n68972), .Y(n68984) );
  NOR2xp33_ASAP7_75t_SL U66423 ( .A(n68642), .B(n68645), .Y(n75099) );
  NAND2xp33_ASAP7_75t_SRAM U66424 ( .A(n69026), .B(n69025), .Y(n69045) );
  OAI21xp33_ASAP7_75t_SRAM U66425 ( .A1(n69097), .A2(n69096), .B(n69095), .Y(
        n69101) );
  INVxp33_ASAP7_75t_SRAM U66426 ( .A(n57477), .Y(n68899) );
  HB1xp67_ASAP7_75t_SL U66427 ( .A(n68803), .Y(n59480) );
  NAND2xp33_ASAP7_75t_SRAM U66428 ( .A(n68828), .B(n68827), .Y(n68852) );
  NOR2xp33_ASAP7_75t_SL U66429 ( .A(n58389), .B(n68833), .Y(n68840) );
  INVxp33_ASAP7_75t_SRAM U66430 ( .A(n53199), .Y(n68833) );
  INVxp33_ASAP7_75t_SRAM U66431 ( .A(n74559), .Y(n74560) );
  INVxp33_ASAP7_75t_SRAM U66432 ( .A(n74554), .Y(n74555) );
  OAI21xp33_ASAP7_75t_SRAM U66433 ( .A1(n69116), .A2(n69241), .B(n68687), .Y(
        n68688) );
  INVxp33_ASAP7_75t_SRAM U66434 ( .A(n74557), .Y(n74561) );
  NOR2xp33_ASAP7_75t_SL U66435 ( .A(n68702), .B(n68703), .Y(n68707) );
  NAND2xp33_ASAP7_75t_SRAM U66436 ( .A(n75276), .B(n68694), .Y(n68703) );
  NAND4xp25_ASAP7_75t_SL U66437 ( .A(n68700), .B(n68699), .C(n68698), .D(
        n69102), .Y(n74563) );
  XOR2xp5_ASAP7_75t_SL U66438 ( .A(n75275), .B(n75274), .Y(n75283) );
  NOR2xp33_ASAP7_75t_SL U66439 ( .A(n68695), .B(n59392), .Y(n59391) );
  NOR2xp33_ASAP7_75t_SL U66440 ( .A(n68668), .B(n69235), .Y(n68651) );
  NOR2xp33_ASAP7_75t_SL U66441 ( .A(n68627), .B(n69227), .Y(n68668) );
  NOR2xp33_ASAP7_75t_SL U66442 ( .A(n57062), .B(n68803), .Y(n68564) );
  NOR2xp33_ASAP7_75t_SL U66443 ( .A(n75108), .B(n75107), .Y(n75137) );
  XOR2xp5_ASAP7_75t_SL U66444 ( .A(n66840), .B(n66708), .Y(n66709) );
  XNOR2xp5_ASAP7_75t_SL U66445 ( .A(n67104), .B(n67038), .Y(n67109) );
  XOR2xp5_ASAP7_75t_SL U66446 ( .A(n67105), .B(n67103), .Y(n67038) );
  INVxp33_ASAP7_75t_SRAM U66447 ( .A(n66845), .Y(n66693) );
  XNOR2xp5_ASAP7_75t_SL U66448 ( .A(n66893), .B(n66689), .Y(n66841) );
  INVxp33_ASAP7_75t_SRAM U66449 ( .A(n66988), .Y(n66846) );
  XNOR2xp5_ASAP7_75t_SL U66450 ( .A(n66865), .B(n58459), .Y(n66866) );
  NOR2xp33_ASAP7_75t_SL U66451 ( .A(n66845), .B(n66844), .Y(n66987) );
  XOR2xp5_ASAP7_75t_SL U66452 ( .A(n67101), .B(n67099), .Y(n67010) );
  XNOR2xp5_ASAP7_75t_SL U66453 ( .A(n67037), .B(n67049), .Y(n67103) );
  NOR2xp33_ASAP7_75t_SL U66454 ( .A(n67213), .B(n67214), .Y(n74554) );
  XOR2xp5_ASAP7_75t_SL U66455 ( .A(n66871), .B(n66872), .Y(n66680) );
  NOR2xp33_ASAP7_75t_SL U66456 ( .A(n66887), .B(n66886), .Y(n66890) );
  INVxp33_ASAP7_75t_SRAM U66457 ( .A(n66888), .Y(n66886) );
  XNOR2xp5_ASAP7_75t_SL U66458 ( .A(n67007), .B(n66854), .Y(n66865) );
  INVxp33_ASAP7_75t_SRAM U66459 ( .A(n67099), .Y(n67102) );
  XNOR2xp5_ASAP7_75t_SL U66460 ( .A(n67008), .B(n67052), .Y(n67099) );
  NAND2xp33_ASAP7_75t_SRAM U66461 ( .A(n67154), .B(n67139), .Y(n58678) );
  XNOR2xp5_ASAP7_75t_SL U66462 ( .A(n67168), .B(n67167), .Y(n67206) );
  XNOR2xp5_ASAP7_75t_SL U66463 ( .A(n67058), .B(n59170), .Y(n67052) );
  NOR2xp33_ASAP7_75t_SL U66464 ( .A(n59446), .B(n66678), .Y(n66679) );
  NOR2xp33_ASAP7_75t_SL U66465 ( .A(n59440), .B(n66751), .Y(n59101) );
  NOR2xp33_ASAP7_75t_SL U66466 ( .A(n58521), .B(n68119), .Y(n59103) );
  NOR2xp33_ASAP7_75t_SL U66467 ( .A(n67137), .B(n67136), .Y(n67194) );
  XNOR2xp5_ASAP7_75t_SL U66468 ( .A(n67125), .B(n67124), .Y(n67137) );
  AO21x1_ASAP7_75t_SL U66469 ( .A1(n58681), .A2(n67131), .B(n58680), .Y(n67196) );
  AOI31xp33_ASAP7_75t_SL U66470 ( .A1(n67090), .A2(n67088), .A3(n67089), .B(
        n67087), .Y(n67131) );
  NOR2xp33_ASAP7_75t_SL U66471 ( .A(n67019), .B(n67018), .Y(n67083) );
  OAI22xp33_ASAP7_75t_SRAM U66472 ( .A1(n59200), .A2(n53315), .B1(n67017), 
        .B2(n59668), .Y(n67019) );
  INVxp33_ASAP7_75t_SRAM U66473 ( .A(n67029), .Y(n67032) );
  NOR2xp33_ASAP7_75t_SL U66474 ( .A(n66862), .B(n66861), .Y(n67029) );
  NOR2xp33_ASAP7_75t_SL U66475 ( .A(n67026), .B(n67025), .Y(n67028) );
  AOI21xp33_ASAP7_75t_SRAM U66476 ( .A1(n57336), .A2(n66882), .B(n67566), .Y(
        n66885) );
  INVxp33_ASAP7_75t_SRAM U66477 ( .A(n67023), .Y(n67026) );
  NOR2xp33_ASAP7_75t_SL U66478 ( .A(n67153), .B(n67152), .Y(n67156) );
  AOI21xp33_ASAP7_75t_SRAM U66479 ( .A1(n67593), .A2(n67741), .B(n67092), .Y(
        n67093) );
  XNOR2xp5_ASAP7_75t_SL U66480 ( .A(n59617), .B(n59668), .Y(n67018) );
  AOI21xp33_ASAP7_75t_SRAM U66481 ( .A1(n57277), .A2(n57107), .B(n66996), .Y(
        n66997) );
  NAND2xp33_ASAP7_75t_SRAM U66482 ( .A(n59641), .B(n67911), .Y(n66858) );
  OAI21xp33_ASAP7_75t_SRAM U66483 ( .A1(n67736), .A2(n57505), .B(n66855), .Y(
        n67001) );
  NOR2xp33_ASAP7_75t_SL U66484 ( .A(n68629), .B(n68630), .Y(n69301) );
  XNOR2xp5_ASAP7_75t_SL U66485 ( .A(n66604), .B(n66603), .Y(n68634) );
  XNOR2xp5_ASAP7_75t_SL U66486 ( .A(n66559), .B(n66290), .Y(n66592) );
  XNOR2xp5_ASAP7_75t_SL U66487 ( .A(n66341), .B(n66339), .Y(n66597) );
  NAND2xp33_ASAP7_75t_SRAM U66488 ( .A(n66542), .B(n75048), .Y(n66323) );
  XNOR2xp5_ASAP7_75t_SL U66489 ( .A(n66588), .B(n66587), .Y(n66601) );
  XNOR2xp5_ASAP7_75t_SL U66490 ( .A(n68635), .B(n66584), .Y(n68629) );
  XNOR2xp5_ASAP7_75t_SL U66491 ( .A(n66583), .B(n66582), .Y(n66584) );
  XOR2xp5_ASAP7_75t_SL U66492 ( .A(n59617), .B(n59670), .Y(n66853) );
  XNOR2xp5_ASAP7_75t_SL U66493 ( .A(n66492), .B(n66460), .Y(n67168) );
  NOR2xp33_ASAP7_75t_SL U66494 ( .A(n66278), .B(n66282), .Y(n66394) );
  NOR2xp33_ASAP7_75t_SL U66495 ( .A(n66277), .B(n66276), .Y(n66282) );
  NOR2xp33_ASAP7_75t_SL U66496 ( .A(n66275), .B(n66274), .Y(n66278) );
  OAI21xp33_ASAP7_75t_SRAM U66497 ( .A1(n76176), .A2(n66479), .B(n66247), .Y(
        n66277) );
  AOI22xp33_ASAP7_75t_SRAM U66498 ( .A1(n66281), .A2(n59635), .B1(n66331), 
        .B2(n57067), .Y(n66395) );
  XNOR2xp5_ASAP7_75t_SL U66499 ( .A(n66440), .B(n66439), .Y(n66529) );
  XNOR2xp5_ASAP7_75t_SL U66500 ( .A(n66438), .B(n66437), .Y(n66440) );
  XNOR2xp5_ASAP7_75t_SL U66501 ( .A(n66392), .B(n66391), .Y(n66437) );
  OAI21xp33_ASAP7_75t_SRAM U66502 ( .A1(n75899), .A2(n68603), .B(n66316), .Y(
        n66317) );
  NAND2xp33_ASAP7_75t_SRAM U66503 ( .A(n75899), .B(n68602), .Y(n66316) );
  XNOR2xp5_ASAP7_75t_SL U66504 ( .A(n66507), .B(n66506), .Y(n66514) );
  INVxp33_ASAP7_75t_SRAM U66505 ( .A(n66498), .Y(n66499) );
  XNOR2xp5_ASAP7_75t_SL U66506 ( .A(n59607), .B(n59647), .Y(n67078) );
  XNOR2xp5_ASAP7_75t_SL U66507 ( .A(n59640), .B(n59647), .Y(n66455) );
  INVxp33_ASAP7_75t_SRAM U66508 ( .A(n66484), .Y(n66485) );
  INVxp33_ASAP7_75t_SRAM U66509 ( .A(n58476), .Y(n66487) );
  XNOR2xp5_ASAP7_75t_SL U66510 ( .A(n66512), .B(n66511), .Y(n66527) );
  XNOR2xp5_ASAP7_75t_SL U66511 ( .A(n66363), .B(n66366), .Y(n66511) );
  AOI31xp33_ASAP7_75t_SL U66512 ( .A1(n59447), .A2(n66369), .A3(n66364), .B(
        n66368), .Y(n66363) );
  NAND2xp33_ASAP7_75t_SRAM U66513 ( .A(n59607), .B(n59666), .Y(n66364) );
  NAND2xp33_ASAP7_75t_SRAM U66514 ( .A(n57292), .B(n59664), .Y(n66369) );
  OAI21xp33_ASAP7_75t_SRAM U66515 ( .A1(n59664), .A2(n67074), .B(n66350), .Y(
        n66346) );
  NAND2xp33_ASAP7_75t_SRAM U66516 ( .A(n57163), .B(n66344), .Y(n66349) );
  XNOR2xp5_ASAP7_75t_SL U66517 ( .A(n66521), .B(n66520), .Y(n66525) );
  NAND2xp33_ASAP7_75t_SRAM U66518 ( .A(n59455), .B(n59670), .Y(n58666) );
  INVxp33_ASAP7_75t_SRAM U66519 ( .A(n66656), .Y(n66419) );
  NAND2xp33_ASAP7_75t_SRAM U66520 ( .A(n66414), .B(n75048), .Y(n66415) );
  INVxp33_ASAP7_75t_SRAM U66521 ( .A(n67643), .Y(n66413) );
  XNOR2xp5_ASAP7_75t_SL U66522 ( .A(n59596), .B(n57398), .Y(n66423) );
  XNOR2xp5_ASAP7_75t_SL U66523 ( .A(n59637), .B(n57101), .Y(n66414) );
  AOI21xp33_ASAP7_75t_SRAM U66524 ( .A1(n75899), .A2(n66399), .B(n57292), .Y(
        n66400) );
  OAI21xp33_ASAP7_75t_SRAM U66525 ( .A1(n59662), .A2(n57505), .B(n66396), .Y(
        n66464) );
  NOR2xp33_ASAP7_75t_SL U66526 ( .A(n66268), .B(n66267), .Y(n66281) );
  NOR2xp33_ASAP7_75t_SL U66527 ( .A(n66473), .B(n59491), .Y(n66252) );
  NOR2xp33_ASAP7_75t_SL U66528 ( .A(n66431), .B(n59612), .Y(n66250) );
  XNOR2xp5_ASAP7_75t_SL U66529 ( .A(n57456), .B(n57505), .Y(n66431) );
  XNOR2xp5_ASAP7_75t_SL U66530 ( .A(n66430), .B(n66429), .Y(n66519) );
  XNOR2xp5_ASAP7_75t_SL U66531 ( .A(n66389), .B(n66388), .Y(n66429) );
  NOR2xp33_ASAP7_75t_SL U66532 ( .A(n66386), .B(n66385), .Y(n66389) );
  NOR2xp33_ASAP7_75t_SL U66533 ( .A(n68119), .B(n66537), .Y(n66385) );
  NAND2xp33_ASAP7_75t_SRAM U66534 ( .A(n75641), .B(n59607), .Y(n66384) );
  NAND2xp33_ASAP7_75t_SRAM U66535 ( .A(n57260), .B(n66379), .Y(n66382) );
  NOR2xp33_ASAP7_75t_SL U66536 ( .A(n75055), .B(n68613), .Y(n68615) );
  NOR2xp33_ASAP7_75t_SL U66537 ( .A(n66579), .B(n66578), .Y(n68616) );
  AO21x1_ASAP7_75t_SL U66538 ( .A1(n66577), .A2(n66576), .B(n66575), .Y(n66578) );
  XNOR2xp5_ASAP7_75t_SL U66539 ( .A(n68596), .B(n66573), .Y(n66579) );
  XNOR2xp5_ASAP7_75t_SL U66540 ( .A(n68607), .B(n68595), .Y(n66573) );
  NAND2xp33_ASAP7_75t_SRAM U66541 ( .A(n59639), .B(n53310), .Y(n66570) );
  NAND2xp33_ASAP7_75t_SRAM U66542 ( .A(n59637), .B(n53221), .Y(n66571) );
  NOR2xp33_ASAP7_75t_SL U66543 ( .A(n66582), .B(n66583), .Y(n68636) );
  XNOR2xp5_ASAP7_75t_SL U66544 ( .A(n66544), .B(n66567), .Y(n66582) );
  OAI21xp33_ASAP7_75t_SRAM U66545 ( .A1(n59641), .A2(n75947), .B(n66377), .Y(
        n66537) );
  XNOR2xp5_ASAP7_75t_SL U66546 ( .A(n66574), .B(n66576), .Y(n66583) );
  AOI22xp33_ASAP7_75t_SRAM U66547 ( .A1(n59635), .A2(n66550), .B1(n66572), 
        .B2(n57067), .Y(n66551) );
  OAI21xp33_ASAP7_75t_SRAM U66548 ( .A1(n58015), .A2(n59637), .B(n66541), .Y(
        n66550) );
  NAND2xp33_ASAP7_75t_SRAM U66549 ( .A(n59637), .B(n75899), .Y(n66541) );
  NOR2xp33_ASAP7_75t_SL U66550 ( .A(n66549), .B(n66548), .Y(n66553) );
  OAI22xp33_ASAP7_75t_SRAM U66551 ( .A1(n66546), .A2(n75036), .B1(n58785), 
        .B2(n67365), .Y(n66549) );
  HB1xp67_ASAP7_75t_SL U66552 ( .A(n59144), .Y(n59142) );
  OAI22xp33_ASAP7_75t_SRAM U66553 ( .A1(n66372), .A2(n75076), .B1(n75032), 
        .B2(n66284), .Y(n66559) );
  AOI22xp33_ASAP7_75t_SRAM U66554 ( .A1(n59635), .A2(n66331), .B1(n66542), 
        .B2(n57067), .Y(n66338) );
  OAI21xp33_ASAP7_75t_SRAM U66555 ( .A1(n59638), .A2(n59648), .B(n66279), .Y(
        n66331) );
  NAND2xp33_ASAP7_75t_SRAM U66556 ( .A(n59637), .B(n68104), .Y(n66279) );
  INVxp33_ASAP7_75t_SRAM U66557 ( .A(n63362), .Y(n63021) );
  NOR2xp33_ASAP7_75t_SL U66558 ( .A(n63259), .B(n63260), .Y(n63279) );
  XNOR2xp5_ASAP7_75t_SL U66559 ( .A(n62893), .B(n62886), .Y(n63299) );
  XNOR2xp5_ASAP7_75t_SL U66560 ( .A(n62906), .B(n62884), .Y(n62886) );
  NOR2xp33_ASAP7_75t_SL U66561 ( .A(n62948), .B(n63343), .Y(n63370) );
  XNOR2xp5_ASAP7_75t_SL U66562 ( .A(n62933), .B(n62932), .Y(n62946) );
  XNOR2xp5_ASAP7_75t_SL U66563 ( .A(n62914), .B(n62840), .Y(n63367) );
  XNOR2xp5_ASAP7_75t_SL U66564 ( .A(n62916), .B(n62915), .Y(n62840) );
  XNOR2xp5_ASAP7_75t_SL U66565 ( .A(n62931), .B(n62821), .Y(n62914) );
  XNOR2xp5_ASAP7_75t_SL U66566 ( .A(n62861), .B(n62860), .Y(n63343) );
  XNOR2xp5_ASAP7_75t_SL U66567 ( .A(n63029), .B(n63028), .Y(n63042) );
  XNOR2xp5_ASAP7_75t_SL U66568 ( .A(n63027), .B(n63026), .Y(n63028) );
  XNOR2xp5_ASAP7_75t_SL U66569 ( .A(n62994), .B(n62993), .Y(n62988) );
  XNOR2xp5_ASAP7_75t_SL U66570 ( .A(n62928), .B(n62927), .Y(n62989) );
  NAND2xp33_ASAP7_75t_SRAM U66571 ( .A(n57178), .B(n75925), .Y(n62800) );
  XNOR2xp5_ASAP7_75t_SL U66572 ( .A(n59512), .B(n59503), .Y(n62879) );
  XNOR2xp5_ASAP7_75t_SL U66573 ( .A(n62972), .B(n62945), .Y(n62991) );
  XNOR2xp5_ASAP7_75t_SL U66574 ( .A(n62973), .B(n62944), .Y(n62945) );
  XNOR2xp5_ASAP7_75t_SL U66575 ( .A(n62987), .B(n62986), .Y(n62993) );
  NAND2xp33_ASAP7_75t_SRAM U66576 ( .A(n59514), .B(n59614), .Y(n62835) );
  NAND2xp33_ASAP7_75t_SRAM U66577 ( .A(n76028), .B(n57180), .Y(n62837) );
  AOI31xp33_ASAP7_75t_SL U66578 ( .A1(n64625), .A2(n58481), .A3(n62942), .B(
        n62941), .Y(n62973) );
  OAI21xp33_ASAP7_75t_SRAM U66579 ( .A1(n59418), .A2(n57178), .B(n62814), .Y(
        n62942) );
  XNOR2xp5_ASAP7_75t_SL U66580 ( .A(n63002), .B(n62969), .Y(n62992) );
  XNOR2xp5_ASAP7_75t_SL U66581 ( .A(n63006), .B(n63005), .Y(n63020) );
  OAI21xp33_ASAP7_75t_SRAM U66582 ( .A1(n58431), .A2(n59595), .B(n62918), .Y(
        n62965) );
  NAND2xp33_ASAP7_75t_SRAM U66583 ( .A(n59504), .B(n67231), .Y(n62920) );
  NOR2xp33_ASAP7_75t_SL U66584 ( .A(n62960), .B(n64642), .Y(n62961) );
  NOR2xp33_ASAP7_75t_SL U66585 ( .A(n62957), .B(n57156), .Y(n62962) );
  XNOR2xp5_ASAP7_75t_SL U66586 ( .A(n63001), .B(n63000), .Y(n63022) );
  XNOR2xp5_ASAP7_75t_SL U66587 ( .A(n62999), .B(n62998), .Y(n63000) );
  XNOR2xp5_ASAP7_75t_SL U66588 ( .A(n62997), .B(n62996), .Y(n63001) );
  XNOR2xp5_ASAP7_75t_SL U66589 ( .A(n58984), .B(n58983), .Y(n63043) );
  NAND2xp33_ASAP7_75t_SRAM U66590 ( .A(n67428), .B(n59620), .Y(n62706) );
  XNOR2xp5_ASAP7_75t_SL U66591 ( .A(n62720), .B(n62705), .Y(n63027) );
  NOR2xp33_ASAP7_75t_SL U66592 ( .A(n63161), .B(n63160), .Y(n63878) );
  NOR2xp33_ASAP7_75t_SL U66593 ( .A(n64745), .B(n64744), .Y(n64750) );
  XOR2xp5_ASAP7_75t_SL U66594 ( .A(n63155), .B(n63087), .Y(n58502) );
  O2A1O1Ixp5_ASAP7_75t_SL U66595 ( .A1(n62624), .A2(n62623), .B(n57110), .C(
        n62622), .Y(n62625) );
  O2A1O1Ixp5_ASAP7_75t_SL U66596 ( .A1(n53300), .A2(n62614), .B(n57186), .C(
        n59556), .Y(n62623) );
  OAI22xp33_ASAP7_75t_SRAM U66597 ( .A1(n57159), .A2(n62643), .B1(n62940), 
        .B2(n57097), .Y(n63031) );
  NAND2xp33_ASAP7_75t_SRAM U66598 ( .A(n75930), .B(n57178), .Y(n62633) );
  NAND2xp33_ASAP7_75t_SRAM U66599 ( .A(n59230), .B(n67909), .Y(n59060) );
  NOR2xp33_ASAP7_75t_SL U66600 ( .A(n62597), .B(n59506), .Y(n62664) );
  NOR2xp33_ASAP7_75t_SL U66601 ( .A(n62770), .B(n62769), .Y(n63072) );
  NAND2xp33_ASAP7_75t_SRAM U66602 ( .A(n67481), .B(n62725), .Y(n62768) );
  NAND2xp33_ASAP7_75t_SRAM U66603 ( .A(n57180), .B(n67585), .Y(n62651) );
  XNOR2xp5_ASAP7_75t_SL U66604 ( .A(n62766), .B(n62765), .Y(n63078) );
  INVxp33_ASAP7_75t_SRAM U66605 ( .A(n63088), .Y(n62766) );
  XNOR2xp5_ASAP7_75t_SL U66606 ( .A(n63054), .B(n62753), .Y(n63049) );
  XNOR2xp5_ASAP7_75t_SL U66607 ( .A(n63053), .B(n63052), .Y(n62753) );
  XNOR2xp5_ASAP7_75t_SL U66608 ( .A(n63062), .B(n62747), .Y(n63053) );
  NOR2xp33_ASAP7_75t_SL U66609 ( .A(n62732), .B(n58361), .Y(n62733) );
  NOR2xp33_ASAP7_75t_SL U66610 ( .A(n57111), .B(n59012), .Y(n62719) );
  XNOR2xp5_ASAP7_75t_SL U66611 ( .A(n59602), .B(n59512), .Y(n62728) );
  NAND2xp33_ASAP7_75t_SRAM U66612 ( .A(n67629), .B(n59615), .Y(n62742) );
  XNOR2xp5_ASAP7_75t_SL U66613 ( .A(n63237), .B(n63150), .Y(n63151) );
  OAI21xp33_ASAP7_75t_SRAM U66614 ( .A1(n64710), .A2(n64709), .B(n64718), .Y(
        n64719) );
  NAND2xp33_ASAP7_75t_SRAM U66615 ( .A(n59340), .B(n67428), .Y(n63095) );
  NAND2xp33_ASAP7_75t_SRAM U66616 ( .A(n68087), .B(n67428), .Y(n62758) );
  XNOR2xp5_ASAP7_75t_SL U66617 ( .A(n63119), .B(n63118), .Y(n63198) );
  XNOR2xp5_ASAP7_75t_SL U66618 ( .A(n63627), .B(n63628), .Y(n63195) );
  OAI21xp33_ASAP7_75t_SRAM U66619 ( .A1(n67906), .A2(n63143), .B(n63065), .Y(
        n63158) );
  NAND2xp33_ASAP7_75t_SRAM U66620 ( .A(n59506), .B(n63084), .Y(n63085) );
  NAND2xp33_ASAP7_75t_SRAM U66621 ( .A(n59505), .B(n57169), .Y(n63086) );
  XNOR2xp5_ASAP7_75t_SL U66622 ( .A(n63639), .B(n63211), .Y(n63212) );
  XNOR2xp5_ASAP7_75t_SL U66623 ( .A(n63641), .B(n58825), .Y(n63873) );
  XNOR2xp5_ASAP7_75t_SL U66624 ( .A(n64063), .B(n63870), .Y(n64017) );
  INVxp33_ASAP7_75t_SRAM U66625 ( .A(n63645), .Y(n63649) );
  NAND2xp33_ASAP7_75t_SRAM U66626 ( .A(n75900), .B(n68101), .Y(n63146) );
  NOR2xp33_ASAP7_75t_SL U66627 ( .A(n59338), .B(n58884), .Y(n59337) );
  INVxp33_ASAP7_75t_SRAM U66628 ( .A(n63149), .Y(n59338) );
  NOR2xp33_ASAP7_75t_SL U66629 ( .A(n59514), .B(n58536), .Y(n62724) );
  NAND2xp33_ASAP7_75t_SRAM U66630 ( .A(n53280), .B(n67463), .Y(n63228) );
  NOR2xp33_ASAP7_75t_SL U66631 ( .A(n63112), .B(n63111), .Y(n63232) );
  NOR2xp33_ASAP7_75t_SL U66632 ( .A(n63110), .B(n59460), .Y(n63111) );
  XNOR2xp5_ASAP7_75t_SL U66633 ( .A(n57024), .B(n63680), .Y(n63795) );
  XNOR2xp5_ASAP7_75t_SL U66634 ( .A(n64711), .B(n64066), .Y(n64092) );
  XNOR2xp5_ASAP7_75t_SL U66635 ( .A(n64065), .B(n64722), .Y(n64066) );
  XNOR2xp5_ASAP7_75t_SL U66636 ( .A(n63637), .B(n63834), .Y(n63849) );
  NAND2xp33_ASAP7_75t_SRAM U66637 ( .A(n59660), .B(n57180), .Y(n63208) );
  XNOR2xp5_ASAP7_75t_SL U66638 ( .A(n63868), .B(n63867), .Y(n64057) );
  XNOR2xp5_ASAP7_75t_SL U66639 ( .A(n64054), .B(n63866), .Y(n63867) );
  O2A1O1Ixp5_ASAP7_75t_SL U66640 ( .A1(n57167), .A2(n59614), .B(n63614), .C(
        n68079), .Y(n63615) );
  NAND2xp33_ASAP7_75t_SRAM U66641 ( .A(n59614), .B(n67569), .Y(n63614) );
  NOR2xp33_ASAP7_75t_SL U66642 ( .A(n63222), .B(n63221), .Y(n63620) );
  NAND2xp33_ASAP7_75t_SRAM U66643 ( .A(n59606), .B(n58431), .Y(n63220) );
  NAND2xp33_ASAP7_75t_SRAM U66644 ( .A(n67343), .B(n67963), .Y(n63217) );
  NOR2xp33_ASAP7_75t_SL U66645 ( .A(n63216), .B(n63215), .Y(n63622) );
  NOR2xp33_ASAP7_75t_SL U66646 ( .A(n63214), .B(n59460), .Y(n63215) );
  NOR2xp33_ASAP7_75t_SL U66647 ( .A(n64718), .B(n59369), .Y(n59367) );
  XNOR2xp5_ASAP7_75t_SL U66648 ( .A(n58467), .B(n66977), .Y(n59005) );
  NOR2xp33_ASAP7_75t_SL U66649 ( .A(n66671), .B(n66690), .Y(n66672) );
  AO21x1_ASAP7_75t_SL U66650 ( .A1(n66737), .A2(n66739), .B(n66738), .Y(n66691) );
  INVxp33_ASAP7_75t_SRAM U66651 ( .A(n67566), .Y(n66657) );
  XOR2xp5_ASAP7_75t_SL U66652 ( .A(n59393), .B(n66835), .Y(n66673) );
  OAI22xp33_ASAP7_75t_SRAM U66653 ( .A1(n66857), .A2(n59440), .B1(n66619), 
        .B2(n59446), .Y(n66687) );
  NOR2xp33_ASAP7_75t_SL U66654 ( .A(n76071), .B(n59639), .Y(n66615) );
  XNOR2xp5_ASAP7_75t_SL U66655 ( .A(n66833), .B(n58529), .Y(n59393) );
  AOI21xp33_ASAP7_75t_SRAM U66656 ( .A1(n66333), .A2(n59648), .B(n66763), .Y(
        n66830) );
  XNOR2xp5_ASAP7_75t_SL U66657 ( .A(n57107), .B(n59607), .Y(n66857) );
  XOR2xp5_ASAP7_75t_SL U66658 ( .A(n68547), .B(n68548), .Y(n59016) );
  XOR2xp5_ASAP7_75t_SL U66659 ( .A(n66775), .B(n66774), .Y(n66776) );
  XNOR2xp5_ASAP7_75t_SL U66660 ( .A(n68460), .B(n68367), .Y(n68445) );
  XOR2xp5_ASAP7_75t_SL U66661 ( .A(n68458), .B(n68459), .Y(n68367) );
  XNOR2xp5_ASAP7_75t_SL U66662 ( .A(n58500), .B(n59267), .Y(n68541) );
  XNOR2xp5_ASAP7_75t_SL U66663 ( .A(n68527), .B(n68526), .Y(n68556) );
  XNOR2xp5_ASAP7_75t_SL U66664 ( .A(n66913), .B(n66914), .Y(n68524) );
  XNOR2xp5_ASAP7_75t_SL U66665 ( .A(n59071), .B(n59075), .Y(n66909) );
  OAI22xp33_ASAP7_75t_SRAM U66666 ( .A1(n66757), .A2(n59440), .B1(n59446), 
        .B2(n66756), .Y(n66814) );
  XNOR2xp5_ASAP7_75t_SL U66667 ( .A(n58919), .B(n59607), .Y(n66756) );
  XNOR2xp5_ASAP7_75t_SL U66668 ( .A(n59602), .B(n59668), .Y(n66667) );
  NOR2xp33_ASAP7_75t_SL U66669 ( .A(n66665), .B(n66664), .Y(n66748) );
  XNOR2xp5_ASAP7_75t_SL U66670 ( .A(n68535), .B(n59320), .Y(n68550) );
  XNOR2xp5_ASAP7_75t_SL U66671 ( .A(n66975), .B(n66974), .Y(n68534) );
  XOR2xp5_ASAP7_75t_SL U66672 ( .A(n66968), .B(n66967), .Y(n58503) );
  OAI21xp33_ASAP7_75t_SRAM U66673 ( .A1(n67839), .A2(n59637), .B(n66631), .Y(
        n66749) );
  NOR2xp33_ASAP7_75t_SL U66674 ( .A(n59641), .B(n75908), .Y(n66729) );
  XNOR2xp5_ASAP7_75t_SL U66675 ( .A(n67432), .B(n59607), .Y(n66755) );
  NOR2xp33_ASAP7_75t_SL U66676 ( .A(n66920), .B(n68361), .Y(n66927) );
  XNOR2xp5_ASAP7_75t_SL U66677 ( .A(n68406), .B(n59150), .Y(n68436) );
  INVxp33_ASAP7_75t_SRAM U66678 ( .A(n68401), .Y(n68403) );
  NOR2xp33_ASAP7_75t_SL U66679 ( .A(n56857), .B(n59191), .Y(n66710) );
  XNOR2xp5_ASAP7_75t_SL U66680 ( .A(n59603), .B(n59670), .Y(n66711) );
  OAI21xp33_ASAP7_75t_SRAM U66681 ( .A1(n66783), .A2(n58884), .B(n66715), .Y(
        n68479) );
  NAND2xp33_ASAP7_75t_SRAM U66682 ( .A(n59283), .B(n59637), .Y(n66630) );
  NOR2xp33_ASAP7_75t_SL U66683 ( .A(n66728), .B(n66727), .Y(n66963) );
  NOR2xp33_ASAP7_75t_SL U66684 ( .A(n59641), .B(n68087), .Y(n66728) );
  NOR2xp33_ASAP7_75t_SL U66685 ( .A(n66961), .B(n66960), .Y(n59288) );
  NAND2xp33_ASAP7_75t_SRAM U66686 ( .A(n67481), .B(n58015), .Y(n66929) );
  NOR2xp33_ASAP7_75t_SL U66687 ( .A(n68364), .B(n68363), .Y(n68366) );
  NOR2xp33_ASAP7_75t_SL U66688 ( .A(n66919), .B(n66918), .Y(n68361) );
  NAND2xp33_ASAP7_75t_SRAM U66689 ( .A(n57078), .B(n67846), .Y(n66916) );
  INVxp33_ASAP7_75t_SRAM U66690 ( .A(n68468), .Y(n68472) );
  INVxp33_ASAP7_75t_SRAM U66691 ( .A(n66623), .Y(n66796) );
  XNOR2xp5_ASAP7_75t_SL U66692 ( .A(n68315), .B(n58636), .Y(n68349) );
  XNOR2xp5_ASAP7_75t_SL U66693 ( .A(n68300), .B(n68299), .Y(n68314) );
  XNOR2xp5_ASAP7_75t_SL U66694 ( .A(n64987), .B(n64986), .Y(n68337) );
  XNOR2xp5_ASAP7_75t_SL U66695 ( .A(n64692), .B(n64691), .Y(n64715) );
  O2A1O1Ixp5_ASAP7_75t_SL U66696 ( .A1(n58383), .A2(n59656), .B(n58759), .C(
        n64685), .Y(n64687) );
  NOR2xp33_ASAP7_75t_SL U66697 ( .A(n63824), .B(n67442), .Y(n63666) );
  NAND2xp33_ASAP7_75t_SRAM U66698 ( .A(n58919), .B(n67428), .Y(n63657) );
  XNOR2xp5_ASAP7_75t_SL U66699 ( .A(n59331), .B(n64344), .Y(n64683) );
  XNOR2xp5_ASAP7_75t_SL U66700 ( .A(n64345), .B(n64346), .Y(n59331) );
  XNOR2xp5_ASAP7_75t_SL U66701 ( .A(n64671), .B(n64672), .Y(n64673) );
  AOI211xp5_ASAP7_75t_SL U66702 ( .A1(n64668), .A2(n64667), .B(n64666), .C(
        n64665), .Y(n64670) );
  INVxp33_ASAP7_75t_SRAM U66703 ( .A(n64664), .Y(n64666) );
  XNOR2xp5_ASAP7_75t_SL U66704 ( .A(n63846), .B(n63845), .Y(n64088) );
  NAND2xp33_ASAP7_75t_SRAM U66705 ( .A(n59595), .B(n75906), .Y(n63209) );
  XNOR2xp5_ASAP7_75t_SL U66706 ( .A(n68275), .B(n68274), .Y(n68295) );
  XNOR2xp5_ASAP7_75t_SL U66707 ( .A(n68291), .B(n68290), .Y(n68301) );
  INVxp33_ASAP7_75t_SRAM U66708 ( .A(n68288), .Y(n68291) );
  XNOR2xp5_ASAP7_75t_SL U66709 ( .A(n59248), .B(n59246), .Y(n64983) );
  XOR2xp5_ASAP7_75t_SL U66710 ( .A(n64871), .B(n58337), .Y(n59246) );
  XNOR2xp5_ASAP7_75t_SL U66711 ( .A(n64546), .B(n64545), .Y(n64547) );
  XNOR2xp5_ASAP7_75t_SL U66712 ( .A(n64454), .B(n58780), .Y(n64672) );
  NAND2xp33_ASAP7_75t_SRAM U66713 ( .A(n67228), .B(n64897), .Y(n63828) );
  NAND2xp33_ASAP7_75t_SRAM U66714 ( .A(n59609), .B(n67264), .Y(n58936) );
  NOR2xp33_ASAP7_75t_SL U66715 ( .A(n59468), .B(n67920), .Y(n63839) );
  NAND2xp33_ASAP7_75t_SRAM U66716 ( .A(n59593), .B(n67962), .Y(n63635) );
  NAND2xp33_ASAP7_75t_SRAM U66717 ( .A(n59505), .B(n53280), .Y(n63863) );
  NAND2xp33_ASAP7_75t_SRAM U66718 ( .A(n57108), .B(n67569), .Y(n63864) );
  NAND2xp33_ASAP7_75t_SRAM U66719 ( .A(n59599), .B(n67914), .Y(n66422) );
  NAND2xp33_ASAP7_75t_SRAM U66720 ( .A(n64418), .B(n64417), .Y(n64420) );
  INVxp33_ASAP7_75t_SRAM U66721 ( .A(n63859), .Y(n63861) );
  NOR2xp33_ASAP7_75t_SL U66722 ( .A(n64022), .B(n59460), .Y(n64023) );
  NOR2xp33_ASAP7_75t_SL U66723 ( .A(n59515), .B(n64380), .Y(n64024) );
  XOR2xp5_ASAP7_75t_SL U66724 ( .A(n64413), .B(n64412), .Y(n64658) );
  XNOR2xp5_ASAP7_75t_SL U66725 ( .A(n64405), .B(n64526), .Y(n64413) );
  XNOR2xp5_ASAP7_75t_SL U66726 ( .A(n65065), .B(n65064), .Y(n68257) );
  XNOR2xp5_ASAP7_75t_SL U66727 ( .A(n64656), .B(n64655), .Y(n64911) );
  XOR2xp5_ASAP7_75t_SL U66728 ( .A(n64654), .B(n64905), .Y(n64655) );
  XNOR2xp5_ASAP7_75t_SL U66729 ( .A(n64946), .B(n64632), .Y(n64912) );
  XNOR2xp5_ASAP7_75t_SL U66730 ( .A(n64542), .B(n64602), .Y(n64543) );
  XNOR2xp5_ASAP7_75t_SL U66731 ( .A(n64404), .B(n64403), .Y(n64526) );
  INVxp33_ASAP7_75t_SRAM U66732 ( .A(n58432), .Y(n64385) );
  NOR2xp33_ASAP7_75t_SL U66733 ( .A(n64380), .B(n57360), .Y(n64381) );
  NOR2xp33_ASAP7_75t_SL U66734 ( .A(n59515), .B(n64379), .Y(n64382) );
  NAND2xp33_ASAP7_75t_SRAM U66735 ( .A(n67911), .B(n67428), .Y(n64070) );
  NOR2xp33_ASAP7_75t_SL U66736 ( .A(n64374), .B(n59067), .Y(n64349) );
  NOR2xp33_ASAP7_75t_SL U66737 ( .A(n57508), .B(n64072), .Y(n64348) );
  AOI31xp33_ASAP7_75t_SL U66738 ( .A1(n63813), .A2(n63812), .A3(n63811), .B(
        n63810), .Y(n64351) );
  NAND2xp33_ASAP7_75t_SRAM U66739 ( .A(n67911), .B(n58439), .Y(n63813) );
  XNOR2xp5_ASAP7_75t_SL U66740 ( .A(n58402), .B(n59511), .Y(n64035) );
  XNOR2xp5_ASAP7_75t_SL U66741 ( .A(n64477), .B(n64361), .Y(n64524) );
  XNOR2xp5_ASAP7_75t_SL U66742 ( .A(n64530), .B(n64375), .Y(n64376) );
  AOI211xp5_ASAP7_75t_SL U66743 ( .A1(n64970), .A2(n64969), .B(n64968), .C(
        n64967), .Y(n64972) );
  NOR2xp33_ASAP7_75t_SL U66744 ( .A(n64944), .B(n64943), .Y(n64997) );
  NAND2xp33_ASAP7_75t_SRAM U66745 ( .A(n59599), .B(n67227), .Y(n63815) );
  NAND2xp33_ASAP7_75t_SRAM U66746 ( .A(n57180), .B(n58753), .Y(n64372) );
  NAND2xp33_ASAP7_75t_SRAM U66747 ( .A(n59505), .B(n57315), .Y(n64399) );
  O2A1O1Ixp5_ASAP7_75t_SL U66748 ( .A1(n59654), .A2(n64390), .B(n59411), .C(
        n59604), .Y(n64391) );
  XNOR2xp5_ASAP7_75t_SL U66749 ( .A(n64614), .B(n64613), .Y(n64944) );
  NAND2xp33_ASAP7_75t_SRAM U66750 ( .A(n59505), .B(n76077), .Y(n64427) );
  NAND2xp33_ASAP7_75t_SRAM U66751 ( .A(n59283), .B(n59466), .Y(n64446) );
  XNOR2xp5_ASAP7_75t_SL U66752 ( .A(n64583), .B(n64893), .Y(n64585) );
  XNOR2xp5_ASAP7_75t_SL U66753 ( .A(n64583), .B(n64508), .Y(n64519) );
  XNOR2xp5_ASAP7_75t_SL U66754 ( .A(n59511), .B(n59599), .Y(n64616) );
  INVxp33_ASAP7_75t_SRAM U66755 ( .A(n64562), .Y(n64491) );
  XNOR2xp5_ASAP7_75t_SL U66756 ( .A(n58996), .B(n64882), .Y(n64907) );
  XOR2xp5_ASAP7_75t_SL U66757 ( .A(n64883), .B(n64878), .Y(n58996) );
  XNOR2xp5_ASAP7_75t_SL U66758 ( .A(n64653), .B(n64652), .Y(n64905) );
  NAND2xp33_ASAP7_75t_SRAM U66759 ( .A(n76028), .B(n67738), .Y(n64608) );
  O2A1O1Ixp5_ASAP7_75t_SL U66760 ( .A1(n59466), .A2(n57167), .B(n64939), .C(
        n59012), .Y(n64633) );
  NOR2xp33_ASAP7_75t_SL U66761 ( .A(n64636), .B(n64635), .Y(n64885) );
  NOR2xp33_ASAP7_75t_SL U66762 ( .A(n59515), .B(n64922), .Y(n64636) );
  AO21x1_ASAP7_75t_SL U66763 ( .A1(n75900), .A2(n59230), .B(n67960), .Y(n64922) );
  XNOR2xp5_ASAP7_75t_SL U66764 ( .A(n59466), .B(n59620), .Y(n64502) );
  XNOR2xp5_ASAP7_75t_SL U66765 ( .A(n59596), .B(n67228), .Y(n64498) );
  XNOR2xp5_ASAP7_75t_SL U66766 ( .A(n64558), .B(n64559), .Y(n64470) );
  XNOR2xp5_ASAP7_75t_SL U66767 ( .A(n59468), .B(n76028), .Y(n64466) );
  AO21x1_ASAP7_75t_SL U66768 ( .A1(n67912), .A2(n64634), .B(n59129), .Y(n64558) );
  NAND2xp33_ASAP7_75t_SRAM U66769 ( .A(n57112), .B(n59659), .Y(n64479) );
  XNOR2xp5_ASAP7_75t_SL U66770 ( .A(n59609), .B(n57315), .Y(n64643) );
  XNOR2xp5_ASAP7_75t_SL U66771 ( .A(n68369), .B(n67755), .Y(n68354) );
  XNOR2xp5_ASAP7_75t_SL U66772 ( .A(n57108), .B(n59667), .Y(n67750) );
  NAND2xp33_ASAP7_75t_SRAM U66773 ( .A(n59634), .B(n67747), .Y(n59078) );
  NAND2xp33_ASAP7_75t_SRAM U66774 ( .A(n59467), .B(n67736), .Y(n67735) );
  NAND2xp33_ASAP7_75t_SRAM U66775 ( .A(n59641), .B(n76049), .Y(n67705) );
  NAND2xp33_ASAP7_75t_SRAM U66776 ( .A(n53207), .B(n67855), .Y(n67703) );
  XOR2xp5_ASAP7_75t_SL U66777 ( .A(n68392), .B(n68393), .Y(n67694) );
  XNOR2xp5_ASAP7_75t_SL U66778 ( .A(n59024), .B(n59001), .Y(n68392) );
  INVxp33_ASAP7_75t_SRAM U66779 ( .A(n67760), .Y(n67662) );
  INVxp33_ASAP7_75t_SRAM U66780 ( .A(n67766), .Y(n67658) );
  INVxp33_ASAP7_75t_SRAM U66781 ( .A(n67759), .Y(n67663) );
  NOR2xp33_ASAP7_75t_SL U66782 ( .A(n58846), .B(n58847), .Y(n67759) );
  XNOR2xp5_ASAP7_75t_SL U66783 ( .A(n67666), .B(n67573), .Y(n67761) );
  XNOR2xp5_ASAP7_75t_SL U66784 ( .A(n67688), .B(n67572), .Y(n67671) );
  NAND2xp33_ASAP7_75t_SRAM U66785 ( .A(n59653), .B(n59169), .Y(n58982) );
  NOR2xp33_ASAP7_75t_SL U66786 ( .A(n67553), .B(n67554), .Y(n67678) );
  XNOR2xp5_ASAP7_75t_SL U66787 ( .A(n67692), .B(n67538), .Y(n67695) );
  XNOR2xp5_ASAP7_75t_SL U66788 ( .A(n67525), .B(n67524), .Y(n67575) );
  NOR2xp33_ASAP7_75t_SL U66789 ( .A(n67518), .B(n75076), .Y(n67540) );
  NAND2xp33_ASAP7_75t_SRAM U66790 ( .A(n67517), .B(n67516), .Y(n67518) );
  XOR2xp5_ASAP7_75t_SL U66791 ( .A(n67544), .B(n67545), .Y(n67525) );
  NOR2xp33_ASAP7_75t_SL U66792 ( .A(n67512), .B(n68383), .Y(n67541) );
  XNOR2xp5_ASAP7_75t_SL U66793 ( .A(n67679), .B(n67507), .Y(n67577) );
  XNOR2xp5_ASAP7_75t_SL U66794 ( .A(n67259), .B(n57303), .Y(n67787) );
  INVxp33_ASAP7_75t_SRAM U66795 ( .A(n67396), .Y(n67397) );
  NOR2xp33_ASAP7_75t_SL U66796 ( .A(n67579), .B(n67578), .Y(n67396) );
  NAND2xp33_ASAP7_75t_SRAM U66797 ( .A(n59145), .B(n59594), .Y(n58478) );
  NOR2xp33_ASAP7_75t_SL U66798 ( .A(n59097), .B(n59636), .Y(n59096) );
  XNOR2xp5_ASAP7_75t_SL U66799 ( .A(n59594), .B(n59667), .Y(n67534) );
  NOR2xp33_ASAP7_75t_SL U66800 ( .A(n59605), .B(n76172), .Y(n67474) );
  NOR2xp33_ASAP7_75t_SL U66801 ( .A(n59502), .B(n59642), .Y(n67557) );
  NAND2xp33_ASAP7_75t_SRAM U66802 ( .A(n67883), .B(n57321), .Y(n67469) );
  NAND2xp33_ASAP7_75t_SRAM U66803 ( .A(n57321), .B(n67457), .Y(n67462) );
  OAI22xp33_ASAP7_75t_SRAM U66804 ( .A1(n67456), .A2(n59440), .B1(n67455), 
        .B2(n59446), .Y(n67497) );
  XNOR2xp5_ASAP7_75t_SL U66805 ( .A(n67655), .B(n59141), .Y(n67659) );
  XNOR2xp5_ASAP7_75t_SL U66806 ( .A(n67520), .B(n67523), .Y(n59141) );
  NOR2xp33_ASAP7_75t_SL U66807 ( .A(n75032), .B(n67747), .Y(n67519) );
  OAI21xp33_ASAP7_75t_SRAM U66808 ( .A1(n76028), .A2(n59642), .B(n67711), .Y(
        n67279) );
  NOR2xp33_ASAP7_75t_SL U66809 ( .A(n57485), .B(n67408), .Y(n67409) );
  INVxp33_ASAP7_75t_SRAM U66810 ( .A(n56986), .Y(n67384) );
  AOI31xp33_ASAP7_75t_SL U66811 ( .A1(n68333), .A2(n68226), .A3(n68225), .B(
        n68331), .Y(n68227) );
  NAND2xp33_ASAP7_75t_SRAM U66812 ( .A(n58851), .B(n67231), .Y(n64925) );
  NAND2xp33_ASAP7_75t_SRAM U66813 ( .A(n59659), .B(n67458), .Y(n64926) );
  INVxp33_ASAP7_75t_SRAM U66814 ( .A(n68213), .Y(n68215) );
  XOR2xp5_ASAP7_75t_SL U66815 ( .A(n68210), .B(n68209), .Y(n68211) );
  XNOR2xp5_ASAP7_75t_SL U66816 ( .A(n68206), .B(n58352), .Y(n58441) );
  XOR2xp5_ASAP7_75t_SL U66817 ( .A(n68196), .B(n68195), .Y(n68197) );
  XNOR2xp5_ASAP7_75t_SL U66818 ( .A(n68185), .B(n68232), .Y(n68186) );
  O2A1O1Ixp5_ASAP7_75t_SL U66819 ( .A1(n62610), .A2(n57119), .B(n58206), .C(
        n58460), .Y(n62690) );
  NAND2xp33_ASAP7_75t_SRAM U66820 ( .A(n59532), .B(n57465), .Y(n64510) );
  NAND2xp33_ASAP7_75t_SRAM U66821 ( .A(n58439), .B(n75947), .Y(n59373) );
  XNOR2xp5_ASAP7_75t_SL U66822 ( .A(n58923), .B(n67352), .Y(n58922) );
  NOR2xp33_ASAP7_75t_SL U66823 ( .A(n58919), .B(n67948), .Y(n67261) );
  AOI21xp33_ASAP7_75t_SRAM U66824 ( .A1(n58384), .A2(n75906), .B(n67240), .Y(
        n67386) );
  NAND2xp33_ASAP7_75t_SRAM U66825 ( .A(n59619), .B(n56986), .Y(n67269) );
  XOR2xp5_ASAP7_75t_SL U66826 ( .A(n59084), .B(n67293), .Y(n67783) );
  NOR2xp33_ASAP7_75t_SL U66827 ( .A(n67906), .B(n67450), .Y(n59377) );
  XNOR2xp5_ASAP7_75t_SL U66828 ( .A(n59503), .B(n59667), .Y(n67450) );
  NOR2xp33_ASAP7_75t_SL U66829 ( .A(n59230), .B(n67826), .Y(n58960) );
  NOR2xp33_ASAP7_75t_SL U66830 ( .A(n59603), .B(n58901), .Y(n65036) );
  NOR2xp33_ASAP7_75t_SL U66831 ( .A(n57111), .B(n65033), .Y(n65037) );
  XNOR2xp5_ASAP7_75t_SL U66832 ( .A(n59607), .B(n75641), .Y(n65033) );
  XNOR2xp5_ASAP7_75t_SL U66833 ( .A(n67800), .B(n67799), .Y(n68070) );
  NAND2xp33_ASAP7_75t_SRAM U66834 ( .A(n67629), .B(n59050), .Y(n58805) );
  NAND2xp33_ASAP7_75t_SRAM U66835 ( .A(n67443), .B(n67967), .Y(n67448) );
  INVxp33_ASAP7_75t_SRAM U66836 ( .A(n67590), .Y(n67591) );
  XNOR2xp5_ASAP7_75t_SL U66837 ( .A(n58468), .B(n67817), .Y(n58628) );
  OR2x2_ASAP7_75t_SL U66838 ( .A(n66243), .B(n66286), .Y(n75958) );
  OAI21xp33_ASAP7_75t_SRAM U66839 ( .A1(n57347), .A2(n74781), .B(n66288), .Y(
        n66243) );
  NOR2xp33_ASAP7_75t_SL U66840 ( .A(n59012), .B(n67335), .Y(n58643) );
  OAI21xp33_ASAP7_75t_SRAM U66841 ( .A1(n67911), .A2(n59508), .B(n67224), .Y(
        n67225) );
  XNOR2xp5_ASAP7_75t_SL U66842 ( .A(n67776), .B(n67775), .Y(n68035) );
  NOR2xp33_ASAP7_75t_SL U66843 ( .A(n67369), .B(n59356), .Y(n67832) );
  NOR2xp33_ASAP7_75t_SL U66844 ( .A(n67583), .B(n67584), .Y(n67834) );
  NAND2xp33_ASAP7_75t_SRAM U66845 ( .A(n59615), .B(n67736), .Y(n67299) );
  NAND2xp33_ASAP7_75t_SRAM U66846 ( .A(n68011), .B(n59475), .Y(n59317) );
  NOR2xp33_ASAP7_75t_SL U66847 ( .A(n67636), .B(n59599), .Y(n59113) );
  NOR2xp33_ASAP7_75t_SL U66848 ( .A(n67629), .B(n53317), .Y(n63083) );
  XNOR2xp5_ASAP7_75t_SL U66849 ( .A(n59594), .B(n75947), .Y(n67608) );
  XNOR2xp5_ASAP7_75t_SL U66850 ( .A(n59617), .B(n67964), .Y(n67824) );
  XNOR2xp5_ASAP7_75t_SL U66851 ( .A(n59512), .B(n59640), .Y(n67852) );
  NOR2xp33_ASAP7_75t_SL U66852 ( .A(n58369), .B(n68233), .Y(n68031) );
  XNOR2xp5_ASAP7_75t_SL U66853 ( .A(n58430), .B(n58926), .Y(n58754) );
  NOR4xp25_ASAP7_75t_SL U66854 ( .A(n59233), .B(n64965), .C(n59236), .D(n62806), .Y(n67806) );
  NOR3xp33_ASAP7_75t_SL U66855 ( .A(n59234), .B(n63836), .C(n59235), .Y(n59233) );
  AOI21xp33_ASAP7_75t_SRAM U66856 ( .A1(n59543), .A2(n57122), .B(n62556), .Y(
        n62559) );
  INVxp33_ASAP7_75t_SRAM U66857 ( .A(n59543), .Y(n77696) );
  XOR2xp5_ASAP7_75t_SL U66858 ( .A(n58873), .B(n58715), .Y(n58430) );
  XNOR2xp5_ASAP7_75t_SL U66859 ( .A(n67984), .B(n59450), .Y(n58873) );
  NOR2xp33_ASAP7_75t_SL U66860 ( .A(n59509), .B(n59190), .Y(n59110) );
  NOR2xp33_ASAP7_75t_SL U66861 ( .A(n59543), .B(n57186), .Y(n62583) );
  XNOR2xp5_ASAP7_75t_SL U66862 ( .A(n67983), .B(n67982), .Y(n68185) );
  AND2x2_ASAP7_75t_SL U66863 ( .A(n59578), .B(n59546), .Y(n58520) );
  NOR3xp33_ASAP7_75t_SL U66864 ( .A(n62591), .B(n62590), .C(n76690), .Y(n62592) );
  NOR2xp33_ASAP7_75t_SL U66865 ( .A(n59079), .B(n62637), .Y(n62638) );
  NOR2xp33_ASAP7_75t_SL U66866 ( .A(n59534), .B(n63653), .Y(n63655) );
  NOR2xp33_ASAP7_75t_SL U66867 ( .A(n57184), .B(n59448), .Y(n59328) );
  NOR2xp33_ASAP7_75t_SL U66868 ( .A(n68098), .B(n67365), .Y(n67366) );
  NOR2xp33_ASAP7_75t_SL U66869 ( .A(n74781), .B(n66634), .Y(n66287) );
  NOR2xp33_ASAP7_75t_SL U66870 ( .A(n59258), .B(n57219), .Y(n59257) );
  NOR2xp33_ASAP7_75t_SL U66871 ( .A(n58504), .B(n59009), .Y(n67900) );
  NOR2xp33_ASAP7_75t_SL U66872 ( .A(n59553), .B(n62671), .Y(n64389) );
  NOR2xp33_ASAP7_75t_SL U66873 ( .A(n59535), .B(n59474), .Y(n58828) );
  NOR2xp33_ASAP7_75t_SL U66874 ( .A(n59532), .B(n59591), .Y(n63806) );
  AND2x2_ASAP7_75t_SL U66875 ( .A(n63808), .B(n59290), .Y(n67971) );
  O2A1O1Ixp5_ASAP7_75t_SL U66876 ( .A1(n59592), .A2(n64930), .B(n57186), .C(
        n59532), .Y(n64931) );
  NOR2xp33_ASAP7_75t_SL U66877 ( .A(n77717), .B(n59654), .Y(n58980) );
  INVxp33_ASAP7_75t_SRAM U66878 ( .A(n59532), .Y(n77715) );
  NOR2xp33_ASAP7_75t_SL U66879 ( .A(n63569), .B(n59654), .Y(n62681) );
  NOR2xp33_ASAP7_75t_SL U66880 ( .A(n59398), .B(n59646), .Y(n64116) );
  NOR2xp33_ASAP7_75t_SL U66881 ( .A(n59544), .B(n64229), .Y(n62599) );
  OAI21xp33_ASAP7_75t_SRAM U66882 ( .A1(n64229), .A2(n57122), .B(n59544), .Y(
        n59326) );
  HB1xp67_ASAP7_75t_SL U66883 ( .A(n64358), .Y(n59472) );
  OAI21xp33_ASAP7_75t_SRAM U66884 ( .A1(n64894), .A2(n64357), .B(n57209), .Y(
        n64365) );
  XNOR2xp5_ASAP7_75t_SL U66885 ( .A(n58919), .B(n59603), .Y(n68014) );
  NOR2xp33_ASAP7_75t_SL U66886 ( .A(n57122), .B(n58925), .Y(n59181) );
  NAND2xp33_ASAP7_75t_SRAM U66887 ( .A(n58206), .B(n59589), .Y(n62608) );
  NOR2xp33_ASAP7_75t_SL U66888 ( .A(n76653), .B(n76627), .Y(n62605) );
  NOR2xp33_ASAP7_75t_SL U66889 ( .A(n64079), .B(n64080), .Y(n59187) );
  NOR2xp33_ASAP7_75t_SL U66890 ( .A(n61910), .B(n61909), .Y(n61932) );
  INVxp33_ASAP7_75t_SRAM U66891 ( .A(n1690), .Y(n77709) );
  AND2x2_ASAP7_75t_SL U66892 ( .A(n59569), .B(n59542), .Y(n60595) );
  NAND2xp33_ASAP7_75t_SRAM U66893 ( .A(n59556), .B(n62614), .Y(n58860) );
  OR2x2_ASAP7_75t_SL U66894 ( .A(n62632), .B(n62631), .Y(n58408) );
  NOR2xp33_ASAP7_75t_SL U66895 ( .A(n59577), .B(n64357), .Y(n64356) );
  NOR2xp33_ASAP7_75t_SL U66896 ( .A(n75081), .B(n75083), .Y(n75079) );
  NOR2xp33_ASAP7_75t_SL U66897 ( .A(n75067), .B(n68610), .Y(n75055) );
  NOR2xp33_ASAP7_75t_SL U66898 ( .A(n59116), .B(n75034), .Y(n68605) );
  NOR2xp33_ASAP7_75t_SL U66899 ( .A(n68119), .B(n68606), .Y(n66569) );
  NOR2xp33_ASAP7_75t_SL U66900 ( .A(n75053), .B(n75052), .Y(n75065) );
  NAND2xp33_ASAP7_75t_SRAM U66901 ( .A(n59664), .B(n75046), .Y(n75051) );
  XNOR2xp5_ASAP7_75t_SL U66902 ( .A(n75064), .B(n75063), .Y(n75082) );
  XOR2xp5_ASAP7_75t_SL U66903 ( .A(n59670), .B(n59638), .Y(n75040) );
  NOR2xp33_ASAP7_75t_SL U66904 ( .A(n59549), .B(n66294), .Y(n59413) );
  NOR2xp33_ASAP7_75t_SL U66905 ( .A(n75848), .B(n66293), .Y(n66294) );
  INVxp33_ASAP7_75t_SRAM U66906 ( .A(n66292), .Y(n66293) );
  NOR2xp33_ASAP7_75t_SL U66907 ( .A(n59576), .B(n66256), .Y(n66261) );
  NOR2xp33_ASAP7_75t_SL U66908 ( .A(n66240), .B(n66239), .Y(n66242) );
  NAND3xp33_ASAP7_75t_SL U66909 ( .A(n60536), .B(n59405), .C(n61646), .Y(
        n66239) );
  AND2x2_ASAP7_75t_SL U66910 ( .A(n59575), .B(n59576), .Y(n61646) );
  NOR2xp33_ASAP7_75t_SL U66911 ( .A(n74776), .B(n61214), .Y(n60536) );
  XOR2xp5_ASAP7_75t_SL U66912 ( .A(n59670), .B(n59640), .Y(n75077) );
  AND2x2_ASAP7_75t_SL U66913 ( .A(n61965), .B(n58443), .Y(n59424) );
  NOR2xp33_ASAP7_75t_SL U66914 ( .A(n74781), .B(n77735), .Y(n66292) );
  AND4x1_ASAP7_75t_SL U66915 ( .A(n61931), .B(n1588), .C(n61964), .D(n61911), 
        .Y(n61965) );
  NOR2xp33_ASAP7_75t_SL U66916 ( .A(n59445), .B(n59566), .Y(n60629) );
  NAND3xp33_ASAP7_75t_SL U66917 ( .A(n2501), .B(n2526), .C(n2473), .Y(n58717)
         );
  NOR3xp33_ASAP7_75t_SL U66918 ( .A(or1200_cpu_or1200_except_n552), .B(
        or1200_cpu_or1200_except_n555), .C(
        or1200_cpu_or1200_except_ex_freeze_prev), .Y(n62010) );
  NOR2xp33_ASAP7_75t_SL U66919 ( .A(n61214), .B(n61206), .Y(n60658) );
  OAI22xp33_ASAP7_75t_SRAM U66920 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_ine), .A2(n74741), .B1(
        or1200_cpu_or1200_fpu_fpu_op_r_1_), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_ine_o), .Y(n74742) );
  OAI22xp33_ASAP7_75t_SRAM U66921 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[30]), .A2(n74741), 
        .B1(or1200_cpu_or1200_fpu_fpu_op_r_1_), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[30]), .Y(
        n74282) );
  OAI22xp33_ASAP7_75t_SRAM U66922 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[25]), .A2(n74741), 
        .B1(or1200_cpu_or1200_fpu_fpu_op_r_1_), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[25]), .Y(
        n74106) );
  OAI22xp33_ASAP7_75t_SRAM U66923 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_post_norm_div_output[26]), .A2(n74741), 
        .B1(or1200_cpu_or1200_fpu_fpu_op_r_1_), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_postnorm_addsub_output_o[26]), .Y(
        n73901) );
  NOR2xp33_ASAP7_75t_SL U66924 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        n72112), .Y(n72126) );
  NOR2xp33_ASAP7_75t_SL U66925 ( .A(n74237), .B(n72585), .Y(n72588) );
  NOR2xp33_ASAP7_75t_SL U66926 ( .A(n66060), .B(n66080), .Y(n66055) );
  NOR2xp33_ASAP7_75t_SL U66927 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[35]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[34]), .Y(n65378) );
  NOR2xp33_ASAP7_75t_SL U66928 ( .A(n71692), .B(n71661), .Y(n71639) );
  NOR3xp33_ASAP7_75t_SL U66929 ( .A(n62194), .B(n62193), .C(n62192), .Y(n62195) );
  NOR2xp33_ASAP7_75t_SL U66930 ( .A(n64802), .B(n64804), .Y(n74076) );
  O2A1O1Ixp5_ASAP7_75t_SL U66931 ( .A1(n73927), .A2(n74608), .B(n73926), .C(
        n73925), .Y(n73928) );
  O2A1O1Ixp5_ASAP7_75t_SL U66932 ( .A1(n61707), .A2(n75226), .B(n61706), .C(
        n61868), .Y(n77108) );
  NOR2xp33_ASAP7_75t_SL U66933 ( .A(n61802), .B(n61801), .Y(n77905) );
  NOR2xp33_ASAP7_75t_SL U66934 ( .A(n61762), .B(n62250), .Y(n77614) );
  O2A1O1Ixp5_ASAP7_75t_SL U66935 ( .A1(n61530), .A2(n75226), .B(n61706), .C(
        n61868), .Y(n75573) );
  O2A1O1Ixp5_ASAP7_75t_SL U66936 ( .A1(n75866), .A2(n75865), .B(n75864), .C(
        n75863), .Y(n75867) );
  OAI22xp33_ASAP7_75t_SRAM U66937 ( .A1(n2499), .A2(n62005), .B1(n2473), .B2(
        n77567), .Y(n9566) );
  XNOR2xp5_ASAP7_75t_SL U66938 ( .A(n2037), .B(or1200_cpu_or1200_except_n658), 
        .Y(n75158) );
  NOR2xp33_ASAP7_75t_SL U66939 ( .A(or1200_cpu_or1200_mult_mac_n383), .B(
        n69163), .Y(n69191) );
  NOR2xp33_ASAP7_75t_SL U66940 ( .A(or1200_cpu_or1200_mult_mac_n171), .B(
        n63501), .Y(n63518) );
  XOR2xp5_ASAP7_75t_SL U66941 ( .A(or1200_cpu_or1200_mult_mac_n295), .B(
        or1200_cpu_or1200_mult_mac_n149), .Y(n63399) );
  NOR2xp33_ASAP7_75t_SL U66942 ( .A(or1200_cpu_or1200_mult_mac_n387), .B(
        n69188), .Y(n69200) );
  NOR3xp33_ASAP7_75t_SL U66943 ( .A(n75129), .B(n75128), .C(n75127), .Y(n75131) );
  NOR2xp33_ASAP7_75t_SL U66944 ( .A(or1200_cpu_or1200_mult_mac_n403), .B(
        n75116), .Y(n75128) );
  NOR2xp33_ASAP7_75t_SL U66945 ( .A(or1200_cpu_or1200_mult_mac_n405), .B(
        n75126), .Y(n75129) );
  OAI22xp33_ASAP7_75t_SRAM U66946 ( .A1(n2517), .A2(n62005), .B1(n2501), .B2(
        n77567), .Y(n9567) );
  NOR2xp33_ASAP7_75t_SL U66947 ( .A(n65354), .B(n65279), .Y(n65283) );
  AOI31xp33_ASAP7_75t_SL U66948 ( .A1(n77676), .A2(n77128), .A3(n77674), .B(
        n61897), .Y(n61898) );
  NAND2xp33_ASAP7_75t_SRAM U66949 ( .A(n75876), .B(n77124), .Y(n61895) );
  AOI22xp33_ASAP7_75t_SRAM U66950 ( .A1(or1200_cpu_or1200_fpu_result_arith[31]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[31]), .Y(
        n61859) );
  AND2x2_ASAP7_75t_SL U66951 ( .A(n73490), .B(n73489), .Y(n73591) );
  AOI211xp5_ASAP7_75t_SL U66952 ( .A1(or1200_cpu_rf_datab[30]), .A2(n57091), 
        .B(n77184), .C(n75757), .Y(n75758) );
  AOI22xp33_ASAP7_75t_SRAM U66953 ( .A1(n59550), .A2(n75735), .B1(n76429), 
        .B2(n75734), .Y(n75742) );
  INVxp33_ASAP7_75t_SRAM U66954 ( .A(n75707), .Y(n75711) );
  NOR2xp33_ASAP7_75t_SL U66955 ( .A(n69840), .B(n70103), .Y(n69639) );
  AOI22xp33_ASAP7_75t_SRAM U66956 ( .A1(n75853), .A2(n63272), .B1(n60965), 
        .B2(n57191), .Y(n60966) );
  NOR4xp25_ASAP7_75t_SL U66957 ( .A(n62108), .B(n61886), .C(n61104), .D(n61880), .Y(n61639) );
  AOI22xp33_ASAP7_75t_SRAM U66958 ( .A1(n64219), .A2(n62279), .B1(n77076), 
        .B2(n61643), .Y(n60959) );
  INVxp33_ASAP7_75t_SRAM U66959 ( .A(n76763), .Y(n60961) );
  NAND2xp33_ASAP7_75t_SRAM U66960 ( .A(n76782), .B(n75323), .Y(n61353) );
  AOI21xp33_ASAP7_75t_SRAM U66961 ( .A1(n60924), .A2(n57641), .B(n60923), .Y(
        n60925) );
  NOR4xp25_ASAP7_75t_SL U66962 ( .A(n61693), .B(n60908), .C(n60907), .D(n58552), .Y(n77588) );
  AOI22xp33_ASAP7_75t_SRAM U66963 ( .A1(n63272), .A2(n77039), .B1(n68846), 
        .B2(n68812), .Y(n60901) );
  NOR2xp33_ASAP7_75t_SL U66964 ( .A(n61030), .B(n62142), .Y(n60723) );
  NAND2xp33_ASAP7_75t_SRAM U66965 ( .A(n64282), .B(n60691), .Y(n76796) );
  AND2x2_ASAP7_75t_SL U66966 ( .A(n60689), .B(n75876), .Y(n77117) );
  AOI21xp33_ASAP7_75t_SRAM U66967 ( .A1(n75518), .A2(n76289), .B(n60673), .Y(
        n60674) );
  OAI22xp33_ASAP7_75t_SRAM U66968 ( .A1(or1200_cpu_or1200_mult_mac_n128), .A2(
        n77058), .B1(n59710), .B2(n76775), .Y(n60673) );
  AOI31xp33_ASAP7_75t_SL U66969 ( .A1(n61436), .A2(n60850), .A3(n60639), .B(
        n76779), .Y(n60640) );
  AOI22xp33_ASAP7_75t_SRAM U66970 ( .A1(n59709), .A2(n64132), .B1(n59708), 
        .B2(n64131), .Y(n64775) );
  NOR4xp25_ASAP7_75t_SL U66971 ( .A(n64838), .B(n75831), .C(n60638), .D(n64783), .Y(n64131) );
  NOR2xp33_ASAP7_75t_SL U66972 ( .A(n57641), .B(n61514), .Y(n61538) );
  NOR2xp33_ASAP7_75t_SL U66973 ( .A(n60642), .B(n61648), .Y(n60618) );
  INVxp33_ASAP7_75t_SRAM U66974 ( .A(n61647), .Y(n60642) );
  NOR2xp33_ASAP7_75t_SL U66975 ( .A(n59493), .B(n63261), .Y(n77041) );
  INVx1_ASAP7_75t_SL U66976 ( .A(n76720), .Y(n61226) );
  INVxp33_ASAP7_75t_SRAM U66977 ( .A(n60819), .Y(n60897) );
  OAI21xp33_ASAP7_75t_SRAM U66978 ( .A1(n61133), .A2(n61845), .B(n60553), .Y(
        n75561) );
  NAND2xp33_ASAP7_75t_SRAM U66979 ( .A(n77623), .B(n61845), .Y(n60553) );
  NOR2xp33_ASAP7_75t_SL U66980 ( .A(n60542), .B(n60576), .Y(n61480) );
  NAND4xp25_ASAP7_75t_SL U66981 ( .A(n12861), .B(n73839), .C(n12863), .D(
        n21879), .Y(n73840) );
  NOR2xp33_ASAP7_75t_SL U66982 ( .A(n73467), .B(n73466), .Y(n73468) );
  AND2x2_ASAP7_75t_SL U66983 ( .A(n77166), .B(n60551), .Y(n58416) );
  NOR2xp33_ASAP7_75t_SL U66984 ( .A(n60369), .B(n61311), .Y(n60725) );
  NAND3xp33_ASAP7_75t_SL U66985 ( .A(n61154), .B(n61028), .C(n2616), .Y(n61311) );
  O2A1O1Ixp5_ASAP7_75t_SL U66986 ( .A1(n74244), .A2(n74243), .B(n74281), .C(
        n74260), .Y(n2870) );
  NAND2xp33_ASAP7_75t_SRAM U66987 ( .A(n59567), .B(n59182), .Y(n73977) );
  NAND2xp33_ASAP7_75t_SRAM U66988 ( .A(n61969), .B(n61968), .Y(n61972) );
  NOR2xp33_ASAP7_75t_SL U66989 ( .A(n59182), .B(n60762), .Y(n60763) );
  NOR2xp33_ASAP7_75t_SL U66990 ( .A(n77164), .B(n60816), .Y(n60551) );
  NOR2xp33_ASAP7_75t_SL U66991 ( .A(n73529), .B(n73530), .Y(n73490) );
  NOR2xp33_ASAP7_75t_SL U66992 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[3]), .B(
        n73888), .Y(n73887) );
  NOR2xp33_ASAP7_75t_SL U66993 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[2]), .B(
        n73890), .Y(n73869) );
  NOR2xp33_ASAP7_75t_SL U66994 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[0]), .B(
        n73866), .Y(n73865) );
  AOI211xp5_ASAP7_75t_SL U66995 ( .A1(n70996), .A2(n71208), .B(n70866), .C(
        n70865), .Y(n71019) );
  XNOR2xp5_ASAP7_75t_SL U66996 ( .A(n75968), .B(n57398), .Y(n76193) );
  NOR2xp33_ASAP7_75t_SL U66997 ( .A(n60577), .B(n60576), .Y(n77848) );
  NOR2xp33_ASAP7_75t_SL U66998 ( .A(n75196), .B(n75189), .Y(n59869) );
  OAI21xp33_ASAP7_75t_SRAM U66999 ( .A1(n59555), .A2(n2145), .B(n59935), .Y(
        n76616) );
  NOR2xp33_ASAP7_75t_SL U67000 ( .A(n74873), .B(n74872), .Y(n74876) );
  NOR2xp33_ASAP7_75t_SL U67001 ( .A(n74750), .B(n74838), .Y(n74165) );
  NOR3xp33_ASAP7_75t_SL U67002 ( .A(n69151), .B(n69144), .C(n69149), .Y(n69157) );
  XNOR2xp5_ASAP7_75t_SL U67003 ( .A(n59607), .B(n59668), .Y(n66545) );
  NOR2xp33_ASAP7_75t_SL U67004 ( .A(n62971), .B(n62970), .Y(n62974) );
  NAND2xp33_ASAP7_75t_SRAM U67005 ( .A(n75901), .B(n67428), .Y(n62954) );
  NAND2xp33_ASAP7_75t_SRAM U67006 ( .A(n75900), .B(n57422), .Y(n63194) );
  XOR2xp5_ASAP7_75t_SL U67007 ( .A(n59173), .B(n66772), .Y(n66821) );
  XNOR2xp5_ASAP7_75t_SL U67008 ( .A(n59617), .B(n75947), .Y(n66726) );
  XNOR2xp5_ASAP7_75t_SL U67009 ( .A(n64532), .B(n64376), .Y(n64525) );
  INVxp33_ASAP7_75t_SRAM U67010 ( .A(n59534), .Y(n77713) );
  NAND2xp33_ASAP7_75t_SRAM U67011 ( .A(n59442), .B(n59712), .Y(n64233) );
  OR2x2_ASAP7_75t_SL U67012 ( .A(n59709), .B(n60860), .Y(n75710) );
  INVxp33_ASAP7_75t_SRAM U67013 ( .A(n59537), .Y(n63251) );
  NAND2xp33_ASAP7_75t_SRAM U67014 ( .A(n75074), .B(n75048), .Y(n75049) );
  NOR2xp33_ASAP7_75t_SL U67015 ( .A(n59387), .B(n61921), .Y(n61908) );
  INVxp33_ASAP7_75t_SRAM U67016 ( .A(n77831), .Y(n77832) );
  O2A1O1Ixp5_ASAP7_75t_SL U67017 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .A2(
        n72485), .B(n72412), .C(n72221), .Y(n72231) );
  OAI22xp33_ASAP7_75t_SRAM U67018 ( .A1(n59706), .A2(n77786), .B1(n57083), 
        .B2(n1277), .Y(n1278) );
  NOR2xp33_ASAP7_75t_SL U67019 ( .A(n71986), .B(n71985), .Y(n72226) );
  O2A1O1Ixp5_ASAP7_75t_SL U67020 ( .A1(n72197), .A2(n72367), .B(n57123), .C(
        n72196), .Y(n72198) );
  O2A1O1Ixp5_ASAP7_75t_SL U67021 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_13_), 
        .A2(n71617), .B(n71616), .C(n71615), .Y(n71618) );
  NOR2xp33_ASAP7_75t_SL U67022 ( .A(n72976), .B(n72963), .Y(n72734) );
  NOR2xp33_ASAP7_75t_SL U67023 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_13_), 
        .Y(n71433) );
  NOR2xp33_ASAP7_75t_SL U67024 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_), 
        .B(n71605), .Y(n71434) );
  NOR2xp33_ASAP7_75t_SL U67025 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_), .B(
        n73042), .Y(n72987) );
  OR2x2_ASAP7_75t_SL U67026 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .Y(
        n72976) );
  NOR3xp33_ASAP7_75t_SL U67027 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_7_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_5_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_6_), .Y(
        n72994) );
  XNOR2xp5_ASAP7_75t_SL U67028 ( .A(or1200_cpu_or1200_mult_mac_n333), .B(
        or1200_cpu_or1200_mult_mac_n187), .Y(n65135) );
  NOR2xp33_ASAP7_75t_SL U67029 ( .A(n74632), .B(n74634), .Y(n76877) );
  OAI22xp33_ASAP7_75t_SRAM U67030 ( .A1(n1476), .A2(n61596), .B1(n1406), .B2(
        n76716), .Y(n61602) );
  O2A1O1Ixp5_ASAP7_75t_SL U67031 ( .A1(n62380), .A2(n62379), .B(n57126), .C(
        n62378), .Y(n62384) );
  AOI22xp33_ASAP7_75t_SRAM U67032 ( .A1(or1200_cpu_or1200_fpu_result_arith[19]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[19]), .Y(
        n74600) );
  OAI22xp33_ASAP7_75t_SRAM U67033 ( .A1(n1143), .A2(n77033), .B1(n1448), .B2(
        n77034), .Y(n74583) );
  AOI22xp33_ASAP7_75t_SRAM U67034 ( .A1(or1200_pic_picmr_19_), .A2(n74582), 
        .B1(n77043), .B2(n74581), .Y(n74586) );
  OAI21xp33_ASAP7_75t_SRAM U67035 ( .A1(or1200_cpu_or1200_mult_mac_n92), .A2(
        n64785), .B(n63585), .Y(n63588) );
  OAI22xp33_ASAP7_75t_SRAM U67036 ( .A1(n76765), .A2(n63570), .B1(n75701), 
        .B2(n75325), .Y(n63576) );
  AOI22xp33_ASAP7_75t_SRAM U67037 ( .A1(n63552), .A2(n74582), .B1(n77043), 
        .B2(n74972), .Y(n63553) );
  OAI22xp33_ASAP7_75t_SRAM U67038 ( .A1(n1450), .A2(n77034), .B1(n1145), .B2(
        n77033), .Y(n63551) );
  AOI211xp5_ASAP7_75t_SL U67039 ( .A1(or1200_cpu_rf_datab[20]), .A2(n57091), 
        .B(n77184), .C(n64156), .Y(n64157) );
  OAI22xp33_ASAP7_75t_SRAM U67040 ( .A1(n1628), .A2(n59679), .B1(n1626), .B2(
        n57074), .Y(n64156) );
  AOI31xp33_ASAP7_75t_SL U67041 ( .A1(n75577), .A2(n58081), .A3(n64127), .B(
        n64126), .Y(n64130) );
  OAI21xp33_ASAP7_75t_SRAM U67042 ( .A1(or1200_cpu_or1200_mult_mac_n327), .A2(
        n75738), .B(n64125), .Y(n64126) );
  AOI22xp33_ASAP7_75t_SRAM U67043 ( .A1(or1200_cpu_or1200_fpu_result_arith[20]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[20]), .Y(
        n64122) );
  NAND2xp33_ASAP7_75t_SRAM U67044 ( .A(n77082), .B(n64107), .Y(n64141) );
  OAI22xp33_ASAP7_75t_SRAM U67045 ( .A1(n1446), .A2(n77034), .B1(n1141), .B2(
        n77033), .Y(n64100) );
  NOR2xp33_ASAP7_75t_SL U67046 ( .A(n63566), .B(n75840), .Y(n64829) );
  OAI22xp33_ASAP7_75t_SRAM U67047 ( .A1(n1362), .A2(n77035), .B1(n1360), .B2(
        n75364), .Y(n75365) );
  OAI22xp33_ASAP7_75t_SRAM U67048 ( .A1(n1452), .A2(n77034), .B1(n1147), .B2(
        n77033), .Y(n75362) );
  AOI211xp5_ASAP7_75t_SL U67049 ( .A1(or1200_cpu_rf_datab[28]), .A2(n57091), 
        .B(n77184), .C(n77183), .Y(n77189) );
  NOR2xp33_ASAP7_75t_SL U67050 ( .A(n64217), .B(n64216), .Y(n75607) );
  OAI22xp33_ASAP7_75t_SRAM U67051 ( .A1(or1200_cpu_or1200_mult_mac_n80), .A2(
        n64785), .B1(n57068), .B2(n64830), .Y(n64789) );
  OAI22xp33_ASAP7_75t_SRAM U67052 ( .A1(n1438), .A2(n77034), .B1(n1133), .B2(
        n77033), .Y(n64760) );
  AOI211xp5_ASAP7_75t_SL U67053 ( .A1(or1200_cpu_rf_datab[24]), .A2(n57091), 
        .B(n77184), .C(n64803), .Y(n64808) );
  OAI22xp33_ASAP7_75t_SRAM U67054 ( .A1(n1608), .A2(n59679), .B1(n57068), .B2(
        n57074), .Y(n64803) );
  NOR2xp33_ASAP7_75t_SL U67055 ( .A(n75872), .B(n76755), .Y(n74594) );
  OAI22xp33_ASAP7_75t_SRAM U67056 ( .A1(n1442), .A2(n77034), .B1(n1137), .B2(
        n77033), .Y(n64277) );
  NAND3xp33_ASAP7_75t_SL U67057 ( .A(or1200_cpu_or1200_mult_mac_n345), .B(
        or1200_cpu_or1200_mult_mac_n287), .C(or1200_cpu_or1200_mult_mac_n295), 
        .Y(n75502) );
  NOR2xp33_ASAP7_75t_SL U67058 ( .A(n76896), .B(n76895), .Y(n76912) );
  NOR2xp33_ASAP7_75t_SL U67059 ( .A(n3310), .B(n73609), .Y(n73541) );
  NOR2xp33_ASAP7_75t_SL U67060 ( .A(n61083), .B(n61082), .Y(n75217) );
  NOR2xp33_ASAP7_75t_SL U67061 ( .A(n69692), .B(n69688), .Y(n69985) );
  NOR2xp33_ASAP7_75t_SL U67062 ( .A(n69685), .B(n70103), .Y(n69692) );
  NOR2xp33_ASAP7_75t_SL U67063 ( .A(n69919), .B(n70103), .Y(n69679) );
  NOR2xp33_ASAP7_75t_SL U67064 ( .A(n69646), .B(n70103), .Y(n69649) );
  XOR2xp5_ASAP7_75t_SL U67065 ( .A(n73366), .B(n73365), .Y(n78220) );
  NOR2xp33_ASAP7_75t_SL U67066 ( .A(n77208), .B(n63713), .Y(n63726) );
  NAND3xp33_ASAP7_75t_SL U67067 ( .A(n2589), .B(n2814), .C(n3078), .Y(n60501)
         );
  NOR2xp33_ASAP7_75t_SL U67068 ( .A(n59576), .B(n61907), .Y(n61986) );
  NAND3xp33_ASAP7_75t_SL U67069 ( .A(n73515), .B(n73774), .C(n73753), .Y(
        n73529) );
  NOR2xp33_ASAP7_75t_SL U67070 ( .A(n73525), .B(n73533), .Y(n73488) );
  NOR2xp33_ASAP7_75t_SL U67071 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[5]), .B(
        n73882), .Y(n73892) );
  INVxp33_ASAP7_75t_SRAM U67072 ( .A(n68740), .Y(n68742) );
  NOR2xp33_ASAP7_75t_SL U67073 ( .A(n70815), .B(n70814), .Y(n70837) );
  NOR2xp33_ASAP7_75t_SL U67074 ( .A(n78408), .B(n71413), .Y(n70902) );
  OAI21xp33_ASAP7_75t_SRAM U67075 ( .A1(n62477), .A2(n59708), .B(n60261), .Y(
        n77918) );
  NOR2xp33_ASAP7_75t_SL U67076 ( .A(n3088), .B(n61318), .Y(n77997) );
  NOR2xp33_ASAP7_75t_SL U67077 ( .A(n60197), .B(n60202), .Y(n60295) );
  INVx1_ASAP7_75t_SL U67078 ( .A(n60207), .Y(n60293) );
  NOR2xp33_ASAP7_75t_SL U67079 ( .A(n1879), .B(n59574), .Y(n75196) );
  NOR2xp33_ASAP7_75t_SL U67080 ( .A(dbg_stb_i), .B(n59941), .Y(n59942) );
  NOR2xp33_ASAP7_75t_SL U67081 ( .A(dbg_stb_i), .B(n76200), .Y(n59939) );
  NOR2xp33_ASAP7_75t_SL U67082 ( .A(dbg_stb_i), .B(n76204), .Y(n59937) );
  NOR2xp33_ASAP7_75t_SL U67083 ( .A(n74834), .B(n66218), .Y(n74164) );
  INVx1_ASAP7_75t_SL U67084 ( .A(n76976), .Y(n74894) );
  NOR2xp33_ASAP7_75t_SL U67085 ( .A(n69301), .B(n69300), .Y(n69302) );
  INVxp33_ASAP7_75t_SRAM U67086 ( .A(n68850), .Y(n68851) );
  NOR3xp33_ASAP7_75t_SL U67087 ( .A(n62974), .B(n62985), .C(n62973), .Y(n62976) );
  AO22x1_ASAP7_75t_SL U67088 ( .A1(n57463), .A2(n66792), .B1(n66791), .B2(
        n67464), .Y(n58486) );
  NAND2xp33_ASAP7_75t_SRAM U67089 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B(
        n70387), .Y(n70532) );
  NOR2xp33_ASAP7_75t_SL U67090 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[32]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[31]), .Y(n65658) );
  AOI31xp33_ASAP7_75t_SL U67091 ( .A1(n74816), .A2(
        or1200_cpu_or1200_fpu_a_is_inf), .A3(or1200_cpu_or1200_fpu_b_is_inf), 
        .B(or1200_cpu_or1200_fpu_fpu_op_r_1_), .Y(n74819) );
  NOR2xp33_ASAP7_75t_SL U67092 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .B(
        n73040), .Y(n73021) );
  NOR2xp33_ASAP7_75t_SL U67093 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_), 
        .B(n71630), .Y(n71497) );
  NOR2xp33_ASAP7_75t_SL U67094 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_35_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_36_), 
        .Y(n71583) );
  NOR2xp33_ASAP7_75t_SL U67095 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_), 
        .Y(n71628) );
  XOR2xp5_ASAP7_75t_SL U67096 ( .A(n78150), .B(n78149), .Y(n78153) );
  NOR2xp33_ASAP7_75t_SL U67097 ( .A(n72891), .B(n72912), .Y(n72933) );
  OR2x2_ASAP7_75t_SL U67098 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_), .Y(n72614) );
  NOR2xp33_ASAP7_75t_SL U67099 ( .A(n70069), .B(n70076), .Y(n2269) );
  AOI211xp5_ASAP7_75t_SL U67100 ( .A1(n61508), .A2(n61875), .B(n75225), .C(
        n61871), .Y(n75588) );
  NOR2xp33_ASAP7_75t_SL U67101 ( .A(n60788), .B(n63574), .Y(n62535) );
  NOR4xp25_ASAP7_75t_SL U67102 ( .A(n60857), .B(n64302), .C(n64837), .D(n64784), .Y(n63583) );
  NOR2xp33_ASAP7_75t_SL U67103 ( .A(n76896), .B(n76900), .Y(n75665) );
  NOR2xp33_ASAP7_75t_SL U67104 ( .A(n63888), .B(n63887), .Y(n65084) );
  OR2x2_ASAP7_75t_SL U67105 ( .A(n75872), .B(n64858), .Y(n75882) );
  NOR2xp33_ASAP7_75t_SL U67106 ( .A(n69937), .B(n70103), .Y(n69681) );
  NOR2xp33_ASAP7_75t_SL U67107 ( .A(n69650), .B(n70103), .Y(n69653) );
  INVxp33_ASAP7_75t_SRAM U67108 ( .A(n69773), .Y(n69610) );
  NOR2xp33_ASAP7_75t_SL U67109 ( .A(n64324), .B(n64282), .Y(n77128) );
  NOR2xp33_ASAP7_75t_SL U67110 ( .A(n76503), .B(n76498), .Y(n76326) );
  XNOR2xp5_ASAP7_75t_SL U67111 ( .A(n74776), .B(n61972), .Y(n64757) );
  NOR2xp33_ASAP7_75t_SL U67112 ( .A(n71229), .B(n71228), .Y(n71376) );
  INVxp33_ASAP7_75t_SRAM U67113 ( .A(n68756), .Y(n68764) );
  NOR2xp33_ASAP7_75t_SL U67114 ( .A(n59881), .B(n60293), .Y(n60194) );
  NOR2xp33_ASAP7_75t_SL U67115 ( .A(dbg_stb_i), .B(n76201), .Y(n59930) );
  NAND2xp33_ASAP7_75t_SRAM U67116 ( .A(n2496), .B(n59568), .Y(n76201) );
  NOR2xp33_ASAP7_75t_SL U67117 ( .A(dbg_stb_i), .B(n59922), .Y(n59923) );
  NOR2xp33_ASAP7_75t_SL U67118 ( .A(n74158), .B(n74055), .Y(n74209) );
  NOR2xp33_ASAP7_75t_SL U67119 ( .A(n69233), .B(n69230), .Y(n69239) );
  XOR2xp5_ASAP7_75t_SL U67120 ( .A(n67166), .B(n67165), .Y(n67167) );
  AOI22xp33_ASAP7_75t_SRAM U67121 ( .A1(n53298), .A2(n66480), .B1(n67861), 
        .B2(n66348), .Y(n66345) );
  NAND2xp33_ASAP7_75t_SRAM U67122 ( .A(n59505), .B(n67850), .Y(n62834) );
  NAND2xp33_ASAP7_75t_SRAM U67123 ( .A(n53219), .B(n62625), .Y(n62626) );
  NOR2xp33_ASAP7_75t_SL U67124 ( .A(n63214), .B(n59515), .Y(n63112) );
  AOI211xp5_ASAP7_75t_SL U67125 ( .A1(n59656), .A2(n67146), .B(n57505), .C(
        n64685), .Y(n64449) );
  NOR2xp33_ASAP7_75t_SL U67126 ( .A(n57181), .B(n62611), .Y(n58889) );
  INVx1_ASAP7_75t_SL U67127 ( .A(n76430), .Y(n66249) );
  INVx1_ASAP7_75t_SL U67128 ( .A(n74817), .Y(n74744) );
  NOR2xp33_ASAP7_75t_SL U67129 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .Y(
        n70386) );
  OAI22xp33_ASAP7_75t_SRAM U67130 ( .A1(n59706), .A2(n77787), .B1(n57083), 
        .B2(n1262), .Y(n1263) );
  O2A1O1Ixp5_ASAP7_75t_SL U67131 ( .A1(n72303), .A2(n72546), .B(n72302), .C(
        n58599), .Y(n72304) );
  NOR2xp33_ASAP7_75t_SL U67132 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_2_), .B(
        n71772), .Y(n72093) );
  AND2x2_ASAP7_75t_SL U67133 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .B(
        n71894), .Y(n58611) );
  NOR2xp33_ASAP7_75t_SL U67134 ( .A(n65595), .B(n66090), .Y(n65654) );
  INVx1_ASAP7_75t_SL U67135 ( .A(n70081), .Y(n69902) );
  NOR2xp33_ASAP7_75t_SL U67136 ( .A(n78349), .B(n70021), .Y(n69808) );
  AOI211xp5_ASAP7_75t_SL U67137 ( .A1(n66022), .A2(n65977), .B(n65923), .C(
        n65922), .Y(n65924) );
  AOI211xp5_ASAP7_75t_SL U67138 ( .A1(n57194), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[10]), .B(n65700), 
        .C(n65699), .Y(n65965) );
  OAI21xp33_ASAP7_75t_SRAM U67139 ( .A1(n65761), .A2(n65808), .B(n65686), .Y(
        n65840) );
  NOR2xp33_ASAP7_75t_SL U67140 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_0_), .B(
        n74814), .Y(n74815) );
  NOR2xp33_ASAP7_75t_SL U67141 ( .A(n72848), .B(n72840), .Y(n72762) );
  NOR2xp33_ASAP7_75t_SL U67142 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_24_), 
        .Y(n71629) );
  NAND2xp5_ASAP7_75t_SL U67143 ( .A(n2456), .B(n2455), .Y(n70530) );
  XNOR2xp5_ASAP7_75t_SL U67144 ( .A(or1200_cpu_or1200_mult_mac_n301), .B(
        or1200_cpu_or1200_mult_mac_n155), .Y(n63353) );
  XNOR2xp5_ASAP7_75t_SL U67145 ( .A(or1200_cpu_or1200_mult_mac_n345), .B(
        or1200_cpu_or1200_mult_mac_n199), .Y(n75020) );
  NOR2xp33_ASAP7_75t_SL U67146 ( .A(n78362), .B(n59626), .Y(n72647) );
  NOR2xp33_ASAP7_75t_SL U67147 ( .A(n1590), .B(n59689), .Y(n64256) );
  AOI22xp33_ASAP7_75t_SRAM U67148 ( .A1(n1470), .A2(n76712), .B1(n76711), .B2(
        n1163), .Y(n62316) );
  AOI211xp5_ASAP7_75t_SL U67149 ( .A1(n77128), .A2(n77643), .B(n60884), .C(
        n60883), .Y(n60885) );
  AOI21xp33_ASAP7_75t_SRAM U67150 ( .A1(n77039), .A2(n63485), .B(n60821), .Y(
        n60822) );
  OAI22xp33_ASAP7_75t_SRAM U67151 ( .A1(n1458), .A2(n77034), .B1(n1153), .B2(
        n77033), .Y(n60821) );
  NOR2xp33_ASAP7_75t_SL U67152 ( .A(n63567), .B(n73941), .Y(n60801) );
  NOR2xp33_ASAP7_75t_SL U67153 ( .A(n1787), .B(n59679), .Y(n76560) );
  AOI211xp5_ASAP7_75t_SL U67154 ( .A1(n77125), .A2(n73933), .B(n61717), .C(
        n61716), .Y(n61738) );
  O2A1O1Ixp5_ASAP7_75t_SL U67155 ( .A1(n3132), .A2(n69344), .B(n57073), .C(
        n62472), .Y(n62474) );
  NOR2xp33_ASAP7_75t_SL U67156 ( .A(n75872), .B(n61346), .Y(n77096) );
  NOR2xp33_ASAP7_75t_SL U67157 ( .A(n61832), .B(n61721), .Y(n62455) );
  NOR2xp33_ASAP7_75t_SL U67158 ( .A(n64205), .B(n64204), .Y(n64215) );
  OAI22xp33_ASAP7_75t_SRAM U67159 ( .A1(or1200_cpu_or1200_except_n652), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n538), .B2(n77032), .Y(n64204)
         );
  OAI22xp33_ASAP7_75t_SRAM U67160 ( .A1(or1200_cpu_or1200_except_n238), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n136), .B2(n57102), .Y(n64205)
         );
  NAND3xp33_ASAP7_75t_SL U67161 ( .A(n69405), .B(n78382), .C(n78373), .Y(
        n69409) );
  NOR2xp33_ASAP7_75t_SL U67162 ( .A(or1200_cpu_or1200_mult_mac_n347), .B(
        n75692), .Y(n76883) );
  NOR2xp33_ASAP7_75t_SL U67163 ( .A(or1200_cpu_or1200_mult_mac_n189), .B(
        n65140), .Y(n65164) );
  NOR2xp33_ASAP7_75t_SL U67164 ( .A(or1200_cpu_or1200_mult_mac_n185), .B(
        n65124), .Y(n65142) );
  NOR2xp33_ASAP7_75t_SL U67165 ( .A(or1200_cpu_or1200_mult_mac_n177), .B(
        n63891), .Y(n64172) );
  NOR2xp33_ASAP7_75t_SL U67166 ( .A(or1200_cpu_or1200_mult_mac_n161), .B(
        n63422), .Y(n63531) );
  NOR2xp33_ASAP7_75t_SL U67167 ( .A(or1200_cpu_or1200_mult_mac_n163), .B(
        n63453), .Y(n63530) );
  NOR2xp33_ASAP7_75t_SL U67168 ( .A(or1200_cpu_or1200_mult_mac_n153), .B(
        n63334), .Y(n63394) );
  NOR2xp33_ASAP7_75t_SL U67169 ( .A(or1200_cpu_or1200_mult_mac_n151), .B(
        n63315), .Y(n63397) );
  NOR2xp33_ASAP7_75t_SL U67170 ( .A(or1200_cpu_or1200_mult_mac_n289), .B(
        n63272), .Y(n63390) );
  NOR2xp33_ASAP7_75t_SL U67171 ( .A(or1200_cpu_or1200_mult_mac_n159), .B(
        n63409), .Y(n63423) );
  INVxp33_ASAP7_75t_SRAM U67172 ( .A(n69052), .Y(n69055) );
  AOI211xp5_ASAP7_75t_SL U67173 ( .A1(n77220), .A2(or1200_cpu_sr_15_), .B(
        n77218), .C(n77146), .Y(or1200_cpu_or1200_except_n253) );
  NOR2xp33_ASAP7_75t_SL U67174 ( .A(n70970), .B(n70974), .Y(n70945) );
  NOR2xp33_ASAP7_75t_SL U67175 ( .A(n74462), .B(n74221), .Y(n70641) );
  NOR2xp33_ASAP7_75t_SL U67176 ( .A(n70045), .B(n70103), .Y(n69705) );
  NOR2xp33_ASAP7_75t_SL U67177 ( .A(n69990), .B(n70103), .Y(n69696) );
  NOR2xp33_ASAP7_75t_SL U67178 ( .A(n69666), .B(n70103), .Y(n69669) );
  O2A1O1Ixp5_ASAP7_75t_SL U67179 ( .A1(n57185), .A2(n73244), .B(n73243), .C(
        n73242), .Y(n73245) );
  O2A1O1Ixp5_ASAP7_75t_SL U67180 ( .A1(n73483), .A2(n59631), .B(n73233), .C(
        n73232), .Y(n73482) );
  O2A1O1Ixp5_ASAP7_75t_SL U67181 ( .A1(n73185), .A2(n57185), .B(n73184), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[13]), .Y(
        n73186) );
  OAI22xp33_ASAP7_75t_SRAM U67182 ( .A1(or1200_cpu_or1200_if_insn_saved[16]), 
        .A2(n61042), .B1(n61152), .B2(n77454), .Y(n60508) );
  AOI22xp33_ASAP7_75t_SRAM U67183 ( .A1(n60686), .A2(n62000), .B1(n60489), 
        .B2(n77566), .Y(n60342) );
  NOR2xp33_ASAP7_75t_SL U67184 ( .A(n1571), .B(n57120), .Y(n61976) );
  XNOR2xp5_ASAP7_75t_SL U67185 ( .A(n75628), .B(n61966), .Y(n64185) );
  NOR2xp33_ASAP7_75t_SL U67186 ( .A(n61321), .B(n62462), .Y(n60774) );
  NAND2xp33_ASAP7_75t_SRAM U67187 ( .A(n57120), .B(n64930), .Y(n61945) );
  AND2x2_ASAP7_75t_SL U67188 ( .A(n74497), .B(n3143), .Y(n74738) );
  AND2x2_ASAP7_75t_SL U67189 ( .A(n60327), .B(n77359), .Y(n78022) );
  AND2x2_ASAP7_75t_SL U67190 ( .A(n60327), .B(n77359), .Y(n59497) );
  NOR2xp33_ASAP7_75t_SL U67191 ( .A(n77833), .B(n60326), .Y(n60327) );
  NOR2xp33_ASAP7_75t_SL U67192 ( .A(n77456), .B(n77359), .Y(n76846) );
  NOR2xp33_ASAP7_75t_SL U67193 ( .A(n57090), .B(n77954), .Y(n60523) );
  NOR2xp33_ASAP7_75t_SL U67194 ( .A(n3121), .B(n77276), .Y(n60426) );
  NOR2xp33_ASAP7_75t_SL U67195 ( .A(n63956), .B(n63944), .Y(n4133) );
  NOR2xp33_ASAP7_75t_SL U67196 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[5]), .B(
        n70589), .Y(n70602) );
  NOR2xp33_ASAP7_75t_SL U67197 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[1]), .B(
        n70572), .Y(n70580) );
  NOR2xp33_ASAP7_75t_SL U67198 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[0]), .B(
        n70570), .Y(n70572) );
  O2A1O1Ixp5_ASAP7_75t_SL U67199 ( .A1(n59526), .A2(n70869), .B(n70845), .C(
        n70847), .Y(n70859) );
  NOR2xp33_ASAP7_75t_SL U67200 ( .A(n76027), .B(n76060), .Y(n76032) );
  NOR2xp33_ASAP7_75t_SL U67201 ( .A(n60175), .B(n57160), .Y(n65193) );
  NOR2xp33_ASAP7_75t_SL U67202 ( .A(n1868), .B(n57124), .Y(n60019) );
  NOR2xp33_ASAP7_75t_SL U67203 ( .A(n59703), .B(n76844), .Y(n59968) );
  NOR3xp33_ASAP7_75t_SL U67204 ( .A(n60669), .B(n60668), .C(n61647), .Y(n75486) );
  XNOR2xp5_ASAP7_75t_SL U67205 ( .A(or1200_dc_top_tag_2_), .B(n77017), .Y(
        n59791) );
  NOR2xp33_ASAP7_75t_SL U67206 ( .A(n59530), .B(n1885), .Y(n69357) );
  NOR2xp33_ASAP7_75t_SL U67207 ( .A(n59944), .B(n60557), .Y(n59946) );
  INVx1_ASAP7_75t_SL U67208 ( .A(n60554), .Y(n62205) );
  OR2x2_ASAP7_75t_SL U67209 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]), .Y(n65425) );
  XNOR2xp5_ASAP7_75t_SL U67210 ( .A(n57151), .B(n59194), .Y(n59193) );
  NAND2xp33_ASAP7_75t_SRAM U67211 ( .A(n59505), .B(n57274), .Y(n62627) );
  XNOR2xp5_ASAP7_75t_SL U67212 ( .A(n59609), .B(n67228), .Y(n62956) );
  XNOR2xp5_ASAP7_75t_SL U67213 ( .A(n67343), .B(n59603), .Y(n63080) );
  AOI22xp33_ASAP7_75t_SRAM U67214 ( .A1(n67635), .A2(n68019), .B1(n57394), 
        .B2(n67242), .Y(n66612) );
  XNOR2xp5_ASAP7_75t_SL U67215 ( .A(n58726), .B(n68289), .Y(n68290) );
  NOR2xp33_ASAP7_75t_SL U67216 ( .A(n67343), .B(n67560), .Y(n58698) );
  INVxp33_ASAP7_75t_SRAM U67217 ( .A(n59578), .Y(n74799) );
  AOI21xp33_ASAP7_75t_SRAM U67218 ( .A1(n58248), .A2(n59555), .B(n59571), .Y(
        n58972) );
  INVxp33_ASAP7_75t_SRAM U67219 ( .A(n59544), .Y(n78004) );
  NAND2xp33_ASAP7_75t_SRAM U67220 ( .A(n59530), .B(n59529), .Y(n65030) );
  AOI22xp33_ASAP7_75t_SRAM U67221 ( .A1(n72347), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_32_), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_), .B2(n72364), .Y(n72101) );
  AOI22xp33_ASAP7_75t_SRAM U67222 ( .A1(n72347), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_36_), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_), .B2(n72364), .Y(n72022) );
  O2A1O1Ixp5_ASAP7_75t_SL U67223 ( .A1(n70086), .A2(n70085), .B(n70166), .C(
        n70084), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[23]) );
  O2A1O1Ixp5_ASAP7_75t_SL U67224 ( .A1(n70018), .A2(n69467), .B(n69466), .C(
        n69465), .Y(n69509) );
  O2A1O1Ixp5_ASAP7_75t_SL U67225 ( .A1(n72882), .A2(n73042), .B(n72881), .C(
        n72880), .Y(n72884) );
  NOR2xp33_ASAP7_75t_SL U67226 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_25_), 
        .Y(n71627) );
  NOR2xp33_ASAP7_75t_SL U67227 ( .A(n78380), .B(n57190), .Y(n72668) );
  NOR2xp33_ASAP7_75t_SL U67228 ( .A(n78360), .B(n59626), .Y(n72653) );
  O2A1O1Ixp5_ASAP7_75t_SL U67229 ( .A1(n61642), .A2(n61641), .B(n57126), .C(
        n61640), .Y(n61660) );
  O2A1O1Ixp5_ASAP7_75t_SL U67230 ( .A1(n61235), .A2(n61234), .B(n57126), .C(
        n61233), .Y(n61240) );
  XNOR2xp5_ASAP7_75t_SL U67231 ( .A(n75815), .B(n75814), .Y(n75881) );
  OR2x2_ASAP7_75t_SL U67232 ( .A(n3117), .B(or1200_cpu_or1200_except_n646), 
        .Y(n65225) );
  OR2x2_ASAP7_75t_SL U67233 ( .A(or1200_cpu_or1200_mult_mac_n359), .B(
        or1200_cpu_or1200_mult_mac_n213), .Y(n68935) );
  XOR2xp5_ASAP7_75t_SL U67234 ( .A(or1200_cpu_or1200_mult_mac_n157), .B(
        or1200_cpu_or1200_mult_mac_n303), .Y(n63426) );
  NAND4xp25_ASAP7_75t_SL U67235 ( .A(n69051), .B(n69050), .C(n69049), .D(
        n69048), .Y(n69064) );
  NOR2xp33_ASAP7_75t_SL U67236 ( .A(n63261), .B(n68810), .Y(n63266) );
  AOI211xp5_ASAP7_75t_SL U67237 ( .A1(or1200_cpu_rf_datab[31]), .A2(n57091), 
        .B(n77184), .C(n61991), .Y(n61992) );
  OAI22xp33_ASAP7_75t_SRAM U67238 ( .A1(n2958), .A2(n59679), .B1(n59582), .B2(
        n59689), .Y(n61991) );
  NOR4xp25_ASAP7_75t_SL U67239 ( .A(n61887), .B(n61886), .C(n61885), .D(n61884), .Y(n77104) );
  NOR4xp25_ASAP7_75t_SL U67240 ( .A(n61883), .B(n61882), .C(n61881), .D(n61880), .Y(n75590) );
  AOI22xp33_ASAP7_75t_SRAM U67241 ( .A1(n75708), .A2(n75890), .B1(n75861), 
        .B2(n77089), .Y(n61879) );
  NOR2xp33_ASAP7_75t_SL U67242 ( .A(or1200_cpu_epcr_31_), .B(n57170), .Y(
        n61843) );
  XNOR2xp5_ASAP7_75t_SL U67243 ( .A(n61837), .B(n75749), .Y(n61902) );
  NAND2xp33_ASAP7_75t_SRAM U67244 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[2]), .B(n73605), 
        .Y(n73600) );
  NOR2xp33_ASAP7_75t_SL U67245 ( .A(n73524), .B(n73523), .Y(n73526) );
  NOR2xp33_ASAP7_75t_SL U67246 ( .A(n75872), .B(n75863), .Y(n75731) );
  NOR2xp33_ASAP7_75t_SL U67247 ( .A(n59709), .B(n60846), .Y(n62371) );
  OR2x2_ASAP7_75t_SL U67248 ( .A(n2567), .B(n2807), .Y(n58607) );
  NOR2xp33_ASAP7_75t_SL U67249 ( .A(n70640), .B(n74459), .Y(n74715) );
  NOR2xp33_ASAP7_75t_SL U67250 ( .A(n70639), .B(n70638), .Y(n74459) );
  NOR2xp33_ASAP7_75t_SL U67251 ( .A(n69958), .B(n69961), .Y(n69964) );
  NOR3xp33_ASAP7_75t_SL U67252 ( .A(n65261), .B(n65260), .C(n65259), .Y(n65320) );
  NOR2xp33_ASAP7_75t_SL U67253 ( .A(n78005), .B(n75863), .Y(n62362) );
  NOR2xp33_ASAP7_75t_SL U67254 ( .A(n59708), .B(n64218), .Y(n76763) );
  NOR2xp33_ASAP7_75t_SL U67255 ( .A(n59709), .B(n75328), .Y(n77076) );
  XNOR2xp5_ASAP7_75t_SL U67256 ( .A(n73246), .B(n73245), .Y(n73471) );
  O2A1O1Ixp5_ASAP7_75t_SL U67257 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[12]), .A2(
        n59630), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[12]), .C(
        n73181), .Y(n73182) );
  OR2x2_ASAP7_75t_SL U67258 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_19_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_18_), .Y(n69404) );
  NOR2xp33_ASAP7_75t_SL U67259 ( .A(n77014), .B(n77016), .Y(n77149) );
  NOR2xp33_ASAP7_75t_SL U67260 ( .A(n59579), .B(n78327), .Y(n74025) );
  INVxp33_ASAP7_75t_SRAM U67261 ( .A(n73990), .Y(n73993) );
  NOR2xp33_ASAP7_75t_SL U67262 ( .A(n73966), .B(n76346), .Y(n74019) );
  OAI21xp33_ASAP7_75t_SRAM U67263 ( .A1(n59528), .A2(n77735), .B(n73965), .Y(
        n76346) );
  NOR2xp33_ASAP7_75t_SL U67264 ( .A(n59582), .B(n76486), .Y(n76427) );
  NOR2xp33_ASAP7_75t_SL U67265 ( .A(n61323), .B(n60776), .Y(n62463) );
  XOR2xp5_ASAP7_75t_SL U67266 ( .A(n61940), .B(n59535), .Y(n75310) );
  NOR2xp33_ASAP7_75t_SL U67267 ( .A(n74121), .B(n75297), .Y(n75298) );
  INVxp33_ASAP7_75t_SRAM U67268 ( .A(n69368), .Y(n69353) );
  AND2x2_ASAP7_75t_SL U67269 ( .A(n77052), .B(n77163), .Y(n69370) );
  NOR2xp33_ASAP7_75t_SL U67270 ( .A(n63700), .B(n63701), .Y(n69352) );
  NOR2xp33_ASAP7_75t_SL U67271 ( .A(n73893), .B(n73892), .Y(n74069) );
  NAND3xp33_ASAP7_75t_SL U67272 ( .A(n78249), .B(n78248), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_2_), 
        .Y(n73857) );
  NAND2xp33_ASAP7_75t_SRAM U67273 ( .A(n59662), .B(n76185), .Y(n76192) );
  AOI211xp5_ASAP7_75t_SL U67274 ( .A1(n59522), .A2(n71219), .B(n70884), .C(
        n70883), .Y(n71046) );
  XNOR2xp5_ASAP7_75t_SL U67275 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_output_o_31_), .Y(
        n74289) );
  NOR2xp33_ASAP7_75t_SL U67276 ( .A(n2779), .B(n60281), .Y(n77354) );
  NOR2xp33_ASAP7_75t_SL U67277 ( .A(n58401), .B(n62149), .Y(n60300) );
  AOI211xp5_ASAP7_75t_SL U67278 ( .A1(n57198), .A2(n60020), .B(n60019), .C(
        n60018), .Y(n60021) );
  AOI211xp5_ASAP7_75t_SL U67279 ( .A1(n57198), .A2(n60005), .B(n60004), .C(
        n60003), .Y(n60006) );
  NOR2xp33_ASAP7_75t_SL U67280 ( .A(n59550), .B(n57124), .Y(n60004) );
  AND2x2_ASAP7_75t_SL U67281 ( .A(n59992), .B(n59991), .Y(n77257) );
  AOI31xp33_ASAP7_75t_SL U67282 ( .A1(n75765), .A2(n59493), .A3(n60306), .B(
        n76503), .Y(n59962) );
  NOR2xp33_ASAP7_75t_SL U67283 ( .A(n60294), .B(n77765), .Y(n60297) );
  OAI22xp33_ASAP7_75t_SRAM U67284 ( .A1(n60421), .A2(n77358), .B1(n2757), .B2(
        or1200_cpu_or1200_if_insn_saved[28]), .Y(n60314) );
  OAI22xp33_ASAP7_75t_SRAM U67285 ( .A1(n60421), .A2(n60321), .B1(n2757), .B2(
        or1200_cpu_or1200_if_insn_saved[26]), .Y(n60322) );
  AOI21xp33_ASAP7_75t_SRAM U67286 ( .A1(n59564), .A2(n2514), .B(dbg_stb_i), 
        .Y(n60223) );
  XNOR2xp5_ASAP7_75t_SL U67287 ( .A(or1200_dc_top_tag_9_), .B(n75423), .Y(
        n59789) );
  NOR2xp33_ASAP7_75t_SL U67288 ( .A(n75439), .B(n59839), .Y(n75423) );
  XNOR2xp5_ASAP7_75t_SL U67289 ( .A(n1921), .B(n59579), .Y(n60207) );
  AND2x2_ASAP7_75t_SL U67290 ( .A(n1882), .B(n59528), .Y(n69366) );
  NOR2xp33_ASAP7_75t_SL U67291 ( .A(n1909), .B(n59563), .Y(n69356) );
  AND2x2_ASAP7_75t_SL U67292 ( .A(n1885), .B(n59530), .Y(n59864) );
  AND2x2_ASAP7_75t_SL U67293 ( .A(n1909), .B(n59563), .Y(n74041) );
  NOR2xp33_ASAP7_75t_SL U67294 ( .A(n1906), .B(n59577), .Y(n75439) );
  NOR2xp33_ASAP7_75t_SL U67295 ( .A(n1924), .B(n59572), .Y(n59850) );
  NOR2xp33_ASAP7_75t_SL U67296 ( .A(n2039), .B(n59560), .Y(n77148) );
  NOR2xp33_ASAP7_75t_SL U67297 ( .A(n2461), .B(n59557), .Y(n76205) );
  XNOR2xp5_ASAP7_75t_SL U67298 ( .A(n59568), .B(n2496), .Y(n76683) );
  AOI211xp5_ASAP7_75t_SL U67299 ( .A1(n76202), .A2(n76199), .B(n76198), .C(
        n76616), .Y(n76613) );
  NOR2xp33_ASAP7_75t_SL U67300 ( .A(n59545), .B(n2157), .Y(n76198) );
  NOR2xp33_ASAP7_75t_SL U67301 ( .A(n2169), .B(n59559), .Y(n76202) );
  NOR2xp33_ASAP7_75t_SL U67302 ( .A(n2544), .B(n59540), .Y(n76546) );
  NOR2xp33_ASAP7_75t_SL U67303 ( .A(n2073), .B(n59570), .Y(n59843) );
  NOR2xp33_ASAP7_75t_SL U67304 ( .A(n2095), .B(n59541), .Y(n76548) );
  NAND2xp33_ASAP7_75t_SRAM U67305 ( .A(n2119), .B(n59569), .Y(n75775) );
  NOR2xp33_ASAP7_75t_SL U67306 ( .A(n75779), .B(n58539), .Y(n75774) );
  AND2x2_ASAP7_75t_SL U67307 ( .A(n2107), .B(n59542), .Y(n58539) );
  NOR2xp33_ASAP7_75t_SL U67308 ( .A(n2107), .B(n59542), .Y(n75779) );
  AND2x2_ASAP7_75t_SL U67309 ( .A(n1903), .B(n59531), .Y(n59855) );
  AND2x2_ASAP7_75t_SL U67310 ( .A(n1897), .B(n59537), .Y(n59821) );
  NOR2xp33_ASAP7_75t_SL U67311 ( .A(n1897), .B(n59537), .Y(n74118) );
  AND2x2_ASAP7_75t_SL U67312 ( .A(n1906), .B(n59577), .Y(n59839) );
  NAND3xp33_ASAP7_75t_SL U67313 ( .A(n61131), .B(n59946), .C(n60548), .Y(
        n60826) );
  AOI31xp33_ASAP7_75t_SL U67314 ( .A1(n60595), .A2(n59934), .A3(n59932), .B(
        n59933), .Y(n60545) );
  AND2x2_ASAP7_75t_SL U67315 ( .A(n2131), .B(n59571), .Y(n59934) );
  AOI31xp33_ASAP7_75t_SL U67316 ( .A1(n2532), .A2(n59565), .A3(n78439), .B(
        n59920), .Y(n77953) );
  OR2x2_ASAP7_75t_SL U67317 ( .A(n74219), .B(n74218), .Y(n77195) );
  XNOR2xp5_ASAP7_75t_SL U67318 ( .A(n66519), .B(n66518), .Y(n66521) );
  NOR2xp33_ASAP7_75t_SL U67319 ( .A(n57108), .B(n62822), .Y(n62824) );
  NAND2xp33_ASAP7_75t_SRAM U67320 ( .A(n75927), .B(n67428), .Y(n62802) );
  NAND2xp33_ASAP7_75t_SRAM U67321 ( .A(n59656), .B(n53219), .Y(n62862) );
  NOR2xp33_ASAP7_75t_SL U67322 ( .A(n67343), .B(n67232), .Y(n62820) );
  XNOR2xp5_ASAP7_75t_SL U67323 ( .A(n63012), .B(n62985), .Y(n62986) );
  NAND2xp33_ASAP7_75t_SRAM U67324 ( .A(n62831), .B(n53219), .Y(n62832) );
  XNOR2xp5_ASAP7_75t_SL U67325 ( .A(n57257), .B(n59511), .Y(n62692) );
  XOR2xp5_ASAP7_75t_SL U67326 ( .A(n66813), .B(n66815), .Y(n59075) );
  NOR2xp33_ASAP7_75t_SL U67327 ( .A(n53251), .B(n59639), .Y(n66664) );
  NAND2xp33_ASAP7_75t_SRAM U67328 ( .A(n59657), .B(n58809), .Y(n68125) );
  NAND2xp33_ASAP7_75t_SRAM U67329 ( .A(n59711), .B(n59441), .Y(n64779) );
  OAI21xp33_ASAP7_75t_SRAM U67330 ( .A1(n53275), .A2(n75894), .B(n75047), .Y(
        n75074) );
  AOI22xp33_ASAP7_75t_SRAM U67331 ( .A1(n72347), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_), 
        .B2(n72364), .Y(n72359) );
  NOR2xp33_ASAP7_75t_SL U67332 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[24]), .Y(n65552) );
  OR2x2_ASAP7_75t_SL U67333 ( .A(n69948), .B(n69557), .Y(n70035) );
  O2A1O1Ixp5_ASAP7_75t_SL U67334 ( .A1(n65398), .A2(n65374), .B(n65373), .C(
        n65372), .Y(n65376) );
  OAI21xp33_ASAP7_75t_SRAM U67335 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_18_), .A2(n59629), .B(
        n72707), .Y(n1646) );
  OAI21xp33_ASAP7_75t_SRAM U67336 ( .A1(n59629), .A2(n73046), .B(n73045), .Y(
        n1722) );
  OAI21xp33_ASAP7_75t_SRAM U67337 ( .A1(n59629), .A2(n72750), .B(n72749), .Y(
        n1771) );
  NOR2xp33_ASAP7_75t_SL U67338 ( .A(n71676), .B(n71638), .Y(n71719) );
  NOR2xp33_ASAP7_75t_SL U67339 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_), 
        .Y(n71568) );
  NOR2xp33_ASAP7_75t_SL U67340 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_0_), .B(n69376), .Y(
        n70281) );
  NOR2xp33_ASAP7_75t_SL U67341 ( .A(n70255), .B(n70502), .Y(n70280) );
  NOR2xp33_ASAP7_75t_SL U67342 ( .A(n70766), .B(n70785), .Y(n70775) );
  OAI22xp33_ASAP7_75t_SRAM U67343 ( .A1(n70522), .A2(n70422), .B1(n57081), 
        .B2(n70045), .Y(n70053) );
  NOR2xp33_ASAP7_75t_SL U67344 ( .A(n1510), .B(n77685), .Y(n77681) );
  NAND2xp33_ASAP7_75t_SRAM U67345 ( .A(n2440), .B(n74662), .Y(n74690) );
  O2A1O1Ixp5_ASAP7_75t_SL U67346 ( .A1(n64794), .A2(n64793), .B(n57126), .C(
        n64792), .Y(n64795) );
  O2A1O1Ixp5_ASAP7_75t_SL U67347 ( .A1(n70158), .A2(n70157), .B(n70172), .C(
        n70156), .Y(n70161) );
  OAI22xp33_ASAP7_75t_SRAM U67348 ( .A1(n70498), .A2(n70422), .B1(n57081), 
        .B2(n70088), .Y(n70096) );
  NOR3xp33_ASAP7_75t_SL U67349 ( .A(n73611), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[3]), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[4]), .Y(n73590)
         );
  NOR4xp25_ASAP7_75t_SL U67350 ( .A(n62351), .B(n62347), .C(n62346), .D(n62350), .Y(n60810) );
  OR2x2_ASAP7_75t_SL U67351 ( .A(or1200_cpu_or1200_except_n494), .B(
        or1200_cpu_or1200_except_n496), .Y(n61651) );
  NAND4xp25_ASAP7_75t_SL U67352 ( .A(n70632), .B(n70631), .C(n70630), .D(
        n70629), .Y(n74461) );
  NOR2xp33_ASAP7_75t_SL U67353 ( .A(n2865), .B(n2854), .Y(n70629) );
  NOR2xp33_ASAP7_75t_SL U67354 ( .A(n1564), .B(n1600), .Y(n70630) );
  NOR2xp33_ASAP7_75t_SL U67355 ( .A(n2009), .B(n2900), .Y(n70631) );
  NOR2xp33_ASAP7_75t_SL U67356 ( .A(n2860), .B(n1582), .Y(n70632) );
  AOI21xp33_ASAP7_75t_SRAM U67357 ( .A1(n69791), .A2(n69789), .B(n69617), .Y(
        n69618) );
  INVxp33_ASAP7_75t_SRAM U67358 ( .A(n69748), .Y(n69609) );
  NOR2xp33_ASAP7_75t_SL U67359 ( .A(n2191), .B(n77567), .Y(n60495) );
  NAND4xp25_ASAP7_75t_SL U67360 ( .A(n2854), .B(n2860), .C(n2900), .D(n2865), 
        .Y(n65259) );
  AND2x2_ASAP7_75t_SL U67361 ( .A(n1600), .B(n2009), .Y(n65258) );
  NAND2xp33_ASAP7_75t_SRAM U67362 ( .A(n59080), .B(n60629), .Y(n60630) );
  NOR2xp33_ASAP7_75t_SL U67363 ( .A(n73415), .B(n73414), .Y(n73438) );
  O2A1O1Ixp5_ASAP7_75t_SL U67364 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[13]), .A2(
        n59631), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[13]), .C(
        n73186), .Y(n73187) );
  NOR2xp33_ASAP7_75t_SL U67365 ( .A(n2616), .B(n57072), .Y(n61153) );
  XNOR2xp5_ASAP7_75t_SL U67366 ( .A(n62466), .B(n62465), .Y(n76300) );
  O2A1O1Ixp5_ASAP7_75t_SL U67367 ( .A1(n59564), .A2(n60979), .B(n60978), .C(
        n60757), .Y(n61236) );
  XNOR2xp5_ASAP7_75t_SL U67368 ( .A(n77717), .B(n61941), .Y(n61943) );
  NOR2xp33_ASAP7_75t_SL U67369 ( .A(n53455), .B(n57397), .Y(n61941) );
  NAND2xp33_ASAP7_75t_SRAM U67370 ( .A(n53251), .B(n76048), .Y(n76052) );
  NOR2xp33_ASAP7_75t_SL U67371 ( .A(n59527), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_), .Y(
        n72519) );
  NOR3xp33_ASAP7_75t_SL U67372 ( .A(n72517), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_0_), .Y(
        n72523) );
  NOR2xp33_ASAP7_75t_SL U67373 ( .A(n76151), .B(n76150), .Y(n76152) );
  NOR2xp33_ASAP7_75t_SL U67374 ( .A(n751), .B(n59703), .Y(n59988) );
  NOR2xp33_ASAP7_75t_SL U67375 ( .A(n61647), .B(n75478), .Y(n75518) );
  NOR2xp33_ASAP7_75t_SL U67376 ( .A(n57407), .B(n53311), .Y(n61647) );
  NOR2xp33_ASAP7_75t_SL U67377 ( .A(n2035), .B(n62008), .Y(n63719) );
  NAND3xp33_ASAP7_75t_SL U67378 ( .A(n60209), .B(n77418), .C(n59706), .Y(
        n61293) );
  NOR2xp33_ASAP7_75t_SL U67379 ( .A(n74856), .B(n74885), .Y(n74857) );
  O2A1O1Ixp5_ASAP7_75t_SL U67380 ( .A1(n58402), .A2(n57456), .B(n67086), .C(
        n67085), .Y(n67087) );
  XNOR2xp5_ASAP7_75t_SL U67381 ( .A(n63233), .B(n63131), .Y(n63196) );
  NOR2xp33_ASAP7_75t_SL U67382 ( .A(n59653), .B(n59509), .Y(n63810) );
  NOR2xp33_ASAP7_75t_SL U67383 ( .A(n59125), .B(n59042), .Y(n58822) );
  NOR2xp33_ASAP7_75t_SL U67384 ( .A(n59264), .B(n59265), .Y(n59260) );
  INVxp33_ASAP7_75t_SRAM U67385 ( .A(n77910), .Y(n77911) );
  OAI22xp33_ASAP7_75t_SRAM U67386 ( .A1(n71953), .A2(n57208), .B1(n71993), 
        .B2(n71890), .Y(n71893) );
  AOI21xp33_ASAP7_75t_SRAM U67387 ( .A1(n65636), .A2(n65635), .B(n65674), .Y(
        n65637) );
  OAI21xp33_ASAP7_75t_SRAM U67388 ( .A1(n65626), .A2(n65625), .B(n65691), .Y(
        n65641) );
  AOI22xp33_ASAP7_75t_SRAM U67389 ( .A1(n65674), .A2(n66154), .B1(n65639), 
        .B2(n65618), .Y(n65650) );
  INVxp33_ASAP7_75t_SRAM U67390 ( .A(n70080), .Y(n70086) );
  INVx1_ASAP7_75t_SL U67391 ( .A(n58421), .Y(n59687) );
  NOR2xp33_ASAP7_75t_SL U67392 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[5]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[6]), .Y(n65479) );
  NOR2xp33_ASAP7_75t_SL U67393 ( .A(n66195), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n63), .Y(n65476) );
  OAI21xp33_ASAP7_75t_SRAM U67394 ( .A1(n65974), .A2(n65896), .B(n65968), .Y(
        n65899) );
  OAI21xp33_ASAP7_75t_SRAM U67395 ( .A1(n66027), .A2(n65921), .B(n65968), .Y(
        n65890) );
  OAI22xp33_ASAP7_75t_SRAM U67396 ( .A1(n65805), .A2(n58582), .B1(n65804), 
        .B2(n58418), .Y(n65806) );
  AOI22xp33_ASAP7_75t_SRAM U67397 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .A2(n57188), 
        .B1(n57187), .B2(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .Y(n65802) );
  AOI22xp33_ASAP7_75t_SRAM U67398 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[44]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .B2(n57194), .Y(n65803) );
  INVxp33_ASAP7_75t_SRAM U67399 ( .A(n70109), .Y(n69492) );
  OAI21xp33_ASAP7_75t_SRAM U67400 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[29]), .A2(n58571), 
        .B(n65798), .Y(n65799) );
  O2A1O1Ixp5_ASAP7_75t_SL U67401 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .A2(n72234), .B(n72212), .C(n71605), .Y(n71610) );
  OAI22xp33_ASAP7_75t_SRAM U67402 ( .A1(n58418), .A2(n65855), .B1(n65857), 
        .B2(n58571), .Y(n65751) );
  OAI22xp33_ASAP7_75t_SRAM U67403 ( .A1(n65854), .A2(n58419), .B1(n65742), 
        .B2(n58582), .Y(n65752) );
  AOI22xp33_ASAP7_75t_SRAM U67404 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[42]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .B2(n57194), .Y(n65741) );
  AOI22xp33_ASAP7_75t_SRAM U67405 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]), .B2(n57194), .Y(n65866) );
  OAI22xp33_ASAP7_75t_SRAM U67406 ( .A1(n58418), .A2(n65857), .B1(n65856), 
        .B2(n58571), .Y(n65861) );
  OAI22xp33_ASAP7_75t_SRAM U67407 ( .A1(n65855), .A2(n58419), .B1(n65854), 
        .B2(n58582), .Y(n65862) );
  OAI22xp33_ASAP7_75t_SRAM U67408 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .A2(n58582), 
        .B1(n65841), .B2(n65777), .Y(n65764) );
  OAI21xp33_ASAP7_75t_SRAM U67409 ( .A1(n65828), .A2(n65850), .B(n65746), .Y(
        n65747) );
  OAI21xp33_ASAP7_75t_SRAM U67410 ( .A1(n65745), .A2(n65841), .B(n65705), .Y(
        n65807) );
  NOR2xp33_ASAP7_75t_SL U67411 ( .A(n73042), .B(n72962), .Y(n72806) );
  NOR2xp33_ASAP7_75t_SL U67412 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_2_), .B(n70502), .Y(
        n70288) );
  NOR2xp33_ASAP7_75t_SL U67413 ( .A(n78243), .B(n78244), .Y(n72964) );
  NOR2xp33_ASAP7_75t_SL U67414 ( .A(n64327), .B(n64329), .Y(n75459) );
  NOR2xp33_ASAP7_75t_SL U67415 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_5_), .Y(
        n74710) );
  INVxp33_ASAP7_75t_SRAM U67416 ( .A(n76977), .Y(n76975) );
  NOR2xp33_ASAP7_75t_SL U67417 ( .A(n69290), .B(n69274), .Y(n69262) );
  NOR2xp33_ASAP7_75t_SL U67418 ( .A(n69242), .B(n69244), .Y(n74115) );
  NOR2xp33_ASAP7_75t_SL U67419 ( .A(n73953), .B(n76266), .Y(n75801) );
  NAND2xp33_ASAP7_75t_SRAM U67420 ( .A(or1200_cpu_esr[15]), .B(n77048), .Y(
        n77049) );
  OAI22xp33_ASAP7_75t_SRAM U67421 ( .A1(n1456), .A2(n77034), .B1(n1151), .B2(
        n77033), .Y(n77037) );
  AOI22xp33_ASAP7_75t_SRAM U67422 ( .A1(n74609), .A2(n75727), .B1(n75736), 
        .B2(n77715), .Y(n74610) );
  NOR2xp33_ASAP7_75t_SL U67423 ( .A(n73953), .B(n76315), .Y(n64152) );
  AOI21xp33_ASAP7_75t_SRAM U67424 ( .A1(n75736), .A2(n77717), .B(n64128), .Y(
        n64129) );
  NOR2xp33_ASAP7_75t_SL U67425 ( .A(n61784), .B(n61783), .Y(n64119) );
  OAI21xp33_ASAP7_75t_SRAM U67426 ( .A1(n59529), .A2(n64237), .B(n64236), .Y(
        n64245) );
  OAI22xp33_ASAP7_75t_SRAM U67427 ( .A1(n76765), .A2(n75350), .B1(n75326), 
        .B2(n75700), .Y(n64224) );
  OAI22xp33_ASAP7_75t_SRAM U67428 ( .A1(n76764), .A2(n75327), .B1(n75326), 
        .B2(n75325), .Y(n75333) );
  OAI21xp33_ASAP7_75t_SRAM U67429 ( .A1(n75239), .A2(n75863), .B(n64230), .Y(
        n75869) );
  NOR4xp25_ASAP7_75t_SL U67430 ( .A(n64112), .B(n64111), .C(n64110), .D(n64109), .Y(n75871) );
  AND2x2_ASAP7_75t_SL U67431 ( .A(n57126), .B(n75518), .Y(n77031) );
  NOR2xp33_ASAP7_75t_SL U67432 ( .A(n73602), .B(n73652), .Y(n73603) );
  NOR2xp33_ASAP7_75t_SL U67433 ( .A(n75212), .B(n75211), .Y(n75269) );
  AOI22xp33_ASAP7_75t_SRAM U67434 ( .A1(n75646), .A2(n75689), .B1(n75406), 
        .B2(n75203), .Y(n75204) );
  NAND3xp33_ASAP7_75t_SL U67435 ( .A(n62288), .B(n62289), .C(n60810), .Y(
        n62348) );
  NOR2xp33_ASAP7_75t_SL U67436 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_3_), .Y(
        n70623) );
  NOR2xp33_ASAP7_75t_SL U67437 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_22_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_4_), .Y(
        n70624) );
  NOR4xp25_ASAP7_75t_SL U67438 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_15_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_21_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_5_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_9_), .Y(
        n70621) );
  NOR4xp25_ASAP7_75t_SL U67439 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_6_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_8_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_12_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_14_), .Y(
        n70622) );
  NOR4xp25_ASAP7_75t_SL U67440 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_16_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_17_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_18_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_19_), .Y(
        n70619) );
  NOR4xp25_ASAP7_75t_SL U67441 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_10_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_13_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_2_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_0_), .Y(
        n70620) );
  NOR4xp25_ASAP7_75t_SL U67442 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_23_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_24_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_25_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_26_), .Y(
        n70636) );
  NOR4xp25_ASAP7_75t_SL U67443 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_30_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_29_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_28_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_27_), .Y(
        n70637) );
  NOR2xp33_ASAP7_75t_SL U67444 ( .A(n69961), .B(n70003), .Y(n69699) );
  OR2x2_ASAP7_75t_SL U67445 ( .A(n75872), .B(n77066), .Y(n75735) );
  AND2x2_ASAP7_75t_SL U67446 ( .A(n57126), .B(n75518), .Y(n59499) );
  O2A1O1Ixp5_ASAP7_75t_SL U67447 ( .A1(n61145), .A2(n60723), .B(n60722), .C(
        n60721), .Y(n60724) );
  NOR2xp33_ASAP7_75t_SL U67448 ( .A(n60622), .B(n61648), .Y(n61856) );
  NOR2xp33_ASAP7_75t_SL U67449 ( .A(n51957), .B(n73848), .Y(n73849) );
  NOR2xp33_ASAP7_75t_SL U67450 ( .A(n73430), .B(n73429), .Y(n73449) );
  NOR2xp33_ASAP7_75t_SL U67451 ( .A(n73421), .B(n73420), .Y(n73429) );
  NOR2xp33_ASAP7_75t_SL U67452 ( .A(n73413), .B(n73412), .Y(n73414) );
  O2A1O1Ixp5_ASAP7_75t_SL U67453 ( .A1(n73304), .A2(n57185), .B(n73303), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[19]), .Y(
        n73305) );
  NOR2xp33_ASAP7_75t_SL U67454 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[8]), .B(
        n59525), .Y(n73197) );
  NOR2xp33_ASAP7_75t_SL U67455 ( .A(n73166), .B(n73165), .Y(n73434) );
  NOR2xp33_ASAP7_75t_SL U67456 ( .A(n73156), .B(n59630), .Y(n73157) );
  NOR2xp33_ASAP7_75t_SL U67457 ( .A(n60369), .B(n57072), .Y(n62146) );
  NAND2xp33_ASAP7_75t_SRAM U67458 ( .A(n1849), .B(n77354), .Y(n60285) );
  NOR3xp33_ASAP7_75t_SL U67459 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_2_), .B(
        or1200_cpu_or1200_fpu_fpu_op_r_0_), .C(
        or1200_cpu_or1200_fpu_fpu_op_r_1_), .Y(n76494) );
  NOR2xp33_ASAP7_75t_SL U67460 ( .A(n76386), .B(n73967), .Y(n76461) );
  NOR2xp33_ASAP7_75t_SL U67461 ( .A(n74017), .B(n74016), .Y(n76405) );
  NAND2xp33_ASAP7_75t_SRAM U67462 ( .A(n59578), .B(n75456), .Y(n76421) );
  XNOR2xp5_ASAP7_75t_SL U67463 ( .A(n76258), .B(n76257), .Y(n76276) );
  NOR2xp33_ASAP7_75t_SL U67464 ( .A(n63547), .B(n75306), .Y(n75307) );
  NOR2xp33_ASAP7_75t_SL U67465 ( .A(n75684), .B(n75683), .Y(n76270) );
  NOR2xp33_ASAP7_75t_SL U67466 ( .A(n75682), .B(n75681), .Y(n75684) );
  NOR2xp33_ASAP7_75t_SL U67467 ( .A(n61954), .B(n61120), .Y(n62497) );
  INVx1_ASAP7_75t_SL U67468 ( .A(n61064), .Y(n77965) );
  AND2x2_ASAP7_75t_SL U67469 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_25_), 
        .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_24_), 
        .Y(n73861) );
  NAND4xp25_ASAP7_75t_SL U67470 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_30_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_), .Y(n73883) );
  OAI21xp33_ASAP7_75t_SRAM U67471 ( .A1(n63695), .A2(n57160), .B(n63694), .Y(
        n63696) );
  AOI22xp33_ASAP7_75t_SRAM U67472 ( .A1(n77448), .A2(n77247), .B1(n61271), 
        .B2(n57198), .Y(n61273) );
  NOR2xp33_ASAP7_75t_SL U67473 ( .A(n70895), .B(n70882), .Y(n70884) );
  NOR2xp33_ASAP7_75t_SL U67474 ( .A(n58315), .B(n71281), .Y(n71332) );
  XOR2xp5_ASAP7_75t_SL U67475 ( .A(n835), .B(n831), .Y(n77798) );
  NAND3xp33_ASAP7_75t_SL U67476 ( .A(n60290), .B(n1494), .C(n1492), .Y(n60299)
         );
  NOR3xp33_ASAP7_75t_SL U67477 ( .A(n1181), .B(n60233), .C(
        or1200_cpu_or1200_except_n679), .Y(n60234) );
  AND2x2_ASAP7_75t_SL U67478 ( .A(n59462), .B(n53311), .Y(n60668) );
  NAND2xp33_ASAP7_75t_SRAM U67479 ( .A(n59438), .B(n57483), .Y(n60615) );
  O2A1O1Ixp5_ASAP7_75t_SL U67480 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_3_), .A2(n77171), 
        .B(n77139), .C(n74903), .Y(n78190) );
  O2A1O1Ixp5_ASAP7_75t_SL U67481 ( .A1(n57398), .A2(n58759), .B(n66251), .C(
        n66431), .Y(n66273) );
  NAND2xp33_ASAP7_75t_SRAM U67482 ( .A(n67850), .B(n59595), .Y(n62782) );
  NOR2xp33_ASAP7_75t_SL U67483 ( .A(n62728), .B(n59515), .Y(n62716) );
  XNOR2xp5_ASAP7_75t_SL U67484 ( .A(n66826), .B(n66769), .Y(n66819) );
  O2A1O1Ixp5_ASAP7_75t_SL U67485 ( .A1(n58508), .A2(n58672), .B(n67490), .C(
        n67609), .Y(n67493) );
  XNOR2xp5_ASAP7_75t_SL U67486 ( .A(n59601), .B(n67964), .Y(n67465) );
  INVxp33_ASAP7_75t_SRAM U67487 ( .A(n77894), .Y(n77895) );
  OAI21xp33_ASAP7_75t_SRAM U67488 ( .A1(n59708), .A2(n77748), .B(n77689), .Y(
        dwb_dat_o[2]) );
  AOI22xp33_ASAP7_75t_SRAM U67489 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[25]), .B1(n57081), 
        .B2(n70525), .Y(n2260) );
  AOI22xp33_ASAP7_75t_SRAM U67490 ( .A1(n70526), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_rmndr[8]), .B1(n57081), 
        .B2(n70515), .Y(n2226) );
  AOI22xp33_ASAP7_75t_SRAM U67491 ( .A1(n73690), .A2(n57204), .B1(n3313), .B2(
        n59632), .Y(n73644) );
  AOI22xp33_ASAP7_75t_SRAM U67492 ( .A1(n3313), .A2(n57217), .B1(n73728), .B2(
        n57205), .Y(n73694) );
  AO21x1_ASAP7_75t_SL U67493 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .A2(
        n72037), .B(n72036), .Y(n72389) );
  AOI22xp33_ASAP7_75t_SRAM U67494 ( .A1(n57217), .A2(n73690), .B1(n3313), .B2(
        n57205), .Y(n73664) );
  AOI22xp33_ASAP7_75t_SRAM U67495 ( .A1(n57217), .A2(n73667), .B1(n73690), 
        .B2(n57205), .Y(n73620) );
  AOI22xp33_ASAP7_75t_SRAM U67496 ( .A1(n3313), .A2(n57204), .B1(n73728), .B2(
        n59632), .Y(n73621) );
  OAI22xp33_ASAP7_75t_SRAM U67497 ( .A1(n71936), .A2(n57123), .B1(n57203), 
        .B2(n71950), .Y(n71868) );
  OAI21xp33_ASAP7_75t_SRAM U67498 ( .A1(n66124), .A2(n65670), .B(n65505), .Y(
        n66109) );
  AOI22xp33_ASAP7_75t_SRAM U67499 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[32]), .A2(n65634), 
        .B1(n65593), .B2(n65670), .Y(n65594) );
  AOI21xp33_ASAP7_75t_SRAM U67500 ( .A1(n65670), .A2(n65600), .B(n65599), .Y(
        n66115) );
  AOI21xp33_ASAP7_75t_SRAM U67501 ( .A1(n65670), .A2(n65628), .B(n65627), .Y(
        n66151) );
  AOI21xp33_ASAP7_75t_SRAM U67502 ( .A1(n65620), .A2(n65670), .B(n65619), .Y(
        n66148) );
  AOI22xp33_ASAP7_75t_SRAM U67503 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]), .A2(n65621), 
        .B1(n65611), .B2(n65670), .Y(n65612) );
  OAI21xp33_ASAP7_75t_SRAM U67504 ( .A1(n65670), .A2(n65569), .B(n65568), .Y(
        n66099) );
  AOI21xp33_ASAP7_75t_SRAM U67505 ( .A1(n63260), .A2(n63259), .B(n63279), .Y(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N3) );
  INVxp33_ASAP7_75t_SRAM U67506 ( .A(n65457), .Y(n65458) );
  INVxp33_ASAP7_75t_SRAM U67507 ( .A(n65545), .Y(n65548) );
  INVxp33_ASAP7_75t_SRAM U67508 ( .A(n65544), .Y(n65549) );
  INVxp33_ASAP7_75t_SRAM U67509 ( .A(n65543), .Y(n65551) );
  AOI21xp33_ASAP7_75t_SRAM U67510 ( .A1(n65808), .A2(n65807), .B(n65806), .Y(
        n65896) );
  OAI22xp33_ASAP7_75t_SRAM U67511 ( .A1(n78357), .A2(n69563), .B1(n78244), 
        .B2(n78365), .Y(n69442) );
  OAI21xp33_ASAP7_75t_SRAM U67512 ( .A1(n59629), .A2(n72811), .B(n72809), .Y(
        n1799) );
  INVxp33_ASAP7_75t_SRAM U67513 ( .A(n71474), .Y(n71475) );
  INVxp33_ASAP7_75t_SRAM U67514 ( .A(n71501), .Y(n71477) );
  AOI22xp33_ASAP7_75t_SRAM U67515 ( .A1(n73030), .A2(n73029), .B1(n73028), 
        .B2(n73027), .Y(n73033) );
  AOI22xp33_ASAP7_75t_SRAM U67516 ( .A1(n73026), .A2(n73025), .B1(n73024), 
        .B2(n73023), .Y(n73034) );
  OAI21xp33_ASAP7_75t_SRAM U67517 ( .A1(n72993), .A2(n72938), .B(n72999), .Y(
        n72832) );
  AOI22xp33_ASAP7_75t_SRAM U67518 ( .A1(n73030), .A2(n72920), .B1(n73028), 
        .B2(n72938), .Y(n72844) );
  OAI21xp33_ASAP7_75t_SRAM U67519 ( .A1(n57081), .A2(n69840), .B(n69839), .Y(
        n69841) );
  OAI21xp33_ASAP7_75t_SRAM U67520 ( .A1(n57081), .A2(n69855), .B(n69854), .Y(
        n69856) );
  INVxp33_ASAP7_75t_SRAM U67521 ( .A(n72920), .Y(n72924) );
  INVxp33_ASAP7_75t_SRAM U67522 ( .A(n72902), .Y(n72903) );
  INVxp33_ASAP7_75t_SRAM U67523 ( .A(n72901), .Y(n72905) );
  INVxp33_ASAP7_75t_SRAM U67524 ( .A(n72609), .Y(n71538) );
  NOR2xp33_ASAP7_75t_SL U67525 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_5_), .B(
        n74674), .Y(n74695) );
  NOR2xp33_ASAP7_75t_SL U67526 ( .A(n74694), .B(n74642), .Y(n74723) );
  AOI22xp33_ASAP7_75t_SRAM U67527 ( .A1(n77696), .A2(n77070), .B1(n61348), 
        .B2(n57191), .Y(n61349) );
  AOI22xp33_ASAP7_75t_SRAM U67528 ( .A1(n61328), .A2(n74582), .B1(n63410), 
        .B2(n77039), .Y(n61330) );
  OAI22xp33_ASAP7_75t_SRAM U67529 ( .A1(or1200_cpu_or1200_mult_mac_n157), .A2(
        n77057), .B1(n77066), .B2(n76442), .Y(n62364) );
  INVxp33_ASAP7_75t_SRAM U67530 ( .A(n62353), .Y(n62363) );
  AOI22xp33_ASAP7_75t_SRAM U67531 ( .A1(or1200_cpu_or1200_fpu_result_arith[8]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[8]), 
        .Y(n62334) );
  AOI22xp33_ASAP7_75t_SRAM U67532 ( .A1(or1200_cpu_or1200_fpu_result_arith[6]), 
        .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[6]), 
        .Y(n62265) );
  OAI22xp33_ASAP7_75t_SRAM U67533 ( .A1(or1200_cpu_or1200_mult_mac_n147), .A2(
        n77057), .B1(n76438), .B2(n77066), .Y(n61529) );
  AOI22xp33_ASAP7_75t_SRAM U67534 ( .A1(n59182), .A2(n76772), .B1(n61425), 
        .B2(n64220), .Y(n61427) );
  OAI21xp33_ASAP7_75t_SRAM U67535 ( .A1(or1200_cpu_or1200_mult_mac_n120), .A2(
        n77058), .B(n61420), .Y(n61421) );
  AOI22xp33_ASAP7_75t_SRAM U67536 ( .A1(n75852), .A2(n61419), .B1(n63325), 
        .B2(n75853), .Y(n61420) );
  AOI22xp33_ASAP7_75t_SRAM U67537 ( .A1(n76768), .A2(n76767), .B1(n76766), 
        .B2(n77075), .Y(n76769) );
  OAI21xp33_ASAP7_75t_SRAM U67538 ( .A1(n1400), .A2(n77035), .B(n76723), .Y(
        n76726) );
  AOI22xp33_ASAP7_75t_SRAM U67539 ( .A1(n76722), .A2(n77039), .B1(n77041), 
        .B2(n76721), .Y(n76723) );
  OAI21xp33_ASAP7_75t_SRAM U67540 ( .A1(or1200_cpu_or1200_mult_mac_n124), .A2(
        n77058), .B(n61197), .Y(n61198) );
  AOI22xp33_ASAP7_75t_SRAM U67541 ( .A1(n75852), .A2(n76455), .B1(n61249), 
        .B2(n75853), .Y(n61197) );
  OAI22xp33_ASAP7_75t_SRAM U67542 ( .A1(n75702), .A2(n62255), .B1(n63577), 
        .B2(n75325), .Y(n61188) );
  AOI22xp33_ASAP7_75t_SRAM U67543 ( .A1(or1200_cpu_or1200_fpu_result_arith[26]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[26]), .Y(
        n64826) );
  OAI21xp33_ASAP7_75t_SRAM U67544 ( .A1(n69373), .A2(n64814), .B(n77082), .Y(
        n64863) );
  AOI22xp33_ASAP7_75t_SRAM U67545 ( .A1(n74582), .A2(n60820), .B1(n69124), 
        .B2(n77041), .Y(n60823) );
  AOI22xp33_ASAP7_75t_SRAM U67546 ( .A1(or1200_cpu_or1200_fpu_result_arith[27]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[27]), .Y(
        n73917) );
  OAI22xp33_ASAP7_75t_SRAM U67547 ( .A1(n1127), .A2(n75818), .B1(n1432), .B2(
        n75817), .Y(n73909) );
  OAI22xp33_ASAP7_75t_SRAM U67548 ( .A1(or1200_cpu_or1200_mult_mac_n98), .A2(
        n77058), .B1(or1200_cpu_or1200_mult_mac_n171), .B2(n77057), .Y(n77059)
         );
  OAI22xp33_ASAP7_75t_SRAM U67549 ( .A1(n63567), .A2(n75838), .B1(n59534), 
        .B2(n63586), .Y(n63568) );
  AOI22xp33_ASAP7_75t_SRAM U67550 ( .A1(or1200_cpu_or1200_fpu_result_arith[16]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[16]), .Y(
        n62526) );
  OAI22xp33_ASAP7_75t_SRAM U67551 ( .A1(or1200_cpu_or1200_mult_mac_n96), .A2(
        n64785), .B1(n57312), .B2(n64830), .Y(n62517) );
  OAI22xp33_ASAP7_75t_SRAM U67552 ( .A1(n1149), .A2(n77033), .B1(n1454), .B2(
        n77034), .Y(n62503) );
  OAI21xp33_ASAP7_75t_SRAM U67553 ( .A1(or1200_cpu_or1200_mult_mac_n311), .A2(
        n75738), .B(n62429), .Y(n62437) );
  AOI22xp33_ASAP7_75t_SRAM U67554 ( .A1(or1200_cpu_or1200_fpu_result_arith[12]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[12]), .Y(
        n62427) );
  NOR2xp33_ASAP7_75t_SL U67555 ( .A(or1200_cpu_or1200_except_n613), .B(n59675), 
        .Y(n77624) );
  OAI21xp33_ASAP7_75t_SRAM U67556 ( .A1(n77623), .A2(n77626), .B(n62421), .Y(
        n77619) );
  OAI22xp33_ASAP7_75t_SRAM U67557 ( .A1(n1157), .A2(n62419), .B1(n1462), .B2(
        n62418), .Y(n62420) );
  NOR4xp25_ASAP7_75t_SL U67558 ( .A(n62417), .B(n62416), .C(n62415), .D(n58565), .Y(n77630) );
  OAI22xp33_ASAP7_75t_SRAM U67559 ( .A1(or1200_cpu_or1200_except_n212), .A2(
        n57170), .B1(or1200_cpu_or1200_except_n162), .B2(n57102), .Y(n62416)
         );
  NOR2xp33_ASAP7_75t_SL U67560 ( .A(or1200_cpu_or1200_except_n428), .B(n59676), 
        .Y(n62417) );
  AOI211xp5_ASAP7_75t_SL U67561 ( .A1(n77125), .A2(n61796), .B(n61795), .C(
        n77122), .Y(n61797) );
  AOI22xp33_ASAP7_75t_SRAM U67562 ( .A1(or1200_cpu_or1200_fpu_result_arith[10]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[10]), .Y(
        n61775) );
  INVxp33_ASAP7_75t_SRAM U67563 ( .A(n61190), .Y(n61193) );
  AOI22xp33_ASAP7_75t_SRAM U67564 ( .A1(n61748), .A2(n74582), .B1(n61777), 
        .B2(n77039), .Y(n61750) );
  AOI22xp33_ASAP7_75t_SRAM U67565 ( .A1(or1200_cpu_or1200_fpu_result_arith[13]), .A2(n77091), .B1(n77090), .B2(or1200_cpu_or1200_fpu_result_conv[13]), .Y(
        n61100) );
  OAI22xp33_ASAP7_75t_SRAM U67566 ( .A1(or1200_cpu_or1200_mult_mac_n102), .A2(
        n64785), .B1(n59539), .B2(n64830), .Y(n61088) );
  NOR2xp33_ASAP7_75t_SL U67567 ( .A(n61358), .B(n62348), .Y(n61763) );
  OAI22xp33_ASAP7_75t_SRAM U67568 ( .A1(or1200_cpu_or1200_except_n616), .A2(
        n59675), .B1(or1200_cpu_or1200_except_n214), .B2(n57170), .Y(n61073)
         );
  AOI22xp33_ASAP7_75t_SRAM U67569 ( .A1(n1155), .A2(n76711), .B1(n76712), .B2(
        n1460), .Y(n61062) );
  NAND2xp33_ASAP7_75t_SRAM U67570 ( .A(n62319), .B(n77638), .Y(n61067) );
  NOR2xp33_ASAP7_75t_SL U67571 ( .A(or1200_cpu_or1200_except_n160), .B(n57102), 
        .Y(n77635) );
  NOR2xp33_ASAP7_75t_SL U67572 ( .A(or1200_cpu_or1200_except_n514), .B(n77032), 
        .Y(n77636) );
  INVxp33_ASAP7_75t_SRAM U67573 ( .A(n62359), .Y(n61347) );
  OAI22xp33_ASAP7_75t_SRAM U67574 ( .A1(n59536), .A2(n76775), .B1(
        or1200_cpu_or1200_mult_mac_n175), .B2(n77057), .Y(n75320) );
  NOR3xp33_ASAP7_75t_SL U67575 ( .A(n75566), .B(n75565), .C(n75564), .Y(n77660) );
  AOI21xp33_ASAP7_75t_SRAM U67576 ( .A1(n77039), .A2(n75557), .B(n75556), .Y(
        n75560) );
  OAI22xp33_ASAP7_75t_SRAM U67577 ( .A1(n1135), .A2(n77033), .B1(n1440), .B2(
        n77034), .Y(n75556) );
  AOI22xp33_ASAP7_75t_SRAM U67578 ( .A1(n64305), .A2(n75727), .B1(n75736), 
        .B2(n74799), .Y(n64306) );
  OAI22xp33_ASAP7_75t_SRAM U67579 ( .A1(n75832), .A2(n59585), .B1(n57215), 
        .B2(n63571), .Y(n60786) );
  OAI22xp33_ASAP7_75t_SRAM U67580 ( .A1(n75890), .A2(n57197), .B1(n57212), 
        .B2(n59645), .Y(n60787) );
  AOI22xp33_ASAP7_75t_SRAM U67581 ( .A1(n77854), .A2(n76903), .B1(n76902), 
        .B2(n57079), .Y(n76908) );
  OAI21xp33_ASAP7_75t_SRAM U67582 ( .A1(n1582), .A2(n65402), .B(n65308), .Y(
        n65270) );
  O2A1O1Ixp5_ASAP7_75t_SL U67583 ( .A1(n73533), .A2(n73532), .B(n73531), .C(
        n73530), .Y(n73594) );
  O2A1O1Ixp5_ASAP7_75t_SL U67584 ( .A1(n73528), .A2(n73527), .B(n73526), .C(
        n73525), .Y(n73532) );
  NOR2xp33_ASAP7_75t_SL U67585 ( .A(n75853), .B(n76751), .Y(n76755) );
  OAI22xp33_ASAP7_75t_SRAM U67586 ( .A1(n59574), .A2(n75714), .B1(n75713), 
        .B2(n76764), .Y(n75715) );
  INVxp33_ASAP7_75t_SRAM U67587 ( .A(n75706), .Y(n75712) );
  OAI21xp33_ASAP7_75t_SRAM U67588 ( .A1(n59442), .A2(n62432), .B(n60798), .Y(
        n75717) );
  NAND2xp33_ASAP7_75t_SRAM U67589 ( .A(n77128), .B(n77663), .Y(n75880) );
  NOR3xp33_ASAP7_75t_SL U67590 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_20_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_7_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_opb_i_11_), .Y(
        n70625) );
  NAND4xp25_ASAP7_75t_SL U67591 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_3_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_0_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_1_), .Y(
        n70634) );
  NAND4xp25_ASAP7_75t_SL U67592 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_6_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_7_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_4_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo3_5_), .Y(
        n70635) );
  AOI21xp33_ASAP7_75t_SRAM U67593 ( .A1(n60344), .A2(n2596), .B(n60725), .Y(
        n60334) );
  AOI22xp33_ASAP7_75t_SRAM U67594 ( .A1(n59492), .A2(n62000), .B1(n62019), 
        .B2(n77566), .Y(n60380) );
  NOR2xp33_ASAP7_75t_SL U67595 ( .A(n59708), .B(n75328), .Y(n62374) );
  OAI22xp33_ASAP7_75t_SRAM U67596 ( .A1(or1200_cpu_or1200_mult_mac_n141), .A2(
        n77057), .B1(n76431), .B2(n77066), .Y(n60646) );
  HB1xp67_ASAP7_75t_SL U67597 ( .A(n59537), .Y(n59486) );
  AOI21xp33_ASAP7_75t_SRAM U67598 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_31_), .A2(n74518), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_0_), .Y(n73838)
         );
  NOR2xp33_ASAP7_75t_SL U67599 ( .A(n77460), .B(n62002), .Y(n60335) );
  INVxp33_ASAP7_75t_SRAM U67600 ( .A(n75439), .Y(n75444) );
  AOI211xp5_ASAP7_75t_SL U67601 ( .A1(n77217), .A2(n77190), .B(n76510), .C(
        n76509), .Y(n76511) );
  INVxp33_ASAP7_75t_SRAM U67602 ( .A(n76383), .Y(n76385) );
  INVxp33_ASAP7_75t_SRAM U67603 ( .A(n76466), .Y(n76380) );
  INVxp33_ASAP7_75t_SRAM U67604 ( .A(n76363), .Y(n76375) );
  INVxp33_ASAP7_75t_SRAM U67605 ( .A(n76353), .Y(n76356) );
  NOR2xp33_ASAP7_75t_SL U67606 ( .A(n2086), .B(n76323), .Y(n76331) );
  INVxp33_ASAP7_75t_SRAM U67607 ( .A(n73971), .Y(n73973) );
  INVxp33_ASAP7_75t_SRAM U67608 ( .A(n59529), .Y(n64241) );
  NOR2xp33_ASAP7_75t_SL U67609 ( .A(n61323), .B(n61322), .Y(n61674) );
  NOR2xp33_ASAP7_75t_SL U67610 ( .A(n61321), .B(n61320), .Y(n61322) );
  AOI21xp33_ASAP7_75t_SRAM U67611 ( .A1(n62676), .A2(n62737), .B(n53455), .Y(
        n60739) );
  NOR2xp33_ASAP7_75t_SL U67612 ( .A(n73887), .B(n73876), .Y(n73875) );
  NOR4xp25_ASAP7_75t_SL U67613 ( .A(n73874), .B(n73873), .C(n73872), .D(n73871), .Y(n74361) );
  NAND4xp25_ASAP7_75t_SL U67614 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_27_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_29_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_), .Y(n73884) );
  OAI21xp33_ASAP7_75t_SRAM U67615 ( .A1(n59556), .A2(n57124), .B(n61166), .Y(
        n61173) );
  OAI22xp33_ASAP7_75t_SRAM U67616 ( .A1(n76591), .A2(n57160), .B1(n1033), .B2(
        n57168), .Y(n61574) );
  NOR2xp33_ASAP7_75t_SL U67617 ( .A(n57090), .B(n61045), .Y(n61050) );
  NAND2xp33_ASAP7_75t_SRAM U67618 ( .A(n59702), .B(
        or1200_cpu_or1200_genpc_pcreg_default[2]), .Y(n63741) );
  NAND2xp33_ASAP7_75t_SRAM U67619 ( .A(n77337), .B(n77348), .Y(n77400) );
  NAND2xp33_ASAP7_75t_SRAM U67620 ( .A(n22057), .B(n60101), .Y(n77346) );
  INVx1_ASAP7_75t_SL U67621 ( .A(n77998), .Y(n77765) );
  O2A1O1Ixp5_ASAP7_75t_SL U67622 ( .A1(n74894), .A2(n74893), .B(n74892), .C(
        n76932), .Y(n74895) );
  NAND2xp33_ASAP7_75t_SRAM U67623 ( .A(n74835), .B(n76956), .Y(n74836) );
  O2A1O1Ixp5_ASAP7_75t_SL U67624 ( .A1(n77193), .A2(n77196), .B(n74886), .C(
        n74885), .Y(n74897) );
  XNOR2xp5_ASAP7_75t_SL U67625 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_0_), .B(n74204), 
        .Y(n74211) );
  NOR2xp33_ASAP7_75t_SL U67626 ( .A(n75096), .B(n75095), .Y(n68647) );
  XNOR2xp5_ASAP7_75t_SL U67627 ( .A(n66395), .B(n66394), .Y(n66442) );
  XNOR2xp5_ASAP7_75t_SL U67628 ( .A(n59637), .B(n57336), .Y(n66572) );
  XNOR2xp5_ASAP7_75t_SL U67629 ( .A(n59638), .B(n57325), .Y(n66542) );
  AOI21xp33_ASAP7_75t_SRAM U67630 ( .A1(n59503), .A2(n67227), .B(n62876), .Y(
        n62878) );
  XNOR2xp5_ASAP7_75t_SL U67631 ( .A(n62871), .B(n62870), .Y(n62872) );
  NAND2xp33_ASAP7_75t_SRAM U67632 ( .A(n59504), .B(n57422), .Y(n62801) );
  NAND2xp33_ASAP7_75t_SRAM U67633 ( .A(n58431), .B(n67428), .Y(n62783) );
  NOR2xp33_ASAP7_75t_SL U67634 ( .A(n67227), .B(n59503), .Y(n62876) );
  NAND2xp33_ASAP7_75t_SRAM U67635 ( .A(n53320), .B(n75901), .Y(n63223) );
  AOI21xp33_ASAP7_75t_SRAM U67636 ( .A1(n59518), .A2(n76057), .B(n59140), .Y(
        n59139) );
  XNOR2xp5_ASAP7_75t_SL U67637 ( .A(n57107), .B(n58383), .Y(n66955) );
  XNOR2xp5_ASAP7_75t_SL U67638 ( .A(n59617), .B(n59647), .Y(n68381) );
  OAI21xp33_ASAP7_75t_SRAM U67639 ( .A1(n57110), .A2(n59459), .B(n68079), .Y(
        n65063) );
  INVxp33_ASAP7_75t_SRAM U67640 ( .A(n67837), .Y(n67838) );
  O2A1O1Ixp5_ASAP7_75t_SL U67641 ( .A1(n59620), .A2(n59239), .B(n57176), .C(
        n67915), .Y(n67917) );
  XNOR2xp5_ASAP7_75t_SL U67642 ( .A(n59638), .B(n59664), .Y(n75073) );
  NAND2xp33_ASAP7_75t_SRAM U67643 ( .A(n59190), .B(n59637), .Y(n75047) );
  INVxp33_ASAP7_75t_SRAM U67644 ( .A(n77913), .Y(n77914) );
  INVxp33_ASAP7_75t_SRAM U67645 ( .A(n77860), .Y(n77861) );
  INVxp33_ASAP7_75t_SRAM U67646 ( .A(n77857), .Y(n77858) );
  INVxp33_ASAP7_75t_SRAM U67647 ( .A(n77891), .Y(n77892) );
  INVxp33_ASAP7_75t_SRAM U67648 ( .A(n77878), .Y(n77879) );
  INVxp33_ASAP7_75t_SRAM U67649 ( .A(n77881), .Y(n77882) );
  INVxp33_ASAP7_75t_SRAM U67650 ( .A(n77907), .Y(n77908) );
  INVxp33_ASAP7_75t_SRAM U67651 ( .A(n77902), .Y(n77903) );
  INVxp33_ASAP7_75t_SRAM U67652 ( .A(n77897), .Y(n77898) );
  INVxp33_ASAP7_75t_SRAM U67653 ( .A(n77886), .Y(n77887) );
  INVxp33_ASAP7_75t_SRAM U67654 ( .A(n77867), .Y(n77868) );
  INVxp33_ASAP7_75t_SRAM U67655 ( .A(n77905), .Y(n77906) );
  AND3x1_ASAP7_75t_SL U67656 ( .A(n77967), .B(n77966), .C(n77965), .Y(n78176)
         );
  NAND2xp33_ASAP7_75t_SRAM U67657 ( .A(n77994), .B(n77993), .Y(n4139) );
  OAI21xp33_ASAP7_75t_SRAM U67658 ( .A1(n59581), .A2(n77748), .B(n77694), .Y(
        dwb_dat_o[7]) );
  OAI21xp33_ASAP7_75t_SRAM U67659 ( .A1(n59556), .A2(n77748), .B(n77693), .Y(
        dwb_dat_o[6]) );
  OAI21xp33_ASAP7_75t_SRAM U67660 ( .A1(n59544), .A2(n77748), .B(n77692), .Y(
        dwb_dat_o[5]) );
  OAI21xp33_ASAP7_75t_SRAM U67661 ( .A1(n59567), .A2(n77748), .B(n77691), .Y(
        dwb_dat_o[4]) );
  OAI21xp33_ASAP7_75t_SRAM U67662 ( .A1(n59558), .A2(n77748), .B(n77690), .Y(
        dwb_dat_o[3]) );
  OAI21xp33_ASAP7_75t_SRAM U67663 ( .A1(n59442), .A2(n77748), .B(n77688), .Y(
        dwb_dat_o[1]) );
  OAI21xp33_ASAP7_75t_SRAM U67664 ( .A1(n59710), .A2(n77748), .B(n77687), .Y(
        dwb_dat_o[0]) );
  AOI21xp33_ASAP7_75t_SRAM U67665 ( .A1(n77735), .A2(n77746), .B(n77734), .Y(
        n4252) );
  OAI22xp33_ASAP7_75t_SRAM U67666 ( .A1(n57500), .A2(n77745), .B1(n59708), 
        .B2(n77744), .Y(n77734) );
  AOI21xp33_ASAP7_75t_SRAM U67667 ( .A1(n77742), .A2(n78005), .B(n77738), .Y(
        n4248) );
  OAI22xp33_ASAP7_75t_SRAM U67668 ( .A1(n1868), .A2(n77741), .B1(n59553), .B2(
        n77745), .Y(n77738) );
  NAND2xp33_ASAP7_75t_SRAM U67669 ( .A(n2607), .B(n77763), .Y(n77725) );
  INVxp33_ASAP7_75t_SRAM U67670 ( .A(n60277), .Y(n60280) );
  OAI21xp33_ASAP7_75t_SRAM U67671 ( .A1(n3084), .A2(n77476), .B(n61999), .Y(
        n9389) );
  AOI22xp33_ASAP7_75t_SRAM U67672 ( .A1(n73743), .A2(n57204), .B1(n73753), 
        .B2(n59632), .Y(n73693) );
  AOI22xp33_ASAP7_75t_SRAM U67673 ( .A1(n73728), .A2(n57204), .B1(n73743), 
        .B2(n59632), .Y(n73665) );
  OAI22xp33_ASAP7_75t_SRAM U67674 ( .A1(n72310), .A2(n57123), .B1(n57203), 
        .B2(n72318), .Y(n72261) );
  OAI22xp33_ASAP7_75t_SRAM U67675 ( .A1(n72350), .A2(n57123), .B1(n57203), 
        .B2(n72313), .Y(n72259) );
  OAI22xp33_ASAP7_75t_SRAM U67676 ( .A1(n72310), .A2(n57127), .B1(n57203), 
        .B2(n72319), .Y(n72292) );
  OAI22xp33_ASAP7_75t_SRAM U67677 ( .A1(n72319), .A2(n57127), .B1(n57203), 
        .B2(n72307), .Y(n72244) );
  OAI22xp33_ASAP7_75t_SRAM U67678 ( .A1(n72306), .A2(n57123), .B1(n57203), 
        .B2(n72253), .Y(n72255) );
  OR3x1_ASAP7_75t_SL U67679 ( .A(n77686), .B(n78166), .C(n77491), .Y(n4318) );
  OAI22xp33_ASAP7_75t_SRAM U67680 ( .A1(n72311), .A2(n57123), .B1(n57203), 
        .B2(n72310), .Y(n72315) );
  OAI22xp33_ASAP7_75t_SRAM U67681 ( .A1(n72317), .A2(n57125), .B1(n57203), 
        .B2(n72316), .Y(n72321) );
  AOI22xp33_ASAP7_75t_SRAM U67682 ( .A1(n72347), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_), 
        .B1(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), .B2(n58447), .Y(n71971) );
  OAI21xp33_ASAP7_75t_SRAM U67683 ( .A1(n65629), .A2(n65832), .B(n65511), .Y(
        n66108) );
  AOI22xp33_ASAP7_75t_SRAM U67684 ( .A1(n66182), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .B2(n66146), 
        .Y(n65505) );
  OAI21xp33_ASAP7_75t_SRAM U67685 ( .A1(n65629), .A2(n65859), .B(n65504), .Y(
        n66104) );
  AOI22xp33_ASAP7_75t_SRAM U67686 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]), .A2(n59562), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .B2(n74206), .Y(n66124) );
  AOI22xp33_ASAP7_75t_SRAM U67687 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[46]), .A2(n59562), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[45]), .B2(n74206), .Y(n65588) );
  OAI21xp33_ASAP7_75t_SRAM U67688 ( .A1(n59562), .A2(n65684), .B(n65510), .Y(
        n65593) );
  OAI21xp33_ASAP7_75t_SRAM U67689 ( .A1(n74206), .A2(n65631), .B(n65512), .Y(
        n65602) );
  OAI22xp33_ASAP7_75t_SRAM U67690 ( .A1(n65831), .A2(n66181), .B1(n65761), 
        .B2(n65653), .Y(n65590) );
  OAI21xp33_ASAP7_75t_SRAM U67691 ( .A1(n59562), .A2(n65761), .B(n65508), .Y(
        n65592) );
  AOI22xp33_ASAP7_75t_SRAM U67692 ( .A1(n66182), .A2(n65644), .B1(n65643), 
        .B2(n66146), .Y(n65645) );
  OAI22xp33_ASAP7_75t_SRAM U67693 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[33]), .A2(n65646), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[32]), .B2(n66181), .Y(n65619) );
  OAI21xp33_ASAP7_75t_SRAM U67694 ( .A1(n65745), .A2(n65646), .B(n66181), .Y(
        n65614) );
  OAI22xp33_ASAP7_75t_SRAM U67695 ( .A1(n65711), .A2(n65653), .B1(n65629), 
        .B2(n65743), .Y(n65615) );
  AOI22xp33_ASAP7_75t_SRAM U67696 ( .A1(n66182), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[20]), .B2(n66146), 
        .Y(n65568) );
  OAI21xp33_ASAP7_75t_SRAM U67697 ( .A1(n74206), .A2(n65583), .B(n65567), .Y(
        n65628) );
  AOI22xp33_ASAP7_75t_SRAM U67698 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[31]), .A2(n59562), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .B2(n74206), .Y(n65620) );
  OAI21xp33_ASAP7_75t_SRAM U67699 ( .A1(n59562), .A2(n65804), .B(n65571), .Y(
        n65611) );
  AOI22xp33_ASAP7_75t_SRAM U67700 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[45]), .A2(n59562), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[44]), .B2(n74206), .Y(n65616) );
  AOI22xp33_ASAP7_75t_SRAM U67701 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[1]), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .B1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[40]), .B2(n74206), 
        .Y(n65562) );
  INVxp33_ASAP7_75t_SRAM U67702 ( .A(n65447), .Y(n65448) );
  OAI21xp33_ASAP7_75t_SRAM U67703 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .A2(n65808), 
        .B(n58582), .Y(n65800) );
  OAI22xp33_ASAP7_75t_SRAM U67704 ( .A1(n748), .A2(n74916), .B1(n59581), .B2(
        n74934), .Y(n74917) );
  INVxp33_ASAP7_75t_SRAM U67705 ( .A(n53614), .Y(n74918) );
  INVxp33_ASAP7_75t_SRAM U67706 ( .A(n59885), .Y(n59888) );
  INVxp33_ASAP7_75t_SRAM U67707 ( .A(n78166), .Y(n77413) );
  INVxp33_ASAP7_75t_SRAM U67708 ( .A(n61293), .Y(n61295) );
  AOI21xp33_ASAP7_75t_SRAM U67709 ( .A1(n77967), .A2(n77481), .B(n3092), .Y(
        n77475) );
  OAI21xp33_ASAP7_75t_SRAM U67710 ( .A1(n78092), .A2(n78091), .B(n78090), .Y(
        n78093) );
  OAI21xp33_ASAP7_75t_SRAM U67711 ( .A1(n78067), .A2(n56829), .B(n78066), .Y(
        n9356) );
  OAI22xp33_ASAP7_75t_SRAM U67712 ( .A1(n77453), .A2(n77452), .B1(n77451), 
        .B2(n77450), .Y(or1200_cpu_or1200_except_n1731) );
  OAI22xp33_ASAP7_75t_SRAM U67713 ( .A1(or1200_cpu_or1200_mult_mac_n233), .A2(
        n76909), .B1(n77019), .B2(n69182), .Y(n69128) );
  OAI22xp33_ASAP7_75t_SRAM U67714 ( .A1(or1200_cpu_or1200_mult_mac_n217), .A2(
        n76909), .B1(n77600), .B2(n69182), .Y(n68952) );
  OAI22xp33_ASAP7_75t_SRAM U67715 ( .A1(or1200_cpu_or1200_mult_mac_n237), .A2(
        n76909), .B1(n76235), .B2(n69182), .Y(n69183) );
  AOI22xp33_ASAP7_75t_SRAM U67716 ( .A1(or1200_cpu_or1200_except_n294), .A2(
        n77437), .B1(n77436), .B2(n77439), .Y(or1200_cpu_or1200_except_n1788)
         );
  OAI22xp33_ASAP7_75t_SRAM U67717 ( .A1(n1821), .A2(n77463), .B1(n59542), .B2(
        n59688), .Y(n61377) );
  OAI21xp33_ASAP7_75t_SRAM U67718 ( .A1(n76978), .A2(n76977), .B(n76976), .Y(
        n76979) );
  INVxp33_ASAP7_75t_SRAM U67719 ( .A(n76934), .Y(n76967) );
  INVxp33_ASAP7_75t_SRAM U67720 ( .A(n76933), .Y(n76969) );
  AOI21xp33_ASAP7_75t_SRAM U67721 ( .A1(n74926), .A2(n74925), .B(n74942), .Y(
        n74932) );
  INVxp33_ASAP7_75t_SRAM U67722 ( .A(n77436), .Y(n74927) );
  INVxp33_ASAP7_75t_SRAM U67723 ( .A(n74935), .Y(n74941) );
  AOI22xp33_ASAP7_75t_SRAM U67724 ( .A1(n69023), .A2(n68812), .B1(n77623), 
        .B2(n61332), .Y(n61329) );
  INVxp33_ASAP7_75t_SRAM U67725 ( .A(n62371), .Y(n62376) );
  AOI22xp33_ASAP7_75t_SRAM U67726 ( .A1(n63411), .A2(n76753), .B1(n64776), 
        .B2(n77060), .Y(n62367) );
  AOI22xp33_ASAP7_75t_SRAM U67727 ( .A1(n64775), .A2(n62363), .B1(n62362), 
        .B2(n62361), .Y(n62370) );
  OAI22xp33_ASAP7_75t_SRAM U67728 ( .A1(or1200_cpu_or1200_mult_mac_n157), .A2(
        n63555), .B1(n62319), .B2(n62323), .Y(n62320) );
  OAI21xp33_ASAP7_75t_SRAM U67729 ( .A1(n59555), .A2(n62276), .B(n62275), .Y(
        n62277) );
  OAI22xp33_ASAP7_75t_SRAM U67730 ( .A1(n62319), .A2(n62242), .B1(
        or1200_cpu_or1200_mult_mac_n153), .B2(n63555), .Y(n62239) );
  AOI21xp33_ASAP7_75t_SRAM U67731 ( .A1(or1200_cpu_or1200_rf_rf_we_allow), 
        .A2(n57144), .B(n77566), .Y(or1200_cpu_or1200_rf_n12) );
  OAI22xp33_ASAP7_75t_SRAM U67732 ( .A1(n59558), .A2(n76775), .B1(
        or1200_cpu_or1200_mult_mac_n122), .B2(n77058), .Y(n61527) );
  AOI21xp33_ASAP7_75t_SRAM U67733 ( .A1(n61500), .A2(n58206), .B(n61499), .Y(
        n61501) );
  AOI22xp33_ASAP7_75t_SRAM U67734 ( .A1(n61495), .A2(n61494), .B1(n61493), 
        .B2(n62374), .Y(n61502) );
  INVxp33_ASAP7_75t_SRAM U67735 ( .A(n61486), .Y(n61487) );
  AOI22xp33_ASAP7_75t_SRAM U67736 ( .A1(n61474), .A2(n74582), .B1(n77043), 
        .B2(n76855), .Y(n61475) );
  OAI21xp33_ASAP7_75t_SRAM U67737 ( .A1(n59563), .A2(n61413), .B(n61412), .Y(
        n61414) );
  AOI22xp33_ASAP7_75t_SRAM U67738 ( .A1(n61411), .A2(n66239), .B1(n62682), 
        .B2(n61635), .Y(n61412) );
  AOI21xp33_ASAP7_75t_SRAM U67739 ( .A1(n77060), .A2(n57214), .B(n76776), .Y(
        n76777) );
  OAI22xp33_ASAP7_75t_SRAM U67740 ( .A1(n59581), .A2(n76775), .B1(n76774), 
        .B2(n77066), .Y(n76776) );
  OAI22xp33_ASAP7_75t_SRAM U67741 ( .A1(or1200_cpu_or1200_mult_mac_n114), .A2(
        n77058), .B1(or1200_cpu_or1200_mult_mac_n155), .B2(n76751), .Y(n76752)
         );
  OAI21xp33_ASAP7_75t_SRAM U67742 ( .A1(n1398), .A2(n76716), .B(n76715), .Y(
        n76727) );
  AOI22xp33_ASAP7_75t_SRAM U67743 ( .A1(n1472), .A2(n76712), .B1(n76711), .B2(
        n1165), .Y(n76714) );
  AOI22xp33_ASAP7_75t_SRAM U67744 ( .A1(n74582), .A2(n61250), .B1(n68849), 
        .B2(n68812), .Y(n61251) );
  AOI22xp33_ASAP7_75t_SRAM U67745 ( .A1(n77623), .A2(n61254), .B1(n61249), 
        .B2(n75368), .Y(n61252) );
  INVxp33_ASAP7_75t_SRAM U67746 ( .A(n62612), .Y(n61211) );
  AOI22xp33_ASAP7_75t_SRAM U67747 ( .A1(n61411), .A2(n61214), .B1(n64839), 
        .B2(n64235), .Y(n61202) );
  OAI21xp33_ASAP7_75t_SRAM U67748 ( .A1(n61201), .A2(n61200), .B(n61199), .Y(
        n61204) );
  AOI21xp33_ASAP7_75t_SRAM U67749 ( .A1(n76772), .A2(n53316), .B(n61198), .Y(
        n61199) );
  OAI22xp33_ASAP7_75t_SRAM U67750 ( .A1(n2561), .A2(n59679), .B1(n59442), .B2(
        n57074), .Y(n61014) );
  OAI22xp33_ASAP7_75t_SRAM U67751 ( .A1(n59528), .A2(n75239), .B1(n75745), 
        .B2(n75702), .Y(n64844) );
  OAI22xp33_ASAP7_75t_SRAM U67752 ( .A1(n77735), .A2(n64835), .B1(n1571), .B2(
        n77097), .Y(n64848) );
  OAI22xp33_ASAP7_75t_SRAM U67753 ( .A1(or1200_cpu_or1200_mult_mac_n106), .A2(
        n77058), .B1(or1200_cpu_or1200_mult_mac_n163), .B2(n76751), .Y(n61719)
         );
  OAI21xp33_ASAP7_75t_SRAM U67754 ( .A1(or1200_cpu_or1200_mult_mac_n106), .A2(
        n61826), .B(n61718), .Y(n61722) );
  AOI21xp33_ASAP7_75t_SRAM U67755 ( .A1(n59712), .A2(n59576), .B(n59442), .Y(
        n61707) );
  OAI21xp33_ASAP7_75t_SRAM U67756 ( .A1(n59540), .A2(n75734), .B(n64830), .Y(
        n61700) );
  OAI22xp33_ASAP7_75t_SRAM U67757 ( .A1(n76764), .A2(n64843), .B1(n75713), 
        .B2(n75710), .Y(n63575) );
  AOI21xp33_ASAP7_75t_SRAM U67758 ( .A1(n64829), .A2(n63569), .B(n63568), .Y(
        n63582) );
  AOI22xp33_ASAP7_75t_SRAM U67759 ( .A1(n75847), .A2(n59712), .B1(n62519), 
        .B2(n75245), .Y(n62520) );
  INVxp33_ASAP7_75t_SRAM U67760 ( .A(n75328), .Y(n62522) );
  INVxp33_ASAP7_75t_SRAM U67761 ( .A(n77081), .Y(n62515) );
  INVxp33_ASAP7_75t_SRAM U67762 ( .A(n61243), .Y(n61244) );
  INVxp33_ASAP7_75t_SRAM U67763 ( .A(n61242), .Y(n61245) );
  INVxp33_ASAP7_75t_SRAM U67764 ( .A(n62333), .Y(n61774) );
  AOI22xp33_ASAP7_75t_SRAM U67765 ( .A1(n62738), .A2(n75736), .B1(n61764), 
        .B2(n75727), .Y(n61765) );
  AOI22xp33_ASAP7_75t_SRAM U67766 ( .A1(n69024), .A2(n68812), .B1(n77623), 
        .B2(n61752), .Y(n61749) );
  OAI22xp33_ASAP7_75t_SRAM U67767 ( .A1(n1386), .A2(n76716), .B1(n61746), .B2(
        n61745), .Y(n61752) );
  OAI22xp33_ASAP7_75t_SRAM U67768 ( .A1(n62418), .A2(n61744), .B1(n62404), 
        .B2(n62419), .Y(n61745) );
  OAI22xp33_ASAP7_75t_SRAM U67769 ( .A1(or1200_cpu_or1200_mult_mac_n181), .A2(
        n75723), .B1(n59567), .B2(n75722), .Y(n64128) );
  OAI21xp33_ASAP7_75t_SRAM U67770 ( .A1(n64116), .A2(n75347), .B(n64115), .Y(
        n64117) );
  INVxp33_ASAP7_75t_SRAM U67771 ( .A(n62444), .Y(n61086) );
  OAI22xp33_ASAP7_75t_SRAM U67772 ( .A1(n62355), .A2(n75324), .B1(n61347), 
        .B2(n75327), .Y(n64225) );
  OAI22xp33_ASAP7_75t_SRAM U67773 ( .A1(n75330), .A2(n75838), .B1(n75329), 
        .B2(n75328), .Y(n75331) );
  OAI22xp33_ASAP7_75t_SRAM U67774 ( .A1(n59442), .A2(n75319), .B1(n77066), 
        .B2(n76450), .Y(n75321) );
  OAI21xp33_ASAP7_75t_SRAM U67775 ( .A1(n59576), .A2(n59442), .B(n57197), .Y(
        n61530) );
  AOI22xp33_ASAP7_75t_SRAM U67776 ( .A1(n77757), .A2(n77116), .B1(n77752), 
        .B2(n77087), .Y(n75571) );
  OAI21xp33_ASAP7_75t_SRAM U67777 ( .A1(n57197), .A2(n76627), .B(n58081), .Y(
        n62423) );
  OAI22xp33_ASAP7_75t_SRAM U67778 ( .A1(n77278), .A2(n59585), .B1(n76653), 
        .B2(n59645), .Y(n62424) );
  AOI22xp33_ASAP7_75t_SRAM U67779 ( .A1(n61438), .A2(n77242), .B1(n59708), 
        .B2(n62518), .Y(n75865) );
  AOI22xp33_ASAP7_75t_SRAM U67780 ( .A1(n75847), .A2(n59387), .B1(n75846), 
        .B2(n57191), .Y(n75859) );
  OAI22xp33_ASAP7_75t_SRAM U67781 ( .A1(n75840), .A2(n59645), .B1(n75839), 
        .B2(n75838), .Y(n75842) );
  AOI21xp33_ASAP7_75t_SRAM U67782 ( .A1(n59586), .A2(n75832), .B(n75831), .Y(
        n75837) );
  AOI22xp33_ASAP7_75t_SRAM U67783 ( .A1(n75847), .A2(n56954), .B1(n64776), 
        .B2(n75245), .Y(n64777) );
  OAI21xp33_ASAP7_75t_SRAM U67784 ( .A1(n59710), .A2(n62604), .B(n62430), .Y(
        n62431) );
  OAI21xp33_ASAP7_75t_SRAM U67785 ( .A1(n59710), .A2(n57641), .B(n59443), .Y(
        n62533) );
  OAI22xp33_ASAP7_75t_SRAM U67786 ( .A1(or1200_cpu_or1200_except_n258), .A2(
        n58547), .B1(n77210), .B2(or1200_cpu_or1200_except_n122), .Y(n77211)
         );
  INVxp33_ASAP7_75t_SRAM U67787 ( .A(n76503), .Y(n75524) );
  INVxp33_ASAP7_75t_SRAM U67788 ( .A(n65344), .Y(n65292) );
  AOI22xp33_ASAP7_75t_SRAM U67789 ( .A1(n77209), .A2(or1200_cpu_to_sr[1]), 
        .B1(n62156), .B2(n77215), .Y(n62157) );
  AOI22xp33_ASAP7_75t_SRAM U67790 ( .A1(n77209), .A2(or1200_cpu_to_sr[2]), 
        .B1(n63764), .B2(n77215), .Y(n63765) );
  OAI22xp33_ASAP7_75t_SRAM U67791 ( .A1(or1200_cpu_or1200_mult_mac_n183), .A2(
        n75723), .B1(n59544), .B2(n75722), .Y(n62114) );
  INVxp33_ASAP7_75t_SRAM U67792 ( .A(n77163), .Y(n77167) );
  OAI21xp33_ASAP7_75t_SRAM U67793 ( .A1(n59563), .A2(n59443), .B(n59585), .Y(
        n61875) );
  OAI21xp33_ASAP7_75t_SRAM U67794 ( .A1(n57377), .A2(n59442), .B(n59712), .Y(
        n61877) );
  AOI22xp33_ASAP7_75t_SRAM U67795 ( .A1(n78327), .A2(n75736), .B1(n61865), 
        .B2(n75727), .Y(n61866) );
  OAI21xp33_ASAP7_75t_SRAM U67796 ( .A1(n78182), .A2(n75735), .B(n61859), .Y(
        n61860) );
  INVxp33_ASAP7_75t_SRAM U67797 ( .A(n73907), .Y(n61847) );
  OAI22xp33_ASAP7_75t_SRAM U67798 ( .A1(n57090), .A2(n77407), .B1(n2589), .B2(
        n77454), .Y(n9572) );
  OAI22xp33_ASAP7_75t_SRAM U67799 ( .A1(n57090), .A2(n77455), .B1(n2616), .B2(
        n77454), .Y(n9571) );
  OAI22xp33_ASAP7_75t_SRAM U67800 ( .A1(n76765), .A2(n75240), .B1(n59575), 
        .B2(n75239), .Y(n75242) );
  INVxp33_ASAP7_75t_SRAM U67801 ( .A(n64229), .Y(n75239) );
  OAI22xp33_ASAP7_75t_SRAM U67802 ( .A1(n76874), .A2(n57197), .B1(n64114), 
        .B2(n59585), .Y(n62121) );
  OAI22xp33_ASAP7_75t_SRAM U67803 ( .A1(n63668), .A2(n63571), .B1(n57209), 
        .B2(n59645), .Y(n62122) );
  OAI22xp33_ASAP7_75t_SRAM U67804 ( .A1(n59530), .A2(n59585), .B1(n64232), 
        .B2(n64231), .Y(n75235) );
  OAI21xp33_ASAP7_75t_SRAM U67805 ( .A1(n78435), .A2(n65244), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_11_), .Y(n65239) );
  OAI22xp33_ASAP7_75t_SRAM U67806 ( .A1(or1200_cpu_or1200_mult_mac_n201), .A2(
        n75723), .B1(n59552), .B2(n75722), .Y(n75724) );
  OAI21xp33_ASAP7_75t_SRAM U67807 ( .A1(n59710), .A2(n57082), .B(n61190), .Y(
        n62432) );
  INVxp33_ASAP7_75t_SRAM U67808 ( .A(n65115), .Y(n65118) );
  AOI21xp33_ASAP7_75t_SRAM U67809 ( .A1(n65313), .A2(n65344), .B(n65297), .Y(
        n65295) );
  OAI21xp33_ASAP7_75t_SRAM U67810 ( .A1(n65289), .A2(n65354), .B(n65308), .Y(
        n65300) );
  OAI21xp33_ASAP7_75t_SRAM U67811 ( .A1(n65353), .A2(n65354), .B(n65308), .Y(
        n65296) );
  AOI21xp33_ASAP7_75t_SRAM U67812 ( .A1(n64229), .A2(n76782), .B(n76772), .Y(
        n61524) );
  AOI22xp33_ASAP7_75t_SRAM U67813 ( .A1(n60945), .A2(n60944), .B1(n64221), 
        .B2(n60943), .Y(n60948) );
  OAI22xp33_ASAP7_75t_SRAM U67814 ( .A1(n59579), .A2(n57197), .B1(n59575), 
        .B2(n59645), .Y(n60942) );
  OAI21xp33_ASAP7_75t_SRAM U67815 ( .A1(n59557), .A2(n75714), .B(n76770), .Y(
        n60939) );
  INVxp33_ASAP7_75t_SRAM U67816 ( .A(n66253), .Y(n61650) );
  OAI22xp33_ASAP7_75t_SRAM U67817 ( .A1(n57210), .A2(n63571), .B1(n57128), 
        .B2(n59645), .Y(n60679) );
  AOI21xp33_ASAP7_75t_SRAM U67818 ( .A1(n59541), .A2(n59710), .B(n59442), .Y(
        n62430) );
  AOI22xp33_ASAP7_75t_SRAM U67819 ( .A1(n60799), .A2(n64229), .B1(n59712), 
        .B2(n76773), .Y(n60634) );
  AOI21xp33_ASAP7_75t_SRAM U67820 ( .A1(n60644), .A2(n60623), .B(n59438), .Y(
        n60624) );
  OAI21xp33_ASAP7_75t_SRAM U67821 ( .A1(n57082), .A2(n60913), .B(n59570), .Y(
        n60656) );
  AOI21xp33_ASAP7_75t_SRAM U67822 ( .A1(n76653), .A2(n59542), .B(n58206), .Y(
        n60913) );
  INVxp33_ASAP7_75t_SRAM U67823 ( .A(n65030), .Y(n60604) );
  INVxp33_ASAP7_75t_SRAM U67824 ( .A(n66240), .Y(n60601) );
  OAI21xp33_ASAP7_75t_SRAM U67825 ( .A1(n60598), .A2(n62609), .B(n60597), .Y(
        n60603) );
  INVxp33_ASAP7_75t_SRAM U67826 ( .A(n60946), .Y(n60616) );
  AOI21xp33_ASAP7_75t_SRAM U67827 ( .A1(n62000), .A2(n60623), .B(n62072), .Y(
        n60371) );
  AOI22xp33_ASAP7_75t_SRAM U67828 ( .A1(n77456), .A2(n77357), .B1(n69332), 
        .B2(n57137), .Y(n69333) );
  INVxp33_ASAP7_75t_SRAM U67829 ( .A(n78067), .Y(n78068) );
  AOI21xp33_ASAP7_75t_SRAM U67830 ( .A1(n59533), .A2(n77713), .B(n76443), .Y(
        n76447) );
  INVxp33_ASAP7_75t_SRAM U67831 ( .A(n76277), .Y(n76306) );
  OAI21xp33_ASAP7_75t_SRAM U67832 ( .A1(n59550), .A2(n66249), .B(n57120), .Y(
        n61905) );
  HB1xp67_ASAP7_75t_SL U67833 ( .A(n59070), .Y(n59069) );
  OAI21xp33_ASAP7_75t_SRAM U67834 ( .A1(n59556), .A2(n61923), .B(n57120), .Y(
        n60766) );
  OAI21xp33_ASAP7_75t_SRAM U67835 ( .A1(n74416), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_20_), 
        .B(n74426), .Y(n74417) );
  OAI22xp33_ASAP7_75t_SRAM U67836 ( .A1(n2713), .A2(n61042), .B1(n3117), .B2(
        n77454), .Y(n60428) );
  INVxp33_ASAP7_75t_SRAM U67837 ( .A(n60422), .Y(n60423) );
  INVxp33_ASAP7_75t_SRAM U67838 ( .A(n60420), .Y(n60427) );
  OAI22xp33_ASAP7_75t_SRAM U67839 ( .A1(or1200_cpu_or1200_except_n212), .A2(
        n58547), .B1(n77295), .B2(n77254), .Y(n63936) );
  OAI22xp33_ASAP7_75t_SRAM U67840 ( .A1(n3057), .A2(n74953), .B1(n76821), .B2(
        n61570), .Y(n61571) );
  OAI22xp33_ASAP7_75t_SRAM U67841 ( .A1(or1200_cpu_or1200_except_n208), .A2(
        n58547), .B1(or1200_cpu_or1200_except_n116), .B2(
        or1200_cpu_or1200_except_n292), .Y(n63690) );
  OAI22xp33_ASAP7_75t_SRAM U67842 ( .A1(n75781), .A2(n59494), .B1(n57500), 
        .B2(n57124), .Y(n63691) );
  OAI22xp33_ASAP7_75t_SRAM U67843 ( .A1(or1200_cpu_or1200_except_n198), .A2(
        n58547), .B1(n77597), .B2(n59494), .Y(n77255) );
  OAI22xp33_ASAP7_75t_SRAM U67844 ( .A1(or1200_cpu_or1200_except_n204), .A2(
        n58547), .B1(n59554), .B2(n57124), .Y(n76829) );
  OAI21xp33_ASAP7_75t_SRAM U67845 ( .A1(n76828), .A2(n59494), .B(n76827), .Y(
        n76830) );
  INVxp33_ASAP7_75t_SRAM U67846 ( .A(n76826), .Y(n76827) );
  INVxp33_ASAP7_75t_SRAM U67847 ( .A(n77250), .Y(n76837) );
  OAI21xp33_ASAP7_75t_SRAM U67848 ( .A1(n60424), .A2(n60421), .B(n60422), .Y(
        n60406) );
  INVxp33_ASAP7_75t_SRAM U67849 ( .A(n60458), .Y(n60455) );
  OAI22xp33_ASAP7_75t_SRAM U67850 ( .A1(or1200_cpu_or1200_except_n194), .A2(
        n58547), .B1(n77591), .B2(n59494), .Y(n61581) );
  OAI21xp33_ASAP7_75t_SRAM U67851 ( .A1(n57086), .A2(n68809), .B(n68904), .Y(
        n58685) );
  OAI21xp33_ASAP7_75t_SRAM U67852 ( .A1(n68758), .A2(n68757), .B(n68756), .Y(
        n68759) );
  AOI22xp33_ASAP7_75t_SRAM U67853 ( .A1(n57198), .A2(n63744), .B1(n77918), 
        .B2(n63743), .Y(n63745) );
  OAI22xp33_ASAP7_75t_SRAM U67854 ( .A1(or1200_cpu_or1200_except_n216), .A2(
        n58547), .B1(n77019), .B2(n59494), .Y(n60160) );
  OAI22xp33_ASAP7_75t_SRAM U67855 ( .A1(or1200_cpu_or1200_except_n224), .A2(
        n58547), .B1(n74984), .B2(n77254), .Y(n60137) );
  OAI22xp33_ASAP7_75t_SRAM U67856 ( .A1(or1200_cpu_or1200_except_n226), .A2(
        n58547), .B1(n74639), .B2(n59494), .Y(n60128) );
  INVxp33_ASAP7_75t_SRAM U67857 ( .A(n77304), .Y(n60101) );
  OAI22xp33_ASAP7_75t_SRAM U67858 ( .A1(or1200_cpu_or1200_except_n218), .A2(
        n58547), .B1(n77646), .B2(n77254), .Y(n60093) );
  OAI22xp33_ASAP7_75t_SRAM U67859 ( .A1(n59547), .A2(n57124), .B1(n75620), 
        .B2(n59494), .Y(n60074) );
  OAI22xp33_ASAP7_75t_SRAM U67860 ( .A1(n59546), .A2(n57124), .B1(n75431), 
        .B2(n77254), .Y(n60063) );
  OAI22xp33_ASAP7_75t_SRAM U67861 ( .A1(or1200_cpu_or1200_except_n232), .A2(
        n58547), .B1(n59578), .B2(n57124), .Y(n60055) );
  OAI22xp33_ASAP7_75t_SRAM U67862 ( .A1(or1200_cpu_or1200_except_n214), .A2(
        n58547), .B1(n77637), .B2(n59494), .Y(n60046) );
  OAI21xp33_ASAP7_75t_SRAM U67863 ( .A1(n67441), .A2(n57456), .B(n67084), .Y(
        n67086) );
  INVxp33_ASAP7_75t_SRAM U67864 ( .A(n67147), .Y(n67148) );
  AOI21xp33_ASAP7_75t_SRAM U67865 ( .A1(n67861), .A2(n59659), .B(n59641), .Y(
        n67094) );
  OAI21xp33_ASAP7_75t_SRAM U67866 ( .A1(n75947), .A2(n68124), .B(n59641), .Y(
        n66246) );
  INVxp33_ASAP7_75t_SRAM U67867 ( .A(n67244), .Y(n66399) );
  OAI21xp33_ASAP7_75t_SRAM U67868 ( .A1(n75899), .A2(n57302), .B(n57292), .Y(
        n66402) );
  AOI21xp33_ASAP7_75t_SRAM U67869 ( .A1(n53298), .A2(n75899), .B(n57078), .Y(
        n66383) );
  AOI22xp33_ASAP7_75t_SRAM U67870 ( .A1(n59476), .A2(n59514), .B1(n59656), 
        .B2(n58424), .Y(n63271) );
  OAI21xp33_ASAP7_75t_SRAM U67871 ( .A1(n67850), .A2(n59476), .B(n62895), .Y(
        n63278) );
  OAI21xp33_ASAP7_75t_SRAM U67872 ( .A1(n76679), .A2(n75922), .B(n57881), .Y(
        n62894) );
  INVxp33_ASAP7_75t_SRAM U67873 ( .A(n62880), .Y(n62883) );
  INVxp33_ASAP7_75t_SRAM U67874 ( .A(n62575), .Y(n62659) );
  INVxp33_ASAP7_75t_SRAM U67875 ( .A(n62658), .Y(n62660) );
  AOI21xp33_ASAP7_75t_SRAM U67876 ( .A1(n59656), .A2(n58402), .B(n63120), .Y(
        n59119) );
  AOI21xp33_ASAP7_75t_SRAM U67877 ( .A1(n59670), .A2(n59606), .B(n58671), .Y(
        n58670) );
  INVxp33_ASAP7_75t_SRAM U67878 ( .A(n66798), .Y(n66799) );
  AOI22xp33_ASAP7_75t_SRAM U67879 ( .A1(n57213), .A2(n59654), .B1(n64026), 
        .B2(n64025), .Y(n64028) );
  INVxp33_ASAP7_75t_SRAM U67880 ( .A(n63808), .Y(n64932) );
  OAI21xp33_ASAP7_75t_SRAM U67881 ( .A1(n57310), .A2(n67536), .B(n67230), .Y(
        n64335) );
  INVxp33_ASAP7_75t_SRAM U67882 ( .A(n64389), .Y(n64390) );
  OAI21xp33_ASAP7_75t_SRAM U67883 ( .A1(n59653), .A2(n68097), .B(n59503), .Y(
        n64421) );
  INVxp33_ASAP7_75t_SRAM U67884 ( .A(n64503), .Y(n64505) );
  INVxp33_ASAP7_75t_SRAM U67885 ( .A(n64924), .Y(n64483) );
  OAI21xp33_ASAP7_75t_SRAM U67886 ( .A1(n58402), .A2(n59200), .B(n59659), .Y(
        n67542) );
  INVxp33_ASAP7_75t_SRAM U67887 ( .A(n68047), .Y(n68075) );
  INVxp33_ASAP7_75t_SRAM U67888 ( .A(n65034), .Y(n65035) );
  OAI21xp33_ASAP7_75t_SRAM U67889 ( .A1(n57347), .A2(n74799), .B(n53229), .Y(
        n64623) );
  INVxp33_ASAP7_75t_SRAM U67890 ( .A(n67354), .Y(n67357) );
  INVxp33_ASAP7_75t_SRAM U67891 ( .A(n67645), .Y(n58899) );
  INVxp33_ASAP7_75t_SRAM U67892 ( .A(n67308), .Y(n67309) );
  OAI21xp33_ASAP7_75t_SRAM U67893 ( .A1(n53316), .A2(n66258), .B(n62637), .Y(
        n62574) );
  INVxp33_ASAP7_75t_SRAM U67894 ( .A(n63172), .Y(n60929) );
  NOR2xp33_ASAP7_75t_SL U67895 ( .A(n77034), .B(n68810), .Y(n75408) );
  INVx1_ASAP7_75t_SL U67896 ( .A(n77675), .Y(n77645) );
  NAND2xp33_ASAP7_75t_SRAM U67897 ( .A(dwb_dat_i[23]), .B(n59696), .Y(n4264)
         );
  NAND2xp33_ASAP7_75t_SRAM U67898 ( .A(dwb_dat_i[21]), .B(n59696), .Y(n4269)
         );
  NAND2xp33_ASAP7_75t_SRAM U67899 ( .A(n78176), .B(n77977), .Y(n4313) );
  NAND2xp33_ASAP7_75t_SRAM U67900 ( .A(n78176), .B(n77980), .Y(n4312) );
  NAND2xp33_ASAP7_75t_SRAM U67901 ( .A(n78176), .B(n77974), .Y(n4314) );
  NAND2xp33_ASAP7_75t_SRAM U67902 ( .A(n78176), .B(n77983), .Y(n4311) );
  NAND2xp33_ASAP7_75t_SRAM U67903 ( .A(dwb_dat_i[19]), .B(n59696), .Y(n4277)
         );
  NAND2xp33_ASAP7_75t_SRAM U67904 ( .A(n78176), .B(n77986), .Y(n4310) );
  NAND2xp33_ASAP7_75t_SRAM U67905 ( .A(n78176), .B(n77992), .Y(n4309) );
  NAND2xp33_ASAP7_75t_SRAM U67906 ( .A(dwb_dat_i[18]), .B(n59696), .Y(n4280)
         );
  NAND2xp33_ASAP7_75t_SRAM U67907 ( .A(n78176), .B(n77968), .Y(n4316) );
  NAND2xp33_ASAP7_75t_SRAM U67908 ( .A(dwb_dat_i[17]), .B(n59696), .Y(n4283)
         );
  NAND2xp33_ASAP7_75t_SRAM U67909 ( .A(n78176), .B(n77971), .Y(n4315) );
  NAND2xp33_ASAP7_75t_SRAM U67910 ( .A(dwb_dat_i[20]), .B(n59696), .Y(n4272)
         );
  NAND2xp33_ASAP7_75t_SRAM U67911 ( .A(dwb_dat_i[16]), .B(n59696), .Y(n4286)
         );
  NAND2xp33_ASAP7_75t_SRAM U67912 ( .A(dwb_dat_i[15]), .B(n59696), .Y(n4289)
         );
  NAND2xp33_ASAP7_75t_SRAM U67913 ( .A(dwb_dat_i[14]), .B(n59696), .Y(n4292)
         );
  NAND2xp33_ASAP7_75t_SRAM U67914 ( .A(dwb_dat_i[13]), .B(n59696), .Y(n4295)
         );
  NAND2xp33_ASAP7_75t_SRAM U67915 ( .A(dwb_dat_i[12]), .B(n59696), .Y(n4298)
         );
  NAND2xp33_ASAP7_75t_SRAM U67916 ( .A(dwb_dat_i[11]), .B(n59696), .Y(n4301)
         );
  NAND2xp33_ASAP7_75t_SRAM U67917 ( .A(dwb_dat_i[9]), .B(n59696), .Y(n4226) );
  NAND2xp33_ASAP7_75t_SRAM U67918 ( .A(dwb_dat_i[8]), .B(n59696), .Y(n4229) );
  NAND2xp33_ASAP7_75t_SRAM U67919 ( .A(or1200_cpu_or1200_rf_addra_last_4_), 
        .B(n77962), .Y(or1200_cpu_or1200_rf_n130) );
  NAND2xp33_ASAP7_75t_SRAM U67920 ( .A(or1200_cpu_or1200_rf_addra_last_0_), 
        .B(n77962), .Y(or1200_cpu_or1200_rf_n142) );
  NAND2xp33_ASAP7_75t_SRAM U67921 ( .A(or1200_cpu_or1200_rf_addra_last_1_), 
        .B(n77962), .Y(or1200_cpu_or1200_rf_n139) );
  NAND2xp33_ASAP7_75t_SRAM U67922 ( .A(or1200_cpu_or1200_rf_addra_last_2_), 
        .B(n77962), .Y(or1200_cpu_or1200_rf_n136) );
  NAND2xp33_ASAP7_75t_SRAM U67923 ( .A(or1200_cpu_or1200_rf_addra_last_3_), 
        .B(n77962), .Y(or1200_cpu_or1200_rf_n133) );
  NAND2xp33_ASAP7_75t_SRAM U67924 ( .A(dwb_dat_i[25]), .B(n59696), .Y(n4255)
         );
  NAND2xp33_ASAP7_75t_SRAM U67925 ( .A(dwb_dat_i[29]), .B(n59696), .Y(n4247)
         );
  NAND2xp33_ASAP7_75t_SRAM U67926 ( .A(dwb_dat_i[26]), .B(n59696), .Y(n4253)
         );
  NAND2xp33_ASAP7_75t_SRAM U67927 ( .A(dwb_dat_i[31]), .B(n59696), .Y(n4241)
         );
  NAND2xp33_ASAP7_75t_SRAM U67928 ( .A(dwb_dat_i[24]), .B(n59696), .Y(n4257)
         );
  NAND2xp33_ASAP7_75t_SRAM U67929 ( .A(dwb_dat_i[30]), .B(n59696), .Y(n4243)
         );
  NAND2xp33_ASAP7_75t_SRAM U67930 ( .A(dwb_dat_i[28]), .B(n59696), .Y(n4249)
         );
  NAND2xp33_ASAP7_75t_SRAM U67931 ( .A(dwb_dat_i[22]), .B(n59696), .Y(n4266)
         );
  NAND2xp33_ASAP7_75t_SRAM U67932 ( .A(dwb_dat_i[2]), .B(n59696), .Y(n4245) );
  NAND2xp33_ASAP7_75t_SRAM U67933 ( .A(dwb_dat_i[3]), .B(n59696), .Y(n4239) );
  NAND2xp33_ASAP7_75t_SRAM U67934 ( .A(dwb_dat_i[0]), .B(n59696), .Y(n4305) );
  NAND2xp33_ASAP7_75t_SRAM U67935 ( .A(dwb_dat_i[10]), .B(n59696), .Y(n4303)
         );
  NAND2xp33_ASAP7_75t_SRAM U67936 ( .A(dwb_dat_i[27]), .B(n59696), .Y(n4251)
         );
  NAND2xp33_ASAP7_75t_SRAM U67937 ( .A(dwb_dat_i[5]), .B(n59696), .Y(n4235) );
  NAND2xp33_ASAP7_75t_SRAM U67938 ( .A(n77833), .B(n77832), .Y(n3645) );
  NAND2xp33_ASAP7_75t_SRAM U67939 ( .A(dwb_dat_i[6]), .B(n59696), .Y(n4233) );
  NAND2xp33_ASAP7_75t_SRAM U67940 ( .A(dwb_dat_i[1]), .B(n59696), .Y(n4274) );
  NAND2xp33_ASAP7_75t_SRAM U67941 ( .A(dwb_dat_i[7]), .B(n59696), .Y(n4231) );
  NAND2xp33_ASAP7_75t_SRAM U67942 ( .A(dwb_dat_i[4]), .B(n59696), .Y(n4237) );
  NAND2xp33_ASAP7_75t_SRAM U67943 ( .A(n77929), .B(n77923), .Y(
        or1200_cpu_or1200_rf_n116) );
  NAND2xp33_ASAP7_75t_SRAM U67944 ( .A(n77957), .B(n77936), .Y(
        or1200_cpu_or1200_rf_n131) );
  NAND2xp33_ASAP7_75t_SRAM U67945 ( .A(n77957), .B(n77942), .Y(
        or1200_cpu_or1200_rf_n134) );
  NAND2xp33_ASAP7_75t_SRAM U67946 ( .A(n77926), .B(n77929), .Y(
        or1200_cpu_or1200_rf_n122) );
  NAND2xp33_ASAP7_75t_SRAM U67947 ( .A(n77957), .B(n77946), .Y(
        or1200_cpu_or1200_rf_n137) );
  NAND2xp33_ASAP7_75t_SRAM U67948 ( .A(n77929), .B(n77865), .Y(
        or1200_cpu_or1200_rf_n60) );
  NAND2xp33_ASAP7_75t_SRAM U67949 ( .A(n77957), .B(n77951), .Y(
        or1200_cpu_or1200_rf_n140) );
  NAND2xp33_ASAP7_75t_SRAM U67950 ( .A(n77930), .B(n77929), .Y(
        or1200_cpu_or1200_rf_n128) );
  NAND2xp33_ASAP7_75t_SRAM U67951 ( .A(n77929), .B(n77914), .Y(
        or1200_cpu_or1200_rf_n104) );
  NAND2xp33_ASAP7_75t_SRAM U67952 ( .A(n77961), .B(n77957), .Y(
        or1200_cpu_or1200_rf_n144) );
  NOR2xp33_ASAP7_75t_SL U67953 ( .A(n78177), .B(n77952), .Y(n77957) );
  NAND2xp33_ASAP7_75t_SRAM U67954 ( .A(n77929), .B(n77912), .Y(
        or1200_cpu_or1200_rf_n102) );
  NAND2xp33_ASAP7_75t_SRAM U67955 ( .A(n77924), .B(n77929), .Y(
        or1200_cpu_or1200_rf_n118) );
  NAND2xp33_ASAP7_75t_SRAM U67956 ( .A(n77929), .B(n77870), .Y(
        or1200_cpu_or1200_rf_n64) );
  NAND2xp33_ASAP7_75t_SRAM U67957 ( .A(n77925), .B(n77929), .Y(
        or1200_cpu_or1200_rf_n120) );
  NAND2xp33_ASAP7_75t_SRAM U67958 ( .A(n77929), .B(n77861), .Y(
        or1200_cpu_or1200_rf_n56) );
  NAND2xp33_ASAP7_75t_SRAM U67959 ( .A(n77929), .B(n77884), .Y(
        or1200_cpu_or1200_rf_n76) );
  NAND2xp33_ASAP7_75t_SRAM U67960 ( .A(n77929), .B(n77921), .Y(
        or1200_cpu_or1200_rf_n112) );
  NAND2xp33_ASAP7_75t_SRAM U67961 ( .A(n77927), .B(n77929), .Y(
        or1200_cpu_or1200_rf_n124) );
  NAND2xp33_ASAP7_75t_SRAM U67962 ( .A(n77929), .B(n77874), .Y(
        or1200_cpu_or1200_rf_n68) );
  NAND2xp33_ASAP7_75t_SRAM U67963 ( .A(n77929), .B(n77858), .Y(
        or1200_cpu_or1200_rf_n54) );
  NAND2xp33_ASAP7_75t_SRAM U67964 ( .A(n77929), .B(n77892), .Y(
        or1200_cpu_or1200_rf_n82) );
  NAND2xp33_ASAP7_75t_SRAM U67965 ( .A(n77929), .B(n77876), .Y(
        or1200_cpu_or1200_rf_n70) );
  NAND2xp33_ASAP7_75t_SRAM U67966 ( .A(n77929), .B(n77855), .Y(
        or1200_cpu_or1200_rf_n52) );
  NAND2xp33_ASAP7_75t_SRAM U67967 ( .A(n77879), .B(n77929), .Y(
        or1200_cpu_or1200_rf_n72) );
  NAND2xp33_ASAP7_75t_SRAM U67968 ( .A(n77929), .B(n77909), .Y(
        or1200_cpu_or1200_rf_n98) );
  NAND2xp33_ASAP7_75t_SRAM U67969 ( .A(n77929), .B(n77863), .Y(
        or1200_cpu_or1200_rf_n58) );
  NAND2xp33_ASAP7_75t_SRAM U67970 ( .A(n77929), .B(n77882), .Y(
        or1200_cpu_or1200_rf_n74) );
  NAND2xp33_ASAP7_75t_SRAM U67971 ( .A(n77929), .B(n77908), .Y(
        or1200_cpu_or1200_rf_n96) );
  NAND2xp33_ASAP7_75t_SRAM U67972 ( .A(n77929), .B(n77903), .Y(
        or1200_cpu_or1200_rf_n90) );
  NAND2xp33_ASAP7_75t_SRAM U67973 ( .A(n77929), .B(n77898), .Y(
        or1200_cpu_or1200_rf_n86) );
  NAND2xp33_ASAP7_75t_SRAM U67974 ( .A(n77929), .B(n77900), .Y(
        or1200_cpu_or1200_rf_n88) );
  NAND2xp33_ASAP7_75t_SRAM U67975 ( .A(n77929), .B(n77915), .Y(
        or1200_cpu_or1200_rf_n106) );
  NAND2xp33_ASAP7_75t_SRAM U67976 ( .A(n77929), .B(n77904), .Y(
        or1200_cpu_or1200_rf_n92) );
  NAND2xp33_ASAP7_75t_SRAM U67977 ( .A(n77929), .B(n77887), .Y(
        or1200_cpu_or1200_rf_n78) );
  NAND2xp33_ASAP7_75t_SRAM U67978 ( .A(n77929), .B(n77919), .Y(
        or1200_cpu_or1200_rf_n110) );
  NAND2xp33_ASAP7_75t_SRAM U67979 ( .A(n77929), .B(n77868), .Y(
        or1200_cpu_or1200_rf_n62) );
  NAND2xp33_ASAP7_75t_SRAM U67980 ( .A(n77929), .B(n77872), .Y(
        or1200_cpu_or1200_rf_n66) );
  NAND2xp33_ASAP7_75t_SRAM U67981 ( .A(n77929), .B(n77917), .Y(
        or1200_cpu_or1200_rf_n108) );
  NAND2xp33_ASAP7_75t_SRAM U67982 ( .A(n77929), .B(n77889), .Y(
        or1200_cpu_or1200_rf_n80) );
  NAND2xp33_ASAP7_75t_SRAM U67983 ( .A(n77929), .B(n77911), .Y(
        or1200_cpu_or1200_rf_n100) );
  NAND2xp33_ASAP7_75t_SRAM U67984 ( .A(n77929), .B(n77906), .Y(
        or1200_cpu_or1200_rf_n94) );
  NAND2xp33_ASAP7_75t_SRAM U67985 ( .A(n77929), .B(n77895), .Y(
        or1200_cpu_or1200_rf_n84) );
  NAND2xp33_ASAP7_75t_SRAM U67986 ( .A(n77931), .B(n77952), .Y(
        or1200_cpu_or1200_rf_n132) );
  NAND2xp33_ASAP7_75t_SRAM U67987 ( .A(n77937), .B(n77928), .Y(
        or1200_cpu_or1200_rf_n121) );
  NAND2xp33_ASAP7_75t_SRAM U67988 ( .A(n59493), .B(n77952), .Y(
        or1200_cpu_or1200_rf_n145) );
  NAND2xp33_ASAP7_75t_SRAM U67989 ( .A(n77943), .B(n77928), .Y(
        or1200_cpu_or1200_rf_n123) );
  NAND2xp33_ASAP7_75t_SRAM U67990 ( .A(n77952), .B(n77965), .Y(
        or1200_cpu_or1200_rf_n141) );
  NAND2xp33_ASAP7_75t_SRAM U67991 ( .A(n77928), .B(n77862), .Y(
        or1200_cpu_or1200_rf_n59) );
  NAND2xp33_ASAP7_75t_SRAM U67992 ( .A(n77928), .B(n77871), .Y(
        or1200_cpu_or1200_rf_n67) );
  NAND2xp33_ASAP7_75t_SRAM U67993 ( .A(n77937), .B(n77952), .Y(
        or1200_cpu_or1200_rf_n135) );
  NAND2xp33_ASAP7_75t_SRAM U67994 ( .A(n77928), .B(n77869), .Y(
        or1200_cpu_or1200_rf_n65) );
  NAND2xp33_ASAP7_75t_SRAM U67995 ( .A(n77928), .B(n77873), .Y(
        or1200_cpu_or1200_rf_n69) );
  NAND2xp33_ASAP7_75t_SRAM U67996 ( .A(n59493), .B(n77928), .Y(
        or1200_cpu_or1200_rf_n129) );
  NAND2xp33_ASAP7_75t_SRAM U67997 ( .A(n77928), .B(n77866), .Y(
        or1200_cpu_or1200_rf_n63) );
  NAND2xp33_ASAP7_75t_SRAM U67998 ( .A(n77928), .B(n77875), .Y(
        or1200_cpu_or1200_rf_n71) );
  NAND2xp33_ASAP7_75t_SRAM U67999 ( .A(n77928), .B(n77854), .Y(
        or1200_cpu_or1200_rf_n53) );
  NAND2xp33_ASAP7_75t_SRAM U68000 ( .A(n77928), .B(n77877), .Y(
        or1200_cpu_or1200_rf_n73) );
  NAND2xp33_ASAP7_75t_SRAM U68001 ( .A(n77928), .B(n77864), .Y(
        or1200_cpu_or1200_rf_n61) );
  NAND2xp33_ASAP7_75t_SRAM U68002 ( .A(n77928), .B(n77856), .Y(
        or1200_cpu_or1200_rf_n55) );
  NAND2xp33_ASAP7_75t_SRAM U68003 ( .A(n77928), .B(n77880), .Y(
        or1200_cpu_or1200_rf_n75) );
  NAND2xp33_ASAP7_75t_SRAM U68004 ( .A(n77928), .B(n77859), .Y(
        or1200_cpu_or1200_rf_n57) );
  NAND2xp33_ASAP7_75t_SRAM U68005 ( .A(n77928), .B(n77883), .Y(
        or1200_cpu_or1200_rf_n77) );
  NAND2xp33_ASAP7_75t_SRAM U68006 ( .A(n77931), .B(n77928), .Y(
        or1200_cpu_or1200_rf_n119) );
  NAND2xp33_ASAP7_75t_SRAM U68007 ( .A(n77928), .B(n77965), .Y(
        or1200_cpu_or1200_rf_n125) );
  NAND2xp33_ASAP7_75t_SRAM U68008 ( .A(n77928), .B(n77885), .Y(
        or1200_cpu_or1200_rf_n79) );
  NAND2xp33_ASAP7_75t_SRAM U68009 ( .A(n77943), .B(n77952), .Y(
        or1200_cpu_or1200_rf_n138) );
  NAND2xp33_ASAP7_75t_SRAM U68010 ( .A(n77928), .B(n77986), .Y(
        or1200_cpu_or1200_rf_n99) );
  NAND2xp33_ASAP7_75t_SRAM U68011 ( .A(n77928), .B(n77888), .Y(
        or1200_cpu_or1200_rf_n81) );
  NAND2xp33_ASAP7_75t_SRAM U68012 ( .A(n77928), .B(n77890), .Y(
        or1200_cpu_or1200_rf_n83) );
  NAND2xp33_ASAP7_75t_SRAM U68013 ( .A(n77928), .B(n77922), .Y(
        or1200_cpu_or1200_rf_n117) );
  NAND2xp33_ASAP7_75t_SRAM U68014 ( .A(n77928), .B(n77893), .Y(
        or1200_cpu_or1200_rf_n85) );
  NAND2xp33_ASAP7_75t_SRAM U68015 ( .A(n77928), .B(n77992), .Y(
        or1200_cpu_or1200_rf_n97) );
  NAND2xp33_ASAP7_75t_SRAM U68016 ( .A(n77928), .B(n77896), .Y(
        or1200_cpu_or1200_rf_n87) );
  NAND2xp33_ASAP7_75t_SRAM U68017 ( .A(n77928), .B(n77977), .Y(
        or1200_cpu_or1200_rf_n105) );
  NAND2xp33_ASAP7_75t_SRAM U68018 ( .A(n77928), .B(n77899), .Y(
        or1200_cpu_or1200_rf_n89) );
  NAND2xp33_ASAP7_75t_SRAM U68019 ( .A(n77928), .B(n77916), .Y(
        or1200_cpu_or1200_rf_n109) );
  NAND2xp33_ASAP7_75t_SRAM U68020 ( .A(n77928), .B(n77901), .Y(
        or1200_cpu_or1200_rf_n91) );
  NAND2xp33_ASAP7_75t_SRAM U68021 ( .A(n77928), .B(n77971), .Y(
        or1200_cpu_or1200_rf_n93) );
  NAND2xp33_ASAP7_75t_SRAM U68022 ( .A(n77928), .B(n77968), .Y(
        or1200_cpu_or1200_rf_n95) );
  NAND2xp33_ASAP7_75t_SRAM U68023 ( .A(n77928), .B(n77983), .Y(
        or1200_cpu_or1200_rf_n101) );
  NAND2xp33_ASAP7_75t_SRAM U68024 ( .A(n77928), .B(n77918), .Y(
        or1200_cpu_or1200_rf_n111) );
  NAND2xp33_ASAP7_75t_SRAM U68025 ( .A(n77928), .B(n77980), .Y(
        or1200_cpu_or1200_rf_n103) );
  NAND2xp33_ASAP7_75t_SRAM U68026 ( .A(n77928), .B(n77920), .Y(
        or1200_cpu_or1200_rf_n113) );
  NAND2xp33_ASAP7_75t_SRAM U68027 ( .A(n77928), .B(n77974), .Y(
        or1200_cpu_or1200_rf_n107) );
  NAND2xp33_ASAP7_75t_SRAM U68028 ( .A(n3105), .B(n78002), .Y(n4230) );
  NAND2xp33_ASAP7_75t_SRAM U68029 ( .A(n77929), .B(n77849), .Y(
        or1200_cpu_or1200_rf_N31) );
  NAND2xp33_ASAP7_75t_SRAM U68030 ( .A(n3105), .B(n59443), .Y(n4273) );
  NAND2xp33_ASAP7_75t_SRAM U68031 ( .A(n3086), .B(n78163), .Y(n78164) );
  NAND2xp33_ASAP7_75t_SRAM U68032 ( .A(n3105), .B(n59709), .Y(n4244) );
  NAND2xp33_ASAP7_75t_SRAM U68033 ( .A(n3105), .B(n57214), .Y(n4238) );
  NAND2xp33_ASAP7_75t_SRAM U68034 ( .A(n3105), .B(n78004), .Y(n4234) );
  NAND2xp33_ASAP7_75t_SRAM U68035 ( .A(n3105), .B(n78005), .Y(n4236) );
  NAND2xp33_ASAP7_75t_SRAM U68036 ( .A(n3105), .B(n59712), .Y(n4304) );
  NAND2xp33_ASAP7_75t_SRAM U68037 ( .A(n3105), .B(n78003), .Y(n4232) );
  NAND2xp33_ASAP7_75t_SRAM U68038 ( .A(or1200_dc_top_from_dcram_31_), .B(
        n77748), .Y(n77747) );
  NAND2xp33_ASAP7_75t_SRAM U68039 ( .A(or1200_dc_top_from_dcram_10_), .B(
        n77748), .Y(n77698) );
  NAND2xp33_ASAP7_75t_SRAM U68040 ( .A(or1200_dc_top_from_dcram_9_), .B(n77748), .Y(n77697) );
  NAND2xp33_ASAP7_75t_SRAM U68041 ( .A(n77696), .B(n77704), .Y(n4225) );
  NAND2xp33_ASAP7_75t_SRAM U68042 ( .A(n77706), .B(n59443), .Y(n4224) );
  NAND2xp33_ASAP7_75t_SRAM U68043 ( .A(or1200_dc_top_from_dcram_8_), .B(n77748), .Y(n77695) );
  NAND2xp33_ASAP7_75t_SRAM U68044 ( .A(n56954), .B(n77704), .Y(n4228) );
  NAND2xp33_ASAP7_75t_SRAM U68045 ( .A(n77706), .B(n59712), .Y(n4227) );
  NAND2xp33_ASAP7_75t_SRAM U68046 ( .A(or1200_dc_top_from_dcram_7_), .B(n77748), .Y(n77694) );
  NAND2xp33_ASAP7_75t_SRAM U68047 ( .A(or1200_dc_top_from_dcram_6_), .B(n77748), .Y(n77693) );
  NAND2xp33_ASAP7_75t_SRAM U68048 ( .A(or1200_dc_top_from_dcram_5_), .B(n77748), .Y(n77692) );
  NAND2xp33_ASAP7_75t_SRAM U68049 ( .A(or1200_dc_top_from_dcram_4_), .B(n77748), .Y(n77691) );
  NAND2xp33_ASAP7_75t_SRAM U68050 ( .A(or1200_dc_top_from_dcram_3_), .B(n77748), .Y(n77690) );
  NAND2xp33_ASAP7_75t_SRAM U68051 ( .A(or1200_dc_top_from_dcram_2_), .B(n77748), .Y(n77689) );
  NAND2xp33_ASAP7_75t_SRAM U68052 ( .A(or1200_dc_top_from_dcram_1_), .B(n77748), .Y(n77688) );
  NAND2xp33_ASAP7_75t_SRAM U68053 ( .A(or1200_dc_top_from_dcram_0_), .B(n77748), .Y(n77687) );
  NOR4xp25_ASAP7_75t_SL U68054 ( .A(n77577), .B(n77576), .C(n77575), .D(n77574), .Y(n77578) );
  NOR4xp25_ASAP7_75t_SL U68055 ( .A(n77573), .B(n77572), .C(n77571), .D(n77570), .Y(n77579) );
  NAND2xp33_ASAP7_75t_SRAM U68056 ( .A(or1200_dc_top_from_dcram_11_), .B(
        n77748), .Y(n77699) );
  NAND2xp33_ASAP7_75t_SRAM U68057 ( .A(n57219), .B(n77704), .Y(n4300) );
  NAND2xp33_ASAP7_75t_SRAM U68058 ( .A(n77706), .B(n57214), .Y(n4299) );
  NAND2xp33_ASAP7_75t_SRAM U68059 ( .A(or1200_dc_top_from_dcram_12_), .B(
        n77748), .Y(n77700) );
  NAND2xp33_ASAP7_75t_SRAM U68060 ( .A(n59387), .B(n77704), .Y(n4297) );
  NAND2xp33_ASAP7_75t_SRAM U68061 ( .A(n77706), .B(n78005), .Y(n4296) );
  NAND2xp33_ASAP7_75t_SRAM U68062 ( .A(or1200_dc_top_from_dcram_13_), .B(
        n77748), .Y(n77702) );
  NAND2xp33_ASAP7_75t_SRAM U68063 ( .A(n77701), .B(n77704), .Y(n4294) );
  NAND2xp33_ASAP7_75t_SRAM U68064 ( .A(n77706), .B(n78004), .Y(n4293) );
  NAND2xp33_ASAP7_75t_SRAM U68065 ( .A(or1200_dc_top_from_dcram_14_), .B(
        n77748), .Y(n77703) );
  NAND2xp33_ASAP7_75t_SRAM U68066 ( .A(n57213), .B(n77704), .Y(n4291) );
  NAND2xp33_ASAP7_75t_SRAM U68067 ( .A(n77706), .B(n78003), .Y(n4290) );
  NAND2xp33_ASAP7_75t_SRAM U68068 ( .A(or1200_dc_top_from_dcram_15_), .B(
        n77748), .Y(n77707) );
  NAND2xp33_ASAP7_75t_SRAM U68069 ( .A(n77705), .B(n77704), .Y(n4288) );
  INVx1_ASAP7_75t_SL U68070 ( .A(n77706), .Y(n77704) );
  NAND2xp33_ASAP7_75t_SRAM U68071 ( .A(n77706), .B(n78002), .Y(n4287) );
  NOR2xp33_ASAP7_75t_SL U68072 ( .A(n77725), .B(n77753), .Y(n77706) );
  NAND2xp33_ASAP7_75t_SRAM U68073 ( .A(or1200_dc_top_from_dcram_16_), .B(
        n77748), .Y(n77710) );
  NAND2xp33_ASAP7_75t_SRAM U68074 ( .A(n59712), .B(n77721), .Y(n4285) );
  NAND2xp33_ASAP7_75t_SRAM U68075 ( .A(n77723), .B(n77709), .Y(n4284) );
  NAND2xp33_ASAP7_75t_SRAM U68076 ( .A(or1200_dc_top_from_dcram_17_), .B(
        n77748), .Y(n77712) );
  NAND2xp33_ASAP7_75t_SRAM U68077 ( .A(n59443), .B(n77721), .Y(n4282) );
  NAND2xp33_ASAP7_75t_SRAM U68078 ( .A(n77723), .B(n77711), .Y(n4281) );
  NAND2xp33_ASAP7_75t_SRAM U68079 ( .A(or1200_dc_top_from_dcram_18_), .B(
        n77748), .Y(n77714) );
  NAND2xp33_ASAP7_75t_SRAM U68080 ( .A(n59709), .B(n77721), .Y(n4279) );
  NAND2xp33_ASAP7_75t_SRAM U68081 ( .A(n77723), .B(n77713), .Y(n4278) );
  NAND2xp33_ASAP7_75t_SRAM U68082 ( .A(or1200_dc_top_from_dcram_19_), .B(
        n77748), .Y(n77716) );
  NAND2xp33_ASAP7_75t_SRAM U68083 ( .A(n57214), .B(n77721), .Y(n4276) );
  NAND2xp33_ASAP7_75t_SRAM U68084 ( .A(n77723), .B(n77715), .Y(n4275) );
  NAND2xp33_ASAP7_75t_SRAM U68085 ( .A(or1200_dc_top_from_dcram_20_), .B(
        n77748), .Y(n77718) );
  NAND2xp33_ASAP7_75t_SRAM U68086 ( .A(n78005), .B(n77721), .Y(n4271) );
  NAND2xp33_ASAP7_75t_SRAM U68087 ( .A(n77723), .B(n77717), .Y(n4270) );
  NAND2xp33_ASAP7_75t_SRAM U68088 ( .A(or1200_dc_top_from_dcram_21_), .B(
        n77748), .Y(n77719) );
  NAND2xp33_ASAP7_75t_SRAM U68089 ( .A(n78004), .B(n77721), .Y(n4268) );
  NAND2xp33_ASAP7_75t_SRAM U68090 ( .A(n77723), .B(n57218), .Y(n4267) );
  NAND2xp33_ASAP7_75t_SRAM U68091 ( .A(or1200_dc_top_from_dcram_22_), .B(
        n77748), .Y(n77720) );
  NAND2xp33_ASAP7_75t_SRAM U68092 ( .A(or1200_dc_top_from_dcram_23_), .B(
        n77748), .Y(n77724) );
  NAND2xp33_ASAP7_75t_SRAM U68093 ( .A(n78002), .B(n77721), .Y(n4263) );
  NAND2xp33_ASAP7_75t_SRAM U68094 ( .A(n77723), .B(n77722), .Y(n4262) );
  NOR2xp33_ASAP7_75t_SL U68095 ( .A(n77754), .B(n77725), .Y(n77723) );
  NAND2xp33_ASAP7_75t_SRAM U68096 ( .A(or1200_dc_top_from_dcram_24_), .B(
        n77748), .Y(n77731) );
  NAND2xp33_ASAP7_75t_SRAM U68097 ( .A(or1200_dc_top_from_dcram_25_), .B(
        n77748), .Y(n77733) );
  NAND2xp33_ASAP7_75t_SRAM U68098 ( .A(or1200_dc_top_from_dcram_30_), .B(
        n77748), .Y(n77743) );
  NAND2xp33_ASAP7_75t_SRAM U68099 ( .A(or1200_dc_top_from_dcram_26_), .B(
        n77748), .Y(n77736) );
  NAND2xp33_ASAP7_75t_SRAM U68100 ( .A(or1200_dc_top_from_dcram_27_), .B(
        n77748), .Y(n77737) );
  NAND2xp33_ASAP7_75t_SRAM U68101 ( .A(or1200_dc_top_from_dcram_28_), .B(
        n77748), .Y(n77739) );
  NAND2xp33_ASAP7_75t_SRAM U68102 ( .A(or1200_dc_top_from_dcram_29_), .B(
        n77748), .Y(n77740) );
  NAND2xp33_ASAP7_75t_SRAM U68103 ( .A(n77751), .B(n77727), .Y(n77745) );
  NOR2xp33_ASAP7_75t_SL U68104 ( .A(n77726), .B(n77728), .Y(n77741) );
  NOR2xp33_ASAP7_75t_SL U68105 ( .A(n77729), .B(n77728), .Y(n77742) );
  NAND2xp33_ASAP7_75t_SRAM U68106 ( .A(n60274), .B(n60273), .Y(n60275) );
  NOR2xp33_ASAP7_75t_SL U68107 ( .A(n61280), .B(n57084), .Y(n60278) );
  AOI211xp5_ASAP7_75t_SL U68108 ( .A1(n833), .A2(n77793), .B(n57084), .C(
        n77803), .Y(n77794) );
  AOI31xp33_ASAP7_75t_SL U68109 ( .A1(n70296), .A2(n69377), .A3(n2451), .B(
        n70477), .Y(n69378) );
  NAND2xp33_ASAP7_75t_SRAM U68110 ( .A(n77418), .B(n77417), .Y(n77419) );
  NOR2xp33_ASAP7_75t_SL U68111 ( .A(clmode_i[1]), .B(clmode_i[0]), .Y(n61280)
         );
  NOR2xp33_ASAP7_75t_SL U68112 ( .A(n27499), .B(n70530), .Y(n70527) );
  NAND2xp33_ASAP7_75t_SRAM U68113 ( .A(n74285), .B(n74284), .Y(n74287) );
  NOR2xp33_ASAP7_75t_SL U68114 ( .A(n2473), .B(n62006), .Y(
        or1200_cpu_or1200_mult_mac_N294) );
  NOR2xp33_ASAP7_75t_SL U68115 ( .A(n53250), .B(n62006), .Y(
        or1200_cpu_or1200_mult_mac_N292) );
  NOR2xp33_ASAP7_75t_SL U68116 ( .A(n2501), .B(n62006), .Y(
        or1200_cpu_or1200_mult_mac_N293) );
  NOR2xp33_ASAP7_75t_SL U68117 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_), .B(n78243), .Y(n52547)
         );
  NOR2xp33_ASAP7_75t_SL U68118 ( .A(n3423), .B(n77759), .Y(n77755) );
  NOR2xp33_ASAP7_75t_SL U68119 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_23_), .B(n78244), .Y(
        n52549) );
  NOR2xp33_ASAP7_75t_SL U68120 ( .A(n59710), .B(n76679), .Y(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N1) );
  NOR2xp33_ASAP7_75t_SL U68121 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_3_), .B(n62055), .Y(n62058) );
  AOI211xp5_ASAP7_75t_SL U68122 ( .A1(n73663), .A2(n73763), .B(n73648), .C(
        n73647), .Y(n73649) );
  NOR2xp33_ASAP7_75t_SL U68123 ( .A(n70405), .B(n70451), .Y(n70366) );
  NOR2xp33_ASAP7_75t_SL U68124 ( .A(n70407), .B(n70406), .Y(n2364) );
  NOR2xp33_ASAP7_75t_SL U68125 ( .A(n74655), .B(n70488), .Y(n70472) );
  NOR2xp33_ASAP7_75t_SL U68126 ( .A(n74513), .B(n2934), .Y(n74516) );
  NOR2xp33_ASAP7_75t_SL U68127 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B(
        n70470), .Y(n70302) );
  NOR2xp33_ASAP7_75t_SL U68128 ( .A(n70535), .B(n70537), .Y(n70550) );
  AOI211xp5_ASAP7_75t_SL U68129 ( .A1(n70545), .A2(n70333), .B(n70332), .C(
        n70331), .Y(n2328) );
  NOR2xp33_ASAP7_75t_SL U68130 ( .A(n70405), .B(n70547), .Y(n70331) );
  NOR2xp33_ASAP7_75t_SL U68131 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .B(
        n70295), .Y(n70401) );
  AOI211xp5_ASAP7_75t_SL U68132 ( .A1(n74686), .A2(n74691), .B(n70329), .C(
        n70328), .Y(n70330) );
  NOR2xp33_ASAP7_75t_SL U68133 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B(
        n70405), .Y(n70545) );
  NOR2xp33_ASAP7_75t_SL U68134 ( .A(n74706), .B(n70388), .Y(n70321) );
  NOR2xp33_ASAP7_75t_SL U68135 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_2_), .B(n62038), .Y(n62039) );
  NOR2xp33_ASAP7_75t_SL U68136 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_1_), .B(n62037), .Y(n62040) );
  NAND2xp33_ASAP7_75t_SRAM U68137 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_0_), .Y(n62037) );
  NOR2xp33_ASAP7_75t_SL U68138 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_0_), .B(n62046), .Y(n62041) );
  NOR2xp33_ASAP7_75t_SL U68139 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_4_), .B(or1200_cpu_or1200_fpu_fpu_arith_s_count_3_), .Y(n62060) );
  NOR2xp33_ASAP7_75t_SL U68140 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_0_), .B(or1200_cpu_or1200_fpu_fpu_arith_s_count_5_), .Y(n62036) );
  NOR2xp33_ASAP7_75t_SL U68141 ( .A(n62054), .B(n62053), .Y(n62056) );
  NAND2xp33_ASAP7_75t_SRAM U68142 ( .A(n70317), .B(n74680), .Y(n70318) );
  NOR2xp33_ASAP7_75t_SL U68143 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .B(
        n70359), .Y(n70387) );
  AOI31xp33_ASAP7_75t_SL U68144 ( .A1(n70475), .A2(n70551), .A3(n70474), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .Y(
        n70375) );
  NOR2xp33_ASAP7_75t_SL U68145 ( .A(n70338), .B(n70337), .Y(n70373) );
  NOR2xp33_ASAP7_75t_SL U68146 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_11_), .B(
        n70440), .Y(n70412) );
  NOR2xp33_ASAP7_75t_SL U68147 ( .A(n70267), .B(n70266), .Y(n70301) );
  NOR2xp33_ASAP7_75t_SL U68148 ( .A(n70300), .B(n70299), .Y(n70339) );
  NAND2xp33_ASAP7_75t_SRAM U68149 ( .A(n70354), .B(n74680), .Y(n70345) );
  NAND2xp33_ASAP7_75t_SRAM U68150 ( .A(n2442), .B(n74680), .Y(n70380) );
  NOR2xp33_ASAP7_75t_SL U68151 ( .A(n70425), .B(n70424), .Y(n70489) );
  NAND2xp33_ASAP7_75t_SRAM U68152 ( .A(n74655), .B(n74680), .Y(n70390) );
  NOR2xp33_ASAP7_75t_SL U68153 ( .A(n58620), .B(n70250), .Y(n70359) );
  NOR2xp33_ASAP7_75t_SL U68154 ( .A(DP_OP_741J1_129_6992_n46), .B(n70540), .Y(
        n70250) );
  NOR2xp33_ASAP7_75t_SL U68155 ( .A(n74706), .B(n70389), .Y(n70450) );
  NAND2xp33_ASAP7_75t_SRAM U68156 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_), .B(
        n74680), .Y(n70314) );
  NOR2xp33_ASAP7_75t_SL U68157 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .B(
        n70536), .Y(n70451) );
  NAND2xp33_ASAP7_75t_SRAM U68158 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .B(
        n74680), .Y(n70355) );
  NOR2xp33_ASAP7_75t_SL U68159 ( .A(n70427), .B(n70426), .Y(n70444) );
  OR2x2_ASAP7_75t_SL U68160 ( .A(n74718), .B(n70272), .Y(n70405) );
  AOI211xp5_ASAP7_75t_SL U68161 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_8_), .A2(
        n74686), .B(n70442), .C(n70441), .Y(n70538) );
  NOR2xp33_ASAP7_75t_SL U68162 ( .A(n70439), .B(n70488), .Y(n70442) );
  NOR2xp33_ASAP7_75t_SL U68163 ( .A(n70402), .B(n74706), .Y(n70539) );
  NOR2xp33_ASAP7_75t_SL U68164 ( .A(n70426), .B(n70383), .Y(n70469) );
  NOR2xp33_ASAP7_75t_SL U68165 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_4_), .B(
        n70537), .Y(n70383) );
  NOR2xp33_ASAP7_75t_SL U68166 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .B(
        n70537), .Y(n70426) );
  NOR2xp33_ASAP7_75t_SL U68167 ( .A(n70459), .B(n70458), .Y(n70544) );
  NAND2xp33_ASAP7_75t_SRAM U68168 ( .A(n74674), .B(n74680), .Y(n70457) );
  NAND2xp33_ASAP7_75t_SRAM U68169 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_7_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_), .Y(
        n70456) );
  NOR2xp33_ASAP7_75t_SL U68170 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .B(
        n70440), .Y(n70445) );
  AOI211xp5_ASAP7_75t_SL U68171 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_), .A2(
        n74686), .B(n70292), .C(n70291), .Y(n70294) );
  NOR2xp33_ASAP7_75t_SL U68172 ( .A(n70317), .B(n70540), .Y(n70292) );
  NOR2xp33_ASAP7_75t_SL U68173 ( .A(n70552), .B(n70540), .Y(n70257) );
  NOR2xp33_ASAP7_75t_SL U68174 ( .A(DP_OP_741J1_129_6992_n46), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_), .Y(
        n70258) );
  NOR2xp33_ASAP7_75t_SL U68175 ( .A(n77499), .B(n77498), .Y(n6739) );
  NOR2xp33_ASAP7_75t_SL U68176 ( .A(n77497), .B(n4318), .Y(n77498) );
  NOR2xp33_ASAP7_75t_SL U68177 ( .A(n77234), .B(n77301), .Y(n2409) );
  NOR2xp33_ASAP7_75t_SL U68178 ( .A(n75455), .B(n77301), .Y(n2950) );
  NOR2xp33_ASAP7_75t_SL U68179 ( .A(n74550), .B(n76985), .Y(n74551) );
  NOR2xp33_ASAP7_75t_SL U68180 ( .A(n74546), .B(n74545), .Y(n74547) );
  NOR4xp25_ASAP7_75t_SL U68181 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_3_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_2_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_5_), .Y(n74541) );
  NOR4xp25_ASAP7_75t_SL U68182 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_7_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_6_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_9_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_10_), .Y(n74542) );
  NOR4xp25_ASAP7_75t_SL U68183 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_12_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_13_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_14_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_15_), .Y(n74543) );
  NOR4xp25_ASAP7_75t_SL U68184 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_16_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_19_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_21_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_20_), .Y(n74544) );
  NOR4xp25_ASAP7_75t_SL U68185 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_22_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_8_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_23_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_0_), .Y(n74539) );
  NOR4xp25_ASAP7_75t_SL U68186 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_11_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_17_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_18_), .Y(n74540) );
  NOR4xp25_ASAP7_75t_SL U68187 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_33_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_32_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_31_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_35_), .Y(n74534) );
  NOR4xp25_ASAP7_75t_SL U68188 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_34_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_36_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_38_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_41_), .Y(n74535) );
  NOR4xp25_ASAP7_75t_SL U68189 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_42_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_39_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_40_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_45_), .Y(n74536) );
  NOR4xp25_ASAP7_75t_SL U68190 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_48_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_47_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_46_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_49_), .Y(n74537) );
  NOR4xp25_ASAP7_75t_SL U68191 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_27_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_37_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_43_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_44_), .Y(n74532) );
  NOR4xp25_ASAP7_75t_SL U68192 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_30_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_29_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_28_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvdnd_i_26_), .Y(n74533) );
  NOR2xp33_ASAP7_75t_SL U68193 ( .A(n2944), .B(n78249), .Y(n74531) );
  NOR2xp33_ASAP7_75t_SL U68194 ( .A(n77234), .B(n74770), .Y(n74757) );
  NOR2xp33_ASAP7_75t_SL U68195 ( .A(n74525), .B(n74524), .Y(n74526) );
  NOR2xp33_ASAP7_75t_SL U68196 ( .A(n74523), .B(n74522), .Y(n74527) );
  NOR2xp33_ASAP7_75t_SL U68197 ( .A(n74521), .B(n74520), .Y(n74528) );
  NAND2xp33_ASAP7_75t_SRAM U68198 ( .A(dwb_adr_o[2]), .B(n77773), .Y(n77775)
         );
  AOI211xp5_ASAP7_75t_SL U68199 ( .A1(n59625), .A2(n72464), .B(n72420), .C(
        n72419), .Y(n72429) );
  NOR2xp33_ASAP7_75t_SL U68200 ( .A(n59622), .B(n72466), .Y(n72420) );
  NOR2xp33_ASAP7_75t_SL U68201 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .B(
        n59705), .Y(n73813) );
  AOI31xp33_ASAP7_75t_SL U68202 ( .A1(n59618), .A2(n59656), .A3(n59514), .B(
        n63271), .Y(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_mult_x_1_n211) );
  AOI211xp5_ASAP7_75t_SL U68203 ( .A1(n72131), .A2(n72396), .B(n72099), .C(
        n72098), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n91) );
  NOR2xp33_ASAP7_75t_SL U68204 ( .A(n72390), .B(n72106), .Y(n72099) );
  AOI211xp5_ASAP7_75t_SL U68205 ( .A1(n73774), .A2(n59705), .B(n73793), .C(
        n73773), .Y(n73775) );
  NOR2xp33_ASAP7_75t_SL U68206 ( .A(n73791), .B(n73830), .Y(n73773) );
  NOR2xp33_ASAP7_75t_SL U68207 ( .A(n57192), .B(n72210), .Y(n72475) );
  NOR2xp33_ASAP7_75t_SL U68208 ( .A(n72216), .B(n72215), .Y(n72473) );
  AOI211xp5_ASAP7_75t_SL U68209 ( .A1(n72131), .A2(n72369), .B(n72130), .C(
        n72129), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n90) );
  AOI211xp5_ASAP7_75t_SL U68210 ( .A1(n72126), .A2(n72125), .B(n72124), .C(
        n72123), .Y(n72128) );
  NOR2xp33_ASAP7_75t_SL U68211 ( .A(n72122), .B(n72121), .Y(n72123) );
  NOR2xp33_ASAP7_75t_SL U68212 ( .A(n72119), .B(n72118), .Y(n72124) );
  NOR2xp33_ASAP7_75t_SL U68213 ( .A(n71991), .B(n71990), .Y(n72233) );
  NAND2xp33_ASAP7_75t_SRAM U68214 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .B(
        n72502), .Y(n72441) );
  AOI211xp5_ASAP7_75t_SL U68215 ( .A1(n72417), .A2(n72493), .B(n72439), .C(
        n72438), .Y(n72449) );
  NOR2xp33_ASAP7_75t_SL U68216 ( .A(n59624), .B(n72436), .Y(n72438) );
  NOR2xp33_ASAP7_75t_SL U68217 ( .A(n72237), .B(n72236), .Y(n72336) );
  NOR2xp33_ASAP7_75t_SL U68218 ( .A(n72434), .B(n72220), .Y(n72478) );
  NOR4xp25_ASAP7_75t_SL U68219 ( .A(n72485), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_3_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .D(
        n71983), .Y(n71988) );
  AOI211xp5_ASAP7_75t_SL U68220 ( .A1(n72093), .A2(n72044), .B(n71981), .C(
        n71980), .Y(n71982) );
  AOI211xp5_ASAP7_75t_SL U68221 ( .A1(n73780), .A2(n73754), .B(n73701), .C(
        n73700), .Y(n73702) );
  NOR2xp33_ASAP7_75t_SL U68222 ( .A(n73684), .B(n73683), .Y(n73815) );
  NOR2xp33_ASAP7_75t_SL U68223 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .B(
        n73751), .Y(n73683) );
  AOI211xp5_ASAP7_75t_SL U68224 ( .A1(n73763), .A2(n73780), .B(n73707), .C(
        n73793), .Y(n73720) );
  NOR2xp33_ASAP7_75t_SL U68225 ( .A(n73706), .B(n59704), .Y(n73707) );
  AOI211xp5_ASAP7_75t_SL U68226 ( .A1(n72105), .A2(n71927), .B(n71767), .C(
        n71766), .Y(n71769) );
  NOR2xp33_ASAP7_75t_SL U68227 ( .A(n72067), .B(n71765), .Y(n71766) );
  AOI211xp5_ASAP7_75t_SL U68228 ( .A1(n58599), .A2(n72459), .B(n72458), .C(
        n72457), .Y(n72460) );
  NOR2xp33_ASAP7_75t_SL U68229 ( .A(n72499), .B(n72456), .Y(n72457) );
  AOI211xp5_ASAP7_75t_SL U68230 ( .A1(n73767), .A2(n59705), .B(n73793), .C(
        n73766), .Y(n73768) );
  NOR2xp33_ASAP7_75t_SL U68231 ( .A(n73635), .B(n73634), .Y(n73704) );
  AOI211xp5_ASAP7_75t_SL U68232 ( .A1(n72387), .A2(n72474), .B(n72386), .C(
        n72385), .Y(n72388) );
  NOR2xp33_ASAP7_75t_SL U68233 ( .A(n72415), .B(n72384), .Y(n72385) );
  NOR2xp33_ASAP7_75t_SL U68234 ( .A(n72355), .B(n72354), .Y(n72383) );
  NOR2xp33_ASAP7_75t_SL U68235 ( .A(n72340), .B(n72339), .Y(n72387) );
  NOR2xp33_ASAP7_75t_SL U68236 ( .A(n73667), .B(n59704), .Y(n73676) );
  AOI31xp33_ASAP7_75t_SL U68237 ( .A1(n73745), .A2(n73686), .A3(n73744), .B(
        n73666), .Y(n73677) );
  NOR2xp33_ASAP7_75t_SL U68238 ( .A(n3310), .B(n59704), .Y(n73629) );
  NOR2xp33_ASAP7_75t_SL U68239 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .B(
        n73698), .Y(n73663) );
  AOI31xp33_ASAP7_75t_SL U68240 ( .A1(n73730), .A2(n73686), .A3(n73729), .B(
        n73622), .Y(n73631) );
  NOR2xp33_ASAP7_75t_SL U68241 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[8]), .B(n59704), .Y(
        n73819) );
  NOR2xp33_ASAP7_75t_SL U68242 ( .A(n73714), .B(n73713), .Y(n73820) );
  NOR2xp33_ASAP7_75t_SL U68243 ( .A(n73710), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .Y(
        n73711) );
  NOR2xp33_ASAP7_75t_SL U68244 ( .A(n72268), .B(n72458), .Y(n72515) );
  NOR2xp33_ASAP7_75t_SL U68245 ( .A(n72267), .B(n72325), .Y(n72469) );
  NOR2xp33_ASAP7_75t_SL U68246 ( .A(n72265), .B(n72264), .Y(n72488) );
  NOR2xp33_ASAP7_75t_SL U68247 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_14_), 
        .B(n72517), .Y(n72349) );
  NOR2xp33_ASAP7_75t_SL U68248 ( .A(n59527), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_), 
        .Y(n72342) );
  NOR2xp33_ASAP7_75t_SL U68249 ( .A(n72495), .B(n58599), .Y(n72131) );
  NOR2xp33_ASAP7_75t_SL U68250 ( .A(n72190), .B(n72189), .Y(n72468) );
  NOR2xp33_ASAP7_75t_SL U68251 ( .A(n73823), .B(n59704), .Y(n73824) );
  NOR2xp33_ASAP7_75t_SL U68252 ( .A(n73758), .B(n73757), .Y(n73826) );
  NOR2xp33_ASAP7_75t_SL U68253 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[7]), .B(n59704), .Y(
        n73821) );
  AOI211xp5_ASAP7_75t_SL U68254 ( .A1(n72534), .A2(n72374), .B(n72373), .C(
        n72372), .Y(n72512) );
  NOR2xp33_ASAP7_75t_SL U68255 ( .A(n59622), .B(n72371), .Y(n72372) );
  NOR2xp33_ASAP7_75t_SL U68256 ( .A(n59623), .B(n72370), .Y(n72373) );
  AOI211xp5_ASAP7_75t_SL U68257 ( .A1(n72242), .A2(n72459), .B(n71920), .C(
        n72020), .Y(n71921) );
  AOI211xp5_ASAP7_75t_SL U68258 ( .A1(n72116), .A2(n72039), .B(n71917), .C(
        n71916), .Y(n72459) );
  NOR2xp33_ASAP7_75t_SL U68259 ( .A(n72085), .B(n72354), .Y(n71917) );
  NOR2xp33_ASAP7_75t_SL U68260 ( .A(n72298), .B(n72482), .Y(n72299) );
  NOR2xp33_ASAP7_75t_SL U68261 ( .A(n72316), .B(n57127), .Y(n72294) );
  NOR2xp33_ASAP7_75t_SL U68262 ( .A(n72308), .B(n57125), .Y(n72296) );
  NOR2xp33_ASAP7_75t_SL U68263 ( .A(n72292), .B(n72291), .Y(n72479) );
  AOI211xp5_ASAP7_75t_SL U68264 ( .A1(n72417), .A2(n72398), .B(n72024), .C(
        n72023), .Y(n72513) );
  NOR2xp33_ASAP7_75t_SL U68265 ( .A(n59623), .B(n72322), .Y(n72024) );
  AOI211xp5_ASAP7_75t_SL U68266 ( .A1(n72192), .A2(n57192), .B(n71939), .C(
        n72020), .Y(n71940) );
  NOR2xp33_ASAP7_75t_SL U68267 ( .A(n72207), .B(n72467), .Y(n71939) );
  NOR2xp33_ASAP7_75t_SL U68268 ( .A(n71761), .B(n71760), .Y(n71992) );
  NOR2xp33_ASAP7_75t_SL U68269 ( .A(n72119), .B(n72025), .Y(n71891) );
  NOR2xp33_ASAP7_75t_SL U68270 ( .A(n59624), .B(n72020), .Y(n71908) );
  NOR2xp33_ASAP7_75t_SL U68271 ( .A(n71829), .B(n71828), .Y(n71830) );
  AOI211xp5_ASAP7_75t_SL U68272 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .A2(
        n71856), .B(n71824), .C(n71823), .Y(n71979) );
  NOR2xp33_ASAP7_75t_SL U68273 ( .A(n72005), .B(n57208), .Y(n71823) );
  NOR2xp33_ASAP7_75t_SL U68274 ( .A(n71994), .B(n58422), .Y(n71824) );
  AOI211xp5_ASAP7_75t_SL U68275 ( .A1(n57192), .A2(n72329), .B(n72020), .C(
        n71959), .Y(n71960) );
  NOR2xp33_ASAP7_75t_SL U68276 ( .A(n71983), .B(n72330), .Y(n71959) );
  NOR2xp33_ASAP7_75t_SL U68277 ( .A(n71859), .B(n71858), .Y(n72009) );
  NAND2xp33_ASAP7_75t_SRAM U68278 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_36_), 
        .Y(n71822) );
  AOI211xp5_ASAP7_75t_SL U68279 ( .A1(n57192), .A2(n72471), .B(n72020), .C(
        n71976), .Y(n71977) );
  NOR2xp33_ASAP7_75t_SL U68280 ( .A(n72207), .B(n72210), .Y(n71976) );
  NOR2xp33_ASAP7_75t_SL U68281 ( .A(n72495), .B(n72325), .Y(n72331) );
  NOR2xp33_ASAP7_75t_SL U68282 ( .A(n71841), .B(n57192), .Y(n72325) );
  NOR2xp33_ASAP7_75t_SL U68283 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .Y(
        n71841) );
  AOI211xp5_ASAP7_75t_SL U68284 ( .A1(n72116), .A2(n72125), .B(n71963), .C(
        n71962), .Y(n71964) );
  NOR2xp33_ASAP7_75t_SL U68285 ( .A(n72085), .B(n72108), .Y(n71962) );
  NOR2xp33_ASAP7_75t_SL U68286 ( .A(n72355), .B(n72118), .Y(n71963) );
  AOI211xp5_ASAP7_75t_SL U68287 ( .A1(n72412), .A2(n72411), .B(n72410), .C(
        n72409), .Y(n72413) );
  AOI211xp5_ASAP7_75t_SL U68288 ( .A1(n72117), .A2(n72116), .B(n72115), .C(
        n72114), .Y(n72397) );
  NOR2xp33_ASAP7_75t_SL U68289 ( .A(n72355), .B(n72108), .Y(n72115) );
  NOR2xp33_ASAP7_75t_SL U68290 ( .A(n59622), .B(n72271), .Y(n72327) );
  NOR2xp33_ASAP7_75t_SL U68291 ( .A(n72004), .B(n72003), .Y(n72275) );
  NOR2xp33_ASAP7_75t_SL U68292 ( .A(n59622), .B(n72435), .Y(n72497) );
  NOR2xp33_ASAP7_75t_SL U68293 ( .A(n59705), .B(n73831), .Y(n73832) );
  NOR2xp33_ASAP7_75t_SL U68294 ( .A(n3337), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .Y(
        n73685) );
  AND2x2_ASAP7_75t_SL U68295 ( .A(n72499), .B(n57192), .Y(n72500) );
  NAND2xp33_ASAP7_75t_SRAM U68296 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_), 
        .B(n72367), .Y(n72247) );
  AOI31xp33_ASAP7_75t_SL U68297 ( .A1(n72324), .A2(n72474), .A3(n72323), .B(
        n72171), .Y(n72174) );
  NOR2xp33_ASAP7_75t_SL U68298 ( .A(n72147), .B(n72118), .Y(n72169) );
  NOR2xp33_ASAP7_75t_SL U68299 ( .A(n72310), .B(n57208), .Y(n71884) );
  NOR2xp33_ASAP7_75t_SL U68300 ( .A(n72351), .B(n71890), .Y(n71887) );
  NOR2xp33_ASAP7_75t_SL U68301 ( .A(n71872), .B(n71871), .Y(n72113) );
  NOR2xp33_ASAP7_75t_SL U68302 ( .A(n59624), .B(n72271), .Y(n72445) );
  NOR2xp33_ASAP7_75t_SL U68303 ( .A(n71852), .B(n71851), .Y(n72158) );
  NAND2xp33_ASAP7_75t_SRAM U68304 ( .A(n72286), .B(n72091), .Y(n71843) );
  NOR2xp33_ASAP7_75t_SL U68305 ( .A(n72284), .B(n72283), .Y(n72289) );
  NOR2xp33_ASAP7_75t_SL U68306 ( .A(n72355), .B(n72059), .Y(n72281) );
  NOR2xp33_ASAP7_75t_SL U68307 ( .A(n59622), .B(n72465), .Y(n72279) );
  NOR2xp33_ASAP7_75t_SL U68308 ( .A(n72244), .B(n72243), .Y(n72466) );
  OR2x2_ASAP7_75t_SL U68309 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .Y(
        n72495) );
  NOR2xp33_ASAP7_75t_SL U68310 ( .A(n71950), .B(n57127), .Y(n72224) );
  NOR2xp33_ASAP7_75t_SL U68311 ( .A(n71821), .B(n71820), .Y(n72137) );
  NOR2xp33_ASAP7_75t_SL U68312 ( .A(n71810), .B(n71809), .Y(n72046) );
  NAND2xp33_ASAP7_75t_SRAM U68313 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_24_), 
        .Y(n71807) );
  NOR2xp33_ASAP7_75t_SL U68314 ( .A(n72136), .B(n72135), .Y(n72303) );
  NOR2xp33_ASAP7_75t_SL U68315 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .B(
        n72006), .Y(n71985) );
  NOR2xp33_ASAP7_75t_SL U68316 ( .A(n72035), .B(n72034), .Y(n72220) );
  NAND2xp33_ASAP7_75t_SRAM U68317 ( .A(n59527), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_), 
        .Y(n72033) );
  NOR2xp33_ASAP7_75t_SL U68318 ( .A(n72134), .B(n72133), .Y(n72337) );
  AOI211xp5_ASAP7_75t_SL U68319 ( .A1(n59625), .A2(n72493), .B(n72257), .C(
        n72256), .Y(n72391) );
  NOR2xp33_ASAP7_75t_SL U68320 ( .A(n72156), .B(n72155), .Y(n72271) );
  NOR2xp33_ASAP7_75t_SL U68321 ( .A(n72199), .B(n72198), .Y(n72435) );
  NOR2xp33_ASAP7_75t_SL U68322 ( .A(n59527), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_), 
        .Y(n72196) );
  NOR2xp33_ASAP7_75t_SL U68323 ( .A(n59622), .B(n72432), .Y(n72257) );
  NOR2xp33_ASAP7_75t_SL U68324 ( .A(n72255), .B(n72254), .Y(n72432) );
  NOR2xp33_ASAP7_75t_SL U68325 ( .A(n59527), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_), 
        .Y(n72293) );
  NOR2xp33_ASAP7_75t_SL U68326 ( .A(n72089), .B(n72088), .Y(n72392) );
  NOR2xp33_ASAP7_75t_SL U68327 ( .A(n71846), .B(n71845), .Y(n72086) );
  NOR2xp33_ASAP7_75t_SL U68328 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_), 
        .Y(n71883) );
  NOR2xp33_ASAP7_75t_SL U68329 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_14_), 
        .B(n71894), .Y(n71882) );
  NOR2xp33_ASAP7_75t_SL U68330 ( .A(n71838), .B(n71837), .Y(n72083) );
  NOR2xp33_ASAP7_75t_SL U68331 ( .A(n72008), .B(n72007), .Y(n72200) );
  NOR2xp33_ASAP7_75t_SL U68332 ( .A(n72367), .B(n72006), .Y(n72007) );
  NOR2xp33_ASAP7_75t_SL U68333 ( .A(n71955), .B(n71954), .Y(n72153) );
  NOR2xp33_ASAP7_75t_SL U68334 ( .A(n71950), .B(n57125), .Y(n71937) );
  NOR2xp33_ASAP7_75t_SL U68335 ( .A(n71780), .B(n71779), .Y(n72064) );
  AOI31xp33_ASAP7_75t_SL U68336 ( .A1(n71778), .A2(n71890), .A3(n71777), .B(
        n71874), .Y(n71779) );
  NOR2xp33_ASAP7_75t_SL U68337 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_), 
        .B(n71899), .Y(n71874) );
  NAND2xp33_ASAP7_75t_SRAM U68338 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .Y(n71777) );
  NOR2xp33_ASAP7_75t_SL U68339 ( .A(n72351), .B(n57208), .Y(n71780) );
  NAND2xp33_ASAP7_75t_SRAM U68340 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_), 
        .Y(n71770) );
  AOI211xp5_ASAP7_75t_SL U68341 ( .A1(n72072), .A2(n72286), .B(n71758), .C(
        n71757), .Y(n72149) );
  NOR2xp33_ASAP7_75t_SL U68342 ( .A(n71755), .B(n71754), .Y(n72068) );
  NOR2xp33_ASAP7_75t_SL U68343 ( .A(n72112), .B(n72059), .Y(n71758) );
  NOR2xp33_ASAP7_75t_SL U68344 ( .A(n71752), .B(n71751), .Y(n72059) );
  OR2x2_ASAP7_75t_SL U68345 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .B(
        n71894), .Y(n58608) );
  NOR2xp33_ASAP7_75t_SL U68346 ( .A(n72143), .B(n72142), .Y(n72245) );
  NOR2xp33_ASAP7_75t_SL U68347 ( .A(n71953), .B(n57125), .Y(n71932) );
  NOR2xp33_ASAP7_75t_SL U68348 ( .A(n72056), .B(n72055), .Y(n72235) );
  NOR2xp33_ASAP7_75t_SL U68349 ( .A(n73742), .B(n73741), .Y(n73825) );
  NOR2xp33_ASAP7_75t_SL U68350 ( .A(n73668), .B(n58619), .Y(n73736) );
  NOR2xp33_ASAP7_75t_SL U68351 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[4]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .Y(
        n73619) );
  NOR2xp33_ASAP7_75t_SL U68352 ( .A(n73727), .B(n73726), .Y(n73822) );
  AOI31xp33_ASAP7_75t_SL U68353 ( .A1(n59632), .A2(n73752), .A3(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[3]), .B(n59705), .Y(
        n73724) );
  NOR2xp33_ASAP7_75t_SL U68354 ( .A(n73752), .B(n73722), .Y(n73723) );
  OR2x2_ASAP7_75t_SL U68355 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[0]), .B(
        n73617), .Y(n58400) );
  OR2x2_ASAP7_75t_SL U68356 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[1]), .B(
        n73641), .Y(n58619) );
  OR2x2_ASAP7_75t_SL U68357 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[1]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[0]), .Y(
        n58423) );
  AOI211xp5_ASAP7_75t_SL U68358 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[0]), .A2(
        n70311), .B(n70221), .C(n70242), .Y(n3162) );
  NOR2xp33_ASAP7_75t_SL U68359 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[5]), .B(
        n70234), .Y(n70224) );
  NOR2xp33_ASAP7_75t_SL U68360 ( .A(n70220), .B(n70219), .Y(n70576) );
  NOR2xp33_ASAP7_75t_SL U68361 ( .A(n70218), .B(n70237), .Y(n70220) );
  NOR2xp33_ASAP7_75t_SL U68362 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[3]), .B(
        n70241), .Y(n70240) );
  NOR2xp33_ASAP7_75t_SL U68363 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[1]), .B(
        n70221), .Y(n70222) );
  NOR2xp33_ASAP7_75t_SL U68364 ( .A(n70217), .B(n70216), .Y(n70232) );
  NOR2xp33_ASAP7_75t_SL U68365 ( .A(n70215), .B(n70214), .Y(n70217) );
  NOR2xp33_ASAP7_75t_SL U68366 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[5]), .B(
        n70233), .Y(n70214) );
  NOR2xp33_ASAP7_75t_SL U68367 ( .A(n72268), .B(n72476), .Y(n72486) );
  NOR2xp33_ASAP7_75t_SL U68368 ( .A(n72241), .B(n57192), .Y(n72268) );
  OR2x2_ASAP7_75t_SL U68369 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_0_), .Y(
        n58422) );
  NAND2xp33_ASAP7_75t_SRAM U68370 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .Y(n72366) );
  NOR2xp33_ASAP7_75t_SL U68371 ( .A(n72315), .B(n72314), .Y(n72509) );
  NOR2xp33_ASAP7_75t_SL U68372 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_13_), 
        .B(n72517), .Y(n72312) );
  NOR2xp33_ASAP7_75t_SL U68373 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_10_), 
        .B(n57123), .Y(n72505) );
  NAND2xp33_ASAP7_75t_SRAM U68374 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_), 
        .B(n58447), .Y(n72358) );
  NOR2xp33_ASAP7_75t_SL U68375 ( .A(n72357), .B(n72356), .Y(n72404) );
  NOR2xp33_ASAP7_75t_SL U68376 ( .A(n72166), .B(n72165), .Y(n72370) );
  NOR2xp33_ASAP7_75t_SL U68377 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .B(n72517), .Y(n71931) );
  NAND2xp33_ASAP7_75t_SRAM U68378 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_42_), 
        .B(n72364), .Y(n71970) );
  NOR2xp33_ASAP7_75t_SL U68379 ( .A(n74581), .B(n77287), .Y(n63769) );
  NOR2xp33_ASAP7_75t_SL U68380 ( .A(n75454), .B(n75766), .Y(n75616) );
  NAND2xp33_ASAP7_75t_SRAM U68381 ( .A(n75453), .B(n75452), .Y(n75454) );
  NOR4xp25_ASAP7_75t_SL U68382 ( .A(n65608), .B(n65607), .C(n65606), .D(n65605), .Y(n65610) );
  NOR2xp33_ASAP7_75t_SL U68383 ( .A(n66120), .B(n65595), .Y(n65596) );
  NOR2xp33_ASAP7_75t_SL U68384 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[8]), .B(n65663), .Y(
        n65581) );
  NAND2xp33_ASAP7_75t_SRAM U68385 ( .A(n75406), .B(n75405), .Y(n75409) );
  AOI211xp5_ASAP7_75t_SL U68386 ( .A1(n66167), .A2(n65536), .B(n65535), .C(
        n65577), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n3) );
  NOR4xp25_ASAP7_75t_SL U68387 ( .A(n65522), .B(n65521), .C(n65520), .D(n65519), .Y(n65536) );
  NAND2xp33_ASAP7_75t_SRAM U68388 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .B(n66146), 
        .Y(n65502) );
  AOI31xp33_ASAP7_75t_SL U68389 ( .A1(n66167), .A2(n66143), .A3(n66142), .B(
        n66141), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n5) );
  NAND2xp33_ASAP7_75t_SRAM U68390 ( .A(n74142), .B(n66135), .Y(n66140) );
  NOR2xp33_ASAP7_75t_SL U68391 ( .A(n66123), .B(n66122), .Y(n66133) );
  NAND2xp33_ASAP7_75t_SRAM U68392 ( .A(n59562), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .Y(n65510) );
  NAND2xp33_ASAP7_75t_SRAM U68393 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]), .B(n74206), 
        .Y(n65512) );
  AOI211xp5_ASAP7_75t_SL U68394 ( .A1(n66182), .A2(n65592), .B(n65591), .C(
        n65590), .Y(n66117) );
  NOR2xp33_ASAP7_75t_SL U68395 ( .A(n65832), .B(n65646), .Y(n65591) );
  NAND2xp33_ASAP7_75t_SRAM U68396 ( .A(n59562), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]), .Y(n65508) );
  NOR2xp33_ASAP7_75t_SL U68397 ( .A(n65580), .B(n65579), .Y(n66114) );
  NOR2xp33_ASAP7_75t_SL U68398 ( .A(n65805), .B(n65646), .Y(n65579) );
  NOR2xp33_ASAP7_75t_SL U68399 ( .A(n65578), .B(n66181), .Y(n65580) );
  AOI31xp33_ASAP7_75t_SL U68400 ( .A1(n66092), .A2(n65657), .A3(n65656), .B(
        n65655), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n2) );
  AOI211xp5_ASAP7_75t_SL U68401 ( .A1(n65650), .A2(n65649), .B(n65648), .C(
        n65647), .Y(n65657) );
  AOI211xp5_ASAP7_75t_SL U68402 ( .A1(n65642), .A2(n66148), .B(n65641), .C(
        n65640), .Y(n65648) );
  AOI211xp5_ASAP7_75t_SL U68403 ( .A1(n65634), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .B(n65633), 
        .C(n65632), .Y(n65636) );
  NAND2xp33_ASAP7_75t_SRAM U68404 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]), .B(n66146), 
        .Y(n65624) );
  NOR2xp33_ASAP7_75t_SL U68405 ( .A(n65615), .B(n65614), .Y(n66149) );
  NOR2xp33_ASAP7_75t_SL U68406 ( .A(n65530), .B(n76976), .Y(n65534) );
  NOR2xp33_ASAP7_75t_SL U68407 ( .A(n66185), .B(n66180), .Y(n66136) );
  NAND2xp33_ASAP7_75t_SRAM U68408 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]), .B(n74206), 
        .Y(n65567) );
  NOR2xp33_ASAP7_75t_SL U68409 ( .A(n65639), .B(n66150), .Y(n66116) );
  NAND2xp33_ASAP7_75t_SRAM U68410 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), .B(n66146), 
        .Y(n65573) );
  NAND2xp33_ASAP7_75t_SRAM U68411 ( .A(n59562), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[39]), .Y(n65571) );
  NOR2xp33_ASAP7_75t_SL U68412 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .B(n65639), .Y(
        n65517) );
  AOI211xp5_ASAP7_75t_SL U68413 ( .A1(n65670), .A2(n65566), .B(n65565), .C(
        n65564), .Y(n66097) );
  NOR2xp33_ASAP7_75t_SL U68414 ( .A(n66089), .B(n65646), .Y(n65564) );
  NOR2xp33_ASAP7_75t_SL U68415 ( .A(n65742), .B(n66181), .Y(n65565) );
  AOI211xp5_ASAP7_75t_SL U68416 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[25]), .A2(n66182), 
        .B(n65576), .C(n65575), .Y(n66094) );
  NOR2xp33_ASAP7_75t_SL U68417 ( .A(n65506), .B(n65674), .Y(n65601) );
  NOR2xp33_ASAP7_75t_SL U68418 ( .A(n74138), .B(n65674), .Y(n66152) );
  NOR2xp33_ASAP7_75t_SL U68419 ( .A(n65501), .B(n65667), .Y(n66092) );
  NOR2xp33_ASAP7_75t_SL U68420 ( .A(n1179), .B(n75397), .Y(n62212) );
  NOR2xp33_ASAP7_75t_SL U68421 ( .A(n1139), .B(n75645), .Y(n75394) );
  NOR2xp33_ASAP7_75t_SL U68422 ( .A(n62207), .B(n75648), .Y(n75397) );
  NOR2xp33_ASAP7_75t_SL U68423 ( .A(n1171), .B(n62224), .Y(n62226) );
  NOR2xp33_ASAP7_75t_SL U68424 ( .A(n75648), .B(n62228), .Y(n62224) );
  NOR2xp33_ASAP7_75t_SL U68425 ( .A(n1143), .B(n64180), .Y(n63917) );
  NOR2xp33_ASAP7_75t_SL U68426 ( .A(n75648), .B(n75396), .Y(n64180) );
  NOR2xp33_ASAP7_75t_SL U68427 ( .A(n66224), .B(n75645), .Y(n75396) );
  AOI31xp33_ASAP7_75t_SL U68428 ( .A1(n74487), .A2(n74488), .A3(n74486), .B(
        n74485), .Y(n74728) );
  NOR4xp25_ASAP7_75t_SL U68429 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_5_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_6_), .D(
        n74484), .Y(n74485) );
  NOR2xp33_ASAP7_75t_SL U68430 ( .A(n74481), .B(n74480), .Y(n74489) );
  NOR4xp25_ASAP7_75t_SL U68431 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_12_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_11_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_10_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_9_), .Y(
        n74477) );
  NOR4xp25_ASAP7_75t_SL U68432 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_16_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_15_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_14_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_13_), .Y(
        n74478) );
  NOR4xp25_ASAP7_75t_SL U68433 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_20_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_19_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_18_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_17_), .Y(
        n74479) );
  NOR4xp25_ASAP7_75t_SL U68434 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_3_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_2_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_1_), .Y(
        n74474) );
  NOR4xp25_ASAP7_75t_SL U68435 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_8_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_7_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_6_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_5_), .Y(
        n74475) );
  NOR4xp25_ASAP7_75t_SL U68436 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_3_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_4_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_0_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_1_), .Y(
        n74486) );
  NOR4xp25_ASAP7_75t_SL U68437 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_2_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_6_), .D(
        n74473), .Y(n74488) );
  NOR4xp25_ASAP7_75t_SL U68438 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_19_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_20_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_21_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_22_), .Y(
        n74470) );
  NOR4xp25_ASAP7_75t_SL U68439 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_15_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_16_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_17_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_18_), .Y(
        n74471) );
  NOR4xp25_ASAP7_75t_SL U68440 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_11_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_12_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_13_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_14_), .Y(
        n74472) );
  NOR4xp25_ASAP7_75t_SL U68441 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_7_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_8_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_9_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_10_), .Y(
        n74467) );
  NOR4xp25_ASAP7_75t_SL U68442 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_3_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_4_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opa_i_5_), .Y(
        n74468) );
  NOR4xp25_ASAP7_75t_SL U68443 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_5_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_6_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_7_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_2_), .Y(
        n74487) );
  NOR2xp33_ASAP7_75t_SL U68444 ( .A(n70686), .B(n59697), .Y(n70694) );
  NOR2xp33_ASAP7_75t_SL U68445 ( .A(n72563), .B(n72562), .Y(n74099) );
  NOR2xp33_ASAP7_75t_SL U68446 ( .A(n72579), .B(n74098), .Y(n72563) );
  NOR4xp25_ASAP7_75t_SL U68447 ( .A(n74252), .B(n74264), .C(n72587), .D(n72586), .Y(n72593) );
  NOR2xp33_ASAP7_75t_SL U68448 ( .A(n72585), .B(n74234), .Y(n74252) );
  NOR2xp33_ASAP7_75t_SL U68449 ( .A(n72584), .B(n74235), .Y(n74234) );
  NOR2xp33_ASAP7_75t_SL U68450 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_5_), .B(
        n72583), .Y(n74232) );
  NOR2xp33_ASAP7_75t_SL U68451 ( .A(n72579), .B(n72578), .Y(n72577) );
  NOR2xp33_ASAP7_75t_SL U68452 ( .A(n74491), .B(n74490), .Y(n74730) );
  NOR2xp33_ASAP7_75t_SL U68453 ( .A(n72575), .B(n72574), .Y(n74490) );
  NOR2xp33_ASAP7_75t_SL U68454 ( .A(n72572), .B(n72571), .Y(n72573) );
  NOR2xp33_ASAP7_75t_SL U68455 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_1_), .Y(
        n72566) );
  NOR2xp33_ASAP7_75t_SL U68456 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_3_), .Y(
        n72567) );
  NOR2xp33_ASAP7_75t_SL U68457 ( .A(n77932), .B(n78177), .Y(n77933) );
  NOR2xp33_ASAP7_75t_SL U68458 ( .A(n66078), .B(n66077), .Y(n66082) );
  NOR2xp33_ASAP7_75t_SL U68459 ( .A(n65480), .B(n65561), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n59) );
  AOI211xp5_ASAP7_75t_SL U68460 ( .A1(n65476), .A2(n65475), .B(n65474), .C(
        n65473), .Y(n65477) );
  NAND2xp33_ASAP7_75t_SRAM U68461 ( .A(n65449), .B(n65448), .Y(n65472) );
  NOR2xp33_ASAP7_75t_SL U68462 ( .A(n65446), .B(n65537), .Y(n65475) );
  NOR2xp33_ASAP7_75t_SL U68463 ( .A(n3086), .B(n78163), .Y(n77480) );
  NOR2xp33_ASAP7_75t_SL U68464 ( .A(n65561), .B(n65560), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n61) );
  NOR2xp33_ASAP7_75t_SL U68465 ( .A(n65743), .B(n65546), .Y(n65547) );
  AOI211xp5_ASAP7_75t_SL U68466 ( .A1(n70083), .A2(n69956), .B(n69955), .C(
        n69954), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[18]) );
  AOI31xp33_ASAP7_75t_SL U68467 ( .A1(n71609), .A2(n72164), .A3(n71586), .B(
        n71585), .Y(n71595) );
  NOR2xp33_ASAP7_75t_SL U68468 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_), 
        .B(n71579), .Y(n71598) );
  AOI211xp5_ASAP7_75t_SL U68469 ( .A1(n71574), .A2(n71573), .B(n71572), .C(
        n71571), .Y(n71575) );
  NOR2xp33_ASAP7_75t_SL U68470 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_1_), 
        .B(n71604), .Y(n71559) );
  NOR2xp33_ASAP7_75t_SL U68471 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .B(n71601), .Y(n71578) );
  AOI211xp5_ASAP7_75t_SL U68472 ( .A1(n70124), .A2(n78329), .B(n69899), .C(
        n70057), .Y(n69725) );
  AOI211xp5_ASAP7_75t_SL U68473 ( .A1(n70149), .A2(n69947), .B(n69946), .C(
        n69945), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[44]) );
  NOR2xp33_ASAP7_75t_SL U68474 ( .A(n69941), .B(n69940), .Y(n69946) );
  NOR2xp33_ASAP7_75t_SL U68475 ( .A(n70078), .B(n69808), .Y(n69810) );
  NOR2xp33_ASAP7_75t_SL U68476 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[1]), .B(n65443), .Y(
        n65662) );
  AOI211xp5_ASAP7_75t_SL U68477 ( .A1(n70083), .A2(n70067), .B(n70066), .C(
        n70065), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[22]) );
  AOI211xp5_ASAP7_75t_SL U68478 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[14]), .B(n69871), .C(n69870), .Y(n70061) );
  NOR2xp33_ASAP7_75t_SL U68479 ( .A(n78428), .B(n69925), .Y(n69870) );
  AOI211xp5_ASAP7_75t_SL U68480 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[18]), .B(n69951), .C(n69950), .Y(n70063) );
  NAND2xp33_ASAP7_75t_SRAM U68481 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]), .B(n70104), .Y(n69949) );
  NOR2xp33_ASAP7_75t_SL U68482 ( .A(n78424), .B(n70054), .Y(n69951) );
  AOI211xp5_ASAP7_75t_SL U68483 ( .A1(n70057), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[19]), .B(n70056), .C(n70055), .Y(n70058) );
  NOR2xp33_ASAP7_75t_SL U68484 ( .A(n78366), .B(n70054), .Y(n70055) );
  AOI211xp5_ASAP7_75t_SL U68485 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[10]), .B(n69814), .C(n69813), .Y(n70059) );
  NOR2xp33_ASAP7_75t_SL U68486 ( .A(n78344), .B(n70054), .Y(n69813) );
  NOR2xp33_ASAP7_75t_SL U68487 ( .A(n69899), .B(n69815), .Y(n69769) );
  NOR2xp33_ASAP7_75t_SL U68488 ( .A(n65445), .B(n65444), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n58) );
  AOI31xp33_ASAP7_75t_SL U68489 ( .A1(n65476), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[11]), .A3(n65792), 
        .B(n65441), .Y(n65442) );
  NOR2xp33_ASAP7_75t_SL U68490 ( .A(n65433), .B(n65432), .Y(n65558) );
  NOR2xp33_ASAP7_75t_SL U68491 ( .A(n65430), .B(n65545), .Y(n65433) );
  NOR4xp25_ASAP7_75t_SL U68492 ( .A(n65445), .B(n65561), .C(n65429), .D(n65428), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n60) );
  NOR2xp33_ASAP7_75t_SL U68493 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]), .B(n65466), 
        .Y(n65434) );
  NAND2xp33_ASAP7_75t_SRAM U68494 ( .A(n65462), .B(n65419), .Y(n65546) );
  NOR2xp33_ASAP7_75t_SL U68495 ( .A(n65418), .B(n65478), .Y(n65429) );
  NOR2xp33_ASAP7_75t_SL U68496 ( .A(n65414), .B(n65461), .Y(n65415) );
  NOR2xp33_ASAP7_75t_SL U68497 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[3]), .B(n66192), .Y(
        n65417) );
  AOI211xp5_ASAP7_75t_SL U68498 ( .A1(n65423), .A2(n65412), .B(n65411), .C(
        n65473), .Y(n65413) );
  NOR2xp33_ASAP7_75t_SL U68499 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[27]), .Y(n65381) );
  NOR2xp33_ASAP7_75t_SL U68500 ( .A(n69902), .B(n70135), .Y(n69798) );
  NOR2xp33_ASAP7_75t_SL U68501 ( .A(n78368), .B(n70054), .Y(n70036) );
  AOI211xp5_ASAP7_75t_SL U68502 ( .A1(n70083), .A2(n70001), .B(n70000), .C(
        n69999), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[20]) );
  AOI211xp5_ASAP7_75t_SL U68503 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[12]), .B(n69844), .C(n69843), .Y(n69997) );
  NOR2xp33_ASAP7_75t_SL U68504 ( .A(n78346), .B(n70054), .Y(n69843) );
  AOI211xp5_ASAP7_75t_SL U68505 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[20]), .B(n69994), .C(n69993), .Y(n69995) );
  NOR2xp33_ASAP7_75t_SL U68506 ( .A(n78356), .B(n70054), .Y(n69993) );
  AOI211xp5_ASAP7_75t_SL U68507 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[8]), .B(n69559), 
        .C(n69558), .Y(n69996) );
  NOR2xp33_ASAP7_75t_SL U68508 ( .A(n78340), .B(n70054), .Y(n69558) );
  AOI211xp5_ASAP7_75t_SL U68509 ( .A1(n70031), .A2(n69932), .B(n69931), .C(
        n69930), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[17]) );
  NOR2xp33_ASAP7_75t_SL U68510 ( .A(n69952), .B(n70041), .Y(n69931) );
  AOI211xp5_ASAP7_75t_SL U68511 ( .A1(n71801), .A2(n71800), .B(n71799), .C(
        n71798), .Y(n71802) );
  NOR2xp33_ASAP7_75t_SL U68512 ( .A(n69578), .B(n69746), .Y(n69792) );
  NOR2xp33_ASAP7_75t_SL U68513 ( .A(n69495), .B(n69494), .Y(n69795) );
  NOR2xp33_ASAP7_75t_SL U68514 ( .A(n70078), .B(n70017), .Y(n69494) );
  NOR2xp33_ASAP7_75t_SL U68515 ( .A(n70118), .B(n69743), .Y(n69495) );
  AOI211xp5_ASAP7_75t_SL U68516 ( .A1(n66022), .A2(n65932), .B(n65899), .C(
        n65898), .Y(n65900) );
  NOR2xp33_ASAP7_75t_SL U68517 ( .A(n65890), .B(n65889), .Y(n65891) );
  AOI211xp5_ASAP7_75t_SL U68518 ( .A1(n69984), .A2(n69983), .B(n69982), .C(
        n69981), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[19]) );
  NOR2xp33_ASAP7_75t_SL U68519 ( .A(n78424), .B(n70104), .Y(n69974) );
  NOR2xp33_ASAP7_75t_SL U68520 ( .A(n70060), .B(n69971), .Y(n69982) );
  NOR2xp33_ASAP7_75t_SL U68521 ( .A(n69903), .B(n69902), .Y(n70031) );
  NOR2xp33_ASAP7_75t_SL U68522 ( .A(n69899), .B(n69898), .Y(n69984) );
  NOR2xp33_ASAP7_75t_SL U68523 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_14_), .B(n70114), .Y(
        n69463) );
  NAND2xp33_ASAP7_75t_SRAM U68524 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_13_), .B(n70112), .Y(
        n69466) );
  NOR2xp33_ASAP7_75t_SL U68525 ( .A(n78347), .B(n69564), .Y(n69457) );
  AOI211xp5_ASAP7_75t_SL U68526 ( .A1(n66024), .A2(n65932), .B(n65810), .C(
        n65809), .Y(n65811) );
  NOR2xp33_ASAP7_75t_SL U68527 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_30_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_30_), .Y(n78224) );
  NOR2xp33_ASAP7_75t_SL U68528 ( .A(n78345), .B(n70021), .Y(n69490) );
  NOR2xp33_ASAP7_75t_SL U68529 ( .A(n70135), .B(n69926), .Y(n69740) );
  NOR2xp33_ASAP7_75t_SL U68530 ( .A(n69899), .B(n69932), .Y(n69741) );
  NOR2xp33_ASAP7_75t_SL U68531 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_18_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_), 
        .Y(n71540) );
  AOI211xp5_ASAP7_75t_SL U68532 ( .A1(n65978), .A2(n65945), .B(n65874), .C(
        n65873), .Y(n65875) );
  AOI211xp5_ASAP7_75t_SL U68533 ( .A1(n65978), .A2(n65977), .B(n65976), .C(
        n65975), .Y(n65979) );
  AOI211xp5_ASAP7_75t_SL U68534 ( .A1(n69515), .A2(n70149), .B(n69454), .C(
        n69453), .Y(or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[48]) );
  NOR2xp33_ASAP7_75t_SL U68535 ( .A(n69941), .B(n69570), .Y(n69453) );
  AOI211xp5_ASAP7_75t_SL U68536 ( .A1(n78431), .A2(n70109), .B(n70114), .C(
        n69467), .Y(n69441) );
  NOR2xp33_ASAP7_75t_SL U68537 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_15_), .B(n70109), .Y(
        n69467) );
  NOR2xp33_ASAP7_75t_SL U68538 ( .A(n59703), .B(n4138), .Y(or1200_immu_top_N10) );
  AOI211xp5_ASAP7_75t_SL U68539 ( .A1(n70038), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[7]), .B(n69778), 
        .C(n69777), .Y(n69971) );
  NOR2xp33_ASAP7_75t_SL U68540 ( .A(n78338), .B(n70054), .Y(n69777) );
  NOR2xp33_ASAP7_75t_SL U68541 ( .A(n78350), .B(n70035), .Y(n69973) );
  NOR2xp33_ASAP7_75t_SL U68542 ( .A(n78337), .B(n69564), .Y(n69450) );
  NOR2xp33_ASAP7_75t_SL U68543 ( .A(n78352), .B(n69564), .Y(n69424) );
  NOR2xp33_ASAP7_75t_SL U68544 ( .A(n59703), .B(n4089), .Y(or1200_immu_top_N9)
         );
  AOI211xp5_ASAP7_75t_SL U68545 ( .A1(n66051), .A2(n65945), .B(n65944), .C(
        n65943), .Y(n65946) );
  NOR2xp33_ASAP7_75t_SL U68546 ( .A(n66002), .B(n66001), .Y(n66003) );
  NOR2xp33_ASAP7_75t_SL U68547 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_17_), .B(n65400), .Y(
        n65372) );
  NOR2xp33_ASAP7_75t_SL U68548 ( .A(n65371), .B(n65401), .Y(n65373) );
  AOI31xp33_ASAP7_75t_SL U68549 ( .A1(n71626), .A2(n71625), .A3(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_3_), 
        .B(n71624), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n132)
         );
  NOR2xp33_ASAP7_75t_SL U68550 ( .A(n71546), .B(n71634), .Y(n71612) );
  NOR2xp33_ASAP7_75t_SL U68551 ( .A(n71545), .B(n71569), .Y(n71634) );
  NOR2xp33_ASAP7_75t_SL U68552 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .B(n72350), .Y(n71617) );
  NOR2xp33_ASAP7_75t_SL U68553 ( .A(n59703), .B(n4134), .Y(or1200_immu_top_N14) );
  NOR2xp33_ASAP7_75t_SL U68554 ( .A(n66040), .B(n66039), .Y(n66073) );
  NOR2xp33_ASAP7_75t_SL U68555 ( .A(n65974), .B(n66075), .Y(n66045) );
  NOR2xp33_ASAP7_75t_SL U68556 ( .A(n66040), .B(n66036), .Y(n66071) );
  AOI211xp5_ASAP7_75t_SL U68557 ( .A1(n66022), .A2(n65954), .B(n65904), .C(
        n65903), .Y(n66083) );
  NOR2xp33_ASAP7_75t_SL U68558 ( .A(n65974), .B(n65962), .Y(n65904) );
  NOR2xp33_ASAP7_75t_SL U68559 ( .A(n65776), .B(n65775), .Y(n65901) );
  NOR2xp33_ASAP7_75t_SL U68560 ( .A(n66027), .B(n65953), .Y(n65895) );
  NOR2xp33_ASAP7_75t_SL U68561 ( .A(n59703), .B(n4136), .Y(or1200_immu_top_N12) );
  NOR2xp33_ASAP7_75t_SL U68562 ( .A(n65972), .B(n66000), .Y(n65860) );
  NOR2xp33_ASAP7_75t_SL U68563 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[35]), .B(n58418), 
        .Y(n65851) );
  NOR2xp33_ASAP7_75t_SL U68564 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[29]), .B(n65830), 
        .Y(n65829) );
  NOR2xp33_ASAP7_75t_SL U68565 ( .A(n70078), .B(n69567), .Y(n69568) );
  AOI211xp5_ASAP7_75t_SL U68566 ( .A1(n70019), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_1_), .B(n69566), .C(
        n69565), .Y(n69569) );
  NOR2xp33_ASAP7_75t_SL U68567 ( .A(n78433), .B(n69564), .Y(n69565) );
  NOR2xp33_ASAP7_75t_SL U68568 ( .A(n71515), .B(n71514), .Y(n71519) );
  NOR2xp33_ASAP7_75t_SL U68569 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_23_), .B(n78244), .Y(n71514)
         );
  NOR2xp33_ASAP7_75t_SL U68570 ( .A(n70118), .B(n69567), .Y(n69824) );
  NOR2xp33_ASAP7_75t_SL U68571 ( .A(n69480), .B(n69479), .Y(n69575) );
  NOR2xp33_ASAP7_75t_SL U68572 ( .A(n70114), .B(n69500), .Y(n69480) );
  NOR2xp33_ASAP7_75t_SL U68573 ( .A(n78431), .B(n70109), .Y(n69475) );
  AND2x2_ASAP7_75t_SL U68574 ( .A(n70112), .B(n69421), .Y(n70018) );
  NOR2xp33_ASAP7_75t_SL U68575 ( .A(n59703), .B(n4090), .Y(or1200_immu_top_N8)
         );
  NAND2xp33_ASAP7_75t_SRAM U68576 ( .A(n65745), .B(n65841), .Y(n65850) );
  NOR2xp33_ASAP7_75t_SL U68577 ( .A(n66049), .B(n66063), .Y(n65955) );
  NOR2xp33_ASAP7_75t_SL U68578 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[11]), .B(n65841), 
        .Y(n65819) );
  NOR2xp33_ASAP7_75t_SL U68579 ( .A(n66060), .B(n65753), .Y(n66028) );
  NAND2xp33_ASAP7_75t_SRAM U68580 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[23]), .B(n65808), 
        .Y(n65757) );
  NOR2xp33_ASAP7_75t_SL U68581 ( .A(n70247), .B(n70246), .Y(n70249) );
  NOR2xp33_ASAP7_75t_SL U68582 ( .A(n69384), .B(n69383), .Y(n70246) );
  NOR2xp33_ASAP7_75t_SL U68583 ( .A(n69382), .B(n69381), .Y(n69384) );
  NOR2xp33_ASAP7_75t_SL U68584 ( .A(n72808), .B(n72847), .Y(n72700) );
  NOR2xp33_ASAP7_75t_SL U68585 ( .A(n59703), .B(n4135), .Y(or1200_immu_top_N13) );
  NOR2xp33_ASAP7_75t_SL U68586 ( .A(n59703), .B(n4133), .Y(or1200_immu_top_N15) );
  NOR2xp33_ASAP7_75t_SL U68587 ( .A(n59703), .B(n4091), .Y(or1200_immu_top_N7)
         );
  NOR2xp33_ASAP7_75t_SL U68588 ( .A(n72962), .B(n72824), .Y(n72691) );
  NOR2xp33_ASAP7_75t_SL U68589 ( .A(n59703), .B(n4093), .Y(or1200_immu_top_N5)
         );
  NOR2xp33_ASAP7_75t_SL U68590 ( .A(n69380), .B(n69381), .Y(n69383) );
  NAND2xp33_ASAP7_75t_SRAM U68591 ( .A(n65711), .B(n65808), .Y(n65849) );
  NAND2xp33_ASAP7_75t_SRAM U68592 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[39]), .B(n65841), 
        .Y(n65705) );
  AOI211xp5_ASAP7_75t_SL U68593 ( .A1(n57193), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[15]), .B(n57188), 
        .C(n65701), .Y(n65703) );
  NAND2xp33_ASAP7_75t_SRAM U68594 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[13]), .B(n65830), 
        .Y(n65781) );
  NOR2xp33_ASAP7_75t_SL U68595 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[12]), .B(n65828), 
        .Y(n65818) );
  NOR2xp33_ASAP7_75t_SL U68596 ( .A(n74142), .B(n76976), .Y(n65690) );
  NAND2xp33_ASAP7_75t_SRAM U68597 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[24]), .B(n65808), 
        .Y(n65686) );
  NAND2xp33_ASAP7_75t_SRAM U68598 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[30]), .B(n65808), 
        .Y(n65682) );
  NOR2xp33_ASAP7_75t_SL U68599 ( .A(n66179), .B(n76976), .Y(n65675) );
  NOR2xp33_ASAP7_75t_SL U68600 ( .A(n74147), .B(n76976), .Y(n65665) );
  AOI31xp33_ASAP7_75t_SL U68601 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_3_), .A2(
        n74919), .A3(n74918), .B(n74917), .Y(n74923) );
  NOR2xp33_ASAP7_75t_SL U68602 ( .A(n59703), .B(n4092), .Y(or1200_immu_top_N6)
         );
  NOR2xp33_ASAP7_75t_SL U68603 ( .A(n71789), .B(n71788), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n106) );
  NOR2xp33_ASAP7_75t_SL U68604 ( .A(or1200_cpu_or1200_fpu_a_is_qnan), .B(
        or1200_cpu_or1200_fpu_b_is_qnan), .Y(n74810) );
  NOR2xp33_ASAP7_75t_SL U68605 ( .A(n74755), .B(n74808), .Y(n74921) );
  NAND2xp33_ASAP7_75t_SRAM U68606 ( .A(n74803), .B(n74802), .Y(n74804) );
  NOR2xp33_ASAP7_75t_SL U68607 ( .A(n74894), .B(n76978), .Y(n74805) );
  NOR4xp25_ASAP7_75t_SL U68608 ( .A(n75890), .B(n57215), .C(n59530), .D(n59573), .Y(n74801) );
  NOR2xp33_ASAP7_75t_SL U68609 ( .A(n77625), .B(n77624), .Y(n77629) );
  NOR2xp33_ASAP7_75t_SL U68610 ( .A(n77773), .B(n77415), .Y(n78265) );
  NOR2xp33_ASAP7_75t_SL U68611 ( .A(n59892), .B(n77762), .Y(n77412) );
  NAND2xp33_ASAP7_75t_SRAM U68612 ( .A(n78368), .B(n59629), .Y(n72708) );
  NOR2xp33_ASAP7_75t_SL U68613 ( .A(n72962), .B(n72839), .Y(n72709) );
  NOR2xp33_ASAP7_75t_SL U68614 ( .A(n77999), .B(n61294), .Y(n59890) );
  NOR2xp33_ASAP7_75t_SL U68615 ( .A(n72990), .B(n72986), .Y(n72988) );
  NAND2xp33_ASAP7_75t_SRAM U68616 ( .A(n72719), .B(n73047), .Y(n72721) );
  NOR2xp33_ASAP7_75t_SL U68617 ( .A(n77607), .B(n77606), .Y(n749) );
  NOR2xp33_ASAP7_75t_SL U68618 ( .A(n77645), .B(n77605), .Y(n77606) );
  AOI31xp33_ASAP7_75t_SL U68619 ( .A1(n72840), .A2(n72839), .A3(n72976), .B(
        n72838), .Y(n72842) );
  NOR2xp33_ASAP7_75t_SL U68620 ( .A(n27477), .B(n70344), .Y(n70343) );
  NOR2xp33_ASAP7_75t_SL U68621 ( .A(n70376), .B(n70419), .Y(n70344) );
  NOR2xp33_ASAP7_75t_SL U68622 ( .A(n27472), .B(n70421), .Y(n70420) );
  NOR2xp33_ASAP7_75t_SL U68623 ( .A(n70478), .B(n70419), .Y(n70421) );
  AOI211xp5_ASAP7_75t_SL U68624 ( .A1(n73007), .A2(n72971), .B(n72963), .C(
        n72823), .Y(n72826) );
  NOR2xp33_ASAP7_75t_SL U68625 ( .A(n73002), .B(n72975), .Y(n72823) );
  NAND2xp33_ASAP7_75t_SRAM U68626 ( .A(n78427), .B(n59629), .Y(n72725) );
  NOR2xp33_ASAP7_75t_SL U68627 ( .A(n71726), .B(n71725), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n119) );
  NOR2xp33_ASAP7_75t_SL U68628 ( .A(n71724), .B(n71788), .Y(n71725) );
  AOI211xp5_ASAP7_75t_SL U68629 ( .A1(n71723), .A2(n71741), .B(n71722), .C(
        n71745), .Y(n71726) );
  NOR2xp33_ASAP7_75t_SL U68630 ( .A(n72879), .B(n73011), .Y(n72784) );
  NOR2xp33_ASAP7_75t_SL U68631 ( .A(n61301), .B(n61300), .Y(n61996) );
  NOR2xp33_ASAP7_75t_SL U68632 ( .A(n77483), .B(n61289), .Y(n61291) );
  NOR2xp33_ASAP7_75t_SL U68633 ( .A(n77469), .B(n61318), .Y(n61301) );
  NOR2xp33_ASAP7_75t_SL U68634 ( .A(n78163), .B(n77471), .Y(n77474) );
  NAND2xp33_ASAP7_75t_SRAM U68635 ( .A(n62204), .B(n61844), .Y(n61303) );
  AOI211xp5_ASAP7_75t_SL U68636 ( .A1(n71491), .A2(n71490), .B(n71489), .C(
        n71488), .Y(n71492) );
  AOI211xp5_ASAP7_75t_SL U68637 ( .A1(n71485), .A2(n71484), .B(n71483), .C(
        n71482), .Y(n71486) );
  NOR2xp33_ASAP7_75t_SL U68638 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_30_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_), 
        .Y(n71467) );
  AOI31xp33_ASAP7_75t_SL U68639 ( .A1(n71744), .A2(n71741), .A3(n71740), .B(
        n71739), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n118) );
  NOR2xp33_ASAP7_75t_SL U68640 ( .A(n71738), .B(n71788), .Y(n71739) );
  AND2x2_ASAP7_75t_SL U68641 ( .A(n77831), .B(n4152), .Y(n58609) );
  NAND2xp33_ASAP7_75t_SRAM U68642 ( .A(n63311), .B(n63310), .Y(n63312) );
  NAND2xp33_ASAP7_75t_SRAM U68643 ( .A(n59629), .B(n73022), .Y(n3338) );
  AOI211xp5_ASAP7_75t_SL U68644 ( .A1(n73021), .A2(n73020), .B(n73019), .C(
        n73018), .Y(n73022) );
  NOR2xp33_ASAP7_75t_SL U68645 ( .A(n73017), .B(n73016), .Y(n73018) );
  NOR2xp33_ASAP7_75t_SL U68646 ( .A(n72694), .B(n72963), .Y(n72695) );
  AOI211xp5_ASAP7_75t_SL U68647 ( .A1(n71747), .A2(n71786), .B(n71746), .C(
        n71745), .Y(n71748) );
  NOR2xp33_ASAP7_75t_SL U68648 ( .A(n73044), .B(n73043), .Y(n73046) );
  NOR2xp33_ASAP7_75t_SL U68649 ( .A(n73042), .B(n73041), .Y(n73043) );
  NOR2xp33_ASAP7_75t_SL U68650 ( .A(n72834), .B(n72833), .Y(n73036) );
  NOR2xp33_ASAP7_75t_SL U68651 ( .A(n72832), .B(n72872), .Y(n72833) );
  NOR2xp33_ASAP7_75t_SL U68652 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_0_), .B(
        n72920), .Y(n72872) );
  NOR2xp33_ASAP7_75t_SL U68653 ( .A(n70502), .B(n69805), .Y(n70516) );
  NOR2xp33_ASAP7_75t_SL U68654 ( .A(n70502), .B(n69736), .Y(n70508) );
  NOR2xp33_ASAP7_75t_SL U68655 ( .A(n70502), .B(n69887), .Y(n70517) );
  NOR2xp33_ASAP7_75t_SL U68656 ( .A(n70502), .B(n69866), .Y(n70495) );
  NOR2xp33_ASAP7_75t_SL U68657 ( .A(n70247), .B(n70481), .Y(n70231) );
  INVx1_ASAP7_75t_SL U68658 ( .A(n75649), .Y(n76890) );
  NOR2xp33_ASAP7_75t_SL U68659 ( .A(n72962), .B(n72978), .Y(n72750) );
  NOR2xp33_ASAP7_75t_SL U68660 ( .A(n71747), .B(n71786), .Y(n71746) );
  NOR2xp33_ASAP7_75t_SL U68661 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_0_), .B(
        n71684), .Y(n71747) );
  NOR2xp33_ASAP7_75t_SL U68662 ( .A(n71720), .B(n71794), .Y(n71798) );
  NOR2xp33_ASAP7_75t_SL U68663 ( .A(n71685), .B(n71791), .Y(n71687) );
  NOR2xp33_ASAP7_75t_SL U68664 ( .A(n71646), .B(n71683), .Y(n71787) );
  NOR2xp33_ASAP7_75t_SL U68665 ( .A(n71671), .B(n71655), .Y(n71683) );
  NOR2xp33_ASAP7_75t_SL U68666 ( .A(n71644), .B(n71657), .Y(n71685) );
  NOR2xp33_ASAP7_75t_SL U68667 ( .A(n71681), .B(n71650), .Y(n71731) );
  NOR2xp33_ASAP7_75t_SL U68668 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_3_), .B(
        n71691), .Y(n71650) );
  NOR2xp33_ASAP7_75t_SL U68669 ( .A(n71733), .B(n71700), .Y(n71681) );
  NOR2xp33_ASAP7_75t_SL U68670 ( .A(n71640), .B(n71639), .Y(n71707) );
  NOR2xp33_ASAP7_75t_SL U68671 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_4_), .B(
        n71695), .Y(n71640) );
  NOR2xp33_ASAP7_75t_SL U68672 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_7_), .B(
        n71673), .Y(n71676) );
  NOR2xp33_ASAP7_75t_SL U68673 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_0_), 
        .Y(n71671) );
  NOR2xp33_ASAP7_75t_SL U68674 ( .A(n71713), .B(n71668), .Y(n71712) );
  NOR2xp33_ASAP7_75t_SL U68675 ( .A(n71664), .B(n71694), .Y(n71666) );
  NOR2xp33_ASAP7_75t_SL U68676 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_4_), .B(
        n71659), .Y(n71660) );
  NOR2xp33_ASAP7_75t_SL U68677 ( .A(n71658), .B(n71657), .Y(n71702) );
  NOR2xp33_ASAP7_75t_SL U68678 ( .A(n71656), .B(n71655), .Y(n71658) );
  NAND2xp33_ASAP7_75t_SRAM U68679 ( .A(n77367), .B(n57160), .Y(n78054) );
  NOR2xp33_ASAP7_75t_SL U68680 ( .A(n72781), .B(n72780), .Y(n72846) );
  NOR2xp33_ASAP7_75t_SL U68681 ( .A(n72999), .B(n72727), .Y(n72813) );
  NOR2xp33_ASAP7_75t_SL U68682 ( .A(n72783), .B(n72782), .Y(n72814) );
  NOR2xp33_ASAP7_75t_SL U68683 ( .A(n72755), .B(n72754), .Y(n72792) );
  NOR2xp33_ASAP7_75t_SL U68684 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), .B(
        n72901), .Y(n72702) );
  NOR2xp33_ASAP7_75t_SL U68685 ( .A(n77659), .B(n77657), .Y(n77658) );
  NOR2xp33_ASAP7_75t_SL U68686 ( .A(n70502), .B(n69819), .Y(n70492) );
  NOR2xp33_ASAP7_75t_SL U68687 ( .A(n70502), .B(n69838), .Y(n70493) );
  NOR2xp33_ASAP7_75t_SL U68688 ( .A(n70502), .B(n69751), .Y(n70509) );
  NAND2xp33_ASAP7_75t_SRAM U68689 ( .A(n57081), .B(n69775), .Y(n70511) );
  NAND2xp33_ASAP7_75t_SRAM U68690 ( .A(n57081), .B(n69723), .Y(n70504) );
  NOR2xp33_ASAP7_75t_SL U68691 ( .A(n69722), .B(n69721), .Y(n69729) );
  NOR2xp33_ASAP7_75t_SL U68692 ( .A(n71458), .B(n71509), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n129) );
  AOI211xp5_ASAP7_75t_SL U68693 ( .A1(n71443), .A2(n71452), .B(n71442), .C(
        n71441), .Y(n71444) );
  NOR2xp33_ASAP7_75t_SL U68694 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_6_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_7_), 
        .Y(n71461) );
  NOR2xp33_ASAP7_75t_SL U68695 ( .A(n71510), .B(n71509), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n126) );
  AOI31xp33_ASAP7_75t_SL U68696 ( .A1(n71491), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .A3(n71581), .B(n71454), .Y(n71457) );
  NOR2xp33_ASAP7_75t_SL U68697 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_), 
        .B(n71591), .Y(n71435) );
  AOI31xp33_ASAP7_75t_SL U68698 ( .A1(n71452), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_), 
        .A3(n71995), .B(n71451), .Y(n71453) );
  NOR2xp33_ASAP7_75t_SL U68699 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_43_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_44_), 
        .Y(n71581) );
  AOI31xp33_ASAP7_75t_SL U68700 ( .A1(n71505), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_17_), 
        .A3(n72318), .B(n71504), .Y(n71507) );
  NAND2xp33_ASAP7_75t_SRAM U68701 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_37_), 
        .B(n72079), .Y(n71495) );
  AOI31xp33_ASAP7_75t_SL U68702 ( .A1(n69963), .A2(n69921), .A3(n59621), .B(
        n69920), .Y(n2281) );
  NOR2xp33_ASAP7_75t_SL U68703 ( .A(n70502), .B(n69917), .Y(n70497) );
  NOR2xp33_ASAP7_75t_SL U68704 ( .A(n70502), .B(n69853), .Y(n70494) );
  NOR2xp33_ASAP7_75t_SL U68705 ( .A(n69849), .B(n69861), .Y(n69852) );
  NOR2xp33_ASAP7_75t_SL U68706 ( .A(n77996), .B(n77766), .Y(n77487) );
  NOR2xp33_ASAP7_75t_SL U68707 ( .A(n69770), .B(n69790), .Y(n69784) );
  NOR2xp33_ASAP7_75t_SL U68708 ( .A(n2455), .B(n70376), .Y(n70384) );
  AOI31xp33_ASAP7_75t_SL U68709 ( .A1(n69969), .A2(n69939), .A3(n59621), .B(
        n69938), .Y(n2279) );
  NOR2xp33_ASAP7_75t_SL U68710 ( .A(n70502), .B(n69935), .Y(n70518) );
  NOR2xp33_ASAP7_75t_SL U68711 ( .A(n62484), .B(n62483), .Y(n62481) );
  NOR2xp33_ASAP7_75t_SL U68712 ( .A(n73009), .B(n72728), .Y(n72732) );
  NOR2xp33_ASAP7_75t_SL U68713 ( .A(n70502), .B(n69718), .Y(n70503) );
  NOR2xp33_ASAP7_75t_SL U68714 ( .A(n69758), .B(n69754), .Y(n69772) );
  NOR2xp33_ASAP7_75t_SL U68715 ( .A(n69749), .B(n69750), .Y(n69754) );
  NOR2xp33_ASAP7_75t_SL U68716 ( .A(n70502), .B(n69753), .Y(n70510) );
  NOR2xp33_ASAP7_75t_SL U68717 ( .A(n70502), .B(n69893), .Y(n70496) );
  NAND2xp33_ASAP7_75t_SRAM U68718 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_20_), .B(n65344), .Y(
        n65336) );
  NOR2xp33_ASAP7_75t_SL U68719 ( .A(n61994), .B(n61993), .Y(n59500) );
  NOR2xp33_ASAP7_75t_SL U68720 ( .A(n61994), .B(n61993), .Y(n78157) );
  NOR2xp33_ASAP7_75t_SL U68721 ( .A(n61994), .B(n61993), .Y(n59501) );
  OR2x2_ASAP7_75t_SL U68722 ( .A(n77767), .B(n77766), .Y(n58399) );
  NOR2xp33_ASAP7_75t_SL U68723 ( .A(n77999), .B(n77468), .Y(n61292) );
  NOR2xp33_ASAP7_75t_SL U68724 ( .A(n3111), .B(n61284), .Y(n61305) );
  NOR2xp33_ASAP7_75t_SL U68725 ( .A(n78165), .B(n61296), .Y(n77767) );
  NAND2xp33_ASAP7_75t_SRAM U68726 ( .A(or1200_dc_top_dirty), .B(n3092), .Y(
        n77769) );
  NOR2xp33_ASAP7_75t_SL U68727 ( .A(n70817), .B(n70818), .Y(n70807) );
  NAND2xp33_ASAP7_75t_SRAM U68728 ( .A(n1492), .B(n62027), .Y(n62028) );
  NOR2xp33_ASAP7_75t_SL U68729 ( .A(n62016), .B(n62015), .Y(n62017) );
  NOR2xp33_ASAP7_75t_SL U68730 ( .A(n2657), .B(n62007), .Y(n62032) );
  NOR2xp33_ASAP7_75t_SL U68731 ( .A(n70502), .B(n69965), .Y(n70519) );
  NOR2xp33_ASAP7_75t_SL U68732 ( .A(n69961), .B(n69959), .Y(n69968) );
  AOI31xp33_ASAP7_75t_SL U68733 ( .A1(n69992), .A2(n70013), .A3(n59621), .B(
        n69991), .Y(n2275) );
  NOR2xp33_ASAP7_75t_SL U68734 ( .A(n70502), .B(n69988), .Y(n70520) );
  AOI211xp5_ASAP7_75t_SL U68735 ( .A1(n59674), .A2(n63495), .B(n63494), .C(
        n63493), .Y(n63496) );
  NOR2xp33_ASAP7_75t_SL U68736 ( .A(n77019), .B(n68787), .Y(n63494) );
  NOR2xp33_ASAP7_75t_SL U68737 ( .A(n72970), .B(n72969), .Y(n72982) );
  AOI211xp5_ASAP7_75t_SL U68738 ( .A1(n72990), .A2(n72951), .B(n73024), .C(
        n72992), .Y(n72959) );
  NOR4xp25_ASAP7_75t_SL U68739 ( .A(n72939), .B(n72938), .C(n72937), .D(n72936), .Y(n72946) );
  NOR2xp33_ASAP7_75t_SL U68740 ( .A(n72916), .B(n72936), .Y(n72918) );
  NAND2xp33_ASAP7_75t_SRAM U68741 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[4]), .B(n73047), 
        .Y(n72831) );
  NAND2xp33_ASAP7_75t_SRAM U68742 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[3]), .B(n73047), 
        .Y(n72843) );
  NOR2xp33_ASAP7_75t_SL U68743 ( .A(n72938), .B(n72937), .Y(n72894) );
  NAND2xp33_ASAP7_75t_SRAM U68744 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[5]), .B(n73047), 
        .Y(n72820) );
  NOR2xp33_ASAP7_75t_SL U68745 ( .A(n78343), .B(n57190), .Y(n72773) );
  NOR2xp33_ASAP7_75t_SL U68746 ( .A(n72916), .B(n72893), .Y(n72934) );
  NAND2xp33_ASAP7_75t_SRAM U68747 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[12]), .B(n73047), .Y(n72752) );
  NOR2xp33_ASAP7_75t_SL U68748 ( .A(n72902), .B(n72889), .Y(n72930) );
  NOR2xp33_ASAP7_75t_SL U68749 ( .A(n72904), .B(n72901), .Y(n72929) );
  NAND2xp33_ASAP7_75t_SRAM U68750 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[17]), .B(n73047), .Y(n72710) );
  NOR2xp33_ASAP7_75t_SL U68751 ( .A(n72885), .B(n72966), .Y(n72887) );
  NOR2xp33_ASAP7_75t_SL U68752 ( .A(n68801), .B(n68800), .Y(n68802) );
  NOR2xp33_ASAP7_75t_SL U68753 ( .A(n63905), .B(n63904), .Y(n63906) );
  NOR2xp33_ASAP7_75t_SL U68754 ( .A(n64169), .B(n63894), .Y(n63897) );
  NOR2xp33_ASAP7_75t_SL U68755 ( .A(n63512), .B(n63515), .Y(n63510) );
  AOI211xp5_ASAP7_75t_SL U68756 ( .A1(n75015), .A2(n77885), .B(n63788), .C(
        n63787), .Y(n63789) );
  NOR2xp33_ASAP7_75t_SL U68757 ( .A(n64172), .B(n63786), .Y(n63903) );
  NOR2xp33_ASAP7_75t_SL U68758 ( .A(n64170), .B(n63785), .Y(n63898) );
  NOR2xp33_ASAP7_75t_SL U68759 ( .A(n64171), .B(n65099), .Y(n63785) );
  NOR2xp33_ASAP7_75t_SL U68760 ( .A(n63888), .B(n63893), .Y(n63770) );
  NOR2xp33_ASAP7_75t_SL U68761 ( .A(n64172), .B(n64170), .Y(n63773) );
  NOR2xp33_ASAP7_75t_SL U68762 ( .A(n65209), .B(n65230), .Y(n65219) );
  NOR2xp33_ASAP7_75t_SL U68763 ( .A(n63423), .B(n63425), .Y(n63417) );
  AOI211xp5_ASAP7_75t_SL U68764 ( .A1(n59674), .A2(n63359), .B(n63358), .C(
        n63357), .Y(n63360) );
  NOR2xp33_ASAP7_75t_SL U68765 ( .A(n77603), .B(n68787), .Y(n63358) );
  NOR2xp33_ASAP7_75t_SL U68766 ( .A(n63400), .B(n63395), .Y(n63356) );
  NOR2xp33_ASAP7_75t_SL U68767 ( .A(n65173), .B(n65130), .Y(n65148) );
  AOI211xp5_ASAP7_75t_SL U68768 ( .A1(n75015), .A2(n77977), .B(n63332), .C(
        n63331), .Y(n63333) );
  NOR2xp33_ASAP7_75t_SL U68769 ( .A(n63321), .B(n63397), .Y(n63328) );
  NOR2xp33_ASAP7_75t_SL U68770 ( .A(n62492), .B(n62491), .Y(n62489) );
  NOR2xp33_ASAP7_75t_SL U68771 ( .A(n75020), .B(n75023), .Y(n75021) );
  AOI211xp5_ASAP7_75t_SL U68772 ( .A1(n72665), .A2(n72664), .B(n72663), .C(
        n72667), .Y(n72666) );
  NOR2xp33_ASAP7_75t_SL U68773 ( .A(n78381), .B(n59626), .Y(n72612) );
  NOR2xp33_ASAP7_75t_SL U68774 ( .A(n78378), .B(n59626), .Y(n72613) );
  AOI211xp5_ASAP7_75t_SL U68775 ( .A1(n72614), .A2(n72619), .B(n72642), .C(
        n72667), .Y(n72615) );
  NOR2xp33_ASAP7_75t_SL U68776 ( .A(n72622), .B(n72667), .Y(n72623) );
  NOR2xp33_ASAP7_75t_SL U68777 ( .A(n78375), .B(n59626), .Y(n72618) );
  NOR2xp33_ASAP7_75t_SL U68778 ( .A(n78371), .B(n59626), .Y(n72627) );
  NOR2xp33_ASAP7_75t_SL U68779 ( .A(n72670), .B(n72669), .Y(n72676) );
  NOR2xp33_ASAP7_75t_SL U68780 ( .A(n72667), .B(n72655), .Y(n72656) );
  NOR2xp33_ASAP7_75t_SL U68781 ( .A(n72672), .B(n72671), .Y(n72673) );
  NOR2xp33_ASAP7_75t_SL U68782 ( .A(n70502), .B(n70011), .Y(n70521) );
  NAND2xp33_ASAP7_75t_SRAM U68783 ( .A(n77448), .B(n77447), .Y(n77453) );
  NOR2xp33_ASAP7_75t_SL U68784 ( .A(n77428), .B(n77459), .Y(n9468) );
  NOR2xp33_ASAP7_75t_SL U68785 ( .A(n63292), .B(n63345), .Y(n63294) );
  NOR2xp33_ASAP7_75t_SL U68786 ( .A(n70053), .B(n70052), .Y(n2271) );
  AOI211xp5_ASAP7_75t_SL U68787 ( .A1(n70051), .A2(n70050), .B(n58553), .C(
        n70070), .Y(n70052) );
  NAND2xp33_ASAP7_75t_SRAM U68788 ( .A(n57081), .B(n70044), .Y(n70522) );
  NOR2xp33_ASAP7_75t_SL U68789 ( .A(n1779), .B(n59680), .Y(n77203) );
  NOR2xp33_ASAP7_75t_SL U68790 ( .A(n69133), .B(n69132), .Y(n69134) );
  NOR2xp33_ASAP7_75t_SL U68791 ( .A(n69335), .B(n74797), .Y(n62069) );
  NOR4xp25_ASAP7_75t_SL U68792 ( .A(n77682), .B(n77681), .C(n77680), .D(n77679), .Y(n77684) );
  NOR4xp25_ASAP7_75t_SL U68793 ( .A(n57144), .B(n77678), .C(n77677), .D(n2966), 
        .Y(n77682) );
  NOR2xp33_ASAP7_75t_SL U68794 ( .A(n75611), .B(n57144), .Y(n75609) );
  NOR2xp33_ASAP7_75t_SL U68795 ( .A(n76673), .B(n61156), .Y(n76671) );
  NOR2xp33_ASAP7_75t_SL U68796 ( .A(n77436), .B(n77433), .Y(n77452) );
  NOR2xp33_ASAP7_75t_SL U68797 ( .A(n77432), .B(n77449), .Y(n77433) );
  NOR2xp33_ASAP7_75t_SL U68798 ( .A(or1200_cpu_or1200_except_n294), .B(n77432), 
        .Y(n77440) );
  AOI211xp5_ASAP7_75t_SL U68799 ( .A1(n70075), .A2(n70074), .B(n58553), .C(
        n70089), .Y(n70076) );
  NOR2xp33_ASAP7_75t_SL U68800 ( .A(n70502), .B(n70068), .Y(n70524) );
  NAND2xp33_ASAP7_75t_SRAM U68801 ( .A(n77278), .B(n57144), .Y(n77283) );
  NAND2xp33_ASAP7_75t_SRAM U68802 ( .A(n76874), .B(n57144), .Y(n76878) );
  NAND2xp33_ASAP7_75t_SRAM U68803 ( .A(n75456), .B(n57144), .Y(n75460) );
  NOR2xp33_ASAP7_75t_SL U68804 ( .A(n57144), .B(n77904), .Y(n76556) );
  NAND2xp33_ASAP7_75t_SRAM U68805 ( .A(n57082), .B(n59695), .Y(n61743) );
  NOR2xp33_ASAP7_75t_SL U68806 ( .A(n74718), .B(n74719), .Y(n74721) );
  NAND2xp33_ASAP7_75t_SRAM U68807 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_1_), .B(
        n74677), .Y(n74678) );
  NOR2xp33_ASAP7_75t_SL U68808 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_17_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_16_), .Y(
        n74689) );
  NOR2xp33_ASAP7_75t_SL U68809 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_20_), .Y(
        n74692) );
  NOR2xp33_ASAP7_75t_SL U68810 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_7_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_6_), .Y(
        n74696) );
  NOR2xp33_ASAP7_75t_SL U68811 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_8_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_9_), .Y(
        n74666) );
  NOR2xp33_ASAP7_75t_SL U68812 ( .A(n61132), .B(n68810), .Y(n77993) );
  NOR2xp33_ASAP7_75t_SL U68813 ( .A(n1938), .B(n76542), .Y(n76543) );
  NAND2xp33_ASAP7_75t_SRAM U68814 ( .A(n76990), .B(n75768), .Y(n75772) );
  NOR2xp33_ASAP7_75t_SL U68815 ( .A(n2785), .B(n75767), .Y(n76990) );
  NOR2xp33_ASAP7_75t_SL U68816 ( .A(n1983), .B(n76538), .Y(n77200) );
  NOR2xp33_ASAP7_75t_SL U68817 ( .A(n77994), .B(n62319), .Y(n62204) );
  NOR2xp33_ASAP7_75t_SL U68818 ( .A(n77033), .B(n68810), .Y(n62199) );
  NOR2xp33_ASAP7_75t_SL U68819 ( .A(n62179), .B(n62178), .Y(n62196) );
  NOR4xp25_ASAP7_75t_SL U68820 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_15_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_4_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_11_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_1_), .Y(n76939)
         );
  NOR4xp25_ASAP7_75t_SL U68821 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_8_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_7_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_12_), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_16_), .Y(n76937)
         );
  NOR2xp33_ASAP7_75t_SL U68822 ( .A(n68951), .B(n68971), .Y(n68969) );
  NOR2xp33_ASAP7_75t_SL U68823 ( .A(n69087), .B(n69195), .Y(n69092) );
  NOR2xp33_ASAP7_75t_SL U68824 ( .A(n69089), .B(n69073), .Y(n69077) );
  NOR2xp33_ASAP7_75t_SL U68825 ( .A(n69091), .B(n69072), .Y(n69073) );
  NOR2xp33_ASAP7_75t_SL U68826 ( .A(n69090), .B(n69106), .Y(n69075) );
  NAND2xp33_ASAP7_75t_SRAM U68827 ( .A(n75832), .B(n57144), .Y(n73957) );
  NOR2xp33_ASAP7_75t_SL U68828 ( .A(n77356), .B(n77454), .Y(n9455) );
  NOR2xp33_ASAP7_75t_SL U68829 ( .A(n70907), .B(n70965), .Y(n70891) );
  NAND2xp33_ASAP7_75t_SRAM U68830 ( .A(n74776), .B(n57144), .Y(n74077) );
  NOR2xp33_ASAP7_75t_SL U68831 ( .A(n74943), .B(n74942), .Y(n74946) );
  NOR2xp33_ASAP7_75t_SL U68832 ( .A(or1200_cpu_or1200_except_n290), .B(n77434), 
        .Y(n77430) );
  NAND2xp33_ASAP7_75t_SRAM U68833 ( .A(or1200_cpu_or1200_except_n288), .B(
        or1200_cpu_or1200_except_n294), .Y(n77434) );
  NOR2xp33_ASAP7_75t_SL U68834 ( .A(or1200_cpu_or1200_except_n292), .B(
        or1200_cpu_or1200_except_n286), .Y(n74933) );
  AOI211xp5_ASAP7_75t_SL U68835 ( .A1(n61643), .A2(n61367), .B(n61366), .C(
        n61365), .Y(n61368) );
  NOR2xp33_ASAP7_75t_SL U68836 ( .A(n75349), .B(n75574), .Y(n61365) );
  AOI211xp5_ASAP7_75t_SL U68837 ( .A1(n62348), .A2(n61358), .B(n75882), .C(
        n61763), .Y(n61359) );
  AOI211xp5_ASAP7_75t_SL U68838 ( .A1(n62371), .A2(n61357), .B(n62372), .C(
        n61356), .Y(n61361) );
  AOI211xp5_ASAP7_75t_SL U68839 ( .A1(n61494), .A2(n64219), .B(n61352), .C(
        n61351), .Y(n61362) );
  NAND2xp33_ASAP7_75t_SRAM U68840 ( .A(n62362), .B(n64225), .Y(n61350) );
  NOR2xp33_ASAP7_75t_SL U68841 ( .A(n1824), .B(n76717), .Y(n61326) );
  AOI211xp5_ASAP7_75t_SL U68842 ( .A1(n62292), .A2(n61663), .B(n61662), .C(
        n61661), .Y(n61664) );
  AOI211xp5_ASAP7_75t_SL U68843 ( .A1(n61658), .A2(n61785), .B(n61657), .C(
        n61656), .Y(n61659) );
  NOR2xp33_ASAP7_75t_SL U68844 ( .A(n61615), .B(n61614), .Y(n61617) );
  NOR2xp33_ASAP7_75t_SL U68845 ( .A(n1499), .B(n61755), .Y(n61607) );
  NOR2xp33_ASAP7_75t_SL U68846 ( .A(n1847), .B(n76717), .Y(n61605) );
  AOI211xp5_ASAP7_75t_SL U68847 ( .A1(n77125), .A2(n62388), .B(n62387), .C(
        n77122), .Y(n62389) );
  NOR2xp33_ASAP7_75t_SL U68848 ( .A(n62422), .B(n62377), .Y(n62378) );
  NAND2xp33_ASAP7_75t_SRAM U68849 ( .A(n62366), .B(n75845), .Y(n62368) );
  AOI211xp5_ASAP7_75t_SL U68850 ( .A1(n62345), .A2(n62344), .B(n62343), .C(
        n62342), .Y(n62386) );
  NOR2xp33_ASAP7_75t_SL U68851 ( .A(n75316), .B(n62341), .Y(n62342) );
  AOI211xp5_ASAP7_75t_SL U68852 ( .A1(n62425), .A2(n62338), .B(n62337), .C(
        n62336), .Y(n62339) );
  AOI211xp5_ASAP7_75t_SL U68853 ( .A1(n62326), .A2(n76735), .B(n62325), .C(
        n62324), .Y(n62328) );
  AOI211xp5_ASAP7_75t_SL U68854 ( .A1(n77041), .A2(n69002), .B(n62321), .C(
        n62320), .Y(n62322) );
  NOR2xp33_ASAP7_75t_SL U68855 ( .A(n1396), .B(n77035), .Y(n62321) );
  NOR2xp33_ASAP7_75t_SL U68856 ( .A(n73953), .B(n76296), .Y(n62297) );
  AOI211xp5_ASAP7_75t_SL U68857 ( .A1(n76748), .A2(n62290), .B(n76746), .C(
        n75882), .Y(n62291) );
  AOI211xp5_ASAP7_75t_SL U68858 ( .A1(n77125), .A2(n64315), .B(n62286), .C(
        n62285), .Y(n62294) );
  AOI211xp5_ASAP7_75t_SL U68859 ( .A1(n62274), .A2(n62273), .B(n62272), .C(
        n62271), .Y(n62281) );
  AOI211xp5_ASAP7_75t_SL U68860 ( .A1(n75727), .A2(n62268), .B(n62267), .C(
        n62266), .Y(n62269) );
  NOR2xp33_ASAP7_75t_SL U68861 ( .A(or1200_cpu_or1200_mult_mac_n153), .B(
        n75723), .Y(n62267) );
  NOR2xp33_ASAP7_75t_SL U68862 ( .A(n62259), .B(n62258), .Y(n62283) );
  NOR2xp33_ASAP7_75t_SL U68863 ( .A(n1963), .B(n76717), .Y(n62236) );
  NOR2xp33_ASAP7_75t_SL U68864 ( .A(n1402), .B(n76716), .Y(n62234) );
  OR2x2_ASAP7_75t_SL U68865 ( .A(n2596), .B(n62071), .Y(n74797) );
  AOI211xp5_ASAP7_75t_SL U68866 ( .A1(n77125), .A2(n74621), .B(n61558), .C(
        n61557), .Y(n61562) );
  AOI211xp5_ASAP7_75t_SL U68867 ( .A1(n61539), .A2(n61538), .B(n61537), .C(
        n61536), .Y(n61540) );
  AOI211xp5_ASAP7_75t_SL U68868 ( .A1(n76749), .A2(n61517), .B(n61516), .C(
        n61515), .Y(n61543) );
  AOI211xp5_ASAP7_75t_SL U68869 ( .A1(n62508), .A2(n76866), .B(n61482), .C(
        n64206), .Y(n61484) );
  AOI211xp5_ASAP7_75t_SL U68870 ( .A1(n77041), .A2(n68864), .B(n61473), .C(
        n61472), .Y(n61476) );
  NOR2xp33_ASAP7_75t_SL U68871 ( .A(n1976), .B(n76717), .Y(n61468) );
  NOR2xp33_ASAP7_75t_SL U68872 ( .A(n61467), .B(n61466), .Y(n61485) );
  NOR4xp25_ASAP7_75t_SL U68873 ( .A(n61458), .B(n61457), .C(n61456), .D(n61455), .Y(n61459) );
  AOI211xp5_ASAP7_75t_SL U68874 ( .A1(n61447), .A2(n61446), .B(n75882), .C(
        n61621), .Y(n61457) );
  AND4x1_ASAP7_75t_SL U68875 ( .A(n61542), .B(n61442), .C(n61441), .D(n61440), 
        .Y(n61443) );
  AOI31xp33_ASAP7_75t_SL U68876 ( .A1(n77060), .A2(n61438), .A3(n57214), .B(
        n61421), .Y(n61422) );
  NOR2xp33_ASAP7_75t_SL U68877 ( .A(n61415), .B(n61414), .Y(n61542) );
  NAND2xp33_ASAP7_75t_SRAM U68878 ( .A(n74776), .B(n64357), .Y(n58912) );
  AOI211xp5_ASAP7_75t_SL U68879 ( .A1(n77623), .A2(n61385), .B(n61384), .C(
        n61383), .Y(n61386) );
  NOR2xp33_ASAP7_75t_SL U68880 ( .A(or1200_cpu_or1200_mult_mac_n213), .B(
        n74587), .Y(n61384) );
  NOR2xp33_ASAP7_75t_SL U68881 ( .A(n76807), .B(n76806), .Y(n77910) );
  AOI211xp5_ASAP7_75t_SL U68882 ( .A1(n77117), .A2(n77087), .B(n76798), .C(
        n76797), .Y(n76799) );
  NOR2xp33_ASAP7_75t_SL U68883 ( .A(n76796), .B(n77604), .Y(n76797) );
  NOR2xp33_ASAP7_75t_SL U68884 ( .A(n62347), .B(n62346), .Y(n76747) );
  NOR2xp33_ASAP7_75t_SL U68885 ( .A(n76744), .B(n77605), .Y(n76807) );
  NOR4xp25_ASAP7_75t_SL U68886 ( .A(n76743), .B(n76742), .C(n76741), .D(n76740), .Y(n77605) );
  AOI211xp5_ASAP7_75t_SL U68887 ( .A1(n76735), .A2(n76734), .B(n76733), .C(
        n76732), .Y(n76738) );
  NOR2xp33_ASAP7_75t_SL U68888 ( .A(or1200_cpu_or1200_except_n270), .B(n76731), 
        .Y(n76732) );
  AOI211xp5_ASAP7_75t_SL U68889 ( .A1(n77623), .A2(n76727), .B(n76726), .C(
        n76725), .Y(n76728) );
  NOR2xp33_ASAP7_75t_SL U68890 ( .A(n1828), .B(n76717), .Y(n76718) );
  NOR2xp33_ASAP7_75t_SL U68891 ( .A(n76744), .B(n77590), .Y(n61262) );
  NOR4xp25_ASAP7_75t_SL U68892 ( .A(n61693), .B(n61261), .C(n61260), .D(n61259), .Y(n77590) );
  AOI211xp5_ASAP7_75t_SL U68893 ( .A1(n77090), .A2(
        or1200_cpu_or1200_fpu_result_conv[2]), .B(n58614), .C(n61230), .Y(
        n61231) );
  AOI211xp5_ASAP7_75t_SL U68894 ( .A1(n61229), .A2(n61228), .B(n75882), .C(
        n62288), .Y(n61230) );
  AOI211xp5_ASAP7_75t_SL U68895 ( .A1(n63282), .A2(n76753), .B(n61217), .C(
        n61216), .Y(n61218) );
  NOR2xp33_ASAP7_75t_SL U68896 ( .A(n75700), .B(n61498), .Y(n61630) );
  NAND2xp33_ASAP7_75t_SRAM U68897 ( .A(n62594), .B(n61209), .Y(n61210) );
  NAND2xp33_ASAP7_75t_SRAM U68898 ( .A(n62262), .B(n77076), .Y(n61194) );
  NOR2xp33_ASAP7_75t_SL U68899 ( .A(n59569), .B(n59712), .Y(n61185) );
  NOR2xp33_ASAP7_75t_SL U68900 ( .A(n59710), .B(n59542), .Y(n61186) );
  NOR2xp33_ASAP7_75t_SL U68901 ( .A(n76770), .B(n63583), .Y(n61189) );
  NAND2xp33_ASAP7_75t_SRAM U68902 ( .A(n59545), .B(n62595), .Y(n61209) );
  AOI211xp5_ASAP7_75t_SL U68903 ( .A1(or1200_cpu_rf_datab[26]), .A2(n57091), 
        .B(n77184), .C(n64867), .Y(n64868) );
  NAND2xp33_ASAP7_75t_SRAM U68904 ( .A(n64840), .B(n75717), .Y(n64841) );
  AOI211xp5_ASAP7_75t_SL U68905 ( .A1(n64821), .A2(
        or1200_cpu_or1200_mult_mac_n193), .B(n73907), .C(n64820), .Y(n64822)
         );
  AOI211xp5_ASAP7_75t_SL U68906 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[26]), 
        .B(n64816), .C(n64815), .Y(n64817) );
  NOR2xp33_ASAP7_75t_SL U68907 ( .A(or1200_cpu_or1200_except_n240), .B(n57170), 
        .Y(n64815) );
  AOI211xp5_ASAP7_75t_SL U68908 ( .A1(or1200_cpu_rf_datab[14]), .A2(n57091), 
        .B(n77028), .C(n77027), .Y(n77029) );
  NOR2xp33_ASAP7_75t_SL U68909 ( .A(n2199), .B(n59679), .Y(n77028) );
  NOR4xp25_ASAP7_75t_SL U68910 ( .A(n60867), .B(n60866), .C(n60865), .D(n60864), .Y(n60868) );
  NOR2xp33_ASAP7_75t_SL U68911 ( .A(n63577), .B(n77101), .Y(n60865) );
  AOI211xp5_ASAP7_75t_SL U68912 ( .A1(n77082), .A2(n60853), .B(n60852), .C(
        n60851), .Y(n60869) );
  NOR2xp33_ASAP7_75t_SL U68913 ( .A(n75316), .B(n64313), .Y(n60851) );
  AOI211xp5_ASAP7_75t_SL U68914 ( .A1(or1200_cpu_spr_dat_rf[14]), .A2(n59686), 
        .B(n60832), .C(n60831), .Y(n60836) );
  AOI211xp5_ASAP7_75t_SL U68915 ( .A1(n77040), .A2(n75144), .B(n60829), .C(
        n60828), .Y(n60830) );
  NOR2xp33_ASAP7_75t_SL U68916 ( .A(or1200_cpu_or1200_except_n516), .B(n76724), 
        .Y(n60828) );
  AOI211xp5_ASAP7_75t_SL U68917 ( .A1(n62274), .A2(n62374), .B(n60802), .C(
        n60801), .Y(n60887) );
  NOR2xp33_ASAP7_75t_SL U68918 ( .A(n59552), .B(n76775), .Y(n60793) );
  NAND2xp33_ASAP7_75t_SRAM U68919 ( .A(n59585), .B(n77060), .Y(n60795) );
  AOI211xp5_ASAP7_75t_SL U68920 ( .A1(or1200_cpu_rf_datab[27]), .A2(n57091), 
        .B(n77184), .C(n75803), .Y(n75804) );
  AOI211xp5_ASAP7_75t_SL U68921 ( .A1(n76768), .A2(n76763), .B(n73939), .C(
        n73938), .Y(n73940) );
  NOR2xp33_ASAP7_75t_SL U68922 ( .A(n64858), .B(n73937), .Y(n73945) );
  AOI31xp33_ASAP7_75t_SL U68923 ( .A1(n73937), .A2(n77112), .A3(n73936), .B(
        n73935), .Y(n73947) );
  AOI211xp5_ASAP7_75t_SL U68924 ( .A1(n75741), .A2(n75832), .B(n73929), .C(
        n73928), .Y(n73930) );
  AOI211xp5_ASAP7_75t_SL U68925 ( .A1(n75823), .A2(n75126), .B(n73909), .C(
        n73908), .Y(n73910) );
  NOR2xp33_ASAP7_75t_SL U68926 ( .A(or1200_cpu_or1200_mult_mac_n195), .B(
        n75819), .Y(n73908) );
  AOI211xp5_ASAP7_75t_SL U68927 ( .A1(or1200_cpu_rf_datab[15]), .A2(n57091), 
        .B(n77135), .C(n77134), .Y(n77136) );
  NOR2xp33_ASAP7_75t_SL U68928 ( .A(n2850), .B(n59679), .Y(n77134) );
  NOR2xp33_ASAP7_75t_SL U68929 ( .A(n77705), .B(n59688), .Y(n77132) );
  NOR2xp33_ASAP7_75t_SL U68930 ( .A(n2037), .B(n76557), .Y(n69345) );
  AOI211xp5_ASAP7_75t_SL U68931 ( .A1(n77125), .A2(n77124), .B(n77123), .C(
        n77122), .Y(n77126) );
  AOI211xp5_ASAP7_75t_SL U68932 ( .A1(n77088), .A2(n77087), .B(n77086), .C(
        n77085), .Y(n77121) );
  NAND2xp33_ASAP7_75t_SRAM U68933 ( .A(n77082), .B(n77081), .Y(n77083) );
  AOI211xp5_ASAP7_75t_SL U68934 ( .A1(n77062), .A2(n77061), .B(n77060), .C(
        n77059), .Y(n77072) );
  AOI211xp5_ASAP7_75t_SL U68935 ( .A1(n77039), .A2(n77038), .B(n77037), .C(
        n77036), .Y(n77046) );
  NOR2xp33_ASAP7_75t_SL U68936 ( .A(n1370), .B(n77035), .Y(n77036) );
  AOI211xp5_ASAP7_75t_SL U68937 ( .A1(or1200_cpu_rf_datab[19]), .A2(n57091), 
        .B(n77184), .C(n74636), .Y(n74637) );
  NOR2xp33_ASAP7_75t_SL U68938 ( .A(n74626), .B(n74625), .Y(n74631) );
  NOR2xp33_ASAP7_75t_SL U68939 ( .A(n74616), .B(n74615), .Y(n74617) );
  NOR4xp25_ASAP7_75t_SL U68940 ( .A(n74614), .B(n74613), .C(n74612), .D(n74611), .Y(n74618) );
  AOI211xp5_ASAP7_75t_SL U68941 ( .A1(n74603), .A2(n57214), .B(n74602), .C(
        n74601), .Y(n74604) );
  NOR2xp33_ASAP7_75t_SL U68942 ( .A(or1200_cpu_or1200_mult_mac_n325), .B(
        n75738), .Y(n74601) );
  AOI211xp5_ASAP7_75t_SL U68943 ( .A1(or1200_cpu_rf_datab[11]), .A2(n57091), 
        .B(n76560), .C(n76559), .Y(n76561) );
  NOR2xp33_ASAP7_75t_SL U68944 ( .A(n61709), .B(n61708), .Y(n61714) );
  NOR4xp25_ASAP7_75t_SL U68945 ( .A(n61496), .B(n61887), .C(n62105), .D(n61729), .Y(n76759) );
  NOR2xp33_ASAP7_75t_SL U68946 ( .A(n61694), .B(n61693), .Y(n61695) );
  AOI211xp5_ASAP7_75t_SL U68947 ( .A1(n76534), .A2(n58554), .B(n61692), .C(
        n61691), .Y(n61696) );
  AOI211xp5_ASAP7_75t_SL U68948 ( .A1(n77623), .A2(n61684), .B(n61683), .C(
        n61682), .Y(n61685) );
  NOR2xp33_ASAP7_75t_SL U68949 ( .A(or1200_cpu_or1200_mult_mac_n227), .B(
        n74587), .Y(n61683) );
  NOR2xp33_ASAP7_75t_SL U68950 ( .A(n1790), .B(n76717), .Y(n61680) );
  AOI211xp5_ASAP7_75t_SL U68951 ( .A1(or1200_cpu_rf_datab[18]), .A2(n57091), 
        .B(n77184), .C(n63603), .Y(n63604) );
  NOR4xp25_ASAP7_75t_SL U68952 ( .A(n63593), .B(n63592), .C(n63591), .D(n63590), .Y(n63594) );
  NOR2xp33_ASAP7_75t_SL U68953 ( .A(n63588), .B(n63587), .Y(n63589) );
  AOI211xp5_ASAP7_75t_SL U68954 ( .A1(or1200_cpu_or1200_except_n524), .A2(
        n75311), .B(n76791), .C(n74593), .Y(n63597) );
  AOI211xp5_ASAP7_75t_SL U68955 ( .A1(n63563), .A2(n63562), .B(n75882), .C(
        n74596), .Y(n63598) );
  AOI211xp5_ASAP7_75t_SL U68956 ( .A1(n77051), .A2(n74983), .B(n63561), .C(
        n63560), .Y(n77651) );
  AOI211xp5_ASAP7_75t_SL U68957 ( .A1(or1200_cpu_rf_datab[16]), .A2(n57091), 
        .B(n77184), .C(n62547), .Y(n62548) );
  AOI211xp5_ASAP7_75t_SL U68958 ( .A1(n75876), .A2(n62544), .B(n62543), .C(
        n62542), .Y(n62545) );
  AOI211xp5_ASAP7_75t_SL U68959 ( .A1(n73921), .A2(n63536), .B(n62528), .C(
        n62527), .Y(n62529) );
  NOR2xp33_ASAP7_75t_SL U68960 ( .A(or1200_cpu_or1200_mult_mac_n319), .B(
        n75738), .Y(n62527) );
  AOI211xp5_ASAP7_75t_SL U68961 ( .A1(n75577), .A2(n62518), .B(n62517), .C(
        n62516), .Y(n62524) );
  AOI211xp5_ASAP7_75t_SL U68962 ( .A1(n62514), .A2(n77113), .B(n75882), .C(
        n75360), .Y(n62543) );
  AOI211xp5_ASAP7_75t_SL U68963 ( .A1(n75368), .A2(n63536), .B(n62505), .C(
        n62504), .Y(n62506) );
  AOI211xp5_ASAP7_75t_SL U68964 ( .A1(or1200_cpu_rf_datab[12]), .A2(n57091), 
        .B(n62474), .C(n62473), .Y(n62475) );
  NOR2xp33_ASAP7_75t_SL U68965 ( .A(n2196), .B(n59679), .Y(n62473) );
  NOR2xp33_ASAP7_75t_SL U68966 ( .A(n59387), .B(n59688), .Y(n62472) );
  NOR2xp33_ASAP7_75t_SL U68967 ( .A(n62469), .B(n76557), .Y(n62470) );
  NOR2xp33_ASAP7_75t_SL U68968 ( .A(n73953), .B(n76300), .Y(n62467) );
  AOI211xp5_ASAP7_75t_SL U68969 ( .A1(n77082), .A2(n62450), .B(n62449), .C(
        n62448), .Y(n62451) );
  NOR2xp33_ASAP7_75t_SL U68970 ( .A(n75316), .B(n64121), .Y(n62448) );
  NOR4xp25_ASAP7_75t_SL U68971 ( .A(n62443), .B(n62442), .C(n62441), .D(n62440), .Y(n62452) );
  NOR2xp33_ASAP7_75t_SL U68972 ( .A(n62422), .B(n64136), .Y(n62443) );
  NOR4xp25_ASAP7_75t_SL U68973 ( .A(n62413), .B(n62412), .C(n62411), .D(n62410), .Y(n62414) );
  NOR2xp33_ASAP7_75t_SL U68974 ( .A(n76729), .B(n77626), .Y(n62412) );
  AOI211xp5_ASAP7_75t_SL U68975 ( .A1(or1200_cpu_rf_datab[10]), .A2(n57091), 
        .B(n61804), .C(n61803), .Y(n61805) );
  NOR2xp33_ASAP7_75t_SL U68976 ( .A(n1804), .B(n59679), .Y(n61804) );
  NOR2xp33_ASAP7_75t_SL U68977 ( .A(n73953), .B(n76302), .Y(n61801) );
  NOR2xp33_ASAP7_75t_SL U68978 ( .A(n76791), .B(n61772), .Y(n61773) );
  NOR4xp25_ASAP7_75t_SL U68979 ( .A(n64111), .B(n64303), .C(n63572), .D(n60859), .Y(n63577) );
  AOI211xp5_ASAP7_75t_SL U68980 ( .A1(n62382), .A2(n77613), .B(n61771), .C(
        n61770), .Y(n61793) );
  NAND2xp33_ASAP7_75t_SRAM U68981 ( .A(n57082), .B(n59586), .Y(n61192) );
  NOR2xp33_ASAP7_75t_SL U68982 ( .A(n61784), .B(n62353), .Y(n62273) );
  NOR2xp33_ASAP7_75t_SL U68983 ( .A(n60797), .B(n64109), .Y(n60789) );
  NOR2xp33_ASAP7_75t_SL U68984 ( .A(n63566), .B(n62447), .Y(n61768) );
  NOR2xp33_ASAP7_75t_SL U68985 ( .A(n62422), .B(n63564), .Y(n61771) );
  NOR2xp33_ASAP7_75t_SL U68986 ( .A(n1807), .B(n76717), .Y(n61747) );
  AOI211xp5_ASAP7_75t_SL U68987 ( .A1(n75876), .A2(n64139), .B(n64138), .C(
        n64137), .Y(n64140) );
  AOI211xp5_ASAP7_75t_SL U68988 ( .A1(n75862), .A2(n75584), .B(n64134), .C(
        n64133), .Y(n64135) );
  AOI211xp5_ASAP7_75t_SL U68989 ( .A1(n64119), .A2(n75833), .B(n64118), .C(
        n64117), .Y(n64120) );
  AOI211xp5_ASAP7_75t_SL U68990 ( .A1(n77039), .A2(n65079), .B(n64100), .C(
        n64099), .Y(n64101) );
  NOR2xp33_ASAP7_75t_SL U68991 ( .A(or1200_cpu_or1200_mult_mac_n245), .B(
        n74587), .Y(n64099) );
  AOI211xp5_ASAP7_75t_SL U68992 ( .A1(or1200_cpu_rf_datab[13]), .A2(n57091), 
        .B(n61129), .C(n61128), .Y(n61130) );
  NOR2xp33_ASAP7_75t_SL U68993 ( .A(n1776), .B(n59679), .Y(n61129) );
  NOR4xp25_ASAP7_75t_SL U68994 ( .A(n61115), .B(n61114), .C(n61113), .D(n61112), .Y(n61116) );
  AOI211xp5_ASAP7_75t_SL U68995 ( .A1(n61109), .A2(n61658), .B(n61108), .C(
        n61107), .Y(n61111) );
  AOI211xp5_ASAP7_75t_SL U68996 ( .A1(n73921), .A2(n63489), .B(n61102), .C(
        n61101), .Y(n61103) );
  NOR2xp33_ASAP7_75t_SL U68997 ( .A(or1200_cpu_or1200_mult_mac_n313), .B(
        n75738), .Y(n61101) );
  AOI211xp5_ASAP7_75t_SL U68998 ( .A1(n75577), .A2(n61357), .B(n61089), .C(
        n61088), .Y(n61091) );
  NOR2xp33_ASAP7_75t_SL U68999 ( .A(n76791), .B(n77080), .Y(n61085) );
  NOR2xp33_ASAP7_75t_SL U69000 ( .A(n76801), .B(n75217), .Y(n61115) );
  AOI211xp5_ASAP7_75t_SL U69001 ( .A1(n77051), .A2(n77224), .B(n61073), .C(
        n61072), .Y(n61074) );
  NOR2xp33_ASAP7_75t_SL U69002 ( .A(n1376), .B(n76716), .Y(n61068) );
  NOR2xp33_ASAP7_75t_SL U69003 ( .A(n1779), .B(n76717), .Y(n61061) );
  AOI211xp5_ASAP7_75t_SL U69004 ( .A1(n75235), .A2(n64235), .B(n64234), .C(
        n64829), .Y(n64236) );
  NAND2xp33_ASAP7_75t_SRAM U69005 ( .A(n59584), .B(n62682), .Y(n63566) );
  AOI211xp5_ASAP7_75t_SL U69006 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[25]), 
        .B(n64207), .C(n64206), .Y(n64214) );
  NOR2xp33_ASAP7_75t_SL U69007 ( .A(n76791), .B(n64814), .Y(n64202) );
  NOR4xp25_ASAP7_75t_SL U69008 ( .A(n75354), .B(n75353), .C(n75352), .D(n75351), .Y(n75355) );
  AOI211xp5_ASAP7_75t_SL U69009 ( .A1(n75342), .A2(n75341), .B(n75340), .C(
        n75339), .Y(n75343) );
  NOR2xp33_ASAP7_75t_SL U69010 ( .A(n76765), .B(n75324), .Y(n75334) );
  AOI211xp5_ASAP7_75t_SL U69011 ( .A1(n75323), .A2(n75322), .B(n75321), .C(
        n75320), .Y(n75345) );
  AOI211xp5_ASAP7_75t_SL U69012 ( .A1(n75368), .A2(n75367), .B(n75366), .C(
        n75365), .Y(n75369) );
  AOI211xp5_ASAP7_75t_SL U69013 ( .A1(or1200_cpu_rf_datab[17]), .A2(n57091), 
        .B(n77184), .C(n75381), .Y(n75385) );
  NOR4xp25_ASAP7_75t_SL U69014 ( .A(n75599), .B(n75598), .C(n75597), .D(n75596), .Y(n75600) );
  NOR2xp33_ASAP7_75t_SL U69015 ( .A(n76796), .B(n77656), .Y(n75599) );
  AOI211xp5_ASAP7_75t_SL U69016 ( .A1(n75585), .A2(n75584), .B(n75583), .C(
        n75582), .Y(n75601) );
  NAND2xp33_ASAP7_75t_SRAM U69017 ( .A(n59711), .B(n59575), .Y(n61706) );
  AOI211xp5_ASAP7_75t_SL U69018 ( .A1(or1200_cpu_rf_datab[23]), .A2(n57091), 
        .B(n77184), .C(n75610), .Y(n75615) );
  AOI211xp5_ASAP7_75t_SL U69019 ( .A1(n75890), .A2(n75869), .B(n75868), .C(
        n75867), .Y(n75873) );
  NOR2xp33_ASAP7_75t_SL U69020 ( .A(n62424), .B(n62423), .Y(n75860) );
  NAND2xp33_ASAP7_75t_SRAM U69021 ( .A(n75855), .B(n76753), .Y(n75856) );
  AOI211xp5_ASAP7_75t_SL U69022 ( .A1(n75845), .A2(n75844), .B(n75843), .C(
        n75842), .Y(n75874) );
  NAND2xp33_ASAP7_75t_SRAM U69023 ( .A(n61481), .B(n61480), .Y(n75826) );
  AOI211xp5_ASAP7_75t_SL U69024 ( .A1(n75823), .A2(n75822), .B(n75821), .C(
        n75820), .Y(n75824) );
  NOR2xp33_ASAP7_75t_SL U69025 ( .A(or1200_cpu_or1200_mult_mac_n197), .B(
        n75819), .Y(n75820) );
  AOI211xp5_ASAP7_75t_SL U69026 ( .A1(n65140), .A2(n75342), .B(n64789), .C(
        n64788), .Y(n64790) );
  NAND2xp33_ASAP7_75t_SRAM U69027 ( .A(n59561), .B(n59587), .Y(n64781) );
  NOR2xp33_ASAP7_75t_SL U69028 ( .A(n59535), .B(n63571), .Y(n64109) );
  NOR2xp33_ASAP7_75t_SL U69029 ( .A(n59531), .B(n59584), .Y(n64111) );
  NAND2xp33_ASAP7_75t_SRAM U69030 ( .A(n77242), .B(n59646), .Y(n64768) );
  NAND2xp33_ASAP7_75t_SRAM U69031 ( .A(n59183), .B(n59583), .Y(n61435) );
  NOR2xp33_ASAP7_75t_SL U69032 ( .A(n61434), .B(n61433), .Y(n61437) );
  NOR2xp33_ASAP7_75t_SL U69033 ( .A(n59557), .B(n59584), .Y(n61433) );
  AOI211xp5_ASAP7_75t_SL U69034 ( .A1(n77039), .A2(n64761), .B(n64760), .C(
        n64759), .Y(n64762) );
  NOR2xp33_ASAP7_75t_SL U69035 ( .A(or1200_cpu_or1200_mult_mac_n253), .B(
        n74587), .Y(n64759) );
  NOR2xp33_ASAP7_75t_SL U69036 ( .A(n64855), .B(n64317), .Y(n64318) );
  AOI211xp5_ASAP7_75t_SL U69037 ( .A1(n75876), .A2(n64315), .B(n64314), .C(
        n74626), .Y(n64323) );
  NOR4xp25_ASAP7_75t_SL U69038 ( .A(n64310), .B(n64309), .C(n64308), .D(n64307), .Y(n64311) );
  NOR2xp33_ASAP7_75t_SL U69039 ( .A(n75745), .B(n77103), .Y(n64308) );
  AOI211xp5_ASAP7_75t_SL U69040 ( .A1(n75705), .A2(n75577), .B(n64297), .C(
        n64296), .Y(n64298) );
  NOR2xp33_ASAP7_75t_SL U69041 ( .A(or1200_cpu_or1200_mult_mac_n185), .B(
        n74606), .Y(n64296) );
  AOI211xp5_ASAP7_75t_SL U69042 ( .A1(n75701), .A2(n59709), .B(n75699), .C(
        n64295), .Y(n64297) );
  NOR2xp33_ASAP7_75t_SL U69043 ( .A(n59563), .B(n59584), .Y(n64784) );
  AOI211xp5_ASAP7_75t_SL U69044 ( .A1(n77659), .A2(n75561), .B(n1510), .C(
        n64284), .Y(n64285) );
  AOI211xp5_ASAP7_75t_SL U69045 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[22]), 
        .B(n64280), .C(n64279), .Y(n64281) );
  NOR2xp33_ASAP7_75t_SL U69046 ( .A(or1200_cpu_or1200_except_n142), .B(n57102), 
        .Y(n64279) );
  OR2x2_ASAP7_75t_SL U69047 ( .A(n60827), .B(n60826), .Y(n76724) );
  NAND2xp33_ASAP7_75t_SRAM U69048 ( .A(n76675), .B(n75453), .Y(n60827) );
  NOR2xp33_ASAP7_75t_SL U69049 ( .A(n73953), .B(n76277), .Y(n64326) );
  AOI211xp5_ASAP7_75t_SL U69050 ( .A1(or1200_cpu_rf_datab[22]), .A2(n57091), 
        .B(n77184), .C(n64328), .Y(n64332) );
  NOR2xp33_ASAP7_75t_SL U69051 ( .A(n70096), .B(n70095), .Y(n2267) );
  AOI211xp5_ASAP7_75t_SL U69052 ( .A1(n70094), .A2(n70093), .B(n58553), .C(
        n70097), .Y(n70095) );
  AOI211xp5_ASAP7_75t_SL U69053 ( .A1(n74733), .A2(n59705), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_0_), 
        .C(n74732), .Y(n74735) );
  NOR2xp33_ASAP7_75t_SL U69054 ( .A(n3310), .B(n73652), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_N190) );
  NOR2xp33_ASAP7_75t_SL U69055 ( .A(n65288), .B(n65331), .Y(n2008) );
  NOR2xp33_ASAP7_75t_SL U69056 ( .A(n65305), .B(n65331), .Y(n1997) );
  NOR2xp33_ASAP7_75t_SL U69057 ( .A(n65285), .B(n65331), .Y(n2003) );
  AOI211xp5_ASAP7_75t_SL U69058 ( .A1(n77217), .A2(n76668), .B(n76667), .C(
        n76666), .Y(or1200_cpu_or1200_except_n283) );
  NOR2xp33_ASAP7_75t_SL U69059 ( .A(n76665), .B(n77143), .Y(n76666) );
  AOI31xp33_ASAP7_75t_SL U69060 ( .A1(n77833), .A2(n77501), .A3(n77503), .B(
        n77402), .Y(iwb_biu_N62) );
  NOR2xp33_ASAP7_75t_SL U69061 ( .A(n70926), .B(n70925), .Y(n70924) );
  NOR2xp33_ASAP7_75t_SL U69062 ( .A(n70937), .B(n58303), .Y(n70926) );
  NAND2xp33_ASAP7_75t_SRAM U69063 ( .A(n75769), .B(n77459), .Y(n61059) );
  NOR2xp33_ASAP7_75t_SL U69064 ( .A(n62013), .B(n75509), .Y(n75512) );
  NOR4xp25_ASAP7_75t_SL U69065 ( .A(n1504), .B(n53614), .C(n75488), .D(n75487), 
        .Y(n75516) );
  NOR4xp25_ASAP7_75t_SL U69066 ( .A(n59543), .B(n59580), .C(n59532), .D(n59554), .Y(n75483) );
  NOR4xp25_ASAP7_75t_SL U69067 ( .A(n59556), .B(n59553), .C(n59539), .D(n59581), .Y(n75484) );
  NOR4xp25_ASAP7_75t_SL U69068 ( .A(n75866), .B(n59708), .C(n59546), .D(n59582), .Y(n75485) );
  NOR4xp25_ASAP7_75t_SL U69069 ( .A(n59544), .B(n59534), .C(n1626), .D(n59536), 
        .Y(n75480) );
  NOR2xp33_ASAP7_75t_SL U69070 ( .A(n57318), .B(n75476), .Y(n75479) );
  AOI211xp5_ASAP7_75t_SL U69071 ( .A1(n65357), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_19_), .B(n65293), .C(
        n65331), .Y(n1633) );
  AOI211xp5_ASAP7_75t_SL U69072 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_19_), .A2(n65368), .B(
        n65354), .C(n65292), .Y(n65293) );
  AOI211xp5_ASAP7_75t_SL U69073 ( .A1(n65357), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_18_), .B(n65291), .C(
        n65331), .Y(n1647) );
  AOI31xp33_ASAP7_75t_SL U69074 ( .A1(n76912), .A2(n57079), .A3(n76911), .B(
        n76910), .Y(n76913) );
  NOR4xp25_ASAP7_75t_SL U69075 ( .A(n76912), .B(n76911), .C(n76900), .D(n59671), .Y(n76898) );
  NOR2xp33_ASAP7_75t_SL U69076 ( .A(n75651), .B(n75653), .Y(n75657) );
  NOR2xp33_ASAP7_75t_SL U69077 ( .A(n62355), .B(n60800), .Y(n61106) );
  AOI211xp5_ASAP7_75t_SL U69078 ( .A1(n75246), .A2(n64217), .B(n62119), .C(
        n62118), .Y(n62120) );
  OR2x2_ASAP7_75t_SL U69079 ( .A(n62418), .B(n77621), .Y(n77034) );
  OR2x2_ASAP7_75t_SL U69080 ( .A(n62419), .B(n77621), .Y(n77033) );
  NOR2xp33_ASAP7_75t_SL U69081 ( .A(n73609), .B(n73601), .Y(n73604) );
  NOR4xp25_ASAP7_75t_SL U69082 ( .A(n77167), .B(n77166), .C(n77165), .D(n77164), .Y(n77237) );
  AOI31xp33_ASAP7_75t_SL U69083 ( .A1(n78173), .A2(n63268), .A3(n63267), .B(
        n63269), .Y(n68813) );
  AOI31xp33_ASAP7_75t_SL U69084 ( .A1(n73616), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[4]), .A3(n73615), 
        .B(n73614), .Y(n1524) );
  NOR2xp33_ASAP7_75t_SL U69085 ( .A(n73872), .B(n73652), .Y(n73614) );
  NOR2xp33_ASAP7_75t_SL U69086 ( .A(n65354), .B(n65271), .Y(n65278) );
  NOR2xp33_ASAP7_75t_SL U69087 ( .A(n59572), .B(n57196), .Y(n61884) );
  NOR2xp33_ASAP7_75t_SL U69088 ( .A(n59538), .B(n57197), .Y(n61887) );
  NOR2xp33_ASAP7_75t_SL U69089 ( .A(n59535), .B(n57197), .Y(n61882) );
  NOR2xp33_ASAP7_75t_SL U69090 ( .A(n61729), .B(n61728), .Y(n61730) );
  NOR2xp33_ASAP7_75t_SL U69091 ( .A(n59540), .B(n57196), .Y(n61729) );
  NOR2xp33_ASAP7_75t_SL U69092 ( .A(n59579), .B(n57196), .Y(n76768) );
  NOR4xp25_ASAP7_75t_SL U69093 ( .A(n61871), .B(n61870), .C(n61869), .D(n61868), .Y(n73942) );
  NOR2xp33_ASAP7_75t_SL U69094 ( .A(n59573), .B(n57196), .Y(n61868) );
  NOR2xp33_ASAP7_75t_SL U69095 ( .A(n59530), .B(n63571), .Y(n61869) );
  NOR2xp33_ASAP7_75t_SL U69096 ( .A(n59529), .B(n57197), .Y(n61871) );
  NAND2xp33_ASAP7_75t_SRAM U69097 ( .A(n59079), .B(n59646), .Y(n61489) );
  NOR2xp33_ASAP7_75t_SL U69098 ( .A(n61724), .B(n61723), .Y(n61727) );
  NOR2xp33_ASAP7_75t_SL U69099 ( .A(n59571), .B(n57196), .Y(n61724) );
  NOR2xp33_ASAP7_75t_SL U69100 ( .A(n59579), .B(n75872), .Y(n61861) );
  AOI211xp5_ASAP7_75t_SL U69101 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[31]), 
        .B(n64207), .C(n61843), .Y(n61849) );
  NOR2xp33_ASAP7_75t_SL U69102 ( .A(n73594), .B(n73616), .Y(n73596) );
  NOR2xp33_ASAP7_75t_SL U69103 ( .A(n73593), .B(n73652), .Y(n73599) );
  AND4x1_ASAP7_75t_SL U69104 ( .A(n73653), .B(n73651), .C(n73581), .D(n73580), 
        .Y(n73584) );
  NOR2xp33_ASAP7_75t_SL U69105 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[1]), .B(n73602), 
        .Y(n73505) );
  NOR2xp33_ASAP7_75t_SL U69106 ( .A(n73962), .B(n74030), .Y(n74039) );
  NOR2xp33_ASAP7_75t_SL U69107 ( .A(n76503), .B(n73961), .Y(n74030) );
  NOR2xp33_ASAP7_75t_SL U69108 ( .A(n2961), .B(n77142), .Y(n73962) );
  NOR2xp33_ASAP7_75t_SL U69109 ( .A(n75781), .B(n58299), .Y(n73958) );
  AOI211xp5_ASAP7_75t_SL U69110 ( .A1(or1200_cpu_rf_datab[29]), .A2(n57091), 
        .B(n77184), .C(n75267), .Y(n75273) );
  NOR2xp33_ASAP7_75t_SL U69111 ( .A(n65329), .B(n65328), .Y(n65388) );
  NOR2xp33_ASAP7_75t_SL U69112 ( .A(n65252), .B(n65251), .Y(n65307) );
  AOI211xp5_ASAP7_75t_SL U69113 ( .A1(n75685), .A2(n75259), .B(n75258), .C(
        n75257), .Y(n75265) );
  NOR4xp25_ASAP7_75t_SL U69114 ( .A(n75254), .B(n75253), .C(n75252), .D(n75251), .Y(n75255) );
  NOR2xp33_ASAP7_75t_SL U69115 ( .A(n76764), .B(n75863), .Y(n77061) );
  NOR2xp33_ASAP7_75t_SL U69116 ( .A(n59560), .B(n63571), .Y(n62105) );
  NOR2xp33_ASAP7_75t_SL U69117 ( .A(n59537), .B(n59584), .Y(n62107) );
  NOR2xp33_ASAP7_75t_SL U69118 ( .A(n75242), .B(n75241), .Y(n75243) );
  NOR2xp33_ASAP7_75t_SL U69119 ( .A(n59541), .B(n63571), .Y(n61510) );
  NOR2xp33_ASAP7_75t_SL U69120 ( .A(n59570), .B(n59584), .Y(n61496) );
  NOR2xp33_ASAP7_75t_SL U69121 ( .A(n59555), .B(n63571), .Y(n61506) );
  NOR2xp33_ASAP7_75t_SL U69122 ( .A(n59569), .B(n59585), .Y(n61509) );
  NAND3xp33_ASAP7_75t_SL U69123 ( .A(n57214), .B(n59708), .C(n59567), .Y(
        n76765) );
  NOR2xp33_ASAP7_75t_SL U69124 ( .A(n59568), .B(n63571), .Y(n61095) );
  NOR2xp33_ASAP7_75t_SL U69125 ( .A(n59557), .B(n57197), .Y(n61096) );
  NOR2xp33_ASAP7_75t_SL U69126 ( .A(n59559), .B(n59585), .Y(n61505) );
  NOR2xp33_ASAP7_75t_SL U69127 ( .A(n75233), .B(n76779), .Y(n75234) );
  NOR2xp33_ASAP7_75t_SL U69128 ( .A(n59710), .B(n75456), .Y(n64232) );
  NOR2xp33_ASAP7_75t_SL U69129 ( .A(n59574), .B(n59584), .Y(n75226) );
  NOR2xp33_ASAP7_75t_SL U69130 ( .A(n75225), .B(n75224), .Y(n75231) );
  NOR2xp33_ASAP7_75t_SL U69131 ( .A(n59528), .B(n63571), .Y(n75225) );
  NOR2xp33_ASAP7_75t_SL U69132 ( .A(n75880), .B(n75269), .Y(n75266) );
  AOI211xp5_ASAP7_75t_SL U69133 ( .A1(n59686), .A2(or1200_cpu_spr_dat_rf[29]), 
        .B(n75207), .C(n75206), .Y(n75210) );
  NOR2xp33_ASAP7_75t_SL U69134 ( .A(or1200_cpu_or1200_except_n128), .B(n57102), 
        .Y(n75206) );
  NAND2xp33_ASAP7_75t_SRAM U69135 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .B(n65245), .Y(
        n65240) );
  NOR2xp33_ASAP7_75t_SL U69136 ( .A(n63362), .B(n63361), .Y(n63445) );
  NOR2xp33_ASAP7_75t_SL U69137 ( .A(n73900), .B(n74260), .Y(n2873) );
  NOR2xp33_ASAP7_75t_SL U69138 ( .A(n60339), .B(n57072), .Y(n60726) );
  AOI211xp5_ASAP7_75t_SL U69139 ( .A1(or1200_ic_top_from_icram[28]), .A2(
        n22057), .B(n77358), .C(n77357), .Y(n77360) );
  AOI211xp5_ASAP7_75t_SL U69140 ( .A1(or1200_ic_top_from_icram[26]), .A2(
        n22057), .B(n60321), .C(n77357), .Y(n60318) );
  NOR2xp33_ASAP7_75t_SL U69141 ( .A(n75753), .B(n75752), .Y(n75754) );
  AOI211xp5_ASAP7_75t_SL U69142 ( .A1(n75751), .A2(n75750), .B(n75882), .C(
        n75749), .Y(n75752) );
  NOR2xp33_ASAP7_75t_SL U69143 ( .A(or1200_cpu_or1200_mult_mac_n301), .B(
        n61828), .Y(n62346) );
  NOR2xp33_ASAP7_75t_SL U69144 ( .A(or1200_cpu_or1200_mult_mac_n303), .B(
        n61828), .Y(n62351) );
  AOI211xp5_ASAP7_75t_SL U69145 ( .A1(n75727), .A2(n75726), .B(n75725), .C(
        n75724), .Y(n75728) );
  AOI211xp5_ASAP7_75t_SL U69146 ( .A1(n76766), .A2(n75717), .B(n75716), .C(
        n75715), .Y(n75718) );
  NOR2xp33_ASAP7_75t_SL U69147 ( .A(n59708), .B(n59558), .Y(n61087) );
  NOR2xp33_ASAP7_75t_SL U69148 ( .A(n59533), .B(n57196), .Y(n63572) );
  NOR2xp33_ASAP7_75t_SL U69149 ( .A(n59486), .B(n57197), .Y(n63574) );
  NAND2xp33_ASAP7_75t_SRAM U69150 ( .A(n75832), .B(n75708), .Y(n75709) );
  NOR2xp33_ASAP7_75t_SL U69151 ( .A(n59576), .B(n57196), .Y(n75707) );
  NOR2xp33_ASAP7_75t_SL U69152 ( .A(n60797), .B(n60796), .Y(n60798) );
  NAND2xp33_ASAP7_75t_SRAM U69153 ( .A(n59711), .B(n59570), .Y(n61190) );
  NOR2xp33_ASAP7_75t_SL U69154 ( .A(n59530), .B(n57197), .Y(n64837) );
  NOR2xp33_ASAP7_75t_SL U69155 ( .A(n59709), .B(n62257), .Y(n75699) );
  NOR2xp33_ASAP7_75t_SL U69156 ( .A(n61184), .B(n60847), .Y(n60848) );
  NOR2xp33_ASAP7_75t_SL U69157 ( .A(n59559), .B(n57197), .Y(n60847) );
  NOR2xp33_ASAP7_75t_SL U69158 ( .A(n59555), .B(n57196), .Y(n61184) );
  NOR2xp33_ASAP7_75t_SL U69159 ( .A(n59568), .B(n57196), .Y(n61183) );
  NOR4xp25_ASAP7_75t_SL U69160 ( .A(n64304), .B(n64303), .C(n64302), .D(n64301), .Y(n75745) );
  NOR2xp33_ASAP7_75t_SL U69161 ( .A(n59561), .B(n57196), .Y(n64302) );
  NOR2xp33_ASAP7_75t_SL U69162 ( .A(n57377), .B(n57197), .Y(n64303) );
  NOR2xp33_ASAP7_75t_SL U69163 ( .A(n59571), .B(n2141), .Y(n60871) );
  NOR2xp33_ASAP7_75t_SL U69164 ( .A(n57214), .B(n62682), .Y(n73916) );
  AOI211xp5_ASAP7_75t_SL U69165 ( .A1(n75823), .A2(
        or1200_cpu_or1200_mult_mac_n265), .B(n75694), .C(n75693), .Y(n75695)
         );
  NOR2xp33_ASAP7_75t_SL U69166 ( .A(n75692), .B(n75819), .Y(n75693) );
  NAND2xp33_ASAP7_75t_SRAM U69167 ( .A(n64209), .B(n64208), .Y(n75817) );
  NOR2xp33_ASAP7_75t_SL U69168 ( .A(n59493), .B(n61845), .Y(n75823) );
  AND2x2_ASAP7_75t_SL U69169 ( .A(n61156), .B(n61060), .Y(n58554) );
  NOR2xp33_ASAP7_75t_SL U69170 ( .A(n77171), .B(n76242), .Y(n52505) );
  NOR2xp33_ASAP7_75t_SL U69171 ( .A(or1200_ic_top_from_icram[16]), .B(n77833), 
        .Y(n60506) );
  NOR2xp33_ASAP7_75t_SL U69172 ( .A(n71279), .B(n71278), .Y(n71277) );
  AOI211xp5_ASAP7_75t_SL U69173 ( .A1(n74258), .A2(n74105), .B(n74104), .C(
        n74260), .Y(n2874) );
  AOI211xp5_ASAP7_75t_SL U69174 ( .A1(n74103), .A2(n74102), .B(n74101), .C(
        n58298), .Y(n74104) );
  NOR2xp33_ASAP7_75t_SL U69175 ( .A(n69957), .B(n70003), .Y(n69959) );
  NOR2xp33_ASAP7_75t_SL U69176 ( .A(n69694), .B(n70528), .Y(n69695) );
  NOR2xp33_ASAP7_75t_SL U69177 ( .A(n69686), .B(n59521), .Y(n69691) );
  NOR2xp33_ASAP7_75t_SL U69178 ( .A(n69684), .B(n69683), .Y(n69957) );
  NOR2xp33_ASAP7_75t_SL U69179 ( .A(n69680), .B(n59520), .Y(n69684) );
  NOR2xp33_ASAP7_75t_SL U69180 ( .A(n69672), .B(n70528), .Y(n69678) );
  NOR2xp33_ASAP7_75t_SL U69181 ( .A(n69667), .B(n59521), .Y(n69668) );
  NOR2xp33_ASAP7_75t_SL U69182 ( .A(n69651), .B(n59520), .Y(n69652) );
  NOR2xp33_ASAP7_75t_SL U69183 ( .A(n69647), .B(n70528), .Y(n69648) );
  NOR2xp33_ASAP7_75t_SL U69184 ( .A(n69855), .B(n70103), .Y(n69645) );
  NOR2xp33_ASAP7_75t_SL U69185 ( .A(n69631), .B(n59521), .Y(n69642) );
  NOR2xp33_ASAP7_75t_SL U69186 ( .A(n69624), .B(n59520), .Y(n69630) );
  NOR2xp33_ASAP7_75t_SL U69187 ( .A(n69802), .B(n69799), .Y(n69637) );
  NOR2xp33_ASAP7_75t_SL U69188 ( .A(n69621), .B(n70528), .Y(n69625) );
  NOR2xp33_ASAP7_75t_SL U69189 ( .A(n69601), .B(n69786), .Y(n69780) );
  NOR2xp33_ASAP7_75t_SL U69190 ( .A(n69584), .B(n70528), .Y(n69585) );
  NOR2xp33_ASAP7_75t_SL U69191 ( .A(n65114), .B(n65113), .Y(n65119) );
  NOR2xp33_ASAP7_75t_SL U69192 ( .A(n2609), .B(n62022), .Y(n62003) );
  AOI211xp5_ASAP7_75t_SL U69193 ( .A1(n76842), .A2(n77262), .B(n76843), .C(
        n59703), .Y(n76838) );
  NAND2xp33_ASAP7_75t_SRAM U69194 ( .A(n62009), .B(n62000), .Y(n61146) );
  NOR2xp33_ASAP7_75t_SL U69195 ( .A(n2616), .B(n77426), .Y(n61139) );
  NOR4xp25_ASAP7_75t_SL U69196 ( .A(n61138), .B(n61137), .C(n62014), .D(n62016), .Y(n61149) );
  NAND2xp33_ASAP7_75t_SRAM U69197 ( .A(n2609), .B(n2172), .Y(n62016) );
  AOI211xp5_ASAP7_75t_SL U69198 ( .A1(n77426), .A2(n61032), .B(n77427), .C(
        n62024), .Y(n61134) );
  AOI211xp5_ASAP7_75t_SL U69199 ( .A1(n76926), .A2(n76584), .B(n76583), .C(
        n76582), .Y(n76586) );
  NOR2xp33_ASAP7_75t_SL U69200 ( .A(or1200_cpu_or1200_except_n404), .B(n63715), 
        .Y(n76582) );
  AOI211xp5_ASAP7_75t_SL U69201 ( .A1(n76926), .A2(n76703), .B(n76702), .C(
        n76701), .Y(n76706) );
  NOR2xp33_ASAP7_75t_SL U69202 ( .A(or1200_cpu_or1200_except_n413), .B(n63715), 
        .Y(n76701) );
  AOI211xp5_ASAP7_75t_SL U69203 ( .A1(n76926), .A2(n77275), .B(n76212), .C(
        n76211), .Y(n76214) );
  NOR2xp33_ASAP7_75t_SL U69204 ( .A(or1200_cpu_or1200_except_n407), .B(n63715), 
        .Y(n76211) );
  AOI211xp5_ASAP7_75t_SL U69205 ( .A1(n76926), .A2(n76252), .B(n76251), .C(
        n76250), .Y(n76255) );
  NOR2xp33_ASAP7_75t_SL U69206 ( .A(or1200_cpu_or1200_except_n419), .B(n63715), 
        .Y(n76250) );
  AOI211xp5_ASAP7_75t_SL U69207 ( .A1(n76926), .A2(n76849), .B(n76645), .C(
        n76644), .Y(n76647) );
  NOR2xp33_ASAP7_75t_SL U69208 ( .A(or1200_cpu_or1200_except_n416), .B(n63715), 
        .Y(n76644) );
  AOI211xp5_ASAP7_75t_SL U69209 ( .A1(n76926), .A2(n76607), .B(n76597), .C(
        n76596), .Y(n76599) );
  NOR2xp33_ASAP7_75t_SL U69210 ( .A(or1200_cpu_or1200_except_n410), .B(n63715), 
        .Y(n76596) );
  AOI211xp5_ASAP7_75t_SL U69211 ( .A1(n76926), .A2(n64165), .B(n64159), .C(
        n64158), .Y(n64161) );
  NOR2xp33_ASAP7_75t_SL U69212 ( .A(or1200_cpu_spr_dat_ppc[20]), .B(n63715), 
        .Y(n64158) );
  AOI211xp5_ASAP7_75t_SL U69213 ( .A1(n76926), .A2(n75421), .B(n75411), .C(
        n75410), .Y(n75413) );
  NOR2xp33_ASAP7_75t_SL U69214 ( .A(or1200_cpu_spr_dat_ppc[21]), .B(n63715), 
        .Y(n75410) );
  AOI211xp5_ASAP7_75t_SL U69215 ( .A1(n76926), .A2(n76534), .B(n76525), .C(
        n76524), .Y(n76527) );
  NOR2xp33_ASAP7_75t_SL U69216 ( .A(or1200_cpu_or1200_except_n425), .B(n63715), 
        .Y(n76524) );
  AOI211xp5_ASAP7_75t_SL U69217 ( .A1(n76926), .A2(n75167), .B(n75166), .C(
        n75165), .Y(n75169) );
  NOR2xp33_ASAP7_75t_SL U69218 ( .A(or1200_cpu_or1200_except_n476), .B(n63715), 
        .Y(n75165) );
  AOI211xp5_ASAP7_75t_SL U69219 ( .A1(n76926), .A2(n65234), .B(n65188), .C(
        n65187), .Y(n65190) );
  NOR2xp33_ASAP7_75t_SL U69220 ( .A(or1200_cpu_spr_dat_ppc[26]), .B(n63715), 
        .Y(n65187) );
  AOI211xp5_ASAP7_75t_SL U69221 ( .A1(n76926), .A2(n74970), .B(n74963), .C(
        n74962), .Y(n74965) );
  NOR2xp33_ASAP7_75t_SL U69222 ( .A(or1200_cpu_or1200_except_n446), .B(n63715), 
        .Y(n74962) );
  AOI211xp5_ASAP7_75t_SL U69223 ( .A1(n76926), .A2(n75153), .B(n75152), .C(
        n75151), .Y(n75155) );
  NOR2xp33_ASAP7_75t_SL U69224 ( .A(or1200_cpu_spr_dat_ppc[27]), .B(n63715), 
        .Y(n75151) );
  AOI211xp5_ASAP7_75t_SL U69225 ( .A1(n76926), .A2(n65218), .B(n65198), .C(
        n65197), .Y(n65200) );
  NOR2xp33_ASAP7_75t_SL U69226 ( .A(or1200_cpu_spr_dat_ppc[24]), .B(n63715), 
        .Y(n65197) );
  NOR2xp33_ASAP7_75t_SL U69227 ( .A(or1200_cpu_or1200_except_n398), .B(n63715), 
        .Y(n76563) );
  AOI211xp5_ASAP7_75t_SL U69228 ( .A1(n76926), .A2(n65222), .B(n65215), .C(
        n65214), .Y(n65217) );
  NOR2xp33_ASAP7_75t_SL U69229 ( .A(or1200_cpu_or1200_except_n467), .B(n63715), 
        .Y(n65214) );
  AOI211xp5_ASAP7_75t_SL U69230 ( .A1(n76926), .A2(n64267), .B(n64261), .C(
        n64260), .Y(n64263) );
  NOR2xp33_ASAP7_75t_SL U69231 ( .A(or1200_cpu_spr_dat_ppc[22]), .B(n63715), 
        .Y(n64260) );
  AOI211xp5_ASAP7_75t_SL U69232 ( .A1(n76926), .A2(n75640), .B(n75634), .C(
        n75633), .Y(n75636) );
  NOR2xp33_ASAP7_75t_SL U69233 ( .A(or1200_cpu_or1200_except_n482), .B(n63715), 
        .Y(n75633) );
  AOI211xp5_ASAP7_75t_SL U69234 ( .A1(n76926), .A2(n75186), .B(n75177), .C(
        n75176), .Y(n75179) );
  NOR2xp33_ASAP7_75t_SL U69235 ( .A(or1200_cpu_spr_dat_ppc[29]), .B(n63715), 
        .Y(n75176) );
  AOI211xp5_ASAP7_75t_SL U69236 ( .A1(n76926), .A2(n63998), .B(n63990), .C(
        n63989), .Y(n63992) );
  NOR2xp33_ASAP7_75t_SL U69237 ( .A(or1200_cpu_or1200_except_n437), .B(n63715), 
        .Y(n63989) );
  AOI211xp5_ASAP7_75t_SL U69238 ( .A1(n76926), .A2(n75546), .B(n75537), .C(
        n75536), .Y(n75539) );
  NOR2xp33_ASAP7_75t_SL U69239 ( .A(or1200_cpu_or1200_except_n461), .B(n63715), 
        .Y(n75536) );
  AOI211xp5_ASAP7_75t_SL U69240 ( .A1(n76926), .A2(n76925), .B(n76924), .C(
        n76923), .Y(n76930) );
  NOR2xp33_ASAP7_75t_SL U69241 ( .A(or1200_cpu_spr_dat_ppc[31]), .B(n63715), 
        .Y(n76923) );
  AOI211xp5_ASAP7_75t_SL U69242 ( .A1(n76926), .A2(n63972), .B(n63971), .C(
        n63970), .Y(n63974) );
  NOR2xp33_ASAP7_75t_SL U69243 ( .A(or1200_cpu_or1200_except_n434), .B(n63715), 
        .Y(n63970) );
  AOI211xp5_ASAP7_75t_SL U69244 ( .A1(n76926), .A2(n76574), .B(n76573), .C(
        n76572), .Y(n76576) );
  NOR2xp33_ASAP7_75t_SL U69245 ( .A(or1200_cpu_or1200_except_n401), .B(n63715), 
        .Y(n76572) );
  AND2x2_ASAP7_75t_SL U69246 ( .A(n65322), .B(n65308), .Y(n65313) );
  AOI211xp5_ASAP7_75t_SL U69247 ( .A1(n77125), .A2(n60987), .B(n60986), .C(
        n60985), .Y(n60988) );
  NOR2xp33_ASAP7_75t_SL U69248 ( .A(n60976), .B(n60975), .Y(n60989) );
  NOR2xp33_ASAP7_75t_SL U69249 ( .A(n60964), .B(n61649), .Y(n61500) );
  NOR2xp33_ASAP7_75t_SL U69250 ( .A(n59537), .B(n63571), .Y(n61880) );
  NOR2xp33_ASAP7_75t_SL U69251 ( .A(n59538), .B(n57196), .Y(n61104) );
  NOR2xp33_ASAP7_75t_SL U69252 ( .A(n59560), .B(n59585), .Y(n61886) );
  NOR2xp33_ASAP7_75t_SL U69253 ( .A(n59572), .B(n57197), .Y(n62108) );
  NOR2xp33_ASAP7_75t_SL U69254 ( .A(n59570), .B(n63571), .Y(n61885) );
  NOR2xp33_ASAP7_75t_SL U69255 ( .A(n61097), .B(n61105), .Y(n60958) );
  NOR2xp33_ASAP7_75t_SL U69256 ( .A(n59540), .B(n57197), .Y(n61105) );
  NOR2xp33_ASAP7_75t_SL U69257 ( .A(n59542), .B(n57196), .Y(n61097) );
  NOR2xp33_ASAP7_75t_SL U69258 ( .A(n59709), .B(n61531), .Y(n62279) );
  NOR2xp33_ASAP7_75t_SL U69259 ( .A(n59529), .B(n57196), .Y(n75236) );
  NOR2xp33_ASAP7_75t_SL U69260 ( .A(n59528), .B(n59585), .Y(n61870) );
  NOR2xp33_ASAP7_75t_SL U69261 ( .A(n59573), .B(n57197), .Y(n75224) );
  NAND2xp33_ASAP7_75t_SRAM U69262 ( .A(n59442), .B(n61488), .Y(n75326) );
  NOR2xp33_ASAP7_75t_SL U69263 ( .A(n60955), .B(n73971), .Y(n61488) );
  NOR2xp33_ASAP7_75t_SL U69264 ( .A(n59712), .B(n59183), .Y(n60955) );
  NOR4xp25_ASAP7_75t_SL U69265 ( .A(n61098), .B(n61723), .C(n61094), .D(n61728), .Y(n61638) );
  NOR2xp33_ASAP7_75t_SL U69266 ( .A(n59569), .B(n63571), .Y(n61728) );
  NOR2xp33_ASAP7_75t_SL U69267 ( .A(n59545), .B(n57196), .Y(n61094) );
  NOR2xp33_ASAP7_75t_SL U69268 ( .A(n59555), .B(n59585), .Y(n61723) );
  NOR2xp33_ASAP7_75t_SL U69269 ( .A(n59571), .B(n57197), .Y(n61098) );
  AOI211xp5_ASAP7_75t_SL U69270 ( .A1(n76749), .A2(n60951), .B(n60950), .C(
        n60949), .Y(n60952) );
  NOR2xp33_ASAP7_75t_SL U69271 ( .A(n59708), .B(n75233), .Y(n64221) );
  NOR2xp33_ASAP7_75t_SL U69272 ( .A(n59576), .B(n59585), .Y(n61873) );
  NOR2xp33_ASAP7_75t_SL U69273 ( .A(n59710), .B(n74776), .Y(n61507) );
  NOR2xp33_ASAP7_75t_SL U69274 ( .A(n59561), .B(n59585), .Y(n61878) );
  NOR2xp33_ASAP7_75t_SL U69275 ( .A(n63571), .B(n75710), .Y(n75708) );
  AOI211xp5_ASAP7_75t_SL U69276 ( .A1(n61492), .A2(n59443), .B(n62106), .C(
        n61883), .Y(n75349) );
  NOR2xp33_ASAP7_75t_SL U69277 ( .A(n59533), .B(n59585), .Y(n61883) );
  NOR2xp33_ASAP7_75t_SL U69278 ( .A(n59535), .B(n57196), .Y(n62106) );
  NOR2xp33_ASAP7_75t_SL U69279 ( .A(n59406), .B(n74806), .Y(n60933) );
  NAND2xp33_ASAP7_75t_SRAM U69280 ( .A(n60945), .B(n59530), .Y(n59406) );
  AOI31xp33_ASAP7_75t_SL U69281 ( .A1(n62760), .A2(n63125), .A3(n75378), .B(
        n60931), .Y(n60932) );
  NAND2xp33_ASAP7_75t_SRAM U69282 ( .A(n59568), .B(n59564), .Y(n60954) );
  NAND2xp33_ASAP7_75t_SRAM U69283 ( .A(n60919), .B(n64357), .Y(n61406) );
  AOI211xp5_ASAP7_75t_SL U69284 ( .A1(n60920), .A2(n61650), .B(n60916), .C(
        n61518), .Y(n60926) );
  NOR2xp33_ASAP7_75t_SL U69285 ( .A(n60818), .B(n60826), .Y(n77040) );
  NOR2xp33_ASAP7_75t_SL U69286 ( .A(n59493), .B(n61248), .Y(n68812) );
  NOR2xp33_ASAP7_75t_SL U69287 ( .A(n59493), .B(n61746), .Y(n61595) );
  NOR2xp33_ASAP7_75t_SL U69288 ( .A(n3071), .B(n61056), .Y(n60714) );
  AOI211xp5_ASAP7_75t_SL U69289 ( .A1(n59538), .A2(n59586), .B(n60679), .C(
        n62532), .Y(n62425) );
  NOR2xp33_ASAP7_75t_SL U69290 ( .A(n62762), .B(n57197), .Y(n62532) );
  NOR2xp33_ASAP7_75t_SL U69291 ( .A(n59709), .B(n62353), .Y(n61494) );
  NOR2xp33_ASAP7_75t_SL U69292 ( .A(n64301), .B(n63573), .Y(n60677) );
  NOR2xp33_ASAP7_75t_SL U69293 ( .A(n59535), .B(n59584), .Y(n63573) );
  NOR2xp33_ASAP7_75t_SL U69294 ( .A(n59531), .B(n63571), .Y(n64301) );
  NOR2xp33_ASAP7_75t_SL U69295 ( .A(n59533), .B(n57197), .Y(n64112) );
  NOR2xp33_ASAP7_75t_SL U69296 ( .A(n57377), .B(n57209), .Y(n60665) );
  NOR2xp33_ASAP7_75t_SL U69297 ( .A(n59537), .B(n75378), .Y(n60666) );
  NOR2xp33_ASAP7_75t_SL U69298 ( .A(n57377), .B(n57196), .Y(n64110) );
  NOR2xp33_ASAP7_75t_SL U69299 ( .A(n59563), .B(n63571), .Y(n64836) );
  NOR2xp33_ASAP7_75t_SL U69300 ( .A(n59561), .B(n57197), .Y(n60664) );
  NOR2xp33_ASAP7_75t_SL U69301 ( .A(n59577), .B(n59584), .Y(n64304) );
  NOR2xp33_ASAP7_75t_SL U69302 ( .A(n59708), .B(n62353), .Y(n61511) );
  NOR2xp33_ASAP7_75t_SL U69303 ( .A(n59567), .B(n57214), .Y(n73923) );
  NOR2xp33_ASAP7_75t_SL U69304 ( .A(n60945), .B(n60663), .Y(n61410) );
  NOR2xp33_ASAP7_75t_SL U69305 ( .A(n60662), .B(n61649), .Y(n60944) );
  NOR2xp33_ASAP7_75t_SL U69306 ( .A(n59569), .B(n57196), .Y(n62356) );
  AOI211xp5_ASAP7_75t_SL U69307 ( .A1(n61538), .A2(n60656), .B(n60652), .C(
        n60651), .Y(n60653) );
  NOR2xp33_ASAP7_75t_SL U69308 ( .A(n60642), .B(n60669), .Y(n62013) );
  NAND2xp33_ASAP7_75t_SRAM U69309 ( .A(n59183), .B(n59586), .Y(n60639) );
  NOR2xp33_ASAP7_75t_SL U69310 ( .A(n76486), .B(n61649), .Y(n61411) );
  NOR2xp33_ASAP7_75t_SL U69311 ( .A(n59530), .B(n57196), .Y(n64783) );
  NOR2xp33_ASAP7_75t_SL U69312 ( .A(n59528), .B(n57197), .Y(n75831) );
  NOR2xp33_ASAP7_75t_SL U69313 ( .A(n59529), .B(n59584), .Y(n64838) );
  NOR2xp33_ASAP7_75t_SL U69314 ( .A(n59579), .B(n63571), .Y(n75482) );
  NOR2xp33_ASAP7_75t_SL U69315 ( .A(n59576), .B(n57197), .Y(n60637) );
  NOR2xp33_ASAP7_75t_SL U69316 ( .A(n59575), .B(n59584), .Y(n75706) );
  NOR2xp33_ASAP7_75t_SL U69317 ( .A(n59708), .B(n57214), .Y(n62359) );
  NOR2xp33_ASAP7_75t_SL U69318 ( .A(n60662), .B(n61206), .Y(n60963) );
  NOR2xp33_ASAP7_75t_SL U69319 ( .A(n60605), .B(n74806), .Y(n60613) );
  NOR2xp33_ASAP7_75t_SL U69320 ( .A(n59555), .B(n58343), .Y(n60916) );
  NAND2xp33_ASAP7_75t_SRAM U69321 ( .A(n76653), .B(n62606), .Y(n60609) );
  NOR2xp33_ASAP7_75t_SL U69322 ( .A(n60603), .B(n60602), .Y(n61519) );
  NOR2xp33_ASAP7_75t_SL U69323 ( .A(n59530), .B(n74806), .Y(n60602) );
  NAND2xp33_ASAP7_75t_SRAM U69324 ( .A(n60601), .B(n66241), .Y(n74806) );
  NOR2xp33_ASAP7_75t_SL U69325 ( .A(n57641), .B(n57639), .Y(n60962) );
  NAND2xp33_ASAP7_75t_SRAM U69326 ( .A(n61242), .B(n61243), .Y(n61746) );
  OR2x2_ASAP7_75t_SL U69327 ( .A(n60558), .B(n60557), .Y(n76717) );
  NOR2xp33_ASAP7_75t_SL U69328 ( .A(n61242), .B(n75561), .Y(n61753) );
  NOR2xp33_ASAP7_75t_SL U69329 ( .A(n77931), .B(n77851), .Y(n60538) );
  NOR4xp25_ASAP7_75t_SL U69330 ( .A(n66239), .B(n60616), .C(n74005), .D(n60537), .Y(n60539) );
  NOR4xp25_ASAP7_75t_SL U69331 ( .A(dbg_adr_i[16]), .B(n78448), .C(n78449), 
        .D(n78450), .Y(n60540) );
  NOR2xp33_ASAP7_75t_SL U69332 ( .A(dbg_adr_i[21]), .B(dbg_adr_i[22]), .Y(
        n78442) );
  NOR2xp33_ASAP7_75t_SL U69333 ( .A(dbg_adr_i[19]), .B(dbg_adr_i[20]), .Y(
        n78443) );
  NOR2xp33_ASAP7_75t_SL U69334 ( .A(dbg_adr_i[25]), .B(dbg_adr_i[26]), .Y(
        n78444) );
  NOR2xp33_ASAP7_75t_SL U69335 ( .A(dbg_adr_i[23]), .B(dbg_adr_i[24]), .Y(
        n78445) );
  NOR2xp33_ASAP7_75t_SL U69336 ( .A(dbg_adr_i[30]), .B(dbg_adr_i[31]), .Y(
        n78446) );
  NOR2xp33_ASAP7_75t_SL U69337 ( .A(dbg_adr_i[27]), .B(dbg_adr_i[28]), .Y(
        n78447) );
  NOR4xp25_ASAP7_75t_SL U69338 ( .A(dbg_adr_i[18]), .B(dbg_adr_i[29]), .C(
        dbg_adr_i[17]), .D(n78439), .Y(n60541) );
  NOR2xp33_ASAP7_75t_SL U69339 ( .A(n74251), .B(n74267), .Y(n2871) );
  NOR4xp25_ASAP7_75t_SL U69340 ( .A(n51955), .B(n73841), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_addsub_s_fract_o_6_), .D(n73840), 
        .Y(n73842) );
  NOR2xp33_ASAP7_75t_SL U69341 ( .A(n73470), .B(n73469), .Y(n73474) );
  NOR2xp33_ASAP7_75t_SL U69342 ( .A(n73368), .B(n73362), .Y(n78221) );
  NOR2xp33_ASAP7_75t_SL U69343 ( .A(n73411), .B(n73410), .Y(n73412) );
  NOR2xp33_ASAP7_75t_SL U69344 ( .A(n73369), .B(n73368), .Y(n73370) );
  NOR2xp33_ASAP7_75t_SL U69345 ( .A(n73361), .B(n73360), .Y(n73368) );
  NOR2xp33_ASAP7_75t_SL U69346 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[22]), .B(
        n74502), .Y(n73336) );
  NOR2xp33_ASAP7_75t_SL U69347 ( .A(n73312), .B(n58284), .Y(n73310) );
  NOR2xp33_ASAP7_75t_SL U69348 ( .A(n73258), .B(n58284), .Y(n73262) );
  NOR2xp33_ASAP7_75t_SL U69349 ( .A(n73241), .B(n59631), .Y(n73242) );
  NOR2xp33_ASAP7_75t_SL U69350 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[0]), .B(
        n74502), .Y(n73232) );
  NOR2xp33_ASAP7_75t_SL U69351 ( .A(n73219), .B(n73382), .Y(n73216) );
  NOR2xp33_ASAP7_75t_SL U69352 ( .A(n73209), .B(n58284), .Y(n73210) );
  NOR2xp33_ASAP7_75t_SL U69353 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[8]), .B(
        n74502), .Y(n73213) );
  NOR2xp33_ASAP7_75t_SL U69354 ( .A(n73194), .B(n73382), .Y(n73196) );
  NOR2xp33_ASAP7_75t_SL U69355 ( .A(n73191), .B(n59630), .Y(n73189) );
  NOR2xp33_ASAP7_75t_SL U69356 ( .A(n73193), .B(n73382), .Y(n73190) );
  NOR2xp33_ASAP7_75t_SL U69357 ( .A(n73434), .B(n73433), .Y(n73176) );
  NAND2xp33_ASAP7_75t_SRAM U69358 ( .A(n73171), .B(n74502), .Y(n73173) );
  NOR2xp33_ASAP7_75t_SL U69359 ( .A(n73171), .B(n73382), .Y(n73170) );
  NOR2xp33_ASAP7_75t_SL U69360 ( .A(n73148), .B(n58284), .Y(n73149) );
  NOR2xp33_ASAP7_75t_SL U69361 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[15]), .B(
        n74502), .Y(n73152) );
  NOR2xp33_ASAP7_75t_SL U69362 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[16]), .B(
        n59525), .Y(n73126) );
  NOR2xp33_ASAP7_75t_SL U69363 ( .A(n73115), .B(n58284), .Y(n73113) );
  NOR2xp33_ASAP7_75t_SL U69364 ( .A(n78328), .B(n73853), .Y(n73852) );
  NOR4xp25_ASAP7_75t_SL U69365 ( .A(n73087), .B(n73134), .C(n73086), .D(n73085), .Y(n73091) );
  AOI211xp5_ASAP7_75t_SL U69366 ( .A1(n73054), .A2(n73053), .B(n73052), .C(
        n73208), .Y(n73055) );
  AOI211xp5_ASAP7_75t_SL U69367 ( .A1(n76926), .A2(n63954), .B(n63717), .C(
        n63716), .Y(n63728) );
  NOR2xp33_ASAP7_75t_SL U69368 ( .A(or1200_cpu_or1200_except_n422), .B(n63715), 
        .Y(n63716) );
  AOI211xp5_ASAP7_75t_SL U69369 ( .A1(n76926), .A2(n64011), .B(n63927), .C(
        n63926), .Y(n63929) );
  NOR2xp33_ASAP7_75t_SL U69370 ( .A(or1200_cpu_spr_dat_ppc[17]), .B(n63715), 
        .Y(n63926) );
  AOI211xp5_ASAP7_75t_SL U69371 ( .A1(n76926), .A2(n64015), .B(n63922), .C(
        n63921), .Y(n63924) );
  NOR2xp33_ASAP7_75t_SL U69372 ( .A(or1200_cpu_spr_dat_ppc[19]), .B(n63715), 
        .Y(n63921) );
  AOI211xp5_ASAP7_75t_SL U69373 ( .A1(n76926), .A2(n64006), .B(n63932), .C(
        n63931), .Y(n63934) );
  NOR2xp33_ASAP7_75t_SL U69374 ( .A(or1200_cpu_or1200_except_n440), .B(n63715), 
        .Y(n63931) );
  NOR2xp33_ASAP7_75t_SL U69375 ( .A(n74360), .B(n74503), .Y(n74364) );
  AOI211xp5_ASAP7_75t_SL U69376 ( .A1(n76926), .A2(n63960), .B(n63959), .C(
        n63958), .Y(n63962) );
  NOR2xp33_ASAP7_75t_SL U69377 ( .A(or1200_cpu_or1200_except_n431), .B(n63715), 
        .Y(n63958) );
  NOR2xp33_ASAP7_75t_SL U69378 ( .A(n63721), .B(n69352), .Y(n77248) );
  AOI211xp5_ASAP7_75t_SL U69379 ( .A1(n76926), .A2(n63949), .B(n63948), .C(
        n63947), .Y(n63951) );
  NOR2xp33_ASAP7_75t_SL U69380 ( .A(or1200_cpu_or1200_except_n428), .B(n63715), 
        .Y(n63947) );
  AOI211xp5_ASAP7_75t_SL U69381 ( .A1(n74937), .A2(n74940), .B(n63709), .C(
        n63708), .Y(n63711) );
  AOI211xp5_ASAP7_75t_SL U69382 ( .A1(n63719), .A2(
        or1200_cpu_or1200_except_n565), .B(n77208), .C(n74924), .Y(n63709) );
  NOR2xp33_ASAP7_75t_SL U69383 ( .A(n76542), .B(n63712), .Y(n74940) );
  NOR2xp33_ASAP7_75t_SL U69384 ( .A(n76663), .B(n57170), .Y(n63704) );
  NOR2xp33_ASAP7_75t_SL U69385 ( .A(n63702), .B(n63701), .Y(n63718) );
  NOR2xp33_ASAP7_75t_SL U69386 ( .A(n62007), .B(n57072), .Y(n62072) );
  NOR2xp33_ASAP7_75t_SL U69387 ( .A(n61140), .B(n60351), .Y(n60490) );
  NOR2xp33_ASAP7_75t_SL U69388 ( .A(n2596), .B(n2814), .Y(n60343) );
  NOR2xp33_ASAP7_75t_SL U69389 ( .A(n74510), .B(n74509), .Y(n1522) );
  AOI211xp5_ASAP7_75t_SL U69390 ( .A1(n74508), .A2(n74507), .B(n74506), .C(
        n74505), .Y(n74509) );
  AOI31xp33_ASAP7_75t_SL U69391 ( .A1(n74502), .A2(n74828), .A3(n74501), .B(
        n74513), .Y(n74511) );
  AOI31xp33_ASAP7_75t_SL U69392 ( .A1(n74500), .A2(n74499), .A3(n74498), .B(
        n74497), .Y(n74513) );
  NOR2xp33_ASAP7_75t_SL U69393 ( .A(n74257), .B(n74254), .Y(n74263) );
  NOR4xp25_ASAP7_75t_SL U69394 ( .A(n77537), .B(n2616), .C(n2464), .D(n60358), 
        .Y(n60359) );
  NOR2xp33_ASAP7_75t_SL U69395 ( .A(n76638), .B(n76637), .Y(n76695) );
  NOR2xp33_ASAP7_75t_SL U69396 ( .A(n77990), .B(n77991), .Y(n77987) );
  NOR2xp33_ASAP7_75t_SL U69397 ( .A(n76995), .B(n76996), .Y(n76994) );
  NOR2xp33_ASAP7_75t_SL U69398 ( .A(n76611), .B(n76862), .Y(n76996) );
  NAND2xp33_ASAP7_75t_SRAM U69399 ( .A(n76204), .B(n76203), .Y(n76995) );
  NOR2xp33_ASAP7_75t_SL U69400 ( .A(n74241), .B(n74254), .Y(n74244) );
  NOR2xp33_ASAP7_75t_SL U69401 ( .A(n60337), .B(n77834), .Y(n60336) );
  AND2x2_ASAP7_75t_SL U69402 ( .A(n57144), .B(n77459), .Y(n62000) );
  NOR2xp33_ASAP7_75t_SL U69403 ( .A(n75779), .B(n77990), .Y(n76549) );
  NOR2xp33_ASAP7_75t_SL U69404 ( .A(n76229), .B(n76228), .Y(n78138) );
  NOR2xp33_ASAP7_75t_SL U69405 ( .A(n77223), .B(n78149), .Y(n78155) );
  NOR2xp33_ASAP7_75t_SL U69406 ( .A(n74737), .B(n74503), .Y(n74306) );
  AOI211xp5_ASAP7_75t_SL U69407 ( .A1(n76494), .A2(n76493), .B(n76492), .C(
        n76491), .Y(n76496) );
  NOR4xp25_ASAP7_75t_SL U69408 ( .A(n76470), .B(n76469), .C(n76468), .D(n76467), .Y(n76471) );
  NOR2xp33_ASAP7_75t_SL U69409 ( .A(n76363), .B(n76357), .Y(n76463) );
  NOR4xp25_ASAP7_75t_SL U69410 ( .A(n76456), .B(n76455), .C(n76454), .D(n76453), .Y(n76457) );
  NOR2xp33_ASAP7_75t_SL U69411 ( .A(n76441), .B(n76440), .Y(n76458) );
  NOR2xp33_ASAP7_75t_SL U69412 ( .A(n73976), .B(n76353), .Y(n76438) );
  NAND2xp33_ASAP7_75t_SRAM U69413 ( .A(n74798), .B(n53229), .Y(n76428) );
  NOR2xp33_ASAP7_75t_SL U69414 ( .A(n76409), .B(n53229), .Y(n76473) );
  NOR2xp33_ASAP7_75t_SL U69415 ( .A(n76387), .B(n76372), .Y(n76373) );
  NOR2xp33_ASAP7_75t_SL U69416 ( .A(n76358), .B(n76357), .Y(n76359) );
  NAND2xp33_ASAP7_75t_SRAM U69417 ( .A(n59564), .B(n59443), .Y(n76350) );
  NAND2xp33_ASAP7_75t_SRAM U69418 ( .A(n59442), .B(n59183), .Y(n60980) );
  NOR2xp33_ASAP7_75t_SL U69419 ( .A(n76346), .B(n76345), .Y(n76347) );
  NOR2xp33_ASAP7_75t_SL U69420 ( .A(n59529), .B(n59576), .Y(n74800) );
  AOI211xp5_ASAP7_75t_SL U69421 ( .A1(n76325), .A2(n76324), .B(n2069), .C(
        n76323), .Y(n76328) );
  NAND2xp33_ASAP7_75t_SRAM U69422 ( .A(n59548), .B(n75832), .Y(n76342) );
  NOR2xp33_ASAP7_75t_SL U69423 ( .A(n59548), .B(n75832), .Y(n74018) );
  NOR2xp33_ASAP7_75t_SL U69424 ( .A(n1588), .B(n64241), .Y(n74016) );
  NOR2xp33_ASAP7_75t_SL U69425 ( .A(n57068), .B(n74776), .Y(n74017) );
  NOR2xp33_ASAP7_75t_SL U69426 ( .A(n59547), .B(n75628), .Y(n76406) );
  AOI211xp5_ASAP7_75t_SL U69427 ( .A1(n59561), .A2(n74799), .B(n74011), .C(
        n74010), .Y(n76400) );
  NOR2xp33_ASAP7_75t_SL U69428 ( .A(n59536), .B(n74005), .Y(n74006) );
  NOR2xp33_ASAP7_75t_SL U69429 ( .A(n59536), .B(n75378), .Y(n75318) );
  NAND2xp33_ASAP7_75t_SRAM U69430 ( .A(n59546), .B(n57209), .Y(n74008) );
  NAND2xp33_ASAP7_75t_SRAM U69431 ( .A(n57377), .B(n77717), .Y(n74013) );
  NOR2xp33_ASAP7_75t_SL U69432 ( .A(n74007), .B(n76395), .Y(n74000) );
  NAND2xp33_ASAP7_75t_SRAM U69433 ( .A(n57312), .B(n63251), .Y(n73999) );
  NAND2xp33_ASAP7_75t_SRAM U69434 ( .A(n59536), .B(n75378), .Y(n76449) );
  NAND2xp33_ASAP7_75t_SRAM U69435 ( .A(n59532), .B(n76874), .Y(n74004) );
  NOR2xp33_ASAP7_75t_SL U69436 ( .A(n57377), .B(n77717), .Y(n74007) );
  NAND2xp33_ASAP7_75t_SRAM U69437 ( .A(n59537), .B(n77709), .Y(n73994) );
  NOR2xp33_ASAP7_75t_SL U69438 ( .A(n77064), .B(n76466), .Y(n73995) );
  NOR2xp33_ASAP7_75t_SL U69439 ( .A(n77063), .B(n76465), .Y(n76378) );
  NOR2xp33_ASAP7_75t_SL U69440 ( .A(n59551), .B(n57210), .Y(n77064) );
  NAND2xp33_ASAP7_75t_SRAM U69441 ( .A(n59538), .B(n77701), .Y(n76381) );
  NAND2xp33_ASAP7_75t_SRAM U69442 ( .A(n59570), .B(n59387), .Y(n73991) );
  NOR2xp33_ASAP7_75t_SL U69443 ( .A(n76444), .B(n73987), .Y(n73988) );
  NAND2xp33_ASAP7_75t_SRAM U69444 ( .A(n59541), .B(n62738), .Y(n73986) );
  NAND2xp33_ASAP7_75t_SRAM U69445 ( .A(n59540), .B(n57219), .Y(n76451) );
  NAND2xp33_ASAP7_75t_SRAM U69446 ( .A(n59542), .B(n77696), .Y(n73985) );
  NAND2xp33_ASAP7_75t_SRAM U69447 ( .A(n59569), .B(n56954), .Y(n76445) );
  NAND2xp33_ASAP7_75t_SRAM U69448 ( .A(n59555), .B(n78003), .Y(n73980) );
  NOR2xp33_ASAP7_75t_SL U69449 ( .A(n59545), .B(n78004), .Y(n76357) );
  NAND2xp33_ASAP7_75t_SRAM U69450 ( .A(n59559), .B(n78005), .Y(n73983) );
  NOR2xp33_ASAP7_75t_SL U69451 ( .A(n73975), .B(n76353), .Y(n76351) );
  NOR2xp33_ASAP7_75t_SL U69452 ( .A(n59558), .B(n59079), .Y(n76353) );
  NOR2xp33_ASAP7_75t_SL U69453 ( .A(n59708), .B(n53316), .Y(n73975) );
  NOR2xp33_ASAP7_75t_SL U69454 ( .A(n59557), .B(n57214), .Y(n73976) );
  NOR2xp33_ASAP7_75t_SL U69455 ( .A(n59568), .B(n59709), .Y(n73974) );
  NAND2xp33_ASAP7_75t_SRAM U69456 ( .A(n59443), .B(n73971), .Y(n73972) );
  NOR4xp25_ASAP7_75t_SL U69457 ( .A(n76389), .B(n73987), .C(n76374), .D(n76444), .Y(n74003) );
  NOR2xp33_ASAP7_75t_SL U69458 ( .A(n59540), .B(n57219), .Y(n76444) );
  NAND2xp33_ASAP7_75t_SRAM U69459 ( .A(n59581), .B(n77278), .Y(n76366) );
  NAND2xp33_ASAP7_75t_SRAM U69460 ( .A(n59556), .B(n76627), .Y(n73970) );
  NOR2xp33_ASAP7_75t_SL U69461 ( .A(n59560), .B(n57213), .Y(n73969) );
  NOR2xp33_ASAP7_75t_SL U69462 ( .A(n59572), .B(n77705), .Y(n77063) );
  NOR2xp33_ASAP7_75t_SL U69463 ( .A(n59538), .B(n77701), .Y(n73990) );
  NOR2xp33_ASAP7_75t_SL U69464 ( .A(n59570), .B(n59387), .Y(n73968) );
  NOR2xp33_ASAP7_75t_SL U69465 ( .A(n73967), .B(n76383), .Y(n73989) );
  NOR2xp33_ASAP7_75t_SL U69466 ( .A(n59541), .B(n62738), .Y(n76383) );
  NOR2xp33_ASAP7_75t_SL U69467 ( .A(n59542), .B(n77696), .Y(n73967) );
  NAND2xp33_ASAP7_75t_SRAM U69468 ( .A(n59554), .B(n76653), .Y(n76442) );
  NOR2xp33_ASAP7_75t_SL U69469 ( .A(n59530), .B(n77730), .Y(n73966) );
  NAND2xp33_ASAP7_75t_SRAM U69470 ( .A(n59547), .B(n75628), .Y(n76334) );
  NOR2xp33_ASAP7_75t_SL U69471 ( .A(n59550), .B(n75740), .Y(n75720) );
  NOR2xp33_ASAP7_75t_SL U69472 ( .A(n59549), .B(n57215), .Y(n76333) );
  NOR4xp25_ASAP7_75t_SL U69473 ( .A(n76314), .B(n76313), .C(n76312), .D(n76311), .Y(n76316) );
  AOI211xp5_ASAP7_75t_SL U69474 ( .A1(n76306), .A2(n76305), .B(n76304), .C(
        n76303), .Y(n76308) );
  NOR4xp25_ASAP7_75t_SL U69475 ( .A(n76299), .B(n76804), .C(n76298), .D(n76297), .Y(n76301) );
  NOR2xp33_ASAP7_75t_SL U69476 ( .A(n76284), .B(n76287), .Y(n76285) );
  NOR2xp33_ASAP7_75t_SL U69477 ( .A(n76279), .B(n76278), .Y(n76287) );
  NOR2xp33_ASAP7_75t_SL U69478 ( .A(n64271), .B(n64270), .Y(n64272) );
  NOR2xp33_ASAP7_75t_SL U69479 ( .A(n76274), .B(n76273), .Y(n76310) );
  NOR2xp33_ASAP7_75t_SL U69480 ( .A(n53455), .B(n57183), .Y(n61977) );
  NOR2xp33_ASAP7_75t_SL U69481 ( .A(n59530), .B(n61972), .Y(n64192) );
  XNOR2xp5_ASAP7_75t_SL U69482 ( .A(n59529), .B(n61971), .Y(n64191) );
  AOI211xp5_ASAP7_75t_SL U69483 ( .A1(n62084), .A2(n62085), .B(n64146), .C(
        n62074), .Y(n61948) );
  NOR2xp33_ASAP7_75t_SL U69484 ( .A(n75848), .B(n66288), .Y(n61979) );
  NOR2xp33_ASAP7_75t_SL U69485 ( .A(n59579), .B(n75476), .Y(n75517) );
  NOR2xp33_ASAP7_75t_SL U69486 ( .A(n57209), .B(n61947), .Y(n62088) );
  NOR2xp33_ASAP7_75t_SL U69487 ( .A(n62310), .B(n62307), .Y(n60773) );
  NOR2xp33_ASAP7_75t_SL U69488 ( .A(n59571), .B(n76280), .Y(n62310) );
  NOR2xp33_ASAP7_75t_SL U69489 ( .A(n76627), .B(n60770), .Y(n76288) );
  NOR2xp33_ASAP7_75t_SL U69490 ( .A(n59069), .B(n53455), .Y(n60769) );
  NOR2xp33_ASAP7_75t_SL U69491 ( .A(n53455), .B(n62588), .Y(n60760) );
  NOR2xp33_ASAP7_75t_SL U69492 ( .A(n59183), .B(n60756), .Y(n60757) );
  NOR2xp33_ASAP7_75t_SL U69493 ( .A(n60667), .B(n75478), .Y(n60752) );
  NAND2xp33_ASAP7_75t_SRAM U69494 ( .A(n74034), .B(n59080), .Y(n60667) );
  NOR2xp33_ASAP7_75t_SL U69495 ( .A(n59565), .B(n59712), .Y(n60844) );
  NOR2xp33_ASAP7_75t_SL U69496 ( .A(n59712), .B(n77242), .Y(n60754) );
  NOR2xp33_ASAP7_75t_SL U69497 ( .A(n59398), .B(n57196), .Y(n64776) );
  NOR2xp33_ASAP7_75t_SL U69498 ( .A(n60740), .B(n60739), .Y(n60741) );
  NOR2xp33_ASAP7_75t_SL U69499 ( .A(n62738), .B(n57120), .Y(n60740) );
  NOR2xp33_ASAP7_75t_SL U69500 ( .A(n57641), .B(n60735), .Y(n61953) );
  NOR2xp33_ASAP7_75t_SL U69501 ( .A(n53455), .B(n63129), .Y(n61919) );
  NOR2xp33_ASAP7_75t_SL U69502 ( .A(n63584), .B(n61929), .Y(n61928) );
  NOR2xp33_ASAP7_75t_SL U69503 ( .A(n53455), .B(n63653), .Y(n61929) );
  NOR2xp33_ASAP7_75t_SL U69504 ( .A(n59533), .B(n77713), .Y(n73998) );
  NOR2xp33_ASAP7_75t_SL U69505 ( .A(n78100), .B(n78101), .Y(n74084) );
  NOR2xp33_ASAP7_75t_SL U69506 ( .A(n78094), .B(n74082), .Y(n78101) );
  NOR2xp33_ASAP7_75t_SL U69507 ( .A(n69351), .B(n69350), .Y(n74943) );
  NOR2xp33_ASAP7_75t_SL U69508 ( .A(n73892), .B(n73885), .Y(n74249) );
  NOR2xp33_ASAP7_75t_SL U69509 ( .A(n74103), .B(n74102), .Y(n74101) );
  NOR2xp33_ASAP7_75t_SL U69510 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[4]), .B(
        n73877), .Y(n73878) );
  NOR2xp33_ASAP7_75t_SL U69511 ( .A(n73877), .B(n73869), .Y(n73876) );
  NOR2xp33_ASAP7_75t_SL U69512 ( .A(n73886), .B(n74255), .Y(n73885) );
  NOR2xp33_ASAP7_75t_SL U69513 ( .A(n60424), .B(n60423), .Y(n60425) );
  NOR2xp33_ASAP7_75t_SL U69514 ( .A(n847), .B(n77260), .Y(n63940) );
  AOI211xp5_ASAP7_75t_SL U69515 ( .A1(n63938), .A2(n77257), .B(n63937), .C(
        n63936), .Y(n63942) );
  NOR2xp33_ASAP7_75t_SL U69516 ( .A(n62477), .B(n59553), .Y(n62478) );
  NOR2xp33_ASAP7_75t_SL U69517 ( .A(n62476), .B(n63935), .Y(n62479) );
  NOR2xp33_ASAP7_75t_SL U69518 ( .A(n59553), .B(n57124), .Y(n63937) );
  NOR2xp33_ASAP7_75t_SL U69519 ( .A(n63935), .B(n57160), .Y(n63956) );
  NOR2xp33_ASAP7_75t_SL U69520 ( .A(n63736), .B(n63735), .Y(n76818) );
  NAND2xp33_ASAP7_75t_SRAM U69521 ( .A(n63729), .B(n77250), .Y(n76816) );
  NOR2xp33_ASAP7_75t_SL U69522 ( .A(n61175), .B(n77269), .Y(n76604) );
  AOI211xp5_ASAP7_75t_SL U69523 ( .A1(n77257), .A2(n61174), .B(n61173), .C(
        n61172), .Y(n61175) );
  NAND2xp33_ASAP7_75t_SRAM U69524 ( .A(n61164), .B(n77250), .Y(n76603) );
  AOI211xp5_ASAP7_75t_SL U69525 ( .A1(n57198), .A2(n74951), .B(n74950), .C(
        n74949), .Y(n74952) );
  AOI211xp5_ASAP7_75t_SL U69526 ( .A1(n63763), .A2(n77257), .B(n63691), .C(
        n63690), .Y(n63692) );
  NOR2xp33_ASAP7_75t_SL U69527 ( .A(n1099), .B(n57168), .Y(n63697) );
  NAND2xp33_ASAP7_75t_SRAM U69528 ( .A(n61275), .B(n77250), .Y(n61276) );
  AOI211xp5_ASAP7_75t_SL U69529 ( .A1(n77258), .A2(n77257), .B(n77256), .C(
        n77255), .Y(n77259) );
  NOR2xp33_ASAP7_75t_SL U69530 ( .A(n59544), .B(n57124), .Y(n77256) );
  NOR2xp33_ASAP7_75t_SL U69531 ( .A(n1044), .B(n57168), .Y(n77274) );
  NOR2xp33_ASAP7_75t_SL U69532 ( .A(n71346), .B(n71345), .Y(n71347) );
  XOR2xp5_ASAP7_75t_SL U69533 ( .A(n57336), .B(n53471), .Y(n76173) );
  NAND2xp33_ASAP7_75t_SRAM U69534 ( .A(n76845), .B(n77367), .Y(n78058) );
  NOR2xp33_ASAP7_75t_SL U69535 ( .A(or1200_immu_top_icpu_adr_default_8_), .B(
        n59703), .Y(n78055) );
  AOI211xp5_ASAP7_75t_SL U69536 ( .A1(n76831), .A2(n77257), .B(n76830), .C(
        n76829), .Y(n76832) );
  NOR2xp33_ASAP7_75t_SL U69537 ( .A(n76822), .B(n76821), .Y(n76823) );
  NAND2xp33_ASAP7_75t_SRAM U69538 ( .A(n59702), .B(n1073), .Y(n76824) );
  NOR2xp33_ASAP7_75t_SL U69539 ( .A(n4054), .B(n76837), .Y(n76843) );
  XOR2xp5_ASAP7_75t_SL U69540 ( .A(n68744), .B(n57341), .Y(n52060) );
  NOR4xp25_ASAP7_75t_SL U69541 ( .A(n61038), .B(n61037), .C(n61051), .D(n61036), .Y(n61039) );
  NOR2xp33_ASAP7_75t_SL U69542 ( .A(n71265), .B(n71264), .Y(n71296) );
  NOR2xp33_ASAP7_75t_SL U69543 ( .A(n70829), .B(n70830), .Y(n70860) );
  NOR2xp33_ASAP7_75t_SL U69544 ( .A(n70758), .B(n58328), .Y(n70761) );
  NOR2xp33_ASAP7_75t_SL U69545 ( .A(n71149), .B(n70885), .Y(n70770) );
  NOR2xp33_ASAP7_75t_SL U69546 ( .A(n71365), .B(n70846), .Y(n70848) );
  NOR2xp33_ASAP7_75t_SL U69547 ( .A(n70971), .B(n70970), .Y(n70972) );
  NOR2xp33_ASAP7_75t_SL U69548 ( .A(n70889), .B(n70888), .Y(n70907) );
  NOR2xp33_ASAP7_75t_SL U69549 ( .A(n71076), .B(n71162), .Y(n70883) );
  NOR2xp33_ASAP7_75t_SL U69550 ( .A(n78404), .B(n71413), .Y(n70990) );
  NOR2xp33_ASAP7_75t_SL U69551 ( .A(n71076), .B(n71148), .Y(n70865) );
  NOR2xp33_ASAP7_75t_SL U69552 ( .A(n70895), .B(n70864), .Y(n70866) );
  NOR2xp33_ASAP7_75t_SL U69553 ( .A(n71335), .B(n71146), .Y(n71152) );
  NOR2xp33_ASAP7_75t_SL U69554 ( .A(n71323), .B(n71322), .Y(n71346) );
  NOR2xp33_ASAP7_75t_SL U69555 ( .A(n70809), .B(n70993), .Y(n70810) );
  NOR2xp33_ASAP7_75t_SL U69556 ( .A(n70656), .B(n70655), .Y(n70657) );
  NOR2xp33_ASAP7_75t_SL U69557 ( .A(n75475), .B(n69334), .Y(n76834) );
  NOR2xp33_ASAP7_75t_SL U69558 ( .A(n60464), .B(n60463), .Y(n60465) );
  NOR2xp33_ASAP7_75t_SL U69559 ( .A(n60406), .B(or1200_cpu_or1200_if_if_bypass), .Y(n60459) );
  NOR2xp33_ASAP7_75t_SL U69560 ( .A(n3132), .B(n78440), .Y(n60464) );
  NOR2xp33_ASAP7_75t_SL U69561 ( .A(n60450), .B(n60451), .Y(n60441) );
  NOR2xp33_ASAP7_75t_SL U69562 ( .A(n77843), .B(n77363), .Y(n77365) );
  NOR2xp33_ASAP7_75t_SL U69563 ( .A(n77835), .B(n77836), .Y(n60443) );
  NOR2xp33_ASAP7_75t_SL U69564 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_2_), .Y(
        n72550) );
  NOR4xp25_ASAP7_75t_SL U69565 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_16_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_17_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_19_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_20_), .Y(
        n72551) );
  NOR4xp25_ASAP7_75t_SL U69566 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_10_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_11_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_13_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_14_), .Y(
        n72552) );
  NOR4xp25_ASAP7_75t_SL U69567 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_4_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_5_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_7_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_8_), .Y(
        n72553) );
  AOI211xp5_ASAP7_75t_SL U69568 ( .A1(n61583), .A2(n77257), .B(n61582), .C(
        n61581), .Y(n61584) );
  NOR2xp33_ASAP7_75t_SL U69569 ( .A(n62477), .B(n59558), .Y(n61579) );
  NOR2xp33_ASAP7_75t_SL U69570 ( .A(n62476), .B(n61578), .Y(n61580) );
  NOR2xp33_ASAP7_75t_SL U69571 ( .A(n59558), .B(n57124), .Y(n61582) );
  NOR2xp33_ASAP7_75t_SL U69572 ( .A(n61578), .B(n57160), .Y(n76581) );
  NOR2xp33_ASAP7_75t_SL U69573 ( .A(n68904), .B(n57086), .Y(n58684) );
  NOR2xp33_ASAP7_75t_SL U69574 ( .A(or1200_cpu_or1200_mult_mac_n20), .B(n57105), .Y(n76139) );
  NOR2xp33_ASAP7_75t_SL U69575 ( .A(n76135), .B(n76134), .Y(n76141) );
  NOR2xp33_ASAP7_75t_SL U69576 ( .A(or1200_cpu_or1200_mult_mac_n16), .B(n57105), .Y(n76154) );
  NOR2xp33_ASAP7_75t_SL U69577 ( .A(n76153), .B(n76152), .Y(n76155) );
  NOR2xp33_ASAP7_75t_SL U69578 ( .A(n76149), .B(n76159), .Y(n76153) );
  NOR2xp33_ASAP7_75t_SL U69579 ( .A(or1200_cpu_or1200_mult_mac_n50), .B(n57105), .Y(n76015) );
  NOR2xp33_ASAP7_75t_SL U69580 ( .A(n76047), .B(n76050), .Y(n76043) );
  NOR2xp33_ASAP7_75t_SL U69581 ( .A(n76034), .B(n76042), .Y(n76035) );
  NOR2xp33_ASAP7_75t_SL U69582 ( .A(n77340), .B(n77347), .Y(n77350) );
  NOR2xp33_ASAP7_75t_SL U69583 ( .A(n835), .B(n77799), .Y(n77509) );
  AOI211xp5_ASAP7_75t_SL U69584 ( .A1(n65220), .A2(n77257), .B(n60179), .C(
        n60178), .Y(n60180) );
  NOR2xp33_ASAP7_75t_SL U69585 ( .A(n62476), .B(n60175), .Y(n60177) );
  NOR2xp33_ASAP7_75t_SL U69586 ( .A(n1588), .B(n57124), .Y(n60179) );
  NOR2xp33_ASAP7_75t_SL U69587 ( .A(n60166), .B(n57160), .Y(n63984) );
  AOI211xp5_ASAP7_75t_SL U69588 ( .A1(n60162), .A2(n77257), .B(n60161), .C(
        n60160), .Y(n60163) );
  NOR2xp33_ASAP7_75t_SL U69589 ( .A(n62477), .B(n59552), .Y(n60158) );
  NOR2xp33_ASAP7_75t_SL U69590 ( .A(n62476), .B(n60166), .Y(n60159) );
  NOR2xp33_ASAP7_75t_SL U69591 ( .A(n59552), .B(n57124), .Y(n60161) );
  NOR2xp33_ASAP7_75t_SL U69592 ( .A(n60154), .B(n57160), .Y(n64096) );
  NOR2xp33_ASAP7_75t_SL U69593 ( .A(n928), .B(n57168), .Y(n60155) );
  NOR2xp33_ASAP7_75t_SL U69594 ( .A(n795), .B(n77260), .Y(n60148) );
  NOR2xp33_ASAP7_75t_SL U69595 ( .A(n60146), .B(n57160), .Y(n74961) );
  NOR2xp33_ASAP7_75t_SL U69596 ( .A(n803), .B(n77260), .Y(n60141) );
  AOI211xp5_ASAP7_75t_SL U69597 ( .A1(n60139), .A2(n77257), .B(n60138), .C(
        n60137), .Y(n60144) );
  NOR2xp33_ASAP7_75t_SL U69598 ( .A(n62477), .B(n59534), .Y(n60135) );
  NOR2xp33_ASAP7_75t_SL U69599 ( .A(n62476), .B(n60146), .Y(n60136) );
  NOR2xp33_ASAP7_75t_SL U69600 ( .A(n59534), .B(n57124), .Y(n60138) );
  NOR2xp33_ASAP7_75t_SL U69601 ( .A(n60134), .B(n57160), .Y(n63920) );
  AOI211xp5_ASAP7_75t_SL U69602 ( .A1(n64013), .A2(n77257), .B(n60129), .C(
        n60128), .Y(n60130) );
  NOR2xp33_ASAP7_75t_SL U69603 ( .A(n62477), .B(n59532), .Y(n60126) );
  NOR2xp33_ASAP7_75t_SL U69604 ( .A(n62476), .B(n60134), .Y(n60127) );
  NOR2xp33_ASAP7_75t_SL U69605 ( .A(n59532), .B(n57124), .Y(n60129) );
  NOR2xp33_ASAP7_75t_SL U69606 ( .A(n811), .B(n77260), .Y(n60115) );
  NOR2xp33_ASAP7_75t_SL U69607 ( .A(n60100), .B(n57160), .Y(n63987) );
  AOI211xp5_ASAP7_75t_SL U69608 ( .A1(n60095), .A2(n77257), .B(n60094), .C(
        n60093), .Y(n60096) );
  NOR2xp33_ASAP7_75t_SL U69609 ( .A(n62477), .B(n59551), .Y(n60091) );
  NOR2xp33_ASAP7_75t_SL U69610 ( .A(n62476), .B(n60100), .Y(n60092) );
  NOR2xp33_ASAP7_75t_SL U69611 ( .A(n59551), .B(n57124), .Y(n60094) );
  NOR2xp33_ASAP7_75t_SL U69612 ( .A(n60081), .B(n57160), .Y(n65191) );
  NOR2xp33_ASAP7_75t_SL U69613 ( .A(n955), .B(n57168), .Y(n60082) );
  AOI211xp5_ASAP7_75t_SL U69614 ( .A1(n75544), .A2(n77257), .B(n60075), .C(
        n60074), .Y(n60076) );
  NOR2xp33_ASAP7_75t_SL U69615 ( .A(n62477), .B(n59547), .Y(n60072) );
  NOR2xp33_ASAP7_75t_SL U69616 ( .A(n62476), .B(n60081), .Y(n60073) );
  NOR2xp33_ASAP7_75t_SL U69617 ( .A(or1200_cpu_or1200_except_n234), .B(n58547), 
        .Y(n60075) );
  NOR2xp33_ASAP7_75t_SL U69618 ( .A(n60069), .B(n57160), .Y(n64258) );
  NOR2xp33_ASAP7_75t_SL U69619 ( .A(n937), .B(n57168), .Y(n60070) );
  AOI211xp5_ASAP7_75t_SL U69620 ( .A1(n75418), .A2(n77257), .B(n60064), .C(
        n60063), .Y(n60065) );
  NOR2xp33_ASAP7_75t_SL U69621 ( .A(n62477), .B(n59546), .Y(n60061) );
  NOR2xp33_ASAP7_75t_SL U69622 ( .A(n62476), .B(n60069), .Y(n60062) );
  NOR2xp33_ASAP7_75t_SL U69623 ( .A(or1200_cpu_or1200_except_n230), .B(n58547), 
        .Y(n60064) );
  NOR2xp33_ASAP7_75t_SL U69624 ( .A(n946), .B(n57168), .Y(n60059) );
  NOR2xp33_ASAP7_75t_SL U69625 ( .A(n60052), .B(n57160), .Y(n63969) );
  AOI211xp5_ASAP7_75t_SL U69626 ( .A1(n63968), .A2(n77257), .B(n60047), .C(
        n60046), .Y(n60048) );
  NOR2xp33_ASAP7_75t_SL U69627 ( .A(n62477), .B(n59539), .Y(n60044) );
  NOR2xp33_ASAP7_75t_SL U69628 ( .A(n62476), .B(n60052), .Y(n60045) );
  NOR2xp33_ASAP7_75t_SL U69629 ( .A(n59539), .B(n57124), .Y(n60047) );
  AOI211xp5_ASAP7_75t_SL U69630 ( .A1(n57198), .A2(n75208), .B(n60011), .C(
        n60010), .Y(n60012) );
  NOR2xp33_ASAP7_75t_SL U69631 ( .A(n59549), .B(n57124), .Y(n60011) );
  AOI211xp5_ASAP7_75t_SL U69632 ( .A1(n59998), .A2(n77257), .B(n59997), .C(
        n59996), .Y(n59999) );
  NOR2xp33_ASAP7_75t_SL U69633 ( .A(n76019), .B(n76018), .Y(n76020) );
  NOR2xp33_ASAP7_75t_SL U69634 ( .A(n76128), .B(n76127), .Y(n76134) );
  NOR2xp33_ASAP7_75t_SL U69635 ( .A(n75959), .B(n75960), .Y(n76177) );
  NOR2xp33_ASAP7_75t_SL U69636 ( .A(n75942), .B(n75941), .Y(n75943) );
  NOR2xp33_ASAP7_75t_SL U69637 ( .A(n75909), .B(n75908), .Y(n76081) );
  NOR2xp33_ASAP7_75t_SL U69638 ( .A(n76065), .B(n75906), .Y(n75907) );
  NOR2xp33_ASAP7_75t_SL U69639 ( .A(n76003), .B(n76002), .Y(n76010) );
  NOR2xp33_ASAP7_75t_SL U69640 ( .A(n60513), .B(n78006), .Y(n60514) );
  NOR2xp33_ASAP7_75t_SL U69641 ( .A(n2721), .B(n78009), .Y(n60515) );
  NOR2xp33_ASAP7_75t_SL U69642 ( .A(n60520), .B(n78006), .Y(n60521) );
  NOR2xp33_ASAP7_75t_SL U69643 ( .A(n2717), .B(n78009), .Y(n60522) );
  NOR2xp33_ASAP7_75t_SL U69644 ( .A(n60450), .B(n60449), .Y(n60453) );
  NOR2xp33_ASAP7_75t_SL U69645 ( .A(n60448), .B(n77954), .Y(n60449) );
  NOR2xp33_ASAP7_75t_SL U69646 ( .A(n3134), .B(n78009), .Y(n60450) );
  NOR2xp33_ASAP7_75t_SL U69647 ( .A(n60434), .B(n78006), .Y(n60437) );
  NOR2xp33_ASAP7_75t_SL U69648 ( .A(n2703), .B(n78009), .Y(n77835) );
  OR2x2_ASAP7_75t_SL U69649 ( .A(n60310), .B(or1200_cpu_or1200_if_if_bypass), 
        .Y(n78009) );
  NOR2xp33_ASAP7_75t_SL U69650 ( .A(n60313), .B(n22057), .Y(n77358) );
  NOR2xp33_ASAP7_75t_SL U69651 ( .A(n60316), .B(n22057), .Y(n60321) );
  NAND2xp33_ASAP7_75t_SRAM U69652 ( .A(n62477), .B(dbg_dat_i[2]), .Y(n60261)
         );
  NOR2xp33_ASAP7_75t_SL U69653 ( .A(n60420), .B(n62149), .Y(n60309) );
  NOR2xp33_ASAP7_75t_SL U69654 ( .A(n2033), .B(n60219), .Y(n60220) );
  NOR2xp33_ASAP7_75t_SL U69655 ( .A(n60200), .B(n62002), .Y(n60201) );
  NOR2xp33_ASAP7_75t_SL U69656 ( .A(n75196), .B(n75191), .Y(n77174) );
  NOR2xp33_ASAP7_75t_SL U69657 ( .A(dwb_err_i), .B(dwb_rty_i), .Y(n59713) );
  NOR4xp25_ASAP7_75t_SL U69658 ( .A(n59845), .B(n59844), .C(n59843), .D(n76546), .Y(n59846) );
  NOR2xp33_ASAP7_75t_SL U69659 ( .A(n59840), .B(n59841), .Y(n59842) );
  NOR2xp33_ASAP7_75t_SL U69660 ( .A(dbg_adr_i[10]), .B(n78439), .Y(n59943) );
  NOR2xp33_ASAP7_75t_SL U69661 ( .A(dbg_adr_i[3]), .B(n78439), .Y(n59940) );
  NOR2xp33_ASAP7_75t_SL U69662 ( .A(dbg_adr_i[4]), .B(n78439), .Y(n59938) );
  NOR4xp25_ASAP7_75t_SL U69663 ( .A(dbg_adr_i[8]), .B(dbg_adr_i[7]), .C(
        dbg_adr_i[9]), .D(n78439), .Y(n59933) );
  NOR2xp33_ASAP7_75t_SL U69664 ( .A(dbg_adr_i[2]), .B(n78439), .Y(n59931) );
  NOR2xp33_ASAP7_75t_SL U69665 ( .A(dbg_adr_i[14]), .B(n78439), .Y(n59928) );
  NOR2xp33_ASAP7_75t_SL U69666 ( .A(dbg_adr_i[15]), .B(n78439), .Y(n59924) );
  NOR2xp33_ASAP7_75t_SL U69667 ( .A(dbg_adr_i[0]), .B(n78439), .Y(n59920) );
  NOR2xp33_ASAP7_75t_SL U69668 ( .A(n60421), .B(n60311), .Y(n69331) );
  NOR2xp33_ASAP7_75t_SL U69669 ( .A(iwb_err_i), .B(iwb_rty_i), .Y(n60272) );
  NOR2xp33_ASAP7_75t_SL U69670 ( .A(n58837), .B(n59449), .Y(n58836) );
  NOR2xp33_ASAP7_75t_SL U69671 ( .A(n58546), .B(n68686), .Y(n58837) );
  NOR2xp33_ASAP7_75t_SL U69672 ( .A(n68914), .B(n68913), .Y(n68918) );
  NOR2xp33_ASAP7_75t_SL U69673 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_17_), .B(n74864), 
        .Y(n74861) );
  AND4x1_ASAP7_75t_SL U69674 ( .A(n52491), .B(n52506), .C(n52504), .D(n52490), 
        .Y(n74914) );
  NOR2xp33_ASAP7_75t_SL U69675 ( .A(n74851), .B(n77171), .Y(n74852) );
  NOR2xp33_ASAP7_75t_SL U69676 ( .A(n76934), .B(n77171), .Y(n74216) );
  NOR2xp33_ASAP7_75t_SL U69677 ( .A(n76970), .B(n77171), .Y(n74873) );
  NOR2xp33_ASAP7_75t_SL U69678 ( .A(n76948), .B(n77171), .Y(n74843) );
  NOR4xp25_ASAP7_75t_SL U69679 ( .A(n76242), .B(n74898), .C(n74897), .D(n74896), .Y(n74910) );
  NOR2xp33_ASAP7_75t_SL U69680 ( .A(n74855), .B(n74885), .Y(n74882) );
  NOR2xp33_ASAP7_75t_SL U69681 ( .A(n76943), .B(n76950), .Y(n74850) );
  AOI211xp5_ASAP7_75t_SL U69682 ( .A1(n74209), .A2(n74208), .B(n74752), .C(
        n74207), .Y(n74210) );
  NOR2xp33_ASAP7_75t_SL U69683 ( .A(n74206), .B(n74205), .Y(n74207) );
  AOI211xp5_ASAP7_75t_SL U69684 ( .A1(n74209), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_1_), .B(n74752), .C(
        n74051), .Y(n74052) );
  NOR2xp33_ASAP7_75t_SL U69685 ( .A(n74050), .B(n74205), .Y(n74051) );
  AOI31xp33_ASAP7_75t_SL U69686 ( .A1(n74203), .A2(n74750), .A3(n74055), .B(
        n74054), .Y(n74057) );
  NOR2xp33_ASAP7_75t_SL U69687 ( .A(n74087), .B(n74190), .Y(n74096) );
  NOR2xp33_ASAP7_75t_SL U69688 ( .A(n76963), .B(n77171), .Y(n74859) );
  NOR2xp33_ASAP7_75t_SL U69689 ( .A(n68683), .B(n58745), .Y(n58744) );
  AOI211xp5_ASAP7_75t_SL U69690 ( .A1(n69229), .A2(n59449), .B(n59251), .C(
        n59250), .Y(n59249) );
  NOR2xp33_ASAP7_75t_SL U69691 ( .A(n69237), .B(n59449), .Y(n59250) );
  NOR2xp33_ASAP7_75t_SL U69692 ( .A(n58887), .B(n59346), .Y(n59341) );
  NOR2xp33_ASAP7_75t_SL U69693 ( .A(n58827), .B(n68662), .Y(n59212) );
  NOR2xp33_ASAP7_75t_SL U69694 ( .A(n69145), .B(n57369), .Y(n69146) );
  AOI31xp33_ASAP7_75t_SL U69695 ( .A1(n68657), .A2(n68656), .A3(n57376), .B(
        n68655), .Y(n68658) );
  NOR2xp33_ASAP7_75t_SL U69696 ( .A(n68654), .B(n69300), .Y(n68659) );
  NOR2xp33_ASAP7_75t_SL U69697 ( .A(n68712), .B(n57474), .Y(n68715) );
  NOR2xp33_ASAP7_75t_SL U69698 ( .A(n75100), .B(n75099), .Y(n75101) );
  NOR2xp33_ASAP7_75t_SL U69699 ( .A(n69119), .B(n58895), .Y(n69098) );
  NOR2xp33_ASAP7_75t_SL U69700 ( .A(n58887), .B(n58886), .Y(n68968) );
  NOR2xp33_ASAP7_75t_SL U69701 ( .A(n68973), .B(n68835), .Y(n68838) );
  NAND2xp33_ASAP7_75t_SRAM U69702 ( .A(n69008), .B(n69014), .Y(n69009) );
  NOR2xp33_ASAP7_75t_SL U69703 ( .A(n57131), .B(n69011), .Y(n69010) );
  NOR2xp33_ASAP7_75t_SL U69704 ( .A(n59383), .B(n69011), .Y(n69014) );
  NOR2xp33_ASAP7_75t_SL U69705 ( .A(n69005), .B(n57475), .Y(n69015) );
  NOR2xp33_ASAP7_75t_SL U69706 ( .A(n69008), .B(n57131), .Y(n69007) );
  NAND3xp33_ASAP7_75t_SL U69707 ( .A(n58189), .B(n58770), .C(n58768), .Y(
        n52003) );
  NOR2xp33_ASAP7_75t_SL U69708 ( .A(n58771), .B(n68710), .Y(n58770) );
  NOR2xp33_ASAP7_75t_SL U69709 ( .A(n68705), .B(n68704), .Y(n68706) );
  NOR2xp33_ASAP7_75t_SL U69710 ( .A(n74558), .B(n58772), .Y(n58771) );
  NOR2xp33_ASAP7_75t_SL U69711 ( .A(n75280), .B(n57474), .Y(n75282) );
  NOR2xp33_ASAP7_75t_SL U69712 ( .A(n75111), .B(n75110), .Y(n75113) );
  NOR2xp33_ASAP7_75t_SL U69713 ( .A(n68860), .B(n68850), .Y(n68577) );
  NOR2xp33_ASAP7_75t_SL U69714 ( .A(n66898), .B(n66897), .Y(n66900) );
  NOR2xp33_ASAP7_75t_SL U69715 ( .A(n67154), .B(n67139), .Y(n58679) );
  XNOR2xp5_ASAP7_75t_SL U69716 ( .A(n57292), .B(n59659), .Y(n66852) );
  XOR2xp5_ASAP7_75t_SL U69717 ( .A(n57107), .B(n57322), .Y(n58521) );
  NOR2xp33_ASAP7_75t_SL U69718 ( .A(n56985), .B(n59636), .Y(n66699) );
  NOR2xp33_ASAP7_75t_SL U69719 ( .A(n67134), .B(n67135), .Y(n58680) );
  NOR2xp33_ASAP7_75t_SL U69720 ( .A(n59454), .B(n67029), .Y(n67035) );
  NOR2xp33_ASAP7_75t_SL U69721 ( .A(n66860), .B(n59649), .Y(n66861) );
  NOR2xp33_ASAP7_75t_SL U69722 ( .A(n66876), .B(n75032), .Y(n66877) );
  NOR2xp33_ASAP7_75t_SL U69723 ( .A(n59641), .B(n57662), .Y(n66878) );
  NOR2xp33_ASAP7_75t_SL U69724 ( .A(n67432), .B(n67712), .Y(n66879) );
  NOR2xp33_ASAP7_75t_SL U69725 ( .A(n57107), .B(n57405), .Y(n66996) );
  NOR2xp33_ASAP7_75t_SL U69726 ( .A(n58919), .B(n59640), .Y(n66998) );
  NOR2xp33_ASAP7_75t_SL U69727 ( .A(n59660), .B(n67712), .Y(n66999) );
  XNOR2xp5_ASAP7_75t_SL U69728 ( .A(n57292), .B(n58753), .Y(n58794) );
  NOR2xp33_ASAP7_75t_SL U69729 ( .A(n67432), .B(n75644), .Y(n66697) );
  NOR2xp33_ASAP7_75t_SL U69730 ( .A(n59649), .B(n66413), .Y(n66324) );
  XNOR2xp5_ASAP7_75t_SL U69731 ( .A(n58919), .B(n75644), .Y(n66876) );
  NOR2xp33_ASAP7_75t_SL U69732 ( .A(n66462), .B(n75032), .Y(n66463) );
  XNOR2xp5_ASAP7_75t_SL U69733 ( .A(n75644), .B(n59659), .Y(n66462) );
  NOR2xp33_ASAP7_75t_SL U69734 ( .A(n66365), .B(n57494), .Y(n66370) );
  NOR2xp33_ASAP7_75t_SL U69735 ( .A(n67276), .B(n59639), .Y(n66458) );
  NOR2xp33_ASAP7_75t_SL U69736 ( .A(n58861), .B(n59637), .Y(n66459) );
  NOR2xp33_ASAP7_75t_SL U69737 ( .A(n59641), .B(n67383), .Y(n66454) );
  NOR2xp33_ASAP7_75t_SL U69738 ( .A(n57491), .B(n59664), .Y(n66483) );
  NOR2xp33_ASAP7_75t_SL U69739 ( .A(n59600), .B(n59662), .Y(n66378) );
  NOR2xp33_ASAP7_75t_SL U69740 ( .A(n67911), .B(n66413), .Y(n66416) );
  XNOR2xp5_ASAP7_75t_SL U69741 ( .A(n57311), .B(n57436), .Y(n66351) );
  NOR2xp33_ASAP7_75t_SL U69742 ( .A(n59440), .B(n66467), .Y(n66354) );
  NOR2xp33_ASAP7_75t_SL U69743 ( .A(n57491), .B(n75947), .Y(n66353) );
  NOR2xp33_ASAP7_75t_SL U69744 ( .A(n59475), .B(n57405), .Y(n66357) );
  NOR2xp33_ASAP7_75t_SL U69745 ( .A(n58753), .B(n67712), .Y(n66360) );
  NOR2xp33_ASAP7_75t_SL U69746 ( .A(n59637), .B(n66758), .Y(n66267) );
  NOR2xp33_ASAP7_75t_SL U69747 ( .A(n59639), .B(n66800), .Y(n66268) );
  NOR2xp33_ASAP7_75t_SL U69748 ( .A(n59516), .B(n75644), .Y(n66255) );
  NOR2xp33_ASAP7_75t_SL U69749 ( .A(n68612), .B(n68611), .Y(n68613) );
  NAND2xp33_ASAP7_75t_SRAM U69750 ( .A(n67881), .B(n75947), .Y(n66538) );
  NOR2xp33_ASAP7_75t_SL U69751 ( .A(n67365), .B(n57405), .Y(n66539) );
  XOR2xp5_ASAP7_75t_SL U69752 ( .A(n59518), .B(n59664), .Y(n66568) );
  NOR2xp33_ASAP7_75t_SL U69753 ( .A(n75899), .B(n75467), .Y(n66547) );
  XNOR2xp5_ASAP7_75t_SL U69754 ( .A(n59518), .B(n57336), .Y(n66284) );
  NOR2xp33_ASAP7_75t_SL U69755 ( .A(n63313), .B(n63292), .Y(n62911) );
  NOR2xp33_ASAP7_75t_SL U69756 ( .A(n59476), .B(n67638), .Y(n62897) );
  NAND2xp33_ASAP7_75t_SRAM U69757 ( .A(n67424), .B(n63271), .Y(n63259) );
  NOR2xp33_ASAP7_75t_SL U69758 ( .A(n62891), .B(n62890), .Y(n62892) );
  AOI211xp5_ASAP7_75t_SL U69759 ( .A1(n59656), .A2(n68097), .B(n62887), .C(
        n57178), .Y(n63280) );
  NOR2xp33_ASAP7_75t_SL U69760 ( .A(n58701), .B(n68090), .Y(n62881) );
  NOR2xp33_ASAP7_75t_SL U69761 ( .A(n67228), .B(n59509), .Y(n62874) );
  NOR2xp33_ASAP7_75t_SL U69762 ( .A(n62947), .B(n63370), .Y(n62913) );
  NOR2xp33_ASAP7_75t_SL U69763 ( .A(n59614), .B(n62822), .Y(n62830) );
  NOR2xp33_ASAP7_75t_SL U69764 ( .A(n75930), .B(n59618), .Y(n62803) );
  NOR2xp33_ASAP7_75t_SL U69765 ( .A(n59656), .B(n67536), .Y(n62845) );
  NOR2xp33_ASAP7_75t_SL U69766 ( .A(n57111), .B(n67535), .Y(n62846) );
  NOR2xp33_ASAP7_75t_SL U69767 ( .A(n75925), .B(n59618), .Y(n62842) );
  NOR2xp33_ASAP7_75t_SL U69768 ( .A(n63362), .B(n63363), .Y(n63045) );
  NOR2xp33_ASAP7_75t_SL U69769 ( .A(n59511), .B(n67918), .Y(n62817) );
  NOR2xp33_ASAP7_75t_SL U69770 ( .A(n64083), .B(n58701), .Y(n62818) );
  NOR2xp33_ASAP7_75t_SL U69771 ( .A(n59504), .B(n67463), .Y(n62819) );
  NOR2xp33_ASAP7_75t_SL U69772 ( .A(n62879), .B(n57097), .Y(n62795) );
  NOR2xp33_ASAP7_75t_SL U69773 ( .A(n57159), .B(n62794), .Y(n62796) );
  NOR2xp33_ASAP7_75t_SL U69774 ( .A(n62935), .B(n62934), .Y(n62936) );
  NOR2xp33_ASAP7_75t_SL U69775 ( .A(n75930), .B(n68090), .Y(n62836) );
  NOR2xp33_ASAP7_75t_SL U69776 ( .A(n57111), .B(n64489), .Y(n62939) );
  NOR2xp33_ASAP7_75t_SL U69777 ( .A(n62977), .B(n57362), .Y(n62941) );
  NOR2xp33_ASAP7_75t_SL U69778 ( .A(n59614), .B(n58701), .Y(n62983) );
  NOR2xp33_ASAP7_75t_SL U69779 ( .A(n59505), .B(n59511), .Y(n62984) );
  NAND3xp33_ASAP7_75t_SL U69780 ( .A(n58410), .B(n68079), .C(n62742), .Y(
        n59307) );
  NOR2xp33_ASAP7_75t_SL U69781 ( .A(n59505), .B(n59513), .Y(n62943) );
  NOR2xp33_ASAP7_75t_SL U69782 ( .A(n58931), .B(n67227), .Y(n58932) );
  NOR2xp33_ASAP7_75t_SL U69783 ( .A(n59609), .B(n62922), .Y(n62923) );
  NOR2xp33_ASAP7_75t_SL U69784 ( .A(n76028), .B(n68090), .Y(n62924) );
  NOR2xp33_ASAP7_75t_SL U69785 ( .A(n57159), .B(n62965), .Y(n62919) );
  NOR2xp33_ASAP7_75t_SL U69786 ( .A(n58440), .B(n59620), .Y(n62955) );
  NOR2xp33_ASAP7_75t_SL U69787 ( .A(n75927), .B(n67918), .Y(n62708) );
  NOR2xp33_ASAP7_75t_SL U69788 ( .A(n58440), .B(n59510), .Y(n62707) );
  XNOR2xp5_ASAP7_75t_SL U69789 ( .A(n63167), .B(n63165), .Y(n58945) );
  NOR2xp33_ASAP7_75t_SL U69790 ( .A(n53283), .B(n59504), .Y(n62603) );
  NOR2xp33_ASAP7_75t_SL U69791 ( .A(n67343), .B(n59615), .Y(n62980) );
  AOI211xp5_ASAP7_75t_SL U69792 ( .A1(n59614), .A2(n62662), .B(n62661), .C(
        n68079), .Y(n62663) );
  NOR2xp33_ASAP7_75t_SL U69793 ( .A(n62662), .B(n57108), .Y(n62661) );
  NOR2xp33_ASAP7_75t_SL U69794 ( .A(n67629), .B(n59615), .Y(n62597) );
  NOR2xp33_ASAP7_75t_SL U69795 ( .A(n53283), .B(n59418), .Y(n62665) );
  NOR2xp33_ASAP7_75t_SL U69796 ( .A(n59615), .B(n67920), .Y(n62666) );
  NOR2xp33_ASAP7_75t_SL U69797 ( .A(n57167), .B(n59509), .Y(n62650) );
  NOR2xp33_ASAP7_75t_SL U69798 ( .A(n62719), .B(n62716), .Y(n62717) );
  NOR2xp33_ASAP7_75t_SL U69799 ( .A(n57167), .B(n59618), .Y(n62702) );
  NOR2xp33_ASAP7_75t_SL U69800 ( .A(n59620), .B(n65043), .Y(n62696) );
  NOR2xp33_ASAP7_75t_SL U69801 ( .A(n59614), .B(n67944), .Y(n62745) );
  NOR2xp33_ASAP7_75t_SL U69802 ( .A(n59505), .B(n67444), .Y(n62746) );
  NOR2xp33_ASAP7_75t_SL U69803 ( .A(n63130), .B(n59618), .Y(n63096) );
  NOR2xp33_ASAP7_75t_SL U69804 ( .A(n75900), .B(n59618), .Y(n62759) );
  NOR2xp33_ASAP7_75t_SL U69805 ( .A(n57111), .B(n67442), .Y(n63089) );
  NOR2xp33_ASAP7_75t_SL U69806 ( .A(n53207), .B(n58508), .Y(n63067) );
  NOR2xp33_ASAP7_75t_SL U69807 ( .A(n59502), .B(n59594), .Y(n62653) );
  NOR2xp33_ASAP7_75t_SL U69808 ( .A(n59503), .B(n68087), .Y(n63064) );
  NAND2xp33_ASAP7_75t_SRAM U69809 ( .A(n59504), .B(n59466), .Y(n63147) );
  XNOR2xp5_ASAP7_75t_SL U69810 ( .A(n57113), .B(n67228), .Y(n58473) );
  NOR2xp33_ASAP7_75t_SL U69811 ( .A(n53315), .B(n63097), .Y(n63099) );
  NOR2xp33_ASAP7_75t_SL U69812 ( .A(n57097), .B(n63114), .Y(n58907) );
  NOR2xp33_ASAP7_75t_SL U69813 ( .A(n58408), .B(n59609), .Y(n59211) );
  NOR2xp33_ASAP7_75t_SL U69814 ( .A(n67432), .B(n59509), .Y(n63207) );
  NAND2xp33_ASAP7_75t_SRAM U69815 ( .A(n59615), .B(n59510), .Y(n63202) );
  NOR2xp33_ASAP7_75t_SL U69816 ( .A(n57108), .B(n75904), .Y(n63204) );
  NOR2xp33_ASAP7_75t_SL U69817 ( .A(n67451), .B(n63679), .Y(n63193) );
  AOI211xp5_ASAP7_75t_SL U69818 ( .A1(n64060), .A2(n64059), .B(n64058), .C(
        n64057), .Y(n64064) );
  NOR2xp33_ASAP7_75t_SL U69819 ( .A(n63852), .B(n63853), .Y(n64058) );
  NOR2xp33_ASAP7_75t_SL U69820 ( .A(n53283), .B(n53251), .Y(n63616) );
  NOR2xp33_ASAP7_75t_SL U69821 ( .A(n57110), .B(n76049), .Y(n63617) );
  NOR2xp33_ASAP7_75t_SL U69822 ( .A(n57706), .B(n63219), .Y(n63222) );
  XNOR2xp5_ASAP7_75t_SL U69823 ( .A(n59609), .B(n76028), .Y(n63224) );
  NOR2xp33_ASAP7_75t_SL U69824 ( .A(n63630), .B(n59515), .Y(n63216) );
  NOR2xp33_ASAP7_75t_SL U69825 ( .A(n58962), .B(n67826), .Y(n66617) );
  NOR2xp33_ASAP7_75t_SL U69826 ( .A(n59508), .B(n59670), .Y(n58669) );
  NOR2xp33_ASAP7_75t_SL U69827 ( .A(n68087), .B(n59637), .Y(n66616) );
  NOR2xp33_ASAP7_75t_SL U69828 ( .A(n75900), .B(n67712), .Y(n66681) );
  NOR2xp33_ASAP7_75t_SL U69829 ( .A(n59175), .B(n68119), .Y(n59174) );
  NOR2xp33_ASAP7_75t_SL U69830 ( .A(n59601), .B(n59647), .Y(n66763) );
  NOR2xp33_ASAP7_75t_SL U69831 ( .A(n58670), .B(n59012), .Y(n66668) );
  NOR2xp33_ASAP7_75t_SL U69832 ( .A(n59456), .B(n59670), .Y(n58671) );
  NOR2xp33_ASAP7_75t_SL U69833 ( .A(n59508), .B(n59662), .Y(n66669) );
  NOR2xp33_ASAP7_75t_SL U69834 ( .A(n67826), .B(n53275), .Y(n66670) );
  NOR2xp33_ASAP7_75t_SL U69835 ( .A(n67585), .B(n67712), .Y(n66622) );
  XOR2xp5_ASAP7_75t_SL U69836 ( .A(n68494), .B(n68519), .Y(n59120) );
  AO21x1_ASAP7_75t_SL U69837 ( .A1(n59122), .A2(n58317), .B(n59121), .Y(n68517) );
  NOR2xp33_ASAP7_75t_SL U69838 ( .A(n68514), .B(n68515), .Y(n59121) );
  NOR2xp33_ASAP7_75t_SL U69839 ( .A(n59510), .B(n59637), .Y(n66665) );
  NOR2xp33_ASAP7_75t_SL U69840 ( .A(n57827), .B(n67408), .Y(n66640) );
  NOR2xp33_ASAP7_75t_SL U69841 ( .A(n59508), .B(n58165), .Y(n66744) );
  NOR2xp33_ASAP7_75t_SL U69842 ( .A(n67826), .B(n59664), .Y(n66745) );
  NOR2xp33_ASAP7_75t_SL U69843 ( .A(n59518), .B(n53520), .Y(n59140) );
  NOR2xp33_ASAP7_75t_SL U69844 ( .A(n67962), .B(n59643), .Y(n59301) );
  NOR2xp33_ASAP7_75t_SL U69845 ( .A(n66829), .B(n66797), .Y(n66723) );
  XNOR2xp5_ASAP7_75t_SL U69846 ( .A(n68436), .B(n68435), .Y(n59027) );
  NOR2xp33_ASAP7_75t_SL U69847 ( .A(n59601), .B(n57101), .Y(n66752) );
  NOR2xp33_ASAP7_75t_SL U69848 ( .A(n66720), .B(n66958), .Y(n66721) );
  NOR2xp33_ASAP7_75t_SL U69849 ( .A(n58962), .B(n66716), .Y(n66718) );
  NOR2xp33_ASAP7_75t_SL U69850 ( .A(n59662), .B(n67580), .Y(n59191) );
  NOR2xp33_ASAP7_75t_SL U69851 ( .A(n59456), .B(n53288), .Y(n66714) );
  NOR2xp33_ASAP7_75t_SL U69852 ( .A(n57322), .B(n76071), .Y(n66727) );
  NOR2xp33_ASAP7_75t_SL U69853 ( .A(n75644), .B(n75904), .Y(n66960) );
  NOR2xp33_ASAP7_75t_SL U69854 ( .A(n59620), .B(n57425), .Y(n66961) );
  NOR2xp33_ASAP7_75t_SL U69855 ( .A(n76049), .B(n59519), .Y(n66959) );
  NOR2xp33_ASAP7_75t_SL U69856 ( .A(n66962), .B(n68119), .Y(n66919) );
  XNOR2xp5_ASAP7_75t_SL U69857 ( .A(n76028), .B(n59637), .Y(n66954) );
  NOR2xp33_ASAP7_75t_SL U69858 ( .A(n57101), .B(n68413), .Y(n68417) );
  NAND2xp33_ASAP7_75t_SRAM U69859 ( .A(n59518), .B(n57260), .Y(n68412) );
  NOR2xp33_ASAP7_75t_SL U69860 ( .A(n59012), .B(n66783), .Y(n66784) );
  NOR2xp33_ASAP7_75t_SL U69861 ( .A(n66799), .B(n57172), .Y(n66802) );
  NOR2xp33_ASAP7_75t_SL U69862 ( .A(n59653), .B(n59618), .Y(n63658) );
  NOR2xp33_ASAP7_75t_SL U69863 ( .A(n67288), .B(n67826), .Y(n63631) );
  NOR2xp33_ASAP7_75t_SL U69864 ( .A(n68285), .B(n68284), .Y(n68287) );
  XOR2xp5_ASAP7_75t_SL U69865 ( .A(n64439), .B(n58778), .Y(n58779) );
  NOR2xp33_ASAP7_75t_SL U69866 ( .A(n59033), .B(n59032), .Y(n59034) );
  NOR2xp33_ASAP7_75t_SL U69867 ( .A(n58701), .B(n67951), .Y(n59032) );
  NOR2xp33_ASAP7_75t_SL U69868 ( .A(n57182), .B(n75930), .Y(n58961) );
  NOR2xp33_ASAP7_75t_SL U69869 ( .A(n59467), .B(n67444), .Y(n63840) );
  AOI211xp5_ASAP7_75t_SL U69870 ( .A1(n59614), .A2(n64028), .B(n64027), .C(
        n68079), .Y(n64029) );
  NOR2xp33_ASAP7_75t_SL U69871 ( .A(n57108), .B(n64028), .Y(n64027) );
  NOR2xp33_ASAP7_75t_SL U69872 ( .A(n57662), .B(n59594), .Y(n64386) );
  NOR2xp33_ASAP7_75t_SL U69873 ( .A(n67432), .B(n68011), .Y(n64441) );
  NOR2xp33_ASAP7_75t_SL U69874 ( .A(n57109), .B(n67569), .Y(n64031) );
  NOR2xp33_ASAP7_75t_SL U69875 ( .A(n59618), .B(n57101), .Y(n64071) );
  AND2x2_ASAP7_75t_SL U69876 ( .A(n59656), .B(n57323), .Y(n64345) );
  NOR2xp33_ASAP7_75t_SL U69877 ( .A(n67432), .B(n67463), .Y(n64334) );
  XNOR2xp5_ASAP7_75t_SL U69878 ( .A(n64473), .B(n64476), .Y(n64361) );
  NOR2xp33_ASAP7_75t_SL U69879 ( .A(n58515), .B(n59660), .Y(n64968) );
  NOR2xp33_ASAP7_75t_SL U69880 ( .A(n57111), .B(n57494), .Y(n64963) );
  NOR2xp33_ASAP7_75t_SL U69881 ( .A(n57101), .B(n59509), .Y(n64362) );
  NOR2xp33_ASAP7_75t_SL U69882 ( .A(n57394), .B(n68090), .Y(n64371) );
  NOR2xp33_ASAP7_75t_SL U69883 ( .A(n68102), .B(n64406), .Y(n64407) );
  NOR2xp33_ASAP7_75t_SL U69884 ( .A(n58440), .B(n67736), .Y(n64919) );
  NOR2xp33_ASAP7_75t_SL U69885 ( .A(n57484), .B(n67841), .Y(n64916) );
  NOR2xp33_ASAP7_75t_SL U69886 ( .A(n57108), .B(n59041), .Y(n64425) );
  NOR2xp33_ASAP7_75t_SL U69887 ( .A(n67911), .B(n65043), .Y(n64423) );
  AOI211xp5_ASAP7_75t_SL U69888 ( .A1(n67833), .A2(n64616), .B(n64474), .C(
        n64473), .Y(n64475) );
  NOR2xp33_ASAP7_75t_SL U69889 ( .A(n57111), .B(n59454), .Y(n64473) );
  NOR2xp33_ASAP7_75t_SL U69890 ( .A(n64501), .B(n59253), .Y(n64474) );
  NOR2xp33_ASAP7_75t_SL U69891 ( .A(n59660), .B(n67632), .Y(n64492) );
  NOR2xp33_ASAP7_75t_SL U69892 ( .A(n57107), .B(n67883), .Y(n64646) );
  XNOR2xp5_ASAP7_75t_SL U69893 ( .A(n65028), .B(n64902), .Y(n65051) );
  NOR2xp33_ASAP7_75t_SL U69894 ( .A(n59618), .B(n59650), .Y(n64650) );
  NOR2xp33_ASAP7_75t_SL U69895 ( .A(n65022), .B(n64569), .Y(n64517) );
  NOR2xp33_ASAP7_75t_SL U69896 ( .A(n65022), .B(n64569), .Y(n64570) );
  NOR2xp33_ASAP7_75t_SL U69897 ( .A(n75912), .B(n57110), .Y(n64490) );
  NOR2xp33_ASAP7_75t_SL U69898 ( .A(n59660), .B(n59297), .Y(n64563) );
  NOR2xp33_ASAP7_75t_SL U69899 ( .A(n64483), .B(n57112), .Y(n64484) );
  NOR2xp33_ASAP7_75t_SL U69900 ( .A(n63674), .B(n59659), .Y(n58849) );
  NOR2xp33_ASAP7_75t_SL U69901 ( .A(n57257), .B(n57244), .Y(n64459) );
  XNOR2xp5_ASAP7_75t_SL U69902 ( .A(n68386), .B(n68384), .Y(n59028) );
  NOR2xp33_ASAP7_75t_SL U69903 ( .A(n68087), .B(n58863), .Y(n58864) );
  NOR2xp33_ASAP7_75t_SL U69904 ( .A(n67675), .B(n67674), .Y(n67676) );
  XNOR2xp5_ASAP7_75t_SL U69905 ( .A(n67569), .B(n57292), .Y(n67570) );
  NOR2xp33_ASAP7_75t_SL U69906 ( .A(n59659), .B(n67560), .Y(n59163) );
  XNOR2xp5_ASAP7_75t_SL U69907 ( .A(n75927), .B(n57436), .Y(n67555) );
  NOR2xp33_ASAP7_75t_SL U69908 ( .A(n57169), .B(n57405), .Y(n67533) );
  NOR2xp33_ASAP7_75t_SL U69909 ( .A(n53303), .B(n59647), .Y(n67513) );
  O2A1O1Ixp5_ASAP7_75t_SL U69910 ( .A1(n67494), .A2(n67493), .B(n67492), .C(
        n67491), .Y(n59358) );
  XNOR2xp5_ASAP7_75t_SL U69911 ( .A(n59598), .B(n58919), .Y(n67290) );
  NAND2xp33_ASAP7_75t_SRAM U69912 ( .A(n67535), .B(n57321), .Y(n67490) );
  NOR2xp33_ASAP7_75t_SL U69913 ( .A(n59664), .B(n59297), .Y(n67257) );
  NOR2xp33_ASAP7_75t_SL U69914 ( .A(n59505), .B(n59666), .Y(n67417) );
  NOR2xp33_ASAP7_75t_SL U69915 ( .A(n59065), .B(n57315), .Y(n59064) );
  NOR2xp33_ASAP7_75t_SL U69916 ( .A(n59041), .B(n67566), .Y(n67388) );
  NOR2xp33_ASAP7_75t_SL U69917 ( .A(n68239), .B(n68238), .Y(n68240) );
  NOR2xp33_ASAP7_75t_SL U69918 ( .A(n59456), .B(n67264), .Y(n64958) );
  NAND2xp33_ASAP7_75t_SRAM U69919 ( .A(n57348), .B(n58402), .Y(n64959) );
  NOR2xp33_ASAP7_75t_SL U69920 ( .A(n59012), .B(n67843), .Y(n64940) );
  NOR2xp33_ASAP7_75t_SL U69921 ( .A(n58992), .B(n63082), .Y(n58991) );
  NOR2xp33_ASAP7_75t_SL U69922 ( .A(n59459), .B(n53283), .Y(n58992) );
  NOR2xp33_ASAP7_75t_SL U69923 ( .A(n59647), .B(n67866), .Y(n65045) );
  NOR2xp33_ASAP7_75t_SL U69924 ( .A(n59596), .B(n58431), .Y(n64499) );
  NOR2xp33_ASAP7_75t_SL U69925 ( .A(n59598), .B(n67288), .Y(n64500) );
  NOR2xp33_ASAP7_75t_SL U69926 ( .A(n59509), .B(n58015), .Y(n65018) );
  NOR2xp33_ASAP7_75t_SL U69927 ( .A(n59352), .B(n59514), .Y(n59335) );
  NAND3xp33_ASAP7_75t_SL U69928 ( .A(n59607), .B(n66860), .C(n59656), .Y(
        n59304) );
  NOR3xp33_ASAP7_75t_SL U69929 ( .A(n67234), .B(n67233), .C(n67232), .Y(n67235) );
  NOR2xp33_ASAP7_75t_SL U69930 ( .A(n57274), .B(n59519), .Y(n67239) );
  NOR2xp33_ASAP7_75t_SL U69931 ( .A(n67359), .B(n59046), .Y(n59047) );
  NOR2xp33_ASAP7_75t_SL U69932 ( .A(n57111), .B(n68119), .Y(n68120) );
  NOR2xp33_ASAP7_75t_SL U69933 ( .A(n59012), .B(n68118), .Y(n68121) );
  NOR2xp33_ASAP7_75t_SL U69934 ( .A(n57108), .B(n57101), .Y(n68083) );
  AOI31xp33_ASAP7_75t_SL U69935 ( .A1(n68098), .A2(n57106), .A3(n68097), .B(
        n58015), .Y(n68099) );
  NOR2xp33_ASAP7_75t_SL U69936 ( .A(n59509), .B(n76172), .Y(n68091) );
  MAJx2_ASAP7_75t_SL U69937 ( .A(n59360), .B(n67984), .C(n58843), .Y(n67804)
         );
  NOR2xp33_ASAP7_75t_SL U69938 ( .A(n67640), .B(n59399), .Y(n67876) );
  NOR2xp33_ASAP7_75t_SL U69939 ( .A(n64623), .B(n59044), .Y(n58718) );
  O2A1O1Ixp5_ASAP7_75t_SL U69940 ( .A1(n59618), .A2(n59664), .B(n67859), .C(
        n67858), .Y(n68130) );
  NOR2xp33_ASAP7_75t_SL U69941 ( .A(n59509), .B(n75962), .Y(n67858) );
  NOR2xp33_ASAP7_75t_SL U69942 ( .A(n53283), .B(n75899), .Y(n67362) );
  NOR2xp33_ASAP7_75t_SL U69943 ( .A(n59609), .B(n58526), .Y(n67355) );
  NOR2xp33_ASAP7_75t_SL U69944 ( .A(n59604), .B(n67383), .Y(n67359) );
  NOR2xp33_ASAP7_75t_SL U69945 ( .A(n59125), .B(n66322), .Y(n59124) );
  NOR2xp33_ASAP7_75t_SL U69946 ( .A(n53303), .B(n67334), .Y(n67336) );
  NOR2xp33_ASAP7_75t_SL U69947 ( .A(n59508), .B(n67333), .Y(n67337) );
  NAND2xp33_ASAP7_75t_SRAM U69948 ( .A(n77713), .B(n57122), .Y(n67332) );
  NOR2xp33_ASAP7_75t_SL U69949 ( .A(n59658), .B(n67328), .Y(n67330) );
  AOI211xp5_ASAP7_75t_SL U69950 ( .A1(n67344), .A2(n67715), .B(n58706), .C(
        n67895), .Y(n59137) );
  NOR2xp33_ASAP7_75t_SL U69951 ( .A(n67346), .B(n53493), .Y(n67349) );
  XNOR2xp5_ASAP7_75t_SL U69952 ( .A(n57322), .B(n57425), .Y(n67435) );
  NOR2xp33_ASAP7_75t_SL U69953 ( .A(n59502), .B(n59352), .Y(n67305) );
  NOR2xp33_ASAP7_75t_SL U69954 ( .A(n75927), .B(n58845), .Y(n67321) );
  NOR2xp33_ASAP7_75t_SL U69955 ( .A(n57272), .B(n59503), .Y(n68007) );
  NOR2xp33_ASAP7_75t_SL U69956 ( .A(n59592), .B(n63674), .Y(n68005) );
  NOR2xp33_ASAP7_75t_SL U69957 ( .A(n53317), .B(n68019), .Y(n68018) );
  XNOR2xp5_ASAP7_75t_SL U69958 ( .A(n59079), .B(n62636), .Y(n63674) );
  NOR2xp33_ASAP7_75t_SL U69959 ( .A(n59012), .B(n67827), .Y(n67828) );
  XOR2xp5_ASAP7_75t_SL U69960 ( .A(n57107), .B(n59468), .Y(n67827) );
  NOR2xp33_ASAP7_75t_SL U69961 ( .A(n58919), .B(n59508), .Y(n67830) );
  NOR2xp33_ASAP7_75t_SL U69962 ( .A(n59381), .B(n67826), .Y(n67831) );
  NOR2xp33_ASAP7_75t_SL U69963 ( .A(n57696), .B(n67962), .Y(n67341) );
  XOR2xp5_ASAP7_75t_SL U69964 ( .A(n58863), .B(n75930), .Y(n58398) );
  NOR2xp33_ASAP7_75t_SL U69965 ( .A(n59598), .B(n67846), .Y(n67584) );
  NOR2xp33_ASAP7_75t_SL U69966 ( .A(n67629), .B(n59649), .Y(n58806) );
  NAND3xp33_ASAP7_75t_SL U69967 ( .A(n62808), .B(n57118), .C(n62807), .Y(
        n76632) );
  NOR2xp33_ASAP7_75t_SL U69968 ( .A(n59545), .B(n64894), .Y(n62593) );
  NAND3xp33_ASAP7_75t_SL U69969 ( .A(n62560), .B(n62559), .C(n59197), .Y(
        n68410) );
  NOR2xp33_ASAP7_75t_SL U69970 ( .A(n59596), .B(n59601), .Y(n67637) );
  NOR2xp33_ASAP7_75t_SL U69971 ( .A(n59546), .B(n63654), .Y(n59210) );
  NOR2xp33_ASAP7_75t_SL U69972 ( .A(n67911), .B(n59605), .Y(n67913) );
  NOR2xp33_ASAP7_75t_SL U69973 ( .A(n59509), .B(n59664), .Y(n67924) );
  NOR2xp33_ASAP7_75t_SL U69974 ( .A(n62579), .B(n62578), .Y(n68096) );
  NOR2xp33_ASAP7_75t_SL U69975 ( .A(n63662), .B(n63661), .Y(n63663) );
  NAND2xp33_ASAP7_75t_SRAM U69976 ( .A(n66258), .B(n63660), .Y(n63662) );
  NOR2xp33_ASAP7_75t_SL U69977 ( .A(n59596), .B(n76049), .Y(n67916) );
  NOR2xp33_ASAP7_75t_SL U69978 ( .A(n67972), .B(n57109), .Y(n67973) );
  NOR3xp33_ASAP7_75t_SL U69979 ( .A(n62589), .B(n59471), .C(n58972), .Y(n58973) );
  NOR2xp33_ASAP7_75t_SL U69980 ( .A(n57128), .B(n59479), .Y(n62700) );
  NOR2xp33_ASAP7_75t_SL U69981 ( .A(n59508), .B(n67959), .Y(n67961) );
  NOR2xp33_ASAP7_75t_SL U69982 ( .A(n58513), .B(n61913), .Y(n59019) );
  NOR2xp33_ASAP7_75t_SL U69983 ( .A(n63249), .B(n53615), .Y(n63252) );
  NOR2xp33_ASAP7_75t_SL U69984 ( .A(n63184), .B(n64353), .Y(n63672) );
  AOI31xp33_ASAP7_75t_SL U69985 ( .A1(n63180), .A2(n63179), .A3(n63178), .B(
        n75378), .Y(n63181) );
  NOR2xp33_ASAP7_75t_SL U69986 ( .A(n62591), .B(n59184), .Y(n63178) );
  NAND2xp33_ASAP7_75t_SRAM U69987 ( .A(n59559), .B(n59568), .Y(n59184) );
  NOR2xp33_ASAP7_75t_SL U69988 ( .A(n59654), .B(n62667), .Y(n62670) );
  NOR2xp33_ASAP7_75t_SL U69989 ( .A(n78003), .B(n59654), .Y(n62657) );
  OR2x2_ASAP7_75t_SL U69990 ( .A(n62630), .B(n62631), .Y(n67444) );
  NAND3xp33_ASAP7_75t_SL U69991 ( .A(n75035), .B(n66263), .C(n66262), .Y(
        n66264) );
  NAND2xp33_ASAP7_75t_SRAM U69992 ( .A(n59641), .B(n57456), .Y(n75070) );
  NOR2xp33_ASAP7_75t_SL U69993 ( .A(n68606), .B(n59116), .Y(n68608) );
  NOR2xp33_ASAP7_75t_SL U69994 ( .A(n53300), .B(n58940), .Y(n58939) );
  NOR2xp33_ASAP7_75t_SL U69995 ( .A(n59574), .B(n53300), .Y(n66310) );
  NOR2xp33_ASAP7_75t_SL U69996 ( .A(n65030), .B(n66240), .Y(n65032) );
  NOR2xp33_ASAP7_75t_SL U69997 ( .A(n75054), .B(n58962), .Y(n75068) );
  NOR2xp33_ASAP7_75t_SL U69998 ( .A(n57398), .B(n59670), .Y(n75466) );
  NOR2xp33_ASAP7_75t_SL U69999 ( .A(n57215), .B(n66253), .Y(n66257) );
  XNOR2xp5_ASAP7_75t_SL U70000 ( .A(n59518), .B(n57456), .Y(n75043) );
  NOR2xp33_ASAP7_75t_SL U70001 ( .A(n65031), .B(n61208), .Y(n66283) );
  NAND3xp33_ASAP7_75t_SL U70002 ( .A(n60629), .B(n59080), .C(n59438), .Y(
        n59324) );
  NAND3xp33_ASAP7_75t_SL U70003 ( .A(n59438), .B(n59464), .C(n59566), .Y(
        n59414) );
  NOR2xp33_ASAP7_75t_SL U70004 ( .A(iwb_dat_i[16]), .B(n78006), .Y(n77956) );
  NOR2xp33_ASAP7_75t_SL U70005 ( .A(dc_en), .B(n61293), .Y(n60211) );
  AND2x2_ASAP7_75t_SL U70006 ( .A(n62567), .B(n62565), .Y(n58403) );
  OR2x2_ASAP7_75t_SL U70007 ( .A(n58497), .B(n59465), .Y(n58405) );
  OR2x2_ASAP7_75t_SL U70008 ( .A(n59348), .B(n59349), .Y(n58406) );
  OR2x2_ASAP7_75t_SL U70009 ( .A(n58537), .B(n64894), .Y(n58407) );
  OR2x2_ASAP7_75t_SL U70010 ( .A(n59592), .B(n58853), .Y(n58409) );
  AO21x1_ASAP7_75t_SL U70011 ( .A1(n75922), .A2(n59615), .B(n62943), .Y(n58410) );
  OR2x2_ASAP7_75t_SL U70012 ( .A(n59456), .B(n59662), .Y(n58411) );
  OR2x2_ASAP7_75t_SL U70013 ( .A(n58990), .B(n59662), .Y(n58412) );
  AO21x1_ASAP7_75t_SL U70014 ( .A1(n58433), .A2(n59709), .B(n67860), .Y(n58414) );
  OR2x2_ASAP7_75t_SL U70015 ( .A(n2757), .B(n57090), .Y(n58415) );
  OR2x2_ASAP7_75t_SL U70016 ( .A(n59167), .B(n74788), .Y(n58420) );
  NOR3xp33_ASAP7_75t_SL U70017 ( .A(n59145), .B(n67607), .C(n57112), .Y(n58425) );
  AND2x2_ASAP7_75t_SL U70018 ( .A(n62567), .B(n62566), .Y(n58426) );
  AND3x1_ASAP7_75t_SL U70019 ( .A(n59571), .B(n59542), .C(n59569), .Y(n58428)
         );
  OR2x2_ASAP7_75t_SL U70020 ( .A(n57112), .B(n59145), .Y(n58432) );
  AND2x2_ASAP7_75t_SL U70021 ( .A(n67537), .B(n59232), .Y(n58436) );
  AND2x2_ASAP7_75t_SL U70022 ( .A(n64078), .B(n59655), .Y(n58437) );
  OR2x2_ASAP7_75t_SL U70023 ( .A(n58486), .B(n66810), .Y(n58438) );
  OR2x2_ASAP7_75t_SL U70024 ( .A(n68838), .B(n68908), .Y(n58442) );
  AND3x1_ASAP7_75t_SL U70025 ( .A(n66292), .B(n59549), .C(n1868), .Y(n58443)
         );
  OR2x2_ASAP7_75t_SL U70026 ( .A(n62568), .B(n62572), .Y(n58444) );
  AND2x2_ASAP7_75t_SL U70027 ( .A(n68674), .B(n69116), .Y(n58445) );
  AND2x2_ASAP7_75t_SL U70028 ( .A(n67746), .B(n57067), .Y(n58446) );
  AND2x2_ASAP7_75t_SL U70029 ( .A(n59617), .B(n75900), .Y(n58449) );
  NOR2xp33_ASAP7_75t_SL U70030 ( .A(n59456), .B(n59659), .Y(n58848) );
  AND2x2_ASAP7_75t_SL U70031 ( .A(n69239), .B(n74113), .Y(n58450) );
  MAJx2_ASAP7_75t_SL U70032 ( .A(n58468), .B(n67817), .C(n67816), .Y(n58455)
         );
  OR2x2_ASAP7_75t_SL U70033 ( .A(n64721), .B(n64718), .Y(n58457) );
  OA21x2_ASAP7_75t_SL U70034 ( .A1(n59183), .A2(n66258), .B(n57448), .Y(n58458) );
  AND2x2_ASAP7_75t_SL U70035 ( .A(n62742), .B(n68079), .Y(n58462) );
  OR2x2_ASAP7_75t_SL U70036 ( .A(n62642), .B(n62641), .Y(n58463) );
  AND2x2_ASAP7_75t_SL U70037 ( .A(n67410), .B(n57827), .Y(n58464) );
  OA21x2_ASAP7_75t_SL U70038 ( .A1(n57243), .A2(n58919), .B(n64440), .Y(n58465) );
  MAJx2_ASAP7_75t_SL U70039 ( .A(n66777), .B(n66653), .C(n66774), .Y(n58467)
         );
  OA21x2_ASAP7_75t_SL U70040 ( .A1(n67361), .A2(n59515), .B(n59201), .Y(n58468) );
  AND2x2_ASAP7_75t_SL U70041 ( .A(n75628), .B(n66244), .Y(n58469) );
  OR2x2_ASAP7_75t_SL U70042 ( .A(n64045), .B(n64046), .Y(n58470) );
  OR2x2_ASAP7_75t_SL U70043 ( .A(n68643), .B(n75096), .Y(n58471) );
  AO21x1_ASAP7_75t_SL U70044 ( .A1(n68333), .A2(n68332), .B(n68331), .Y(n58472) );
  AND2x2_ASAP7_75t_SL U70045 ( .A(n76429), .B(n59589), .Y(n58474) );
  AND2x2_ASAP7_75t_SL U70046 ( .A(n67430), .B(n67429), .Y(n58475) );
  OR2x2_ASAP7_75t_SL U70047 ( .A(n62953), .B(n62952), .Y(n58477) );
  AO21x1_ASAP7_75t_SL U70048 ( .A1(n68008), .A2(n56827), .B(n59475), .Y(n58479) );
  AND2x2_ASAP7_75t_SL U70049 ( .A(n59257), .B(n61908), .Y(n58480) );
  AO21x1_ASAP7_75t_SL U70050 ( .A1(n67736), .A2(n67607), .B(n67606), .Y(n58482) );
  AND2x2_ASAP7_75t_SL U70051 ( .A(n59505), .B(n59615), .Y(n58483) );
  OR2x2_ASAP7_75t_SL U70052 ( .A(n69294), .B(n69295), .Y(n58485) );
  AND2x2_ASAP7_75t_SL U70053 ( .A(n1868), .B(n59655), .Y(n58487) );
  OR2x2_ASAP7_75t_SL U70054 ( .A(n61921), .B(n58632), .Y(n58489) );
  AND2x2_ASAP7_75t_SL U70055 ( .A(n59605), .B(n67971), .Y(n58490) );
  OR2x2_ASAP7_75t_SL U70056 ( .A(n67944), .B(n67463), .Y(n58493) );
  MAJx2_ASAP7_75t_SL U70057 ( .A(n68207), .B(n68205), .C(n58352), .Y(n58495)
         );
  OR2x2_ASAP7_75t_SL U70058 ( .A(n64617), .B(n57209), .Y(n58496) );
  AO21x1_ASAP7_75t_SL U70059 ( .A1(n62606), .A2(n62605), .B(n62604), .Y(n58497) );
  XOR2xp5_ASAP7_75t_SL U70060 ( .A(n75901), .B(n75438), .Y(n58498) );
  OR2x2_ASAP7_75t_SL U70061 ( .A(n59125), .B(n64920), .Y(n58501) );
  AND2x2_ASAP7_75t_SL U70062 ( .A(n67899), .B(n75906), .Y(n58504) );
  OR2x2_ASAP7_75t_SL U70063 ( .A(n67337), .B(n67336), .Y(n58505) );
  AND2x2_ASAP7_75t_SL U70064 ( .A(n67343), .B(n53613), .Y(n58506) );
  OR2x2_ASAP7_75t_SL U70065 ( .A(n59301), .B(n66729), .Y(n58507) );
  OR2x2_ASAP7_75t_SL U70066 ( .A(n57272), .B(n67326), .Y(n58508) );
  MAJx2_ASAP7_75t_SL U70067 ( .A(n68531), .B(n68532), .C(n68533), .Y(n58511)
         );
  AND2x2_ASAP7_75t_SL U70068 ( .A(n57501), .B(n64538), .Y(n58512) );
  OR2x2_ASAP7_75t_SL U70069 ( .A(n77701), .B(n61921), .Y(n58513) );
  AO21x1_ASAP7_75t_SL U70070 ( .A1(n57122), .A2(n77696), .B(n67625), .Y(n58514) );
  OR2x2_ASAP7_75t_SL U70071 ( .A(n64966), .B(n57108), .Y(n58515) );
  OR2x2_ASAP7_75t_SL U70072 ( .A(n66860), .B(n59670), .Y(n58516) );
  AO21x1_ASAP7_75t_SL U70073 ( .A1(n53274), .A2(n67979), .B(n58488), .Y(n58518) );
  AND2x2_ASAP7_75t_SL U70074 ( .A(n58919), .B(n67951), .Y(n58519) );
  OA21x2_ASAP7_75t_SL U70075 ( .A1(n58887), .A2(n68973), .B(n68837), .Y(n58522) );
  OR2x2_ASAP7_75t_SL U70076 ( .A(n58928), .B(n58929), .Y(n58523) );
  OR2x2_ASAP7_75t_SL U70077 ( .A(n57068), .B(n67357), .Y(n58526) );
  AND2x2_ASAP7_75t_SL U70078 ( .A(n69040), .B(n69039), .Y(n58527) );
  OR2x2_ASAP7_75t_SL U70079 ( .A(n62709), .B(n62708), .Y(n58528) );
  MAJx2_ASAP7_75t_SL U70080 ( .A(n66626), .B(n66627), .C(n66628), .Y(n58529)
         );
  OA21x2_ASAP7_75t_SL U70081 ( .A1(n57165), .A2(n66535), .B(n59143), .Y(n58530) );
  AND2x2_ASAP7_75t_SL U70082 ( .A(n57177), .B(n59660), .Y(n58531) );
  OR2x2_ASAP7_75t_SL U70083 ( .A(n69240), .B(n69241), .Y(n58533) );
  OR2x2_ASAP7_75t_SL U70084 ( .A(n66860), .B(n59662), .Y(n58534) );
  AND2x2_ASAP7_75t_SL U70085 ( .A(n57448), .B(n53316), .Y(n58535) );
  OR2x2_ASAP7_75t_SL U70086 ( .A(n62722), .B(n62723), .Y(n58536) );
  AND2x2_ASAP7_75t_SL U70087 ( .A(n77242), .B(n59183), .Y(n58537) );
  AND2x2_ASAP7_75t_SL U70088 ( .A(n69115), .B(n69122), .Y(n58538) );
  AND2x2_ASAP7_75t_SL U70089 ( .A(or1200_ic_top_from_icram[22]), .B(n53436), 
        .Y(n58540) );
  AND2x2_ASAP7_75t_SL U70090 ( .A(n68924), .B(n68926), .Y(n58541) );
  OR2x2_ASAP7_75t_SL U70091 ( .A(n62806), .B(n59236), .Y(n58542) );
  OR3x1_ASAP7_75t_SL U70092 ( .A(n69115), .B(n69119), .C(n69114), .Y(n58543)
         );
  AO22x1_ASAP7_75t_SL U70093 ( .A1(n59701), .A2(n76581), .B1(n76580), .B2(
        n53440), .Y(n58545) );
  OA211x2_ASAP7_75t_SL U70094 ( .A1(n77667), .A2(n75880), .B(n75879), .C(
        n75878), .Y(n58548) );
  OA211x2_ASAP7_75t_SL U70095 ( .A1(n75357), .A2(n75602), .B(n75356), .C(
        n75355), .Y(n58549) );
  AND3x1_ASAP7_75t_SL U70096 ( .A(n74289), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_23_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_1_), .Y(
        n58550) );
  AND2x2_ASAP7_75t_SL U70097 ( .A(n2009), .B(n65318), .Y(n58551) );
  AND2x2_ASAP7_75t_SL U70098 ( .A(or1200_cpu_spr_dat_rf[1]), .B(n77848), .Y(
        n58552) );
  OR2x2_ASAP7_75t_SL U70099 ( .A(n58553), .B(n70046), .Y(n58555) );
  OR2x2_ASAP7_75t_SL U70100 ( .A(n2979), .B(n57074), .Y(n58556) );
  OR3x1_ASAP7_75t_SL U70101 ( .A(n62103), .B(n62102), .C(n62101), .Y(n58557)
         );
  AND2x2_ASAP7_75t_SL U70102 ( .A(n74937), .B(n74936), .Y(n58559) );
  AND2x2_ASAP7_75t_SL U70103 ( .A(n76842), .B(n57100), .Y(n58560) );
  AO22x1_ASAP7_75t_SL U70104 ( .A1(n59700), .A2(iwb_adr_o[25]), .B1(n57084), 
        .B2(icbiu_adr_ic_word[25]), .Y(n58561) );
  AO22x1_ASAP7_75t_SL U70105 ( .A1(n59700), .A2(iwb_adr_o[29]), .B1(n57084), 
        .B2(icbiu_adr_ic_word[29]), .Y(n58562) );
  AO22x1_ASAP7_75t_SL U70106 ( .A1(n59700), .A2(iwb_adr_o[27]), .B1(n57084), 
        .B2(icbiu_adr_ic_word[27]), .Y(n58563) );
  AO22x1_ASAP7_75t_SL U70107 ( .A1(n59700), .A2(iwb_adr_o[28]), .B1(n57084), 
        .B2(icbiu_adr_ic_word[28]), .Y(n58564) );
  AO22x1_ASAP7_75t_SL U70108 ( .A1(or1200_cpu_spr_dat_rf[12]), .A2(n59686), 
        .B1(n77587), .B2(n75532), .Y(n58565) );
  OA21x2_ASAP7_75t_SL U70109 ( .A1(n75648), .A2(n62394), .B(n62400), .Y(n58566) );
  AND2x2_ASAP7_75t_SL U70110 ( .A(n76520), .B(n57100), .Y(n58567) );
  AND2x2_ASAP7_75t_SL U70111 ( .A(n69635), .B(n69634), .Y(n58568) );
  OR2x2_ASAP7_75t_SL U70112 ( .A(n58665), .B(n59670), .Y(n58569) );
  OA21x2_ASAP7_75t_SL U70113 ( .A1(n59891), .A2(n61294), .B(n77686), .Y(n58570) );
  AND2x2_ASAP7_75t_SL U70114 ( .A(n78243), .B(n78244), .Y(n58572) );
  OR2x2_ASAP7_75t_SL U70115 ( .A(n77943), .B(n60545), .Y(n58574) );
  OA21x2_ASAP7_75t_SL U70116 ( .A1(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_28_), .A2(n78360), .B(n72605), .Y(n58575) );
  OA21x2_ASAP7_75t_SL U70117 ( .A1(n65972), .A2(n66026), .B(n65877), .Y(n58576) );
  AO22x1_ASAP7_75t_SL U70118 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .A2(n57193), 
        .B1(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[18]), .B2(n57194), .Y(n58578) );
  OA21x2_ASAP7_75t_SL U70119 ( .A1(n69831), .A2(n69818), .B(n69837), .Y(n58579) );
  AO22x1_ASAP7_75t_SL U70120 ( .A1(n59706), .A2(dwb_adr_o[26]), .B1(n57083), 
        .B2(sbbiu_adr_sb[26]), .Y(n58580) );
  AO22x1_ASAP7_75t_SL U70121 ( .A1(n59706), .A2(dwb_adr_o[28]), .B1(n57083), 
        .B2(sbbiu_adr_sb[28]), .Y(n58581) );
  OA21x2_ASAP7_75t_SL U70122 ( .A1(n70118), .A2(n70017), .B(n70077), .Y(n58583) );
  AO22x1_ASAP7_75t_SL U70123 ( .A1(n59706), .A2(dwb_adr_o[27]), .B1(n57083), 
        .B2(sbbiu_adr_sb[27]), .Y(n58584) );
  AO22x1_ASAP7_75t_SL U70124 ( .A1(n59706), .A2(dwb_adr_o[29]), .B1(n57083), 
        .B2(sbbiu_adr_sb[29]), .Y(n58585) );
  AO22x1_ASAP7_75t_SL U70125 ( .A1(n59706), .A2(dwb_adr_o[20]), .B1(n57083), 
        .B2(sbbiu_adr_sb[20]), .Y(n58586) );
  OA21x2_ASAP7_75t_SL U70126 ( .A1(n59533), .A2(n63660), .B(n60932), .Y(n58587) );
  OA21x2_ASAP7_75t_SL U70127 ( .A1(n59569), .A2(n59442), .B(n63571), .Y(n58589) );
  AO22x1_ASAP7_75t_SL U70128 ( .A1(n59706), .A2(dwb_adr_o[19]), .B1(n57083), 
        .B2(sbbiu_adr_sb[19]), .Y(n58590) );
  OA21x2_ASAP7_75t_SL U70129 ( .A1(n75871), .A2(n77078), .B(n75870), .Y(n58591) );
  AO22x1_ASAP7_75t_SL U70130 ( .A1(n59706), .A2(dwb_adr_o[25]), .B1(n57083), 
        .B2(sbbiu_adr_sb[25]), .Y(n58593) );
  AO22x1_ASAP7_75t_SL U70131 ( .A1(n59706), .A2(dwb_adr_o[15]), .B1(n57083), 
        .B2(sbbiu_adr_sb[15]), .Y(n58594) );
  OR2x2_ASAP7_75t_SL U70132 ( .A(n74164), .B(n74163), .Y(n58595) );
  AO22x1_ASAP7_75t_SL U70133 ( .A1(n59706), .A2(dwb_adr_o[17]), .B1(n57083), 
        .B2(sbbiu_adr_sb[17]), .Y(n58596) );
  AO21x1_ASAP7_75t_SL U70134 ( .A1(n66225), .A2(n1137), .B(n75648), .Y(n58597)
         );
  OR2x2_ASAP7_75t_SL U70135 ( .A(n59492), .B(n74029), .Y(n58598) );
  AO22x1_ASAP7_75t_SL U70136 ( .A1(n59706), .A2(dwb_adr_o[14]), .B1(n57083), 
        .B2(sbbiu_adr_sb[14]), .Y(n58602) );
  AO22x1_ASAP7_75t_SL U70137 ( .A1(n59706), .A2(dwb_adr_o[23]), .B1(n57083), 
        .B2(sbbiu_adr_sb[23]), .Y(n58603) );
  AO22x1_ASAP7_75t_SL U70138 ( .A1(n59706), .A2(dwb_adr_o[22]), .B1(n57083), 
        .B2(sbbiu_adr_sb[22]), .Y(n58605) );
  OA21x2_ASAP7_75t_SL U70139 ( .A1(n71568), .A2(n71480), .B(n71479), .Y(n58606) );
  AO22x1_ASAP7_75t_SL U70140 ( .A1(n59706), .A2(dwb_adr_o[12]), .B1(n57083), 
        .B2(sbbiu_adr_sb[12]), .Y(n58610) );
  AND2x2_ASAP7_75t_SL U70141 ( .A(n61033), .B(n61134), .Y(n58613) );
  AO22x1_ASAP7_75t_SL U70142 ( .A1(n77082), .A2(n76681), .B1(
        or1200_cpu_or1200_fpu_result_arith[2]), .B2(n77091), .Y(n58614) );
  AND2x2_ASAP7_75t_SL U70143 ( .A(n72097), .B(n72096), .Y(n58615) );
  AND2x2_ASAP7_75t_SL U70144 ( .A(or1200_cpu_or1200_rf_rf_we_allow), .B(n75518), .Y(n58616) );
  AND2x2_ASAP7_75t_SL U70145 ( .A(or1200_cpu_or1200_except_n658), .B(n2037), 
        .Y(n58618) );
  AND2x2_ASAP7_75t_SL U70146 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_), .B(
        n74680), .Y(n58620) );
  OA21x2_ASAP7_75t_SL U70147 ( .A1(n69369), .A2(n77208), .B(n74938), .Y(n58621) );
  AND3x1_ASAP7_75t_SL U70148 ( .A(n73671), .B(n73670), .C(n73669), .Y(n58623)
         );
  AND2x2_ASAP7_75t_SL U70149 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_count_3_), 
        .B(n62061), .Y(n58624) );
  AND2x2_ASAP7_75t_SL U70150 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_rmode_i_1_), .B(
        n74289), .Y(n58625) );
  OR2x2_ASAP7_75t_SL U70151 ( .A(or1200_cpu_or1200_except_n571), .B(n1737), 
        .Y(n58626) );
  AND4x1_ASAP7_75t_SL U70152 ( .A(n77853), .B(n77852), .C(n77851), .D(n77850), 
        .Y(n77928) );
  NAND3xp33_ASAP7_75t_SL U70153 ( .A(n59484), .B(n57111), .C(n59518), .Y(
        n67878) );
  XOR2xp5_ASAP7_75t_SL U70154 ( .A(n68313), .B(n68314), .Y(n58636) );
  MAJx2_ASAP7_75t_SL U70155 ( .A(n67656), .B(n67655), .C(n67254), .Y(n67274)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70156 ( .A1(n59466), .A2(n59381), .B(n67926), .C(
        n57637), .Y(n67927) );
  MAJIxp5_ASAP7_75t_SL U70157 ( .A(n58348), .B(n68146), .C(n58368), .Y(n68198)
         );
  NOR2xp33_ASAP7_75t_SL U70158 ( .A(n58654), .B(n60613), .Y(n60654) );
  XNOR2xp5_ASAP7_75t_SL U70159 ( .A(n67784), .B(n67785), .Y(n59083) );
  MAJIxp5_ASAP7_75t_SL U70160 ( .A(n67779), .B(n67778), .C(n67777), .Y(n67785)
         );
  MAJIxp5_ASAP7_75t_SL U70161 ( .A(n67313), .B(n57419), .C(n67835), .Y(n67778)
         );
  XOR2xp5_ASAP7_75t_SL U70162 ( .A(n67297), .B(n67296), .Y(n58661) );
  A2O1A1Ixp33_ASAP7_75t_SL U70163 ( .A1(n59463), .A2(n58672), .B(n66718), .C(
        n66717), .Y(n66958) );
  O2A1O1Ixp5_ASAP7_75t_SL U70164 ( .A1(or1200_cpu_or1200_mult_mac_n6), .A2(
        n76191), .B(n75966), .C(n58672), .Y(n76190) );
  AO21x1_ASAP7_75t_SL U70165 ( .A1(n69116), .A2(n58881), .B(n58774), .Y(n69103) );
  A2O1A1Ixp33_ASAP7_75t_SL U70166 ( .A1(n68973), .A2(n59342), .B(n58685), .C(
        n58683), .Y(n52013) );
  NAND3xp33_ASAP7_75t_SL U70167 ( .A(n59345), .B(n68809), .C(n59343), .Y(
        n76879) );
  XNOR2xp5_ASAP7_75t_SL U70168 ( .A(n58689), .B(n67398), .Y(n59222) );
  MAJIxp5_ASAP7_75t_SL U70169 ( .A(n65014), .B(n65013), .C(n58690), .Y(n68279)
         );
  XNOR2xp5_ASAP7_75t_SL U70170 ( .A(n67993), .B(n67994), .Y(n67998) );
  O2A1O1Ixp5_ASAP7_75t_SL U70171 ( .A1(n67831), .A2(n67830), .B(n67829), .C(
        n67828), .Y(n67994) );
  XNOR2xp5_ASAP7_75t_SL U70172 ( .A(n67622), .B(n67623), .Y(n58694) );
  XNOR2xp5_ASAP7_75t_SL U70173 ( .A(n59511), .B(n57630), .Y(n62794) );
  XOR2xp5_ASAP7_75t_SL U70174 ( .A(n59511), .B(n59637), .Y(n67246) );
  XNOR2xp5_ASAP7_75t_SL U70175 ( .A(n58383), .B(n59511), .Y(n64497) );
  XOR2xp5_ASAP7_75t_SL U70176 ( .A(n59603), .B(n59511), .Y(n62750) );
  XOR2xp5_ASAP7_75t_SL U70177 ( .A(n59511), .B(n75996), .Y(n75992) );
  XNOR2xp5_ASAP7_75t_SL U70178 ( .A(n59303), .B(n58705), .Y(n58948) );
  XOR2xp5_ASAP7_75t_SL U70179 ( .A(n68202), .B(n59313), .Y(n58705) );
  MAJIxp5_ASAP7_75t_SL U70180 ( .A(n63153), .B(n63154), .C(n63155), .Y(n63201)
         );
  XNOR2xp5_ASAP7_75t_SL U70181 ( .A(n67175), .B(n67174), .Y(n67176) );
  MAJIxp5_ASAP7_75t_SL U70182 ( .A(n67155), .B(n67156), .C(n58710), .Y(n67174)
         );
  NOR2xp33_ASAP7_75t_SL U70183 ( .A(n59350), .B(n66800), .Y(n66676) );
  MAJIxp5_ASAP7_75t_SL U70184 ( .A(n58723), .B(n68525), .C(n66943), .Y(n68542)
         );
  MAJIxp5_ASAP7_75t_SL U70185 ( .A(n58734), .B(n64436), .C(n64437), .Y(n64674)
         );
  MAJIxp5_ASAP7_75t_SL U70186 ( .A(n68145), .B(n68142), .C(n53503), .Y(n68569)
         );
  XNOR2xp5_ASAP7_75t_SL U70187 ( .A(n58742), .B(n68177), .Y(n58741) );
  XNOR2xp5_ASAP7_75t_SL U70188 ( .A(n67178), .B(n67189), .Y(n58751) );
  XNOR2xp5_ASAP7_75t_SL U70189 ( .A(n67091), .B(n67131), .Y(n67186) );
  MAJx2_ASAP7_75t_SL U70190 ( .A(n59202), .B(n68445), .C(n68446), .Y(n68515)
         );
  MAJIxp5_ASAP7_75t_SL U70191 ( .A(n58781), .B(n58782), .C(n68353), .Y(n59202)
         );
  MAJx2_ASAP7_75t_SL U70192 ( .A(n68385), .B(n68384), .C(n68386), .Y(n68448)
         );
  AND2x2_ASAP7_75t_SL U70193 ( .A(n57325), .B(n58785), .Y(n66318) );
  OR2x2_ASAP7_75t_SL U70194 ( .A(n58408), .B(n57179), .Y(n58790) );
  MAJIxp5_ASAP7_75t_SL U70195 ( .A(n68202), .B(n68203), .C(n58796), .Y(n68190)
         );
  NAND3xp33_ASAP7_75t_SL U70196 ( .A(n58797), .B(n61920), .C(n61964), .Y(
        n61969) );
  OA21x2_ASAP7_75t_SL U70197 ( .A1(n59636), .A2(n58799), .B(n58798), .Y(n66739) );
  A2O1A1Ixp33_ASAP7_75t_SL U70198 ( .A1(n66241), .A2(n65032), .B(n59528), .C(
        n66301), .Y(n58810) );
  A2O1A1Ixp33_ASAP7_75t_SL U70199 ( .A1(n62913), .A2(n63366), .B(n57044), .C(
        n58477), .Y(n58815) );
  XOR2xp5_ASAP7_75t_SL U70200 ( .A(n63792), .B(n58823), .Y(n63684) );
  MAJIxp5_ASAP7_75t_SL U70201 ( .A(n63642), .B(n63643), .C(n63644), .Y(n63790)
         );
  MAJIxp5_ASAP7_75t_SL U70202 ( .A(n63198), .B(n63196), .C(n63197), .Y(n63642)
         );
  XNOR2xp5_ASAP7_75t_SL U70203 ( .A(n63850), .B(n63851), .Y(n58825) );
  OAI211xp5_ASAP7_75t_SL U70204 ( .A1(n58836), .A2(n58838), .B(n58835), .C(
        n58833), .Y(n52000) );
  NAND4xp25_ASAP7_75t_SL U70205 ( .A(n74113), .B(n59457), .C(n59252), .D(
        n58834), .Y(n58833) );
  NAND3xp33_ASAP7_75t_SL U70206 ( .A(n58839), .B(n58546), .C(n68686), .Y(
        n58835) );
  A2O1A1Ixp33_ASAP7_75t_SL U70207 ( .A1(n75470), .A2(n58881), .B(n58842), .C(
        n58840), .Y(n58841) );
  OR2x2_ASAP7_75t_SL U70208 ( .A(n58850), .B(n59659), .Y(n76133) );
  A2O1A1Ixp33_ASAP7_75t_SL U70209 ( .A1(n57180), .A2(n58851), .B(n64071), .C(
        n64070), .Y(n64347) );
  NOR3xp33_ASAP7_75t_SL U70210 ( .A(n64740), .B(n64741), .C(n58855), .Y(n58854) );
  XNOR2xp5_ASAP7_75t_SL U70211 ( .A(n57505), .B(n58861), .Y(n66957) );
  XNOR2xp5_ASAP7_75t_SL U70212 ( .A(n76028), .B(n58863), .Y(n67443) );
  XNOR2xp5_ASAP7_75t_SL U70213 ( .A(n58863), .B(n67911), .Y(n66619) );
  XNOR2xp5_ASAP7_75t_SL U70214 ( .A(n58863), .B(n67944), .Y(n67319) );
  XOR2xp5_ASAP7_75t_SL U70215 ( .A(n59283), .B(n58865), .Y(n59282) );
  NOR3xp33_ASAP7_75t_SL U70216 ( .A(n77314), .B(n77504), .C(n59157), .Y(n77799) );
  AOI211xp5_ASAP7_75t_SL U70217 ( .A1(n69160), .A2(n58538), .B(n58869), .C(
        n58868), .Y(n52012) );
  O2A1O1Ixp5_ASAP7_75t_SL U70218 ( .A1(n58871), .A2(n59659), .B(n67542), .C(
        n67541), .Y(n67543) );
  XNOR2xp5_ASAP7_75t_SL U70219 ( .A(n58877), .B(n63197), .Y(n58876) );
  MAJIxp5_ASAP7_75t_SL U70220 ( .A(n63138), .B(n63136), .C(n63137), .Y(n63197)
         );
  XNOR2xp5_ASAP7_75t_SL U70221 ( .A(n63818), .B(n63819), .Y(n63680) );
  AND2x2_ASAP7_75t_SL U70222 ( .A(n67902), .B(n67864), .Y(n67452) );
  XNOR2xp5_ASAP7_75t_SL U70223 ( .A(n63141), .B(n63140), .Y(n58888) );
  OR2x2_ASAP7_75t_SL U70224 ( .A(n58889), .B(n62685), .Y(n64920) );
  MAJIxp5_ASAP7_75t_SL U70225 ( .A(n68295), .B(n68296), .C(n68294), .Y(n68313)
         );
  OA21x2_ASAP7_75t_SL U70226 ( .A1(n57219), .A2(n62670), .B(n62672), .Y(n58892) );
  OR2x2_ASAP7_75t_SL U70227 ( .A(n59110), .B(n59109), .Y(n67805) );
  NAND3xp33_ASAP7_75t_SL U70228 ( .A(n58900), .B(n59656), .C(n58899), .Y(
        n58898) );
  AND3x1_ASAP7_75t_SL U70229 ( .A(n76430), .B(n58353), .C(n59550), .Y(n58908)
         );
  XNOR2xp5_ASAP7_75t_SL U70230 ( .A(n58414), .B(n59640), .Y(n58913) );
  A2O1A1Ixp33_ASAP7_75t_SL U70231 ( .A1(n75954), .A2(n59664), .B(
        or1200_cpu_or1200_mult_mac_n8), .C(n53275), .Y(n75955) );
  NAND3xp33_ASAP7_75t_SL U70232 ( .A(n67536), .B(n58920), .C(n58919), .Y(
        n64440) );
  OR2x2_ASAP7_75t_SL U70233 ( .A(n60737), .B(n62629), .Y(n62581) );
  AO31x2_ASAP7_75t_SL U70234 ( .A1(n68730), .A2(n59386), .A3(n59385), .B(
        n59384), .Y(n69117) );
  NAND3xp33_ASAP7_75t_SL U70235 ( .A(n66311), .B(n66312), .C(n58939), .Y(
        n66313) );
  MAJIxp5_ASAP7_75t_SL U70236 ( .A(n63109), .B(n58947), .C(n58502), .Y(n63163)
         );
  NOR3xp33_ASAP7_75t_SL U70237 ( .A(n69114), .B(n69235), .C(n68668), .Y(n58958) );
  NOR2xp33_ASAP7_75t_SL U70238 ( .A(n68648), .B(n58956), .Y(n68652) );
  XNOR2xp5_ASAP7_75t_SL U70239 ( .A(n75894), .B(n75930), .Y(n67746) );
  XNOR2xp5_ASAP7_75t_SL U70240 ( .A(n57257), .B(n59670), .Y(n66934) );
  XNOR2xp5_ASAP7_75t_SL U70241 ( .A(n59598), .B(n59670), .Y(n66473) );
  O2A1O1Ixp5_ASAP7_75t_SL U70242 ( .A1(n67601), .A2(n58962), .B(n67372), .C(
        n67371), .Y(n67612) );
  O2A1O1Ixp5_ASAP7_75t_SL U70243 ( .A1(n58478), .A2(n58962), .B(n58975), .C(
        n67609), .Y(n58974) );
  MAJx2_ASAP7_75t_SL U70244 ( .A(n58964), .B(n58459), .C(n66865), .Y(n67101)
         );
  NOR2xp33_ASAP7_75t_SL U70245 ( .A(n67561), .B(n59453), .Y(n59306) );
  OA21x2_ASAP7_75t_SL U70246 ( .A1(n62566), .A2(n62565), .B(n62567), .Y(n64504) );
  XNOR2xp5_ASAP7_75t_SL U70247 ( .A(n68454), .B(n68455), .Y(n58976) );
  MAJIxp5_ASAP7_75t_SL U70248 ( .A(n59068), .B(n67689), .C(n67688), .Y(n68357)
         );
  XOR2xp5_ASAP7_75t_SL U70249 ( .A(n62734), .B(n62731), .Y(n58983) );
  XOR2xp5_ASAP7_75t_SL U70250 ( .A(n58510), .B(n62754), .Y(n58985) );
  MAJIxp5_ASAP7_75t_SL U70251 ( .A(n63032), .B(n63031), .C(n63030), .Y(n62756)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70252 ( .A1(n59618), .A2(n53275), .B(n67925), .C(
        n67924), .Y(n67977) );
  MAJIxp5_ASAP7_75t_SL U70253 ( .A(n64907), .B(n64909), .C(n64908), .Y(n64993)
         );
  MAJIxp5_ASAP7_75t_SL U70254 ( .A(n67763), .B(n58346), .C(n67664), .Y(n68581)
         );
  MAJIxp5_ASAP7_75t_SL U70255 ( .A(n67668), .B(n67669), .C(n56833), .Y(n68393)
         );
  MAJIxp5_ASAP7_75t_SL U70256 ( .A(n67667), .B(n67665), .C(n67666), .Y(n68394)
         );
  MAJIxp5_ASAP7_75t_SL U70257 ( .A(n67577), .B(n67527), .C(n67526), .Y(n67666)
         );
  XOR2xp5_ASAP7_75t_SL U70258 ( .A(n68395), .B(n68397), .Y(n59001) );
  O2A1O1Ixp5_ASAP7_75t_SL U70259 ( .A1(n67963), .A2(n59504), .B(n63147), .C(
        n59012), .Y(n63148) );
  O2A1O1Ixp5_ASAP7_75t_SL U70260 ( .A1(n59606), .A2(n57274), .B(n63220), .C(
        n59012), .Y(n63221) );
  O2A1O1Ixp5_ASAP7_75t_SL U70261 ( .A1(n59466), .A2(n75903), .B(n64446), .C(
        n59012), .Y(n64447) );
  O2A1O1Ixp5_ASAP7_75t_SL U70262 ( .A1(n53303), .A2(n53275), .B(n58411), .C(
        n59012), .Y(n66743) );
  A2O1A1Ixp33_ASAP7_75t_SL U70263 ( .A1(n64401), .A2(n67288), .B(n63631), .C(
        n59012), .Y(n63632) );
  XOR2xp5_ASAP7_75t_SL U70264 ( .A(n68544), .B(n68543), .Y(n59013) );
  AND2x2_ASAP7_75t_SL U70265 ( .A(n58511), .B(n68550), .Y(n59014) );
  OR2x2_ASAP7_75t_SL U70266 ( .A(n58511), .B(n68550), .Y(n59015) );
  AND3x1_ASAP7_75t_SL U70267 ( .A(n61932), .B(n61930), .C(n61931), .Y(n59018)
         );
  AO21x1_ASAP7_75t_SL U70268 ( .A1(n59024), .A2(n59022), .B(n59023), .Y(n68427) );
  MAJIxp5_ASAP7_75t_SL U70269 ( .A(n59021), .B(n68428), .C(n68429), .Y(n68493)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70270 ( .A1(n59203), .A2(n68430), .B(n58364), .C(
        n59026), .Y(n59025) );
  NAND3xp33_ASAP7_75t_SL U70271 ( .A(n68431), .B(n68432), .C(n68434), .Y(
        n59026) );
  MAJIxp5_ASAP7_75t_SL U70272 ( .A(n68492), .B(n68491), .C(n68493), .Y(n68519)
         );
  NOR2xp33_ASAP7_75t_SL U70273 ( .A(n67962), .B(n59601), .Y(n67385) );
  AND2x2_ASAP7_75t_SL U70274 ( .A(n77722), .B(n74787), .Y(n64951) );
  NOR4xp25_ASAP7_75t_SL U70275 ( .A(n67838), .B(n59055), .C(n53207), .D(n59596), .Y(n67840) );
  NOR2xp33_ASAP7_75t_SL U70276 ( .A(n68336), .B(n59294), .Y(n59056) );
  XNOR2xp5_ASAP7_75t_SL U70277 ( .A(n67657), .B(n59279), .Y(n59058) );
  MAJIxp5_ASAP7_75t_SL U70278 ( .A(n59061), .B(n68049), .C(n68050), .Y(n68051)
         );
  NOR2xp33_ASAP7_75t_SL U70279 ( .A(n59062), .B(n68804), .Y(n59344) );
  AND2x2_ASAP7_75t_SL U70280 ( .A(n59066), .B(n68325), .Y(n68331) );
  OR2x2_ASAP7_75t_SL U70281 ( .A(n59066), .B(n68325), .Y(n68333) );
  O2A1O1Ixp5_ASAP7_75t_SL U70282 ( .A1(n59556), .A2(n57120), .B(n60766), .C(
        n59069), .Y(n60770) );
  NAND3xp33_ASAP7_75t_SL U70283 ( .A(n60644), .B(n59080), .C(n62561), .Y(
        n61858) );
  A2O1A1Ixp33_ASAP7_75t_SL U70284 ( .A1(n61336), .A2(n57318), .B(n59080), .C(
        n60670), .Y(n60620) );
  MAJIxp5_ASAP7_75t_SL U70285 ( .A(n59266), .B(n68352), .C(n59081), .Y(n68579)
         );
  MAJIxp5_ASAP7_75t_SL U70286 ( .A(n68037), .B(n68035), .C(n68036), .Y(n68038)
         );
  MAJIxp5_ASAP7_75t_SL U70287 ( .A(n66908), .B(n59085), .C(n66910), .Y(n68547)
         );
  XNOR2xp5_ASAP7_75t_SL U70288 ( .A(n66778), .B(n66779), .Y(n59086) );
  XNOR2xp5_ASAP7_75t_SL U70289 ( .A(n64585), .B(n64584), .Y(n59087) );
  OR2x2_ASAP7_75t_SL U70290 ( .A(n67109), .B(n67110), .Y(n69147) );
  MAJIxp5_ASAP7_75t_SL U70291 ( .A(n67324), .B(n67325), .C(n67783), .Y(n59131)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70292 ( .A1(n67395), .A2(n67394), .B(n67393), .C(
        n67396), .Y(n67790) );
  NAND3xp33_ASAP7_75t_SL U70293 ( .A(n58429), .B(n67397), .C(n58370), .Y(
        n59093) );
  NOR3xp33_ASAP7_75t_SL U70294 ( .A(n67379), .B(n67378), .C(n59114), .Y(n67380) );
  OR2x2_ASAP7_75t_SL U70295 ( .A(n58464), .B(n66640), .Y(n66651) );
  A2O1A1Ixp33_ASAP7_75t_SL U70296 ( .A1(n57108), .A2(n67432), .B(n64397), .C(
        n59506), .Y(n64398) );
  XNOR2xp5_ASAP7_75t_SL U70297 ( .A(n59602), .B(n67736), .Y(n67473) );
  OR3x1_ASAP7_75t_SL U70298 ( .A(n59662), .B(n66860), .C(n59142), .Y(n59143)
         );
  XNOR2xp5_ASAP7_75t_SL U70299 ( .A(n68375), .B(n68373), .Y(n67745) );
  XOR2xp5_ASAP7_75t_SL U70300 ( .A(n68471), .B(n68468), .Y(n59151) );
  MAJIxp5_ASAP7_75t_SL U70301 ( .A(n64708), .B(n64706), .C(n64707), .Y(n64714)
         );
  XNOR2xp5_ASAP7_75t_SL U70302 ( .A(n59152), .B(n59153), .Y(n64724) );
  XOR2xp5_ASAP7_75t_SL U70303 ( .A(n64721), .B(n64722), .Y(n59152) );
  NAND3xp33_ASAP7_75t_SL U70304 ( .A(n59596), .B(n67837), .C(n59436), .Y(
        n59169) );
  XOR2xp5_ASAP7_75t_SL U70305 ( .A(n67005), .B(n67056), .Y(n59170) );
  AND2x2_ASAP7_75t_SL U70306 ( .A(n59555), .B(n59588), .Y(n62804) );
  XOR2xp5_ASAP7_75t_SL U70307 ( .A(n66771), .B(n66770), .Y(n59173) );
  MAJIxp5_ASAP7_75t_SL U70308 ( .A(n68042), .B(n68043), .C(n68045), .Y(n68054)
         );
  MAJIxp5_ASAP7_75t_SL U70309 ( .A(n67940), .B(n67648), .C(n67942), .Y(n68045)
         );
  AO31x2_ASAP7_75t_SL U70310 ( .A1(n64081), .A2(n57271), .A3(n77709), .B(
        n59187), .Y(n76091) );
  OR2x2_ASAP7_75t_SL U70311 ( .A(n57122), .B(n63129), .Y(n64081) );
  OR2x2_ASAP7_75t_SL U70312 ( .A(n59605), .B(n67909), .Y(n67580) );
  OR2x2_ASAP7_75t_SL U70313 ( .A(n59193), .B(n66705), .Y(n66988) );
  XNOR2xp5_ASAP7_75t_SL U70314 ( .A(n66874), .B(n66875), .Y(n59194) );
  MAJIxp5_ASAP7_75t_SL U70315 ( .A(n64964), .B(n64963), .C(n64962), .Y(n65002)
         );
  AOI211xp5_ASAP7_75t_SL U70316 ( .A1(n69308), .A2(n68662), .B(n59212), .C(
        n59213), .Y(n51988) );
  MAJIxp5_ASAP7_75t_SL U70317 ( .A(n66614), .B(n59237), .C(n66736), .Y(n66833)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70318 ( .A1(n58512), .A2(n64537), .B(n64600), .C(
        n57154), .Y(n59240) );
  XOR2xp5_ASAP7_75t_SL U70319 ( .A(n57058), .B(n68467), .Y(n68478) );
  NAND3xp33_ASAP7_75t_SL U70320 ( .A(n62768), .B(n62767), .C(n59456), .Y(
        n62773) );
  OR2x2_ASAP7_75t_SL U70321 ( .A(n59656), .B(n59605), .Y(n62725) );
  XNOR2xp5_ASAP7_75t_SL U70322 ( .A(n58393), .B(n64872), .Y(n59248) );
  O2A1O1Ixp5_ASAP7_75t_SL U70323 ( .A1(n67717), .A2(n67716), .B(n67715), .C(
        n67714), .Y(n68385) );
  NAND3xp33_ASAP7_75t_SL U70324 ( .A(n59259), .B(n59423), .C(n58480), .Y(
        n59261) );
  XOR2xp5_ASAP7_75t_SL U70325 ( .A(n68556), .B(n68555), .Y(n59267) );
  MAJIxp5_ASAP7_75t_SL U70326 ( .A(n68498), .B(n68497), .C(n68499), .Y(n68529)
         );
  MAJIxp5_ASAP7_75t_SL U70327 ( .A(n68448), .B(n68449), .C(n68447), .Y(n68499)
         );
  OR2x2_ASAP7_75t_SL U70328 ( .A(n75106), .B(n75080), .Y(n59273) );
  NAND3xp33_ASAP7_75t_SL U70329 ( .A(n59102), .B(n67705), .C(n67706), .Y(
        n59293) );
  OR2x2_ASAP7_75t_SL U70330 ( .A(n76049), .B(n59641), .Y(n67706) );
  A2O1A1Ixp33_ASAP7_75t_SL U70331 ( .A1(n56827), .A2(n68010), .B(n57104), .C(
        n68009), .Y(n59315) );
  MAJIxp5_ASAP7_75t_SL U70332 ( .A(n67659), .B(n67661), .C(n67660), .Y(n67757)
         );
  MAJIxp5_ASAP7_75t_SL U70333 ( .A(n67654), .B(n67653), .C(n67652), .Y(n67661)
         );
  XOR2xp5_ASAP7_75t_SL U70334 ( .A(n58511), .B(n68550), .Y(n68536) );
  MAJIxp5_ASAP7_75t_SL U70335 ( .A(n68500), .B(n68501), .C(n68502), .Y(n68535)
         );
  OR2x2_ASAP7_75t_SL U70336 ( .A(n77730), .B(n64648), .Y(n67356) );
  NAND3xp33_ASAP7_75t_SL U70337 ( .A(n57333), .B(n59438), .C(n59336), .Y(
        n60669) );
  OR2x2_ASAP7_75t_SL U70338 ( .A(n75897), .B(n68098), .Y(n59407) );
  NAND3xp33_ASAP7_75t_SL U70339 ( .A(n59361), .B(n56838), .C(n62577), .Y(
        n62578) );
  O2A1O1Ixp5_ASAP7_75t_SL U70340 ( .A1(n68263), .A2(n68262), .B(n68261), .C(
        n68260), .Y(n59363) );
  AND2x2_ASAP7_75t_SL U70341 ( .A(n59364), .B(n64047), .Y(n59369) );
  XOR2xp5_ASAP7_75t_SL U70342 ( .A(n68167), .B(n68166), .Y(n59372) );
  O2A1O1Ixp5_ASAP7_75t_SL U70343 ( .A1(n75947), .A2(n58440), .B(n59373), .C(
        n65018), .Y(n68166) );
  NAND3xp33_ASAP7_75t_SL U70344 ( .A(n59382), .B(n68916), .C(n68972), .Y(
        n59386) );
  OR2x2_ASAP7_75t_SL U70345 ( .A(n68517), .B(n68516), .Y(n68972) );
  NAND3xp33_ASAP7_75t_SL U70346 ( .A(n69029), .B(n69028), .C(n69026), .Y(
        n59384) );
  OR2x2_ASAP7_75t_SL U70347 ( .A(n66261), .B(n66270), .Y(n66280) );
  AND2x2_ASAP7_75t_SL U70348 ( .A(n59398), .B(n59646), .Y(n61438) );
  O2A1O1Ixp5_ASAP7_75t_SL U70349 ( .A1(n64343), .A2(n64342), .B(n64341), .C(
        n59410), .Y(n64431) );
  XNOR2xp5_ASAP7_75t_SL U70350 ( .A(n58863), .B(n59662), .Y(n59417) );
  OA21x2_ASAP7_75t_SL U70351 ( .A1(n59419), .A2(n62657), .B(n62656), .Y(n59418) );
  HB1xp67_ASAP7_75t_SL U70352 ( .A(dbg_is_o[0]), .Y(dbg_is_o[1]) );
  NOR2xp33_ASAP7_75t_SL U70353 ( .A(n67230), .B(n53288), .Y(n67238) );
  NOR2xp33_ASAP7_75t_SL U70354 ( .A(n57365), .B(n68104), .Y(n66380) );
  XNOR2xp5_ASAP7_75t_SL U70355 ( .A(n63836), .B(n63835), .Y(n63837) );
  NOR2xp33_ASAP7_75t_SL U70356 ( .A(n59641), .B(n66758), .Y(n66359) );
  O2A1O1Ixp5_ASAP7_75t_SL U70357 ( .A1(n59618), .A2(n76028), .B(n62837), .C(
        n62836), .Y(n62934) );
  NOR2xp33_ASAP7_75t_SL U70358 ( .A(n59434), .B(n68740), .Y(n68739) );
  NOR2xp33_ASAP7_75t_SL U70359 ( .A(n68078), .B(n59659), .Y(n68082) );
  NAND2xp33_ASAP7_75t_SRAM U70360 ( .A(n58384), .B(n67736), .Y(n66855) );
  NOR2xp33_ASAP7_75t_SL U70361 ( .A(n58383), .B(n68087), .Y(n67240) );
  AND2x2_ASAP7_75t_SL U70362 ( .A(n77242), .B(n57117), .Y(n59476) );
  AOI31xp33_ASAP7_75t_SL U70363 ( .A1(n66315), .A2(n66314), .A3(n66313), .B(
        n75033), .Y(n68408) );
  NOR2xp33_ASAP7_75t_SL U70364 ( .A(n66806), .B(n66805), .Y(n66807) );
  NOR2xp33_ASAP7_75t_SL U70365 ( .A(n76028), .B(n65043), .Y(n62979) );
  AOI211xp5_ASAP7_75t_SL U70366 ( .A1(n57110), .A2(n76028), .B(n62743), .C(
        n68079), .Y(n62744) );
  NOR2xp33_ASAP7_75t_SL U70367 ( .A(n76028), .B(n67866), .Y(n62585) );
  NOR2xp33_ASAP7_75t_SL U70368 ( .A(n76028), .B(n59615), .Y(n62743) );
  NOR4xp25_ASAP7_75t_SL U70369 ( .A(n57500), .B(n59552), .C(n59551), .D(n57312), .Y(n75481) );
  NOR2xp33_ASAP7_75t_SL U70370 ( .A(n68158), .B(n59453), .Y(n68089) );
  NOR2xp33_ASAP7_75t_SL U70371 ( .A(n57333), .B(n60642), .Y(n60625) );
  NOR2xp33_ASAP7_75t_SL U70372 ( .A(n57333), .B(n60615), .Y(n60645) );
  AOI31xp33_ASAP7_75t_SL U70373 ( .A1(n68744), .A2(n59434), .A3(n68742), .B(
        n68741), .Y(n68747) );
  AND2x2_ASAP7_75t_SL U70374 ( .A(n77833), .B(n77359), .Y(n59495) );
  AND2x2_ASAP7_75t_SL U70375 ( .A(n77833), .B(n77359), .Y(n59496) );
  OR2x2_ASAP7_75t_SL U70376 ( .A(n77414), .B(n3100), .Y(n61281) );
  NAND3xp33_ASAP7_75t_SL U70377 ( .A(n76615), .B(n59716), .C(n76200), .Y(
        n59717) );
  O2A1O1Ixp5_ASAP7_75t_SL U70378 ( .A1(n76859), .A2(n76861), .B(n76860), .C(
        n59717), .Y(n59718) );
  OR2x2_ASAP7_75t_SL U70379 ( .A(n2131), .B(n59571), .Y(n76636) );
  NAND3xp33_ASAP7_75t_SL U70380 ( .A(n59722), .B(n75774), .C(n75775), .Y(
        n59847) );
  A2O1A1Ixp33_ASAP7_75t_SL U70381 ( .A1(n75777), .A2(n75778), .B(n59847), .C(
        n59725), .Y(n59726) );
  OR2x2_ASAP7_75t_SL U70382 ( .A(n1888), .B(n59561), .Y(n59764) );
  XNOR2xp5_ASAP7_75t_SL U70383 ( .A(or1200_dc_top_tag_11_), .B(n75618), .Y(
        n59730) );
  XNOR2xp5_ASAP7_75t_SL U70384 ( .A(n59731), .B(n59730), .Y(n59736) );
  XNOR2xp5_ASAP7_75t_SL U70385 ( .A(n59734), .B(n59733), .Y(n59735) );
  AO21x1_ASAP7_75t_SL U70386 ( .A1(n59737), .A2(n59866), .B(n75196), .Y(n59739) );
  XNOR2xp5_ASAP7_75t_SL U70387 ( .A(n59739), .B(n59738), .Y(n59744) );
  AO21x1_ASAP7_75t_SL U70388 ( .A1(n59740), .A2(n59926), .B(n77148), .Y(n59742) );
  XNOR2xp5_ASAP7_75t_SL U70389 ( .A(or1200_dc_top_tag_3_), .B(n77147), .Y(
        n59741) );
  XNOR2xp5_ASAP7_75t_SL U70390 ( .A(n59742), .B(n59741), .Y(n59743) );
  NOR3xp33_ASAP7_75t_SL U70391 ( .A(n59745), .B(n59744), .C(n59743), .Y(n59786) );
  OR2x2_ASAP7_75t_SL U70392 ( .A(n1903), .B(n59531), .Y(n59856) );
  NOR3xp33_ASAP7_75t_SL U70393 ( .A(n59747), .B(or1200_dc_top_tag_8_), .C(
        n59794), .Y(n59746) );
  O2A1O1Ixp5_ASAP7_75t_SL U70394 ( .A1(n59794), .A2(n59747), .B(
        or1200_dc_top_tag_8_), .C(n59746), .Y(n59759) );
  OR2x2_ASAP7_75t_SL U70395 ( .A(n1891), .B(n57377), .Y(n59852) );
  OR2x2_ASAP7_75t_SL U70396 ( .A(n1876), .B(n59576), .Y(n59775) );
  OR2x2_ASAP7_75t_SL U70397 ( .A(n1882), .B(n59528), .Y(n59865) );
  O2A1O1Ixp5_ASAP7_75t_SL U70398 ( .A1(n59759), .A2(n59758), .B(n59757), .C(
        n59756), .Y(n59785) );
  OR2x2_ASAP7_75t_SL U70399 ( .A(n1912), .B(n59529), .Y(n59798) );
  NOR3xp33_ASAP7_75t_SL U70400 ( .A(n59762), .B(n69362), .C(
        or1200_dc_top_tag_14_), .Y(n59761) );
  O2A1O1Ixp5_ASAP7_75t_SL U70401 ( .A1(n69362), .A2(n59762), .B(
        or1200_dc_top_tag_14_), .C(n59761), .Y(n59771) );
  AO21x1_ASAP7_75t_SL U70402 ( .A1(n59765), .A2(n75441), .B(n75439), .Y(n59766) );
  O2A1O1Ixp5_ASAP7_75t_SL U70403 ( .A1(n59771), .A2(n69365), .B(n59770), .C(
        n59769), .Y(n59784) );
  NOR3xp33_ASAP7_75t_SL U70404 ( .A(n59773), .B(n75189), .C(
        or1200_dc_top_tag_16_), .Y(n59772) );
  O2A1O1Ixp5_ASAP7_75t_SL U70405 ( .A1(n59773), .A2(n75189), .B(
        or1200_dc_top_tag_16_), .C(n59772), .Y(n59782) );
  XNOR2xp5_ASAP7_75t_SL U70406 ( .A(n60207), .B(n59779), .Y(n59780) );
  O2A1O1Ixp5_ASAP7_75t_SL U70407 ( .A1(n59782), .A2(n77174), .B(n59781), .C(
        n59780), .Y(n59783) );
  NAND4xp25_ASAP7_75t_SL U70408 ( .A(n59786), .B(n59785), .C(n59784), .D(
        n59783), .Y(n59835) );
  XNOR2xp5_ASAP7_75t_SL U70409 ( .A(n59790), .B(n59789), .Y(n59805) );
  OR2x2_ASAP7_75t_SL U70410 ( .A(n2056), .B(n59538), .Y(n77015) );
  XNOR2xp5_ASAP7_75t_SL U70411 ( .A(n59792), .B(n59791), .Y(n59804) );
  OR2x2_ASAP7_75t_SL U70412 ( .A(n1894), .B(n59533), .Y(n74122) );
  XNOR2xp5_ASAP7_75t_SL U70413 ( .A(n59796), .B(n59795), .Y(n59803) );
  XNOR2xp5_ASAP7_75t_SL U70414 ( .A(n59801), .B(n59800), .Y(n59802) );
  NAND4xp25_ASAP7_75t_SL U70415 ( .A(n59805), .B(n59804), .C(n59803), .D(
        n59802), .Y(n59834) );
  NOR3xp33_ASAP7_75t_SL U70416 ( .A(n59807), .B(or1200_dc_top_tag_12_), .C(
        n69356), .Y(n59806) );
  XNOR2xp5_ASAP7_75t_SL U70417 ( .A(n74043), .B(n59808), .Y(n59832) );
  NAND3xp33_ASAP7_75t_SL U70418 ( .A(n59812), .B(n59813), .C(n59811), .Y(
        n59810) );
  A2O1A1Ixp33_ASAP7_75t_SL U70419 ( .A1(n59813), .A2(n59812), .B(n59811), .C(
        n59810), .Y(n59814) );
  XNOR2xp5_ASAP7_75t_SL U70420 ( .A(n77223), .B(n59814), .Y(n59831) );
  NAND3xp33_ASAP7_75t_SL U70421 ( .A(n59819), .B(n59817), .C(n59818), .Y(
        n59816) );
  A2O1A1Ixp33_ASAP7_75t_SL U70422 ( .A1(n59819), .A2(n59818), .B(n59817), .C(
        n59816), .Y(n59820) );
  XNOR2xp5_ASAP7_75t_SL U70423 ( .A(n74982), .B(n59820), .Y(n59830) );
  NAND3xp33_ASAP7_75t_SL U70424 ( .A(n59826), .B(n59825), .C(n59824), .Y(
        n59823) );
  A2O1A1Ixp33_ASAP7_75t_SL U70425 ( .A1(n59826), .A2(n59825), .B(n59824), .C(
        n59823), .Y(n59827) );
  XNOR2xp5_ASAP7_75t_SL U70426 ( .A(n59828), .B(n59827), .Y(n59829) );
  NAND4xp25_ASAP7_75t_SL U70427 ( .A(n59832), .B(n59831), .C(n59830), .D(
        n59829), .Y(n59833) );
  NOR3xp33_ASAP7_75t_SL U70428 ( .A(n59835), .B(n59834), .C(n59833), .Y(n59836) );
  A2O1A1Ixp33_ASAP7_75t_SL U70429 ( .A1(n77292), .A2(n77293), .B(
        or1200_dc_top_tag_0_), .C(n59836), .Y(n59837) );
  NAND3xp33_ASAP7_75t_SL U70430 ( .A(n75442), .B(n78090), .C(n69355), .Y(
        n69363) );
  NAND3xp33_ASAP7_75t_SL U70431 ( .A(n75673), .B(n60198), .C(n60207), .Y(
        n59874) );
  OR2x2_ASAP7_75t_SL U70432 ( .A(n3109), .B(n3107), .Y(n60192) );
  OR2x2_ASAP7_75t_SL U70433 ( .A(n3092), .B(n77473), .Y(n77410) );
  OR2x2_ASAP7_75t_SL U70434 ( .A(n60192), .B(n4320), .Y(n60583) );
  NAND4xp25_ASAP7_75t_SL U70435 ( .A(n61998), .B(n3084), .C(n3111), .D(n77763), 
        .Y(n78000) );
  NAND2xp5_ASAP7_75t_SL U70436 ( .A(dc_en), .B(n78000), .Y(n59878) );
  NAND3xp33_ASAP7_75t_SL U70437 ( .A(n59877), .B(n78184), .C(n61317), .Y(
        n59885) );
  NAND4xp25_ASAP7_75t_SL U70438 ( .A(n60583), .B(n60199), .C(n60191), .D(
        n77429), .Y(n59880) );
  NOR3xp33_ASAP7_75t_SL U70439 ( .A(n75673), .B(n59886), .C(n60196), .Y(n59882) );
  NAND3xp33_ASAP7_75t_SL U70440 ( .A(n59884), .B(n60213), .C(n60212), .Y(
        n61294) );
  O2A1O1Ixp5_ASAP7_75t_SL U70441 ( .A1(n59888), .A2(n61289), .B(n61290), .C(
        n59887), .Y(n59889) );
  OR2x2_ASAP7_75t_SL U70442 ( .A(n3074), .B(n77410), .Y(n77686) );
  OR2x2_ASAP7_75t_SL U70443 ( .A(or1200_cpu_or1200_except_n552), .B(
        or1200_cpu_or1200_except_n555), .Y(n62568) );
  A2O1A1Ixp33_ASAP7_75t_SL U70444 ( .A1(n56968), .A2(n62570), .B(n62568), .C(
        n1753), .Y(n62002) );
  O2A1O1Ixp5_ASAP7_75t_SL U70445 ( .A1(n59925), .A2(n62002), .B(n77581), .C(
        n64282), .Y(n61131) );
  OR2x2_ASAP7_75t_SL U70446 ( .A(dbg_adr_i[13]), .B(n78439), .Y(n59929) );
  NAND3xp33_ASAP7_75t_SL U70447 ( .A(n75687), .B(n60549), .C(n77966), .Y(
        n59944) );
  NAND3xp33_ASAP7_75t_SL U70448 ( .A(n61243), .B(n60552), .C(n77994), .Y(
        n60559) );
  OAI31xp33_ASAP7_75t_SL U70449 ( .A1(n59965), .A2(n77370), .A3(n59964), .B(
        n60317), .Y(n59966) );
  A2O1A1Ixp33_ASAP7_75t_SL U70450 ( .A1(n77621), .A2(n59972), .B(n62319), .C(
        n61248), .Y(n77663) );
  NAND3xp33_ASAP7_75t_SL U70451 ( .A(n59989), .B(n60002), .C(n751), .Y(n60000)
         );
  OR2x2_ASAP7_75t_SL U70452 ( .A(n75143), .B(n77210), .Y(n60017) );
  A2O1A1Ixp33_ASAP7_75t_SL U70453 ( .A1(n60001), .A2(n60000), .B(n76821), .C(
        n59999), .Y(n77382) );
  XNOR2xp5_ASAP7_75t_SL U70454 ( .A(n60002), .B(n60014), .Y(n60008) );
  A2O1A1Ixp33_ASAP7_75t_SL U70455 ( .A1(n60008), .A2(n74956), .B(n60007), .C(
        n57100), .Y(n4097) );
  A2O1A1Ixp33_ASAP7_75t_SL U70456 ( .A1(n60015), .A2(n60014), .B(n60013), .C(
        n57100), .Y(n4099) );
  A2O1A1Ixp33_ASAP7_75t_SL U70457 ( .A1(n60024), .A2(n60023), .B(n60022), .C(
        n57100), .Y(n4101) );
  A2O1A1Ixp33_ASAP7_75t_SL U70458 ( .A1(n60030), .A2(n60029), .B(n60028), .C(
        n57100), .Y(n4103) );
  A2O1A1Ixp33_ASAP7_75t_SL U70459 ( .A1(n60036), .A2(n60035), .B(n60034), .C(
        n57100), .Y(n4106) );
  XNOR2xp5_ASAP7_75t_SL U70460 ( .A(n773), .B(icqmem_adr_qmem[26]), .Y(n60089)
         );
  OAI211xp5_ASAP7_75t_SL U70461 ( .A1(n57068), .A2(n57124), .B(n60038), .C(
        n60037), .Y(n60039) );
  A2O1A1Ixp33_ASAP7_75t_SL U70462 ( .A1(n60040), .A2(n74956), .B(n60039), .C(
        n57100), .Y(n4110) );
  XNOR2xp5_ASAP7_75t_SL U70463 ( .A(n781), .B(icqmem_adr_qmem[24]), .Y(n60088)
         );
  OR2x2_ASAP7_75t_SL U70464 ( .A(n1084), .B(n59703), .Y(n61268) );
  A2O1A1Ixp33_ASAP7_75t_SL U70465 ( .A1(n60050), .A2(n60049), .B(n60156), .C(
        n60048), .Y(n60051) );
  XOR2xp5_ASAP7_75t_SL U70466 ( .A(icqmem_adr_qmem[13]), .B(n825), .Y(n60086)
         );
  OAI211xp5_ASAP7_75t_SL U70467 ( .A1(n60054), .A2(n60053), .B(n60079), .C(
        n60174), .Y(n60057) );
  OAI211xp5_ASAP7_75t_SL U70468 ( .A1(n3003), .A2(n74953), .B(n60057), .C(
        n60056), .Y(n60058) );
  XOR2xp5_ASAP7_75t_SL U70469 ( .A(icqmem_adr_qmem[22]), .B(n789), .Y(n60085)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70470 ( .A1(n60147), .A2(n60067), .B(n60066), .C(
        n60065), .Y(n60068) );
  XOR2xp5_ASAP7_75t_SL U70471 ( .A(n793), .B(icqmem_adr_qmem[21]), .Y(n60084)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70472 ( .A1(n60079), .A2(n60078), .B(n60077), .C(
        n60076), .Y(n60080) );
  XOR2xp5_ASAP7_75t_SL U70473 ( .A(icqmem_adr_qmem[23]), .B(n785), .Y(n60083)
         );
  NAND4xp25_ASAP7_75t_SL U70474 ( .A(n60086), .B(n60085), .C(n60084), .D(
        n60083), .Y(n60087) );
  NOR3xp33_ASAP7_75t_SL U70475 ( .A(n60089), .B(n60088), .C(n60087), .Y(n60186) );
  NAND3xp33_ASAP7_75t_SL U70476 ( .A(n60156), .B(n74956), .C(n60157), .Y(
        n60098) );
  A2O1A1Ixp33_ASAP7_75t_SL U70477 ( .A1(n60098), .A2(n60097), .B(n60116), .C(
        n60096), .Y(n60099) );
  XOR2xp5_ASAP7_75t_SL U70478 ( .A(icqmem_adr_qmem[15]), .B(n817), .Y(n60107)
         );
  OAI211xp5_ASAP7_75t_SL U70479 ( .A1(n61162), .A2(n77429), .B(n60107), .C(
        n60106), .Y(n60123) );
  OAI211xp5_ASAP7_75t_SL U70480 ( .A1(n3018), .A2(n74953), .B(n60112), .C(
        n60111), .Y(n60113) );
  XNOR2xp5_ASAP7_75t_SL U70481 ( .A(n809), .B(icqmem_adr_qmem[17]), .Y(n60122)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70482 ( .A1(n60116), .A2(n74956), .B(n60115), .C(
        n60114), .Y(n60119) );
  OAI211xp5_ASAP7_75t_SL U70483 ( .A1(n3021), .A2(n74953), .B(n60119), .C(
        n60118), .Y(n60120) );
  XNOR2xp5_ASAP7_75t_SL U70484 ( .A(n813), .B(icqmem_adr_qmem[16]), .Y(n60121)
         );
  NOR3xp33_ASAP7_75t_SL U70485 ( .A(n60123), .B(n60122), .C(n60121), .Y(n60185) );
  A2O1A1Ixp33_ASAP7_75t_SL U70486 ( .A1(n60132), .A2(n60131), .B(n60149), .C(
        n60130), .Y(n60133) );
  XNOR2xp5_ASAP7_75t_SL U70487 ( .A(n801), .B(icqmem_adr_qmem[19]), .Y(n60170)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70488 ( .A1(n60142), .A2(n74956), .B(n60141), .C(
        n60140), .Y(n60143) );
  A2O1A1Ixp33_ASAP7_75t_SL U70489 ( .A1(n60149), .A2(n74956), .B(n60148), .C(
        n60147), .Y(n60152) );
  OAI211xp5_ASAP7_75t_SL U70490 ( .A1(n3009), .A2(n74953), .B(n60152), .C(
        n60151), .Y(n60153) );
  XNOR2xp5_ASAP7_75t_SL U70491 ( .A(n797), .B(icqmem_adr_qmem[20]), .Y(n60168)
         );
  XNOR2xp5_ASAP7_75t_SL U70492 ( .A(n60157), .B(n60156), .Y(n60164) );
  XNOR2xp5_ASAP7_75t_SL U70493 ( .A(n821), .B(icqmem_adr_qmem[14]), .Y(n60167)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70494 ( .A1(n775), .A2(n60182), .B(n60181), .C(
        n60180), .Y(n65192) );
  OR2x2_ASAP7_75t_SL U70495 ( .A(n3105), .B(n61287), .Y(n61999) );
  NOR3xp33_ASAP7_75t_SL U70496 ( .A(n60202), .B(n60194), .C(n60197), .Y(n60195) );
  NAND3xp33_ASAP7_75t_SL U70497 ( .A(n61999), .B(n60199), .C(n60294), .Y(
        n60203) );
  A2O1A1Ixp33_ASAP7_75t_SL U70498 ( .A1(n53449), .A2(n60207), .B(n60206), .C(
        n60205), .Y(n60219) );
  NOR3xp33_ASAP7_75t_SL U70499 ( .A(n60219), .B(n60305), .C(n77208), .Y(n60215) );
  NAND3xp33_ASAP7_75t_SL U70500 ( .A(n60668), .B(n60644), .C(n62561), .Y(
        n76327) );
  AND2x2_ASAP7_75t_SL U70501 ( .A(dbg_stb_i), .B(dbg_adr_i[1]), .Y(n60224) );
  A2O1A1Ixp33_ASAP7_75t_SL U70502 ( .A1(n73963), .A2(n78260), .B(
        or1200_cpu_to_sr[1]), .C(n60234), .Y(n75767) );
  NAND3xp33_ASAP7_75t_SL U70503 ( .A(n60258), .B(n60257), .C(n60256), .Y(
        n60259) );
  NAND3xp33_ASAP7_75t_SL U70504 ( .A(n75770), .B(n2798), .C(n75769), .Y(n74936) );
  OR2x2_ASAP7_75t_SL U70505 ( .A(n77501), .B(n22057), .Y(n60287) );
  AND3x1_ASAP7_75t_SL U70506 ( .A(n62148), .B(or1200_cpu_or1200_except_n116), 
        .C(n60300), .Y(n60303) );
  NAND3xp33_ASAP7_75t_SL U70507 ( .A(n57160), .B(or1200_cpu_or1200_except_n116), .C(n3119), .Y(n60420) );
  OR2x2_ASAP7_75t_SL U70508 ( .A(n3121), .B(n59703), .Y(n77368) );
  INVx1_ASAP7_75t_SL U70509 ( .A(iwb_dat_i[28]), .Y(n60313) );
  OA21x2_ASAP7_75t_SL U70510 ( .A1(n60315), .A2(n77954), .B(n60314), .Y(n77839) );
  INVx1_ASAP7_75t_SL U70511 ( .A(iwb_dat_i[26]), .Y(n60316) );
  OR2x2_ASAP7_75t_SL U70512 ( .A(n60421), .B(n60325), .Y(n69330) );
  OA21x2_ASAP7_75t_SL U70513 ( .A1(n60323), .A2(n77954), .B(n60322), .Y(n61037) );
  INVx1_ASAP7_75t_SL U70514 ( .A(iwb_dat_i[27]), .Y(n60331) );
  AND2x2_ASAP7_75t_SL U70515 ( .A(n77833), .B(n77359), .Y(n78021) );
  NAND3xp33_ASAP7_75t_SL U70516 ( .A(n61136), .B(n61145), .C(n2609), .Y(n60722) );
  AO21x1_ASAP7_75t_SL U70517 ( .A1(n60722), .A2(n60333), .B(n60501), .Y(n60341) );
  AND3x1_ASAP7_75t_SL U70518 ( .A(n61155), .B(n60369), .C(n61028), .Y(n60360)
         );
  OR3x1_ASAP7_75t_SL U70519 ( .A(n77426), .B(n2616), .C(n61145), .Y(n62022) );
  OAI211xp5_ASAP7_75t_SL U70520 ( .A1(n60350), .A2(n77379), .B(n60349), .C(
        n60348), .Y(n9603) );
  NOR3xp33_ASAP7_75t_SL U70521 ( .A(n62144), .B(n61154), .C(n77426), .Y(n60491) );
  OAI211xp5_ASAP7_75t_SL U70522 ( .A1(n60357), .A2(n77379), .B(n60356), .C(
        n60355), .Y(n9602) );
  NAND3xp33_ASAP7_75t_SL U70523 ( .A(n60360), .B(n62142), .C(n61145), .Y(
        n60361) );
  OAI211xp5_ASAP7_75t_SL U70524 ( .A1(n60368), .A2(n77379), .B(n60367), .C(
        n60366), .Y(n9605) );
  NAND3xp33_ASAP7_75t_SL U70525 ( .A(n62142), .B(n61312), .C(n61028), .Y(
        n60503) );
  OAI211xp5_ASAP7_75t_SL U70526 ( .A1(n3390), .A2(n60382), .B(n60372), .C(
        n60371), .Y(n9239) );
  OAI211xp5_ASAP7_75t_SL U70527 ( .A1(n60378), .A2(n77379), .B(n60377), .C(
        n60376), .Y(n9604) );
  NAND3xp33_ASAP7_75t_SL U70528 ( .A(n61155), .B(n77425), .C(n60379), .Y(
        n60381) );
  OAI211xp5_ASAP7_75t_SL U70529 ( .A1(n2517), .A2(n60382), .B(n60381), .C(
        n60380), .Y(n9238) );
  OAI211xp5_ASAP7_75t_SL U70530 ( .A1(n60388), .A2(n77379), .B(n60387), .C(
        n60386), .Y(n9598) );
  OAI211xp5_ASAP7_75t_SL U70531 ( .A1(n60394), .A2(n77379), .B(n60393), .C(
        n60392), .Y(n9597) );
  OAI211xp5_ASAP7_75t_SL U70532 ( .A1(n60400), .A2(n77379), .B(n60399), .C(
        n60398), .Y(n9596) );
  AOI21xp5_ASAP7_75t_SL U70533 ( .A1(n59495), .A2(iwb_dat_i[22]), .B(n60405), 
        .Y(n2698) );
  A2O1A1Ixp33_ASAP7_75t_SL U70534 ( .A1(n77376), .A2(n62469), .B(n60408), .C(
        n60407), .Y(n60409) );
  OAI211xp5_ASAP7_75t_SL U70535 ( .A1(n60415), .A2(n77379), .B(n60414), .C(
        n60413), .Y(n9582) );
  NAND2xp5_ASAP7_75t_SL U70536 ( .A(iwb_dat_i[21]), .B(n59495), .Y(n60419) );
  A2O1A1Ixp33_ASAP7_75t_SL U70537 ( .A1(n60427), .A2(n76847), .B(n60426), .C(
        n60425), .Y(n60431) );
  INVx1_ASAP7_75t_SL U70538 ( .A(iwb_dat_i[30]), .Y(n60434) );
  OR2x2_ASAP7_75t_SL U70539 ( .A(n60437), .B(n60436), .Y(or1200_cpu_rf_rdb) );
  INVx1_ASAP7_75t_SL U70540 ( .A(iwb_dat_i[31]), .Y(n77424) );
  OR2x2_ASAP7_75t_SL U70541 ( .A(n60442), .B(n77954), .Y(n77837) );
  INVx1_ASAP7_75t_SL U70542 ( .A(iwb_dat_i[29]), .Y(n77406) );
  NOR3xp33_ASAP7_75t_SL U70543 ( .A(n60454), .B(n77843), .C(or1200_cpu_rf_rdb), 
        .Y(n77394) );
  NOR3xp33_ASAP7_75t_SL U70544 ( .A(n77841), .B(n60456), .C(n60455), .Y(n60467) );
  A2O1A1Ixp33_ASAP7_75t_SL U70545 ( .A1(n77394), .A2(n60467), .B(n77834), .C(
        n60457), .Y(n60470) );
  NAND3xp33_ASAP7_75t_SL U70546 ( .A(n61037), .B(n77839), .C(n60459), .Y(
        n60461) );
  NAND4xp25_ASAP7_75t_SL U70547 ( .A(or1200_cpu_rf_rdb), .B(n77839), .C(n60459), .D(n61045), .Y(n60460) );
  A2O1A1Ixp33_ASAP7_75t_SL U70548 ( .A1(n61046), .A2(n60461), .B(n77363), .C(
        n60460), .Y(n60466) );
  A2O1A1Ixp33_ASAP7_75t_SL U70549 ( .A1(n60468), .A2(n60467), .B(n60466), .C(
        n60465), .Y(n60469) );
  OAI211xp5_ASAP7_75t_SL U70550 ( .A1(n60476), .A2(n77379), .B(n60475), .C(
        n60474), .Y(n9576) );
  INVx1_ASAP7_75t_SL U70551 ( .A(or1200_cpu_rf_addrb[4]), .Y(n60477) );
  INVx1_ASAP7_75t_SL U70552 ( .A(or1200_cpu_rf_addrb[0]), .Y(n60478) );
  INVx1_ASAP7_75t_SL U70553 ( .A(or1200_cpu_rf_addrb[3]), .Y(n60479) );
  OAI211xp5_ASAP7_75t_SL U70554 ( .A1(n60485), .A2(n77379), .B(n60484), .C(
        n60483), .Y(n9581) );
  INVx1_ASAP7_75t_SL U70555 ( .A(or1200_cpu_rf_addrb[1]), .Y(n60487) );
  INVx1_ASAP7_75t_SL U70556 ( .A(or1200_cpu_rf_addrb[2]), .Y(n60488) );
  NAND3xp33_ASAP7_75t_SL U70557 ( .A(n61155), .B(n62142), .C(n61028), .Y(
        n60499) );
  NOR3xp33_ASAP7_75t_SL U70558 ( .A(n60492), .B(n60491), .C(n60490), .Y(n60493) );
  INVx1_ASAP7_75t_SL U70559 ( .A(iwb_dat_i[16]), .Y(n60510) );
  A2O1A1Ixp33_ASAP7_75t_SL U70560 ( .A1(n77833), .A2(n60510), .B(n60506), .C(
        n77359), .Y(n60507) );
  NOR3xp33_ASAP7_75t_SL U70561 ( .A(n77954), .B(or1200_ic_top_from_icram[16]), 
        .C(n57090), .Y(n60509) );
  INVx1_ASAP7_75t_SL U70562 ( .A(iwb_dat_i[17]), .Y(n60513) );
  INVx1_ASAP7_75t_SL U70563 ( .A(iwb_dat_i[19]), .Y(n60520) );
  INVx1_ASAP7_75t_SL U70564 ( .A(iwb_dat_i[20]), .Y(n60528) );
  OAI222xp33_ASAP7_75t_SL U70565 ( .A1(n60529), .A2(n77954), .B1(n78009), .B2(
        n2715), .C1(n78006), .C2(n60528), .Y(n77936) );
  INVx1_ASAP7_75t_SL U70566 ( .A(iwb_dat_i[18]), .Y(n60533) );
  OAI222xp33_ASAP7_75t_SL U70567 ( .A1(n60534), .A2(n77954), .B1(n78009), .B2(
        n2719), .C1(n78006), .C2(n60533), .Y(n77946) );
  NAND4xp25_ASAP7_75t_SL U70568 ( .A(n59563), .B(n59579), .C(n59537), .D(
        n78439), .Y(n60537) );
  A2O1A1Ixp33_ASAP7_75t_SL U70569 ( .A1(n60541), .A2(n60540), .B(n60539), .C(
        n60538), .Y(n60542) );
  NAND3xp33_ASAP7_75t_SL U70570 ( .A(n61480), .B(n60556), .C(n60543), .Y(
        n61342) );
  OR2x2_ASAP7_75t_SL U70571 ( .A(n60834), .B(n60557), .Y(n64283) );
  AND2x2_ASAP7_75t_SL U70572 ( .A(n76720), .B(n60575), .Y(n76735) );
  OR2x2_ASAP7_75t_SL U70573 ( .A(n62205), .B(n60559), .Y(n63261) );
  OAI211xp5_ASAP7_75t_SL U70574 ( .A1(n62319), .A2(n60566), .B(n60565), .C(
        n60564), .Y(n60567) );
  NAND3xp33_ASAP7_75t_SL U70575 ( .A(n77166), .B(n60574), .C(n60573), .Y(
        n60817) );
  OR3x1_ASAP7_75t_SL U70576 ( .A(n61693), .B(n60581), .C(n60580), .Y(n77584)
         );
  OR2x2_ASAP7_75t_SL U70577 ( .A(n2567), .B(n60685), .Y(n64324) );
  OAI211xp5_ASAP7_75t_SL U70578 ( .A1(n62254), .A2(n62377), .B(n60594), .C(
        n60593), .Y(n62544) );
  NAND3xp33_ASAP7_75t_SL U70579 ( .A(n62612), .B(n59540), .C(n57128), .Y(
        n60597) );
  OR3x1_ASAP7_75t_SL U70580 ( .A(n60916), .B(n60606), .C(n77242), .Y(n60612)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70581 ( .A1(n64114), .A2(n59531), .B(n63668), .C(
        n59535), .Y(n60610) );
  NAND3xp33_ASAP7_75t_SL U70582 ( .A(n63179), .B(n59572), .C(n63176), .Y(
        n60608) );
  A2O1A1Ixp33_ASAP7_75t_SL U70583 ( .A1(n59486), .A2(n60610), .B(n63249), .C(
        n60609), .Y(n60611) );
  OR2x2_ASAP7_75t_SL U70584 ( .A(n60615), .B(n59445), .Y(n61648) );
  OR3x1_ASAP7_75t_SL U70585 ( .A(n61214), .B(n57215), .C(n76486), .Y(n60662)
         );
  AND2x2_ASAP7_75t_SL U70586 ( .A(n60668), .B(n60645), .Y(n60672) );
  OR2x2_ASAP7_75t_SL U70587 ( .A(n59545), .B(n59584), .Y(n60849) );
  AND2x2_ASAP7_75t_SL U70588 ( .A(n60627), .B(n76782), .Y(n75322) );
  A2O1A1Ixp33_ASAP7_75t_SL U70589 ( .A1(n62276), .A2(n60634), .B(n59565), .C(
        n60633), .Y(n60652) );
  OR2x2_ASAP7_75t_SL U70590 ( .A(n59558), .B(n59567), .Y(n75866) );
  OR2x2_ASAP7_75t_SL U70591 ( .A(n59568), .B(n57197), .Y(n61436) );
  OR2x2_ASAP7_75t_SL U70592 ( .A(n59557), .B(n63571), .Y(n60850) );
  OAI211xp5_ASAP7_75t_SL U70593 ( .A1(n61531), .A2(n60650), .B(n60649), .C(
        n60648), .Y(n60651) );
  A2O1A1Ixp33_ASAP7_75t_SL U70594 ( .A1(n61519), .A2(n60654), .B(n61526), .C(
        n60653), .Y(n60696) );
  NAND3xp33_ASAP7_75t_SL U70595 ( .A(n66257), .B(n61521), .C(n75740), .Y(
        n61409) );
  OR2x2_ASAP7_75t_SL U70596 ( .A(n59542), .B(n59584), .Y(n60863) );
  NAND3xp33_ASAP7_75t_SL U70597 ( .A(n76782), .B(n59567), .C(n57214), .Y(
        n75328) );
  A2O1A1Ixp33_ASAP7_75t_SL U70598 ( .A1(n60922), .A2(n60675), .B(n61428), .C(
        n60674), .Y(n60676) );
  OR2x2_ASAP7_75t_SL U70599 ( .A(n59486), .B(n59645), .Y(n62534) );
  NAND3xp33_ASAP7_75t_SL U70600 ( .A(n60678), .B(n60677), .C(n62534), .Y(
        n62344) );
  OAI211xp5_ASAP7_75t_SL U70601 ( .A1(n62422), .A2(n62341), .B(n60693), .C(
        n60692), .Y(n60694) );
  O2A1O1Ixp5_ASAP7_75t_SL U70602 ( .A1(n60696), .A2(n60695), .B(n57126), .C(
        n60694), .Y(n60697) );
  OAI211xp5_ASAP7_75t_SL U70603 ( .A1(n64796), .A2(n61241), .B(n60698), .C(
        n60697), .Y(n60699) );
  XOR2xp5_ASAP7_75t_SL U70604 ( .A(n2076), .B(n2664), .Y(n60708) );
  XOR2xp5_ASAP7_75t_SL U70605 ( .A(n2042), .B(n2678), .Y(n60707) );
  XOR2xp5_ASAP7_75t_SL U70606 ( .A(n2059), .B(n2671), .Y(n60709) );
  A2O1A1Ixp33_ASAP7_75t_SL U70607 ( .A1(or1200_cpu_rf_dataa_0_), .A2(n61056), 
        .B(n60714), .C(n60728), .Y(n60715) );
  AO21x1_ASAP7_75t_SL U70608 ( .A1(n60717), .A2(n3390), .B(n69341), .Y(n77462)
         );
  NAND3xp33_ASAP7_75t_SL U70609 ( .A(n57500), .B(n59580), .C(n59553), .Y(
        n60732) );
  OR2x2_ASAP7_75t_SL U70610 ( .A(n60732), .B(n60737), .Y(n61913) );
  O2A1O1Ixp5_ASAP7_75t_SL U70611 ( .A1(n59539), .A2(n60778), .B(n60734), .C(
        n67311), .Y(n60735) );
  OR2x2_ASAP7_75t_SL U70612 ( .A(n53455), .B(n62671), .Y(n60777) );
  A2O1A1Ixp33_ASAP7_75t_SL U70613 ( .A1(n61673), .A2(n61676), .B(n60776), .C(
        n60746), .Y(n62462) );
  O2A1O1Ixp5_ASAP7_75t_SL U70614 ( .A1(n59708), .A2(n57120), .B(n60750), .C(
        n64776), .Y(n60758) );
  XNOR2xp5_ASAP7_75t_SL U70615 ( .A(n53316), .B(n60758), .Y(n61237) );
  O2A1O1Ixp5_ASAP7_75t_SL U70616 ( .A1(n60765), .A2(n61397), .B(n60764), .C(
        n60763), .Y(n60767) );
  XNOR2xp5_ASAP7_75t_SL U70617 ( .A(n78002), .B(n60769), .Y(n76280) );
  XNOR2xp5_ASAP7_75t_SL U70618 ( .A(n59569), .B(n60772), .Y(n62307) );
  A2O1A1Ixp33_ASAP7_75t_SL U70619 ( .A1(n62308), .A2(n62296), .B(n62309), .C(
        n60773), .Y(n62313) );
  XNOR2xp5_ASAP7_75t_SL U70620 ( .A(n59542), .B(n60775), .Y(n61323) );
  OR2x2_ASAP7_75t_SL U70621 ( .A(n59387), .B(n60778), .Y(n60782) );
  XNOR2xp5_ASAP7_75t_SL U70622 ( .A(n59553), .B(n60779), .Y(n60780) );
  OR2x2_ASAP7_75t_SL U70623 ( .A(n60787), .B(n60786), .Y(n64834) );
  AND2x2_ASAP7_75t_SL U70624 ( .A(n60789), .B(n62535), .Y(n62256) );
  NAND3xp33_ASAP7_75t_SL U70625 ( .A(n60799), .B(n76486), .C(n60791), .Y(
        n61854) );
  OAI211xp5_ASAP7_75t_SL U70626 ( .A1(n62256), .A2(n76779), .B(n60795), .C(
        n60794), .Y(n60802) );
  OAI31xp33_ASAP7_75t_SL U70627 ( .A1(n62454), .A2(n61829), .A3(n61833), .B(
        n60814), .Y(n60815) );
  A2O1A1Ixp33_ASAP7_75t_SL U70628 ( .A1(n61829), .A2(n62454), .B(n60815), .C(
        n61735), .Y(n60886) );
  OR2x2_ASAP7_75t_SL U70629 ( .A(n60817), .B(n60816), .Y(n76731) );
  OAI211xp5_ASAP7_75t_SL U70630 ( .A1(n1372), .A2(n75364), .B(n60823), .C(
        n60822), .Y(n60829) );
  OR2x2_ASAP7_75t_SL U70631 ( .A(n60840), .B(n60839), .Y(n75747) );
  XOR2xp5_ASAP7_75t_SL U70632 ( .A(n77021), .B(n77080), .Y(n60853) );
  OR2x2_ASAP7_75t_SL U70633 ( .A(n75872), .B(n60846), .Y(n74607) );
  NAND3xp33_ASAP7_75t_SL U70634 ( .A(n60850), .B(n60849), .C(n60848), .Y(
        n62257) );
  NAND3xp33_ASAP7_75t_SL U70635 ( .A(n61697), .B(n61699), .C(n60855), .Y(
        n60856) );
  OR2x2_ASAP7_75t_SL U70636 ( .A(n59529), .B(n63571), .Y(n75836) );
  OR2x2_ASAP7_75t_SL U70637 ( .A(n59541), .B(n59645), .Y(n61191) );
  OR2x2_ASAP7_75t_SL U70638 ( .A(n75702), .B(n75863), .Y(n75838) );
  OR2x2_ASAP7_75t_SL U70639 ( .A(n75872), .B(n75838), .Y(n77093) );
  OAI211xp5_ASAP7_75t_SL U70640 ( .A1(n62253), .A2(n62422), .B(n60869), .C(
        n60868), .Y(n60870) );
  AO21x1_ASAP7_75t_SL U70641 ( .A1(n77125), .A2(n75747), .B(n60870), .Y(n60884) );
  NAND3xp33_ASAP7_75t_SL U70642 ( .A(n61856), .B(n60872), .C(n60871), .Y(
        n77065) );
  A2O1A1Ixp33_ASAP7_75t_SL U70643 ( .A1(n60887), .A2(n60886), .B(n75872), .C(
        n60885), .Y(n60888) );
  A2O1A1Ixp33_ASAP7_75t_SL U70644 ( .A1(n62762), .A2(n57144), .B(n77243), .C(
        n77024), .Y(n60889) );
  OAI211xp5_ASAP7_75t_SL U70645 ( .A1(n60896), .A2(n77379), .B(n60895), .C(
        n60894), .Y(n9601) );
  OR2x2_ASAP7_75t_SL U70646 ( .A(n64209), .B(n61746), .Y(n61597) );
  OAI211xp5_ASAP7_75t_SL U70647 ( .A1(or1200_cpu_or1200_except_n282), .A2(
        n76731), .B(n60906), .C(n60905), .Y(n60908) );
  NAND4xp25_ASAP7_75t_SL U70648 ( .A(n61538), .B(n57200), .C(n61212), .D(
        n60913), .Y(n60973) );
  A2O1A1Ixp33_ASAP7_75t_SL U70649 ( .A1(n59577), .A2(n60922), .B(n61428), .C(
        n60921), .Y(n60923) );
  A2O1A1Ixp33_ASAP7_75t_SL U70650 ( .A1(n60926), .A2(n61406), .B(n61526), .C(
        n60925), .Y(n60927) );
  OR2x2_ASAP7_75t_SL U70651 ( .A(n57197), .B(n75710), .Y(n75714) );
  AND2x2_ASAP7_75t_SL U70652 ( .A(n59709), .B(n73923), .Y(n75861) );
  AO21x1_ASAP7_75t_SL U70653 ( .A1(n59710), .A2(n59563), .B(n59442), .Y(n64231) );
  A2O1A1Ixp33_ASAP7_75t_SL U70654 ( .A1(n75708), .A2(n59182), .B(n60939), .C(
        n60938), .Y(n60940) );
  OAI211xp5_ASAP7_75t_SL U70655 ( .A1(n62275), .A2(n75348), .B(n60941), .C(
        n60940), .Y(n60950) );
  OR2x2_ASAP7_75t_SL U70656 ( .A(n59568), .B(n59584), .Y(n61491) );
  NAND3xp33_ASAP7_75t_SL U70657 ( .A(n61215), .B(n60946), .C(n74005), .Y(
        n60947) );
  OAI211xp5_ASAP7_75t_SL U70658 ( .A1(n76779), .A2(n61491), .B(n60948), .C(
        n60947), .Y(n60949) );
  A2O1A1Ixp33_ASAP7_75t_SL U70659 ( .A1(n58587), .A2(n60953), .B(n61526), .C(
        n60952), .Y(n60976) );
  OR3x1_ASAP7_75t_SL U70660 ( .A(n61783), .B(n59709), .C(n75326), .Y(n60960)
         );
  OR2x2_ASAP7_75t_SL U70661 ( .A(n59541), .B(n59584), .Y(n61731) );
  NAND3xp33_ASAP7_75t_SL U70662 ( .A(n60958), .B(n61731), .C(n60957), .Y(
        n61643) );
  OAI211xp5_ASAP7_75t_SL U70663 ( .A1(n61638), .A2(n60961), .B(n60960), .C(
        n60959), .Y(n60971) );
  NAND3xp33_ASAP7_75t_SL U70664 ( .A(n61429), .B(n60963), .C(n60962), .Y(
        n60964) );
  NOR3xp33_ASAP7_75t_SL U70665 ( .A(n60971), .B(n60970), .C(n60969), .Y(n60972) );
  A2O1A1Ixp33_ASAP7_75t_SL U70666 ( .A1(n59545), .A2(n60974), .B(n60973), .C(
        n60972), .Y(n60975) );
  OAI211xp5_ASAP7_75t_SL U70667 ( .A1(n77586), .A2(n76796), .B(n60984), .C(
        n60983), .Y(n60985) );
  A2O1A1Ixp33_ASAP7_75t_SL U70668 ( .A1(n61182), .A2(n60989), .B(n75872), .C(
        n60988), .Y(n60990) );
  A2O1A1Ixp33_ASAP7_75t_SL U70669 ( .A1(n77588), .A2(n60992), .B(n76744), .C(
        n60991), .Y(n77921) );
  OAI211xp5_ASAP7_75t_SL U70670 ( .A1(n61017), .A2(n77137), .B(n61016), .C(
        n61015), .Y(n9638) );
  OAI211xp5_ASAP7_75t_SL U70671 ( .A1(n61021), .A2(n77137), .B(n61020), .C(
        n61019), .Y(n9639) );
  OAI211xp5_ASAP7_75t_SL U70672 ( .A1(n61027), .A2(n77379), .B(n61026), .C(
        n61025), .Y(n9599) );
  OR2x2_ASAP7_75t_SL U70673 ( .A(n3078), .B(n61142), .Y(n61147) );
  NOR3xp33_ASAP7_75t_SL U70674 ( .A(n61048), .B(n77397), .C(n61047), .Y(n61049) );
  A2O1A1Ixp33_ASAP7_75t_SL U70675 ( .A1(n61052), .A2(n61051), .B(n61050), .C(
        n61049), .Y(n61053) );
  AO21x1_ASAP7_75t_SL U70676 ( .A1(n62008), .A2(n76720), .B(n61061), .Y(n61084) );
  NAND3xp33_ASAP7_75t_SL U70677 ( .A(n61067), .B(n61677), .C(n61062), .Y(
        n77632) );
  OR3x1_ASAP7_75t_SL U70678 ( .A(n77636), .B(n77635), .C(n61063), .Y(n61119)
         );
  AND2x2_ASAP7_75t_SL U70679 ( .A(n76739), .B(n61342), .Y(n61618) );
  O2A1O1Ixp5_ASAP7_75t_SL U70680 ( .A1(n61069), .A2(n61068), .B(n61067), .C(
        n61066), .Y(n61070) );
  OAI211xp5_ASAP7_75t_SL U70681 ( .A1(or1200_cpu_or1200_except_n258), .A2(
        n76731), .B(n61071), .C(n61070), .Y(n61072) );
  A2O1A1Ixp33_ASAP7_75t_SL U70682 ( .A1(n61086), .A2(n77288), .B(n77227), .C(
        n61085), .Y(n61092) );
  AND2x2_ASAP7_75t_SL U70683 ( .A(n64840), .B(n75731), .Y(n75577) );
  A2O1A1Ixp33_ASAP7_75t_SL U70684 ( .A1(n77097), .A2(n77701), .B(n77096), .C(
        n57641), .Y(n61090) );
  NAND4xp25_ASAP7_75t_SL U70685 ( .A(n61093), .B(n61092), .C(n61091), .D(
        n61090), .Y(n61114) );
  OAI211xp5_ASAP7_75t_SL U70686 ( .A1(n75327), .A2(n77078), .B(n61111), .C(
        n61110), .Y(n61113) );
  OAI211xp5_ASAP7_75t_SL U70687 ( .A1(n75882), .A2(n61117), .B(n62459), .C(
        n61116), .Y(n61118) );
  AO21x1_ASAP7_75t_SL U70688 ( .A1(n57073), .A2(n77900), .B(n61123), .Y(n1777)
         );
  NAND3xp33_ASAP7_75t_SL U70689 ( .A(n61153), .B(n61135), .C(n62022), .Y(
        n61151) );
  NAND4xp25_ASAP7_75t_SL U70690 ( .A(n76809), .B(n74796), .C(n69335), .D(n2122), .Y(n61138) );
  NAND3xp33_ASAP7_75t_SL U70691 ( .A(n61136), .B(n2110), .C(n2499), .Y(n61137)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70692 ( .A1(n3078), .A2(n62024), .B(n77427), .C(
        n61140), .Y(n61141) );
  NAND3xp33_ASAP7_75t_SL U70693 ( .A(n61143), .B(n61142), .C(n61141), .Y(
        n61144) );
  A2O1A1Ixp33_ASAP7_75t_SL U70694 ( .A1(n61147), .A2(n62070), .B(n57093), .C(
        n61146), .Y(n61148) );
  OAI31xp33_ASAP7_75t_SL U70695 ( .A1(n69334), .A2(n3426), .A3(n75475), .B(
        n59702), .Y(n61163) );
  OR2x2_ASAP7_75t_SL U70696 ( .A(n62477), .B(n59556), .Y(n4061) );
  OR2x2_ASAP7_75t_SL U70697 ( .A(n61167), .B(n63741), .Y(n61577) );
  NAND3xp33_ASAP7_75t_SL U70698 ( .A(n74956), .B(
        or1200_cpu_or1200_genpc_pcreg_default[5]), .C(n61169), .Y(n61170) );
  OR2x2_ASAP7_75t_SL U70699 ( .A(n59584), .B(n59571), .Y(n62357) );
  AND2x2_ASAP7_75t_SL U70700 ( .A(n61187), .B(n62357), .Y(n62255) );
  OR2x2_ASAP7_75t_SL U70701 ( .A(n59567), .B(n62355), .Y(n75325) );
  OAI211xp5_ASAP7_75t_SL U70702 ( .A1(n61193), .A2(n62533), .B(n61192), .C(
        n61191), .Y(n62262) );
  A2O1A1Ixp33_ASAP7_75t_SL U70703 ( .A1(n61196), .A2(n61195), .B(n61498), .C(
        n61194), .Y(n61205) );
  NAND3xp33_ASAP7_75t_SL U70704 ( .A(n61521), .B(n57424), .C(n62761), .Y(
        n61426) );
  OR2x2_ASAP7_75t_SL U70705 ( .A(n75710), .B(n75863), .Y(n75835) );
  NOR3xp33_ASAP7_75t_SL U70706 ( .A(n61205), .B(n61204), .C(n61203), .Y(n61223) );
  A2O1A1Ixp33_ASAP7_75t_SL U70707 ( .A1(n59560), .A2(n61212), .B(n61211), .C(
        n61210), .Y(n61213) );
  OR2x2_ASAP7_75t_SL U70708 ( .A(n59709), .B(n75866), .Y(n75700) );
  NOR3xp33_ASAP7_75t_SL U70709 ( .A(n61531), .B(n59708), .C(n75729), .Y(n61216) );
  NAND3xp33_ASAP7_75t_SL U70710 ( .A(n61220), .B(n61219), .C(n61218), .Y(
        n61221) );
  OAI211xp5_ASAP7_75t_SL U70711 ( .A1(n61225), .A2(n61224), .B(n61223), .C(
        n61222), .Y(n61234) );
  OAI211xp5_ASAP7_75t_SL U70712 ( .A1(n62284), .A2(n63565), .B(n61232), .C(
        n61231), .Y(n61233) );
  OAI211xp5_ASAP7_75t_SL U70713 ( .A1(n64853), .A2(n61241), .B(n61240), .C(
        n61239), .Y(n61263) );
  OR2x2_ASAP7_75t_SL U70714 ( .A(n64209), .B(n61248), .Y(n63555) );
  OAI211xp5_ASAP7_75t_SL U70715 ( .A1(or1200_cpu_or1200_except_n492), .A2(
        n76724), .B(n61252), .C(n61251), .Y(n61253) );
  OAI211xp5_ASAP7_75t_SL U70716 ( .A1(n61267), .A2(n77137), .B(n61266), .C(
        n61265), .Y(n9637) );
  OR2x2_ASAP7_75t_SL U70717 ( .A(n62477), .B(n59543), .Y(n4049) );
  NAND3xp33_ASAP7_75t_SL U70718 ( .A(n61274), .B(n61273), .C(n61272), .Y(
        n76520) );
  OR2x2_ASAP7_75t_SL U70719 ( .A(n61280), .B(n57083), .Y(n77416) );
  AND2x2_ASAP7_75t_SL U70720 ( .A(n78165), .B(n77996), .Y(n77488) );
  AND2x2_ASAP7_75t_SL U70721 ( .A(n77765), .B(n61292), .Y(n61304) );
  OR2x2_ASAP7_75t_SL U70722 ( .A(n78163), .B(n77473), .Y(n77483) );
  O2A1O1Ixp5_ASAP7_75t_SL U70723 ( .A1(n61295), .A2(n77413), .B(n3088), .C(
        n61294), .Y(n77469) );
  O2A1O1Ixp5_ASAP7_75t_SL U70724 ( .A1(n61312), .A2(n61311), .B(n61310), .C(
        n3392), .Y(n61313) );
  AO21x1_ASAP7_75t_SL U70725 ( .A1(n61327), .A2(n76720), .B(n61326), .Y(n77610) );
  OAI211xp5_ASAP7_75t_SL U70726 ( .A1(or1200_cpu_or1200_except_n506), .A2(
        n76724), .B(n61330), .C(n61329), .Y(n61331) );
  OR3x1_ASAP7_75t_SL U70727 ( .A(n61341), .B(n61340), .C(n61339), .Y(n61345)
         );
  OAI211xp5_ASAP7_75t_SL U70728 ( .A1(n75348), .A2(n62447), .B(n61350), .C(
        n61349), .Y(n61351) );
  A2O1A1Ixp33_ASAP7_75t_SL U70729 ( .A1(n61362), .A2(n61361), .B(n75872), .C(
        n61360), .Y(n61372) );
  OR3x1_ASAP7_75t_SL U70730 ( .A(n61372), .B(n61371), .C(n61370), .Y(n61373)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70731 ( .A1(n61387), .A2(n76729), .B(n77595), .C(
        n61386), .Y(n61389) );
  OAI211xp5_ASAP7_75t_SL U70732 ( .A1(or1200_cpu_or1200_except_n589), .A2(
        n59675), .B(n61392), .C(n61391), .Y(n61395) );
  OR3x1_ASAP7_75t_SL U70733 ( .A(n61395), .B(n61394), .C(n61393), .Y(n77596)
         );
  OR2x2_ASAP7_75t_SL U70734 ( .A(n61404), .B(n61403), .Y(n75877) );
  AO21x1_ASAP7_75t_SL U70735 ( .A1(n75890), .A2(n57506), .B(n61405), .Y(n61523) );
  OAI211xp5_ASAP7_75t_SL U70736 ( .A1(n64131), .A2(n61424), .B(n61423), .C(
        n61422), .Y(n61431) );
  OAI211xp5_ASAP7_75t_SL U70737 ( .A1(n61429), .A2(n61428), .B(n61427), .C(
        n61426), .Y(n61430) );
  NOR3xp33_ASAP7_75t_SL U70738 ( .A(n61432), .B(n61431), .C(n61430), .Y(n61442) );
  NAND3xp33_ASAP7_75t_SL U70739 ( .A(n61437), .B(n61436), .C(n61435), .Y(
        n62518) );
  OR2x2_ASAP7_75t_SL U70740 ( .A(n61447), .B(n61446), .Y(n61624) );
  XOR2xp5_ASAP7_75t_SL U70741 ( .A(or1200_cpu_or1200_except_n494), .B(
        or1200_cpu_or1200_except_n496), .Y(n61452) );
  OAI211xp5_ASAP7_75t_SL U70742 ( .A1(n62284), .A2(n64121), .B(n61454), .C(
        n61453), .Y(n61455) );
  OAI211xp5_ASAP7_75t_SL U70743 ( .A1(n76295), .A2(n73953), .B(n61460), .C(
        n61459), .Y(n61461) );
  AO21x1_ASAP7_75t_SL U70744 ( .A1(n61469), .A2(n76720), .B(n61468), .Y(n61556) );
  NAND3xp33_ASAP7_75t_SL U70745 ( .A(n61595), .B(n77623), .C(n61470), .Y(
        n61471) );
  OAI211xp5_ASAP7_75t_SL U70746 ( .A1(or1200_cpu_or1200_except_n494), .A2(
        n76724), .B(n61476), .C(n61475), .Y(n61477) );
  NAND3xp33_ASAP7_75t_SL U70747 ( .A(n61485), .B(n61484), .C(n61483), .Y(
        n77593) );
  NAND3xp33_ASAP7_75t_SL U70748 ( .A(n61491), .B(n61490), .C(n61489), .Y(
        n77062) );
  OR2x2_ASAP7_75t_SL U70749 ( .A(n59442), .B(n59577), .Y(n64780) );
  OAI31xp33_ASAP7_75t_SL U70750 ( .A1(n76759), .A2(n76765), .A3(n61498), .B(
        n61497), .Y(n61499) );
  OAI211xp5_ASAP7_75t_SL U70751 ( .A1(n61503), .A2(n73941), .B(n61502), .C(
        n61501), .Y(n61516) );
  OR2x2_ASAP7_75t_SL U70752 ( .A(n59545), .B(n57197), .Y(n61726) );
  OAI31xp33_ASAP7_75t_SL U70753 ( .A1(n61506), .A2(n61505), .A3(n61504), .B(
        n75845), .Y(n61513) );
  OR2x2_ASAP7_75t_SL U70754 ( .A(n59542), .B(n57197), .Y(n61732) );
  OAI211xp5_ASAP7_75t_SL U70755 ( .A1(n63176), .A2(n61514), .B(n61513), .C(
        n61512), .Y(n61515) );
  NOR3xp33_ASAP7_75t_SL U70756 ( .A(n61526), .B(n61525), .C(n62615), .Y(n61528) );
  NOR3xp33_ASAP7_75t_SL U70757 ( .A(n61529), .B(n61528), .C(n61527), .Y(n61535) );
  NOR3xp33_ASAP7_75t_SL U70758 ( .A(n61531), .B(n59708), .C(n77106), .Y(n61532) );
  NAND4xp25_ASAP7_75t_SL U70759 ( .A(n61543), .B(n61542), .C(n61541), .D(
        n61540), .Y(n61552) );
  OR2x2_ASAP7_75t_SL U70760 ( .A(n61551), .B(n61550), .Y(n73933) );
  OAI211xp5_ASAP7_75t_SL U70761 ( .A1(n61628), .A2(n74619), .B(n61555), .C(
        n61554), .Y(n61558) );
  NAND3xp33_ASAP7_75t_SL U70762 ( .A(n61563), .B(n61562), .C(n61561), .Y(
        n61564) );
  OR2x2_ASAP7_75t_SL U70763 ( .A(n62477), .B(n59567), .Y(n4070) );
  A2O1A1Ixp33_ASAP7_75t_SL U70764 ( .A1(
        or1200_cpu_or1200_genpc_pcreg_default[4]), .A2(n59701), .B(n61569), 
        .C(n77251), .Y(n61570) );
  AND2x2_ASAP7_75t_SL U70765 ( .A(n61586), .B(n57100), .Y(n76580) );
  OAI211xp5_ASAP7_75t_SL U70766 ( .A1(n61594), .A2(n77379), .B(n61593), .C(
        n61592), .Y(n9600) );
  OR3x1_ASAP7_75t_SL U70767 ( .A(n61602), .B(n61601), .C(n61600), .Y(n61609)
         );
  NAND4xp25_ASAP7_75t_SL U70768 ( .A(n61613), .B(n61612), .C(n61611), .D(
        n61610), .Y(n61614) );
  OAI211xp5_ASAP7_75t_SL U70769 ( .A1(n77943), .A2(n61618), .B(n61617), .C(
        n61616), .Y(n77599) );
  OR2x2_ASAP7_75t_SL U70770 ( .A(n59708), .B(n75872), .Y(n61784) );
  NAND4xp25_ASAP7_75t_SL U70771 ( .A(n61655), .B(n61654), .C(n61653), .D(
        n61652), .Y(n61656) );
  OAI211xp5_ASAP7_75t_SL U70772 ( .A1(n77598), .A2(n76796), .B(n61660), .C(
        n61659), .Y(n61661) );
  OAI211xp5_ASAP7_75t_SL U70773 ( .A1(n73953), .A2(n76293), .B(n61665), .C(
        n61664), .Y(n61666) );
  OAI211xp5_ASAP7_75t_SL U70774 ( .A1(n77913), .A2(n77137), .B(n61670), .C(
        n61669), .Y(n9634) );
  A2O1A1Ixp33_ASAP7_75t_SL U70775 ( .A1(n61686), .A2(n76729), .B(n77616), .C(
        n61685), .Y(n61687) );
  OAI211xp5_ASAP7_75t_SL U70776 ( .A1(or1200_cpu_or1200_except_n262), .A2(
        n76731), .B(n61690), .C(n61689), .Y(n61691) );
  A2O1A1Ixp33_ASAP7_75t_SL U70777 ( .A1(n61701), .A2(n64835), .B(n61700), .C(
        n57219), .Y(n61702) );
  OAI211xp5_ASAP7_75t_SL U70778 ( .A1(n61772), .A2(n76553), .B(n62444), .C(
        n77082), .Y(n61711) );
  OAI211xp5_ASAP7_75t_SL U70779 ( .A1(n75588), .A2(n77107), .B(n61711), .C(
        n61710), .Y(n61712) );
  NAND3xp33_ASAP7_75t_SL U70780 ( .A(n61715), .B(n61714), .C(n61713), .Y(
        n61716) );
  A2O1A1Ixp33_ASAP7_75t_SL U70781 ( .A1(n61722), .A2(n61721), .B(n62455), .C(
        n61720), .Y(n61736) );
  NAND3xp33_ASAP7_75t_SL U70782 ( .A(n61727), .B(n61726), .C(n61725), .Y(
        n77056) );
  NAND3xp33_ASAP7_75t_SL U70783 ( .A(n61732), .B(n61731), .C(n61730), .Y(
        n77089) );
  A2O1A1Ixp33_ASAP7_75t_SL U70784 ( .A1(n61736), .A2(n61735), .B(n61734), .C(
        n57126), .Y(n61737) );
  NAND3xp33_ASAP7_75t_SL U70785 ( .A(n62459), .B(n61738), .C(n61737), .Y(
        n61739) );
  A2O1A1Ixp33_ASAP7_75t_SL U70786 ( .A1(n77467), .A2(n61743), .B(n76556), .C(
        n61742), .Y(n9659) );
  AO21x1_ASAP7_75t_SL U70787 ( .A1(n75764), .A2(n76720), .B(n61747), .Y(n77613) );
  OAI211xp5_ASAP7_75t_SL U70788 ( .A1(or1200_cpu_or1200_except_n422), .A2(
        n59676), .B(n61758), .C(n61757), .Y(n61761) );
  OR3x1_ASAP7_75t_SL U70789 ( .A(n61761), .B(n61760), .C(n61759), .Y(n61762)
         );
  OR2x2_ASAP7_75t_SL U70790 ( .A(n75872), .B(n76779), .Y(n77099) );
  OAI211xp5_ASAP7_75t_SL U70791 ( .A1(n62256), .A2(n62332), .B(n61766), .C(
        n61765), .Y(n61767) );
  OAI211xp5_ASAP7_75t_SL U70792 ( .A1(or1200_cpu_or1200_mult_mac_n307), .A2(
        n75738), .B(n61779), .C(n61778), .Y(n61780) );
  A2O1A1Ixp33_ASAP7_75t_SL U70793 ( .A1(n77097), .A2(n62738), .B(n77096), .C(
        n58206), .Y(n61787) );
  NAND4xp25_ASAP7_75t_SL U70794 ( .A(n61789), .B(n61788), .C(n61787), .D(
        n61786), .Y(n61790) );
  OAI211xp5_ASAP7_75t_SL U70795 ( .A1(n75882), .A2(n61794), .B(n61793), .C(
        n61792), .Y(n61795) );
  XNOR2xp5_ASAP7_75t_SL U70796 ( .A(n61800), .B(n61799), .Y(n76302) );
  NAND4xp25_ASAP7_75t_SL U70797 ( .A(n61824), .B(n61823), .C(n74597), .D(
        n64319), .Y(n61825) );
  NAND4xp25_ASAP7_75t_SL U70798 ( .A(n61831), .B(n62456), .C(n61830), .D(
        n61829), .Y(n61834) );
  OR3x1_ASAP7_75t_SL U70799 ( .A(n61834), .B(n61833), .C(n61832), .Y(n61835)
         );
  OR2x2_ASAP7_75t_SL U70800 ( .A(n75567), .B(n75568), .Y(n75605) );
  OR2x2_ASAP7_75t_SL U70801 ( .A(or1200_cpu_or1200_except_n542), .B(n73905), 
        .Y(n75884) );
  NAND3xp33_ASAP7_75t_SL U70802 ( .A(n61840), .B(or1200_cpu_or1200_except_n550), .C(n75686), .Y(n61899) );
  AND2x2_ASAP7_75t_SL U70803 ( .A(n59493), .B(n64208), .Y(n75689) );
  OAI211xp5_ASAP7_75t_SL U70804 ( .A1(n75819), .A2(n68814), .B(n61847), .C(
        n61846), .Y(n61848) );
  NAND3xp33_ASAP7_75t_SL U70805 ( .A(n64208), .B(n1426), .C(n64209), .Y(n77674) );
  NAND3xp33_ASAP7_75t_SL U70806 ( .A(n61856), .B(n61855), .C(n57210), .Y(
        n61857) );
  NAND3xp33_ASAP7_75t_SL U70807 ( .A(n76782), .B(n64229), .C(n61861), .Y(
        n61862) );
  OAI211xp5_ASAP7_75t_SL U70808 ( .A1(n59551), .A2(n75722), .B(n61863), .C(
        n61862), .Y(n61864) );
  OAI211xp5_ASAP7_75t_SL U70809 ( .A1(or1200_cpu_or1200_mult_mac_n349), .A2(
        n75738), .B(n61867), .C(n61866), .Y(n61894) );
  NOR3xp33_ASAP7_75t_SL U70810 ( .A(n61890), .B(n61889), .C(n61888), .Y(n61891) );
  NOR3xp33_ASAP7_75t_SL U70811 ( .A(n61894), .B(n61893), .C(n61892), .Y(n61896) );
  NAND3xp33_ASAP7_75t_SL U70812 ( .A(n62134), .B(n61896), .C(n61895), .Y(
        n61897) );
  A2O1A1Ixp33_ASAP7_75t_SL U70813 ( .A1(n61900), .A2(n61899), .B(n76791), .C(
        n61898), .Y(n61901) );
  XNOR2xp5_ASAP7_75t_SL U70814 ( .A(n59582), .B(n61903), .Y(n75476) );
  XNOR2xp5_ASAP7_75t_SL U70815 ( .A(n59576), .B(n61907), .Y(n75679) );
  XNOR2xp5_ASAP7_75t_SL U70816 ( .A(n57215), .B(n61985), .Y(n75260) );
  XNOR2xp5_ASAP7_75t_SL U70817 ( .A(n77709), .B(n61919), .Y(n61939) );
  NAND3xp33_ASAP7_75t_SL U70818 ( .A(n58707), .B(n59536), .C(n59534), .Y(
        n61922) );
  NAND3xp33_ASAP7_75t_SL U70819 ( .A(n61923), .B(n58707), .C(n59536), .Y(
        n61924) );
  O2A1O1Ixp5_ASAP7_75t_SL U70820 ( .A1(n77713), .A2(n61927), .B(n61926), .C(
        n63668), .Y(n63543) );
  OR2x2_ASAP7_75t_SL U70821 ( .A(n59533), .B(n59534), .Y(n63584) );
  XNOR2xp5_ASAP7_75t_SL U70822 ( .A(n59536), .B(n61933), .Y(n61940) );
  XNOR2xp5_ASAP7_75t_SL U70823 ( .A(n59537), .B(n61939), .Y(n62500) );
  XNOR2xp5_ASAP7_75t_SL U70824 ( .A(n59532), .B(n61945), .Y(n61946) );
  O2A1O1Ixp5_ASAP7_75t_SL U70825 ( .A1(n61956), .A2(n62080), .B(n61948), .C(
        n61957), .Y(n61949) );
  NAND3xp33_ASAP7_75t_SL U70826 ( .A(n62077), .B(n62076), .C(n61961), .Y(
        n64186) );
  XNOR2xp5_ASAP7_75t_SL U70827 ( .A(n59561), .B(n61962), .Y(n64271) );
  A2O1A1Ixp33_ASAP7_75t_SL U70828 ( .A1(n64506), .A2(n77730), .B(n53455), .C(
        n61967), .Y(n61968) );
  NAND3xp33_ASAP7_75t_SL U70829 ( .A(n64191), .B(n64189), .C(n64757), .Y(
        n61970) );
  O2A1O1Ixp5_ASAP7_75t_SL U70830 ( .A1(n61975), .A2(n64186), .B(n64193), .C(
        n61974), .Y(n64813) );
  XNOR2xp5_ASAP7_75t_SL U70831 ( .A(n75832), .B(n61982), .Y(n73950) );
  A2O1A1Ixp33_ASAP7_75t_SL U70832 ( .A1(n64813), .A2(n64812), .B(n75809), .C(
        n61984), .Y(n75261) );
  OR2x2_ASAP7_75t_SL U70833 ( .A(n62477), .B(n57500), .Y(n4045) );
  AND2x2_ASAP7_75t_SL U70834 ( .A(n3111), .B(n61998), .Y(n77476) );
  A2O1A1Ixp33_ASAP7_75t_SL U70835 ( .A1(n62024), .A2(n62023), .B(n62022), .C(
        n62021), .Y(n62031) );
  NAND3xp33_ASAP7_75t_SL U70836 ( .A(n62025), .B(
        or1200_cpu_or1200_mult_mac_n285), .C(or1200_cpu_or1200_mult_mac_n139), 
        .Y(n62026) );
  OR2x2_ASAP7_75t_SL U70837 ( .A(or1200_cpu_or1200_fpu_fpu_op_r_2_), .B(
        or1200_cpu_or1200_fpu_fpu_op_r_3_), .Y(n74754) );
  OR2x2_ASAP7_75t_SL U70838 ( .A(n2579), .B(n74754), .Y(n2457) );
  NAND3xp33_ASAP7_75t_SL U70839 ( .A(n78437), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_1_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_s_count_2_), .Y(n62044) );
  O2A1O1Ixp5_ASAP7_75t_SL U70840 ( .A1(n62045), .A2(n62044), .B(n62043), .C(
        n62042), .Y(n62065) );
  OR2x2_ASAP7_75t_SL U70841 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_state), .B(
        or1200_cpu_or1200_fpu_fpu_arith_s_start_i), .Y(n62067) );
  A2O1A1Ixp33_ASAP7_75t_SL U70842 ( .A1(n62059), .A2(n62058), .B(n58624), .C(
        n62057), .Y(n2203) );
  AO21x1_ASAP7_75t_SL U70843 ( .A1(n78245), .A2(n62065), .B(n62064), .Y(n2208)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70844 ( .A1(n62068), .A2(n78245), .B(
        or1200_cpu_or1200_fpu_fpu_arith_done), .C(n62067), .Y(n2201) );
  NAND3xp33_ASAP7_75t_SL U70845 ( .A(n62095), .B(n62094), .C(n62093), .Y(
        n62092) );
  A2O1A1Ixp33_ASAP7_75t_SL U70846 ( .A1(n62095), .A2(n62094), .B(n62093), .C(
        n62092), .Y(n76320) );
  XOR2xp5_ASAP7_75t_SL U70847 ( .A(n64316), .B(n64321), .Y(n62138) );
  A2O1A1Ixp33_ASAP7_75t_SL U70848 ( .A1(n73923), .A2(n62110), .B(n62109), .C(
        n75731), .Y(n62112) );
  A2O1A1Ixp33_ASAP7_75t_SL U70849 ( .A1(n77097), .A2(n57209), .B(n75736), .C(
        n57218), .Y(n62111) );
  OAI211xp5_ASAP7_75t_SL U70850 ( .A1(or1200_cpu_or1200_mult_mac_n329), .A2(
        n75738), .B(n62112), .C(n62111), .Y(n62119) );
  OR2x2_ASAP7_75t_SL U70851 ( .A(n62122), .B(n62121), .Y(n75240) );
  NOR3xp33_ASAP7_75t_SL U70852 ( .A(n62126), .B(n62125), .C(n62124), .Y(n62127) );
  NAND3xp33_ASAP7_75t_SL U70853 ( .A(n3078), .B(n2071), .C(n2037), .Y(n62143)
         );
  NOR3xp33_ASAP7_75t_SL U70854 ( .A(n62145), .B(n62144), .C(n62143), .Y(n62147) );
  OR2x2_ASAP7_75t_SL U70855 ( .A(n62151), .B(n63712), .Y(n62154) );
  AND2x2_ASAP7_75t_SL U70856 ( .A(n62508), .B(n77163), .Y(n76707) );
  OR2x2_ASAP7_75t_SL U70857 ( .A(n62155), .B(n77209), .Y(n76507) );
  NAND4xp25_ASAP7_75t_SL U70858 ( .A(n62173), .B(n62172), .C(n62171), .D(
        n62170), .Y(n62179) );
  NAND4xp25_ASAP7_75t_SL U70859 ( .A(n62177), .B(n62176), .C(n62175), .D(
        n62174), .Y(n62178) );
  NAND3xp33_ASAP7_75t_SL U70860 ( .A(n62197), .B(n62196), .C(n62195), .Y(
        n62202) );
  A2O1A1Ixp33_ASAP7_75t_SL U70861 ( .A1(n62201), .A2(n75691), .B(n62202), .C(
        n62198), .Y(n62200) );
  OR3x1_ASAP7_75t_SL U70862 ( .A(n68810), .B(n75818), .C(n62206), .Y(n62209)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70863 ( .A1(n1179), .A2(n75645), .B(n62212), .C(
        n62211), .Y(n9275) );
  XOR2xp5_ASAP7_75t_SL U70864 ( .A(n1177), .B(n1179), .Y(n62213) );
  A2O1A1Ixp33_ASAP7_75t_SL U70865 ( .A1(n1175), .A2(n62218), .B(n62217), .C(
        n62216), .Y(n9273) );
  A2O1A1Ixp33_ASAP7_75t_SL U70866 ( .A1(n62222), .A2(n62221), .B(n62220), .C(
        n62224), .Y(n62223) );
  A2O1A1Ixp33_ASAP7_75t_SL U70867 ( .A1(n1171), .A2(n62227), .B(n62226), .C(
        n62225), .Y(n9271) );
  OR2x2_ASAP7_75t_SL U70868 ( .A(n62477), .B(n59544), .Y(n4066) );
  A2O1A1Ixp33_ASAP7_75t_SL U70869 ( .A1(n62233), .A2(n62232), .B(n62303), .C(
        n62231), .Y(n9270) );
  NOR3xp33_ASAP7_75t_SL U70870 ( .A(n62240), .B(n62239), .C(n62238), .Y(n62241) );
  A2O1A1Ixp33_ASAP7_75t_SL U70871 ( .A1(n62242), .A2(n76729), .B(n77601), .C(
        n62241), .Y(n62243) );
  OAI211xp5_ASAP7_75t_SL U70872 ( .A1(or1200_cpu_or1200_except_n272), .A2(
        n76731), .B(n62246), .C(n62245), .Y(n62249) );
  OR3x1_ASAP7_75t_SL U70873 ( .A(n62249), .B(n62248), .C(n62247), .Y(n62251)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70874 ( .A1(n77097), .A2(n76627), .B(n75736), .C(
        n78003), .Y(n62261) );
  OAI211xp5_ASAP7_75t_SL U70875 ( .A1(n62263), .A2(n76619), .B(n76792), .C(
        n77082), .Y(n62264) );
  OAI211xp5_ASAP7_75t_SL U70876 ( .A1(n76433), .A2(n75735), .B(n62265), .C(
        n62264), .Y(n62266) );
  NAND4xp25_ASAP7_75t_SL U70877 ( .A(n62283), .B(n62282), .C(n62281), .D(
        n62280), .Y(n62286) );
  AND2x2_ASAP7_75t_SL U70878 ( .A(n62289), .B(n62288), .Y(n76746) );
  OAI211xp5_ASAP7_75t_SL U70879 ( .A1(n76744), .A2(n77602), .B(n62294), .C(
        n62293), .Y(n62298) );
  OAI211xp5_ASAP7_75t_SL U70880 ( .A1(n76628), .A2(n77137), .B(n62301), .C(
        n62300), .Y(n9633) );
  OAI211xp5_ASAP7_75t_SL U70881 ( .A1(n62303), .A2(n62302), .B(n62397), .C(
        n75030), .Y(n62304) );
  OR2x2_ASAP7_75t_SL U70882 ( .A(n62477), .B(n59581), .Y(n4057) );
  AO21x1_ASAP7_75t_SL U70883 ( .A1(n62305), .A2(n75648), .B(n62401), .Y(n62394) );
  A2O1A1Ixp33_ASAP7_75t_SL U70884 ( .A1(n1165), .A2(n62397), .B(n62394), .C(
        n62306), .Y(n9268) );
  A2O1A1Ixp33_ASAP7_75t_SL U70885 ( .A1(n62323), .A2(n76729), .B(n62381), .C(
        n62322), .Y(n62324) );
  OAI211xp5_ASAP7_75t_SL U70886 ( .A1(or1200_cpu_or1200_except_n601), .A2(
        n59675), .B(n62328), .C(n62327), .Y(n62331) );
  NOR3xp33_ASAP7_75t_SL U70887 ( .A(n62331), .B(n62330), .C(n62329), .Y(n77609) );
  OAI211xp5_ASAP7_75t_SL U70888 ( .A1(n76795), .A2(n76851), .B(n62333), .C(
        n77082), .Y(n62335) );
  OAI211xp5_ASAP7_75t_SL U70889 ( .A1(n75735), .A2(n76445), .B(n62335), .C(
        n62334), .Y(n62336) );
  NAND4xp25_ASAP7_75t_SL U70890 ( .A(n62370), .B(n62369), .C(n62368), .D(
        n62367), .Y(n62380) );
  NAND4xp25_ASAP7_75t_SL U70891 ( .A(n62386), .B(n62385), .C(n62384), .D(
        n62383), .Y(n62387) );
  OAI211xp5_ASAP7_75t_SL U70892 ( .A1(n76654), .A2(n77137), .B(n62393), .C(
        n62392), .Y(n9631) );
  OR2x2_ASAP7_75t_SL U70893 ( .A(n62477), .B(n59554), .Y(n4053) );
  A2O1A1Ixp33_ASAP7_75t_SL U70894 ( .A1(n1163), .A2(n62396), .B(n58566), .C(
        n62395), .Y(n9267) );
  OR3x1_ASAP7_75t_SL U70895 ( .A(n1161), .B(n1165), .C(n1163), .Y(n63909) );
  A2O1A1Ixp33_ASAP7_75t_SL U70896 ( .A1(n62401), .A2(n62400), .B(n62399), .C(
        n62398), .Y(n62402) );
  OR2x2_ASAP7_75t_SL U70897 ( .A(n75648), .B(n62483), .Y(n62482) );
  OR2x2_ASAP7_75t_SL U70898 ( .A(n62477), .B(n59580), .Y(n4041) );
  A2O1A1Ixp33_ASAP7_75t_SL U70899 ( .A1(n1183), .A2(n62407), .B(n62482), .C(
        n62406), .Y(n9264) );
  NAND3xp33_ASAP7_75t_SL U70900 ( .A(n75731), .B(n62433), .C(n75862), .Y(
        n62435) );
  A2O1A1Ixp33_ASAP7_75t_SL U70901 ( .A1(n77097), .A2(n57128), .B(n75736), .C(
        n59387), .Y(n62434) );
  OAI211xp5_ASAP7_75t_SL U70902 ( .A1(or1200_cpu_or1200_mult_mac_n104), .A2(
        n64785), .B(n62435), .C(n62434), .Y(n62436) );
  NOR3xp33_ASAP7_75t_SL U70903 ( .A(n62438), .B(n62437), .C(n62436), .Y(n62439) );
  XOR2xp5_ASAP7_75t_SL U70904 ( .A(or1200_cpu_or1200_except_n512), .B(n62444), 
        .Y(n62450) );
  OAI211xp5_ASAP7_75t_SL U70905 ( .A1(n77626), .A2(n76796), .B(n62452), .C(
        n62451), .Y(n62453) );
  OAI211xp5_ASAP7_75t_SL U70906 ( .A1(n62456), .A2(n62455), .B(n62454), .C(
        n77112), .Y(n62457) );
  AND3x1_ASAP7_75t_SL U70907 ( .A(n62459), .B(n62458), .C(n62457), .Y(n62460)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70908 ( .A1(n77630), .A2(n62461), .B(n76744), .C(
        n62460), .Y(n62468) );
  A2O1A1Ixp33_ASAP7_75t_SL U70909 ( .A1(n62482), .A2(n62484), .B(n62481), .C(
        n62480), .Y(n9263) );
  A2O1A1Ixp33_ASAP7_75t_SL U70910 ( .A1(n62488), .A2(n62487), .B(n62491), .C(
        n62486), .Y(n9262) );
  AO21x1_ASAP7_75t_SL U70911 ( .A1(n75649), .A2(n77896), .B(n62490), .Y(n9261)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70912 ( .A1(n62496), .A2(n62495), .B(n62549), .C(
        n62494), .Y(n9260) );
  AO21x1_ASAP7_75t_SL U70913 ( .A1(n69163), .A2(n77041), .B(n62503), .Y(n62505) );
  NAND3xp33_ASAP7_75t_SL U70914 ( .A(n62511), .B(n62510), .C(n62509), .Y(
        n62512) );
  A2O1A1Ixp33_ASAP7_75t_SL U70915 ( .A1(n62522), .A2(n64775), .B(n62521), .C(
        n57126), .Y(n62523) );
  OAI211xp5_ASAP7_75t_SL U70916 ( .A1(n62525), .A2(n77078), .B(n62524), .C(
        n62523), .Y(n62539) );
  OAI211xp5_ASAP7_75t_SL U70917 ( .A1(n62531), .A2(n75587), .B(n62530), .C(
        n62529), .Y(n62538) );
  NOR3xp33_ASAP7_75t_SL U70918 ( .A(n62539), .B(n62538), .C(n62537), .Y(n62540) );
  OAI211xp5_ASAP7_75t_SL U70919 ( .A1(n77649), .A2(n76744), .B(n75358), .C(
        n62545), .Y(n62546) );
  A2O1A1Ixp33_ASAP7_75t_SL U70920 ( .A1(n1149), .A2(n62552), .B(n62551), .C(
        n62550), .Y(n9259) );
  NAND3xp33_ASAP7_75t_SL U70921 ( .A(n67251), .B(n75903), .C(n57178), .Y(
        n62584) );
  A2O1A1Ixp33_ASAP7_75t_SL U70922 ( .A1(n76028), .A2(n57422), .B(n62585), .C(
        n62584), .Y(n62586) );
  A2O1A1Ixp33_ASAP7_75t_SL U70923 ( .A1(n62595), .A2(n62594), .B(n59545), .C(
        n66244), .Y(n62596) );
  O2A1O1Ixp5_ASAP7_75t_SL U70924 ( .A1(n59614), .A2(n75925), .B(n62628), .C(
        n68079), .Y(n62602) );
  O2A1O1Ixp5_ASAP7_75t_SL U70925 ( .A1(n62980), .A2(n62603), .B(n62664), .C(
        n62602), .Y(n63016) );
  NAND3xp33_ASAP7_75t_SL U70926 ( .A(n62606), .B(n62605), .C(n62604), .Y(
        n62607) );
  MAJIxp5_ASAP7_75t_SL U70927 ( .A(n63018), .B(n63016), .C(n63014), .Y(n63032)
         );
  NAND3xp33_ASAP7_75t_SL U70928 ( .A(n66258), .B(n59079), .C(n62637), .Y(
        n62639) );
  XNOR2xp5_ASAP7_75t_SL U70929 ( .A(n59609), .B(n67343), .Y(n62693) );
  O2A1O1Ixp5_ASAP7_75t_SL U70930 ( .A1(n59618), .A2(n67585), .B(n62651), .C(
        n62650), .Y(n63075) );
  XNOR2xp5_ASAP7_75t_SL U70931 ( .A(n62773), .B(n63075), .Y(n62652) );
  O2A1O1Ixp5_ASAP7_75t_SL U70932 ( .A1(n62666), .A2(n62665), .B(n62664), .C(
        n62663), .Y(n62775) );
  XNOR2xp5_ASAP7_75t_SL U70933 ( .A(n62775), .B(n62774), .Y(n62680) );
  O2A1O1Ixp5_ASAP7_75t_SL U70934 ( .A1(n59479), .A2(n59592), .B(n57128), .C(
        n62700), .Y(n62701) );
  A2O1A1Ixp33_ASAP7_75t_SL U70935 ( .A1(n59510), .A2(n58439), .B(n62707), .C(
        n62706), .Y(n62997) );
  XNOR2xp5_ASAP7_75t_SL U70936 ( .A(n62730), .B(n62729), .Y(n62731) );
  MAJIxp5_ASAP7_75t_SL U70937 ( .A(n63044), .B(n57473), .C(n63043), .Y(n63482)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70938 ( .A1(n62746), .A2(n62745), .B(n58462), .C(
        n62744), .Y(n63060) );
  XNOR2xp5_ASAP7_75t_SL U70939 ( .A(n63059), .B(n63060), .Y(n62747) );
  XNOR2xp5_ASAP7_75t_SL U70940 ( .A(n63055), .B(n63056), .Y(n62752) );
  MAJIxp5_ASAP7_75t_SL U70941 ( .A(n62756), .B(n58510), .C(n62755), .Y(n63050)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U70942 ( .A1(n75900), .A2(n57180), .B(n62759), .C(
        n62758), .Y(n63088) );
  MAJIxp5_ASAP7_75t_SL U70943 ( .A(n62777), .B(n62776), .C(n62775), .Y(n63077)
         );
  XNOR2xp5_ASAP7_75t_SL U70944 ( .A(n62778), .B(n63077), .Y(n62779) );
  XNOR2xp5_ASAP7_75t_SL U70945 ( .A(n63050), .B(n63051), .Y(n62780) );
  O2A1O1Ixp5_ASAP7_75t_SL U70946 ( .A1(n63068), .A2(n62876), .B(n62782), .C(
        n67609), .Y(n62791) );
  O2A1O1Ixp5_ASAP7_75t_SL U70947 ( .A1(n62792), .A2(n62791), .B(n62790), .C(
        n62789), .Y(n62861) );
  A2O1A1Ixp33_ASAP7_75t_SL U70948 ( .A1(n75930), .A2(n57180), .B(n62803), .C(
        n62802), .Y(n62829) );
  XOR2xp5_ASAP7_75t_SL U70949 ( .A(n62829), .B(n62824), .Y(n62809) );
  XNOR2xp5_ASAP7_75t_SL U70950 ( .A(n62823), .B(n62809), .Y(n62858) );
  MAJIxp5_ASAP7_75t_SL U70951 ( .A(n62812), .B(n62811), .C(n62810), .Y(n63368)
         );
  XNOR2xp5_ASAP7_75t_SL U70952 ( .A(n62929), .B(n62930), .Y(n62821) );
  A2O1A1Ixp33_ASAP7_75t_SL U70953 ( .A1(n62830), .A2(n62829), .B(n62828), .C(
        n62827), .Y(n62916) );
  XNOR2xp5_ASAP7_75t_SL U70954 ( .A(n67228), .B(n59614), .Y(n62831) );
  A2O1A1Ixp33_ASAP7_75t_SL U70955 ( .A1(n62835), .A2(n62834), .B(n62833), .C(
        n62832), .Y(n62937) );
  XNOR2xp5_ASAP7_75t_SL U70956 ( .A(n62838), .B(n62934), .Y(n62839) );
  NAND3xp33_ASAP7_75t_SL U70957 ( .A(n58424), .B(n59565), .C(n62880), .Y(
        n62841) );
  A2O1A1Ixp33_ASAP7_75t_SL U70958 ( .A1(n75925), .A2(n57180), .B(n62842), .C(
        n62841), .Y(n62869) );
  O2A1O1Ixp5_ASAP7_75t_SL U70959 ( .A1(n62846), .A2(n62845), .B(n57159), .C(
        n62844), .Y(n62871) );
  XNOR2xp5_ASAP7_75t_SL U70960 ( .A(n59511), .B(n59503), .Y(n62848) );
  A2O1A1Ixp33_ASAP7_75t_SL U70961 ( .A1(n62855), .A2(n62854), .B(n62853), .C(
        n62852), .Y(n62948) );
  XNOR2xp5_ASAP7_75t_SL U70962 ( .A(n53458), .B(n62856), .Y(n62859) );
  XNOR2xp5_ASAP7_75t_SL U70963 ( .A(n62859), .B(n62858), .Y(n62860) );
  XNOR2xp5_ASAP7_75t_SL U70964 ( .A(n62869), .B(n62868), .Y(n62873) );
  XNOR2xp5_ASAP7_75t_SL U70965 ( .A(n62873), .B(n62872), .Y(n62905) );
  O2A1O1Ixp5_ASAP7_75t_SL U70966 ( .A1(n59618), .A2(n62883), .B(n62882), .C(
        n62881), .Y(n62907) );
  A2O1A1Ixp33_ASAP7_75t_SL U70967 ( .A1(n63298), .A2(n63297), .B(n63296), .C(
        n62899), .Y(n62900) );
  MAJIxp5_ASAP7_75t_SL U70968 ( .A(n62917), .B(n62915), .C(n62916), .Y(n62953)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70969 ( .A1(n64083), .A2(n59504), .B(n62920), .C(
        n62919), .Y(n62968) );
  O2A1O1Ixp5_ASAP7_75t_SL U70970 ( .A1(n59618), .A2(n53261), .B(n62925), .C(
        n62924), .Y(n62967) );
  XNOR2xp5_ASAP7_75t_SL U70971 ( .A(n62926), .B(n62967), .Y(n62927) );
  MAJIxp5_ASAP7_75t_SL U70972 ( .A(n62931), .B(n62930), .C(n62929), .Y(n62990)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70973 ( .A1(n62939), .A2(n62938), .B(n62937), .C(
        n62936), .Y(n62972) );
  XNOR2xp5_ASAP7_75t_SL U70974 ( .A(n62970), .B(n62971), .Y(n62944) );
  A2O1A1Ixp33_ASAP7_75t_SL U70975 ( .A1(n59620), .A2(n58439), .B(n62955), .C(
        n62954), .Y(n63007) );
  XNOR2xp5_ASAP7_75t_SL U70976 ( .A(n57109), .B(n67227), .Y(n62960) );
  MAJIxp5_ASAP7_75t_SL U70977 ( .A(n62968), .B(n62966), .C(n62967), .Y(n63003)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70978 ( .A1(n62985), .A2(n62974), .B(n62973), .C(
        n62972), .Y(n62975) );
  A2O1A1Ixp33_ASAP7_75t_SL U70979 ( .A1(n76028), .A2(n64424), .B(n62979), .C(
        n62978), .Y(n63011) );
  O2A1O1Ixp5_ASAP7_75t_SL U70980 ( .A1(n59504), .A2(n57108), .B(n62981), .C(
        n68079), .Y(n62982) );
  O2A1O1Ixp5_ASAP7_75t_SL U70981 ( .A1(n62984), .A2(n62983), .B(n58462), .C(
        n62982), .Y(n63012) );
  MAJIxp5_ASAP7_75t_SL U70982 ( .A(n62990), .B(n62991), .C(n62989), .Y(n63362)
         );
  MAJIxp5_ASAP7_75t_SL U70983 ( .A(n63013), .B(n63012), .C(n63011), .Y(n63034)
         );
  MAJIxp5_ASAP7_75t_SL U70984 ( .A(n63024), .B(n63023), .C(n63022), .Y(n63476)
         );
  MAJIxp5_ASAP7_75t_SL U70985 ( .A(n63035), .B(n63033), .C(n63034), .Y(n63040)
         );
  XNOR2xp5_ASAP7_75t_SL U70986 ( .A(n63040), .B(n63036), .Y(n63037) );
  MAJIxp5_ASAP7_75t_SL U70987 ( .A(n63042), .B(n63041), .C(n63040), .Y(n63047)
         );
  MAJIxp5_ASAP7_75t_SL U70988 ( .A(n63062), .B(n63061), .C(n63060), .Y(n63141)
         );
  NAND3xp33_ASAP7_75t_SL U70989 ( .A(n63210), .B(n64625), .C(n58481), .Y(
        n63065) );
  XNOR2xp5_ASAP7_75t_SL U70990 ( .A(n63157), .B(n58350), .Y(n63071) );
  MAJIxp5_ASAP7_75t_SL U70991 ( .A(n63078), .B(n63077), .C(n63076), .Y(n63109)
         );
  XNOR2xp5_ASAP7_75t_SL U70992 ( .A(n53317), .B(n75901), .Y(n63084) );
  XNOR2xp5_ASAP7_75t_SL U70993 ( .A(n59511), .B(n59606), .Y(n63149) );
  A2O1A1Ixp33_ASAP7_75t_SL U70994 ( .A1(n63094), .A2(n57347), .B(n63192), .C(
        n63673), .Y(n63835) );
  A2O1A1Ixp33_ASAP7_75t_SL U70995 ( .A1(n63130), .A2(n57180), .B(n63096), .C(
        n63095), .Y(n63137) );
  OAI211xp5_ASAP7_75t_SL U70996 ( .A1(n58207), .A2(n63188), .B(n63251), .C(
        n59588), .Y(n63185) );
  XNOR2xp5_ASAP7_75t_SL U70997 ( .A(n63234), .B(n63646), .Y(n63131) );
  MAJIxp5_ASAP7_75t_SL U70998 ( .A(n63142), .B(n63141), .C(n63140), .Y(n63166)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U70999 ( .A1(n75900), .A2(n67601), .B(n63146), .C(
        n63145), .Y(n63236) );
  MAJIxp5_ASAP7_75t_SL U71000 ( .A(n63164), .B(n58382), .C(n63162), .Y(n63686)
         );
  MAJIxp5_ASAP7_75t_SL U71001 ( .A(n63166), .B(n63167), .C(n63168), .Y(n63609)
         );
  NAND3xp33_ASAP7_75t_SL U71002 ( .A(n63183), .B(n67227), .C(n67738), .Y(
        n63802) );
  NAND3xp33_ASAP7_75t_SL U71003 ( .A(n63190), .B(n53291), .C(n63827), .Y(
        n63627) );
  O2A1O1Ixp5_ASAP7_75t_SL U71004 ( .A1(n75900), .A2(n67866), .B(n63194), .C(
        n63193), .Y(n63628) );
  MAJIxp5_ASAP7_75t_SL U71005 ( .A(n63201), .B(n63200), .C(n63199), .Y(n63626)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71006 ( .A1(n63205), .A2(n63204), .B(n68081), .C(
        n63203), .Y(n63640) );
  O2A1O1Ixp5_ASAP7_75t_SL U71007 ( .A1(n59618), .A2(n59660), .B(n63208), .C(
        n63207), .Y(n63639) );
  A2O1A1Ixp33_ASAP7_75t_SL U71008 ( .A1(n59508), .A2(n67343), .B(n63218), .C(
        n63217), .Y(n63219) );
  XNOR2xp5_ASAP7_75t_SL U71009 ( .A(n63620), .B(n63621), .Y(n63225) );
  XNOR2xp5_ASAP7_75t_SL U71010 ( .A(n63626), .B(n63227), .Y(n63608) );
  MAJIxp5_ASAP7_75t_SL U71011 ( .A(n63232), .B(n63231), .C(n63230), .Y(n63652)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71012 ( .A1(n63647), .A2(n63235), .B(n63646), .C(
        n63645), .Y(n63651) );
  MAJIxp5_ASAP7_75t_SL U71013 ( .A(n63238), .B(n63237), .C(n63236), .Y(n63650)
         );
  OAI211xp5_ASAP7_75t_SL U71014 ( .A1(n63879), .A2(n63244), .B(n64743), .C(
        n63256), .Y(n63687) );
  OAI222xp33_ASAP7_75t_SL U71015 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n108), .B1(n76633), .B2(n58720), .C1(n57105), .C2(or1200_cpu_or1200_mult_mac_n106), .Y(or1200_cpu_or1200_mult_mac_n1549)
         );
  OAI222xp33_ASAP7_75t_SL U71016 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n106), .B1(n76633), .B2(n59604), .C1(n57105), .C2(or1200_cpu_or1200_mult_mac_n104), .Y(or1200_cpu_or1200_mult_mac_n1548)
         );
  OAI222xp33_ASAP7_75t_SL U71017 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n104), .B1(n76633), .B2(n59508), .C1(n57105), .C2(or1200_cpu_or1200_mult_mac_n102), .Y(n52047) );
  OAI222xp33_ASAP7_75t_SL U71018 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n102), .B1(n76633), .B2(n67963), .C1(n57105), .C2(or1200_cpu_or1200_mult_mac_n100), .Y(n14249) );
  OAI222xp33_ASAP7_75t_SL U71019 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n98), .B1(n76633), .B2(n59477), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n96), .Y(
        or1200_cpu_or1200_mult_mac_n1544) );
  O2A1O1Ixp5_ASAP7_75t_SL U71020 ( .A1(n63252), .A2(n57119), .B(n63251), .C(
        n63250), .Y(n63659) );
  OAI222xp33_ASAP7_75t_SL U71021 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n96), .B1(n76633), .B2(n63659), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n94), .Y(n14251) );
  XOR2xp5_ASAP7_75t_SL U71022 ( .A(n63258), .B(n58306), .Y(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N17) );
  NAND3xp33_ASAP7_75t_SL U71023 ( .A(n63265), .B(
        or1200_cpu_or1200_mult_mac_n269), .C(or1200_cpu_or1200_mult_mac_n273), 
        .Y(n63262) );
  OR2x2_ASAP7_75t_SL U71024 ( .A(or1200_cpu_or1200_mult_mac_n289), .B(
        or1200_cpu_or1200_mult_mac_n143), .Y(n63375) );
  OR2x2_ASAP7_75t_SL U71025 ( .A(or1200_cpu_or1200_mult_mac_n291), .B(
        or1200_cpu_or1200_mult_mac_n145), .Y(n63307) );
  AO21x1_ASAP7_75t_SL U71026 ( .A1(n63339), .A2(n63316), .B(n63338), .Y(n63318) );
  A2O1A1Ixp33_ASAP7_75t_SL U71027 ( .A1(or1200_cpu_or1200_mult_mac_n295), .A2(
        n63325), .B(n63324), .C(n63323), .Y(n63384) );
  A2O1A1Ixp33_ASAP7_75t_SL U71028 ( .A1(n63342), .A2(n63373), .B(n63379), .C(
        n63341), .Y(n63352) );
  XNOR2xp5_ASAP7_75t_SL U71029 ( .A(n63356), .B(n63351), .Y(n63359) );
  AO21x1_ASAP7_75t_SL U71030 ( .A1(n63376), .A2(n63352), .B(n63371), .Y(n63355) );
  OAI211xp5_ASAP7_75t_SL U71031 ( .A1(n63375), .A2(n63374), .B(n63373), .C(
        n63378), .Y(n63381) );
  A2O1A1Ixp33_ASAP7_75t_SL U71032 ( .A1(n63383), .A2(n63382), .B(n63381), .C(
        n63380), .Y(n63461) );
  NAND3xp33_ASAP7_75t_SL U71033 ( .A(n63391), .B(n63390), .C(n63389), .Y(
        n63392) );
  NAND3xp33_ASAP7_75t_SL U71034 ( .A(n63398), .B(n63393), .C(n63392), .Y(
        n63403) );
  XOR2xp5_ASAP7_75t_SL U71035 ( .A(n63417), .B(n63414), .Y(n63420) );
  XNOR2xp5_ASAP7_75t_SL U71036 ( .A(n63417), .B(n63416), .Y(n63418) );
  XNOR2xp5_ASAP7_75t_SL U71037 ( .A(n63437), .B(n63436), .Y(n63438) );
  OAI211xp5_ASAP7_75t_SL U71038 ( .A1(n63522), .A2(n63441), .B(n63454), .C(
        n57080), .Y(n63442) );
  OAI211xp5_ASAP7_75t_SL U71039 ( .A1(or1200_cpu_or1200_mult_mac_n163), .A2(
        n76889), .B(n63443), .C(n63442), .Y(or1200_cpu_or1200_mult_mac_n1582)
         );
  AND2x2_ASAP7_75t_SL U71040 ( .A(n63520), .B(n63506), .Y(n63462) );
  XOR2xp5_ASAP7_75t_SL U71041 ( .A(n63462), .B(n63467), .Y(n63465) );
  NAND3xp33_ASAP7_75t_SL U71042 ( .A(n63461), .B(n63460), .C(n63459), .Y(
        n65087) );
  XOR2xp5_ASAP7_75t_SL U71043 ( .A(n63462), .B(n63468), .Y(n63463) );
  XOR2xp5_ASAP7_75t_SL U71044 ( .A(n63470), .B(n63484), .Y(n63473) );
  XOR2xp5_ASAP7_75t_SL U71045 ( .A(n63470), .B(n63469), .Y(n63471) );
  MAJIxp5_ASAP7_75t_SL U71046 ( .A(n63480), .B(n63479), .C(n63478), .Y(n76226)
         );
  AND2x2_ASAP7_75t_SL U71047 ( .A(n63504), .B(n63503), .Y(n63508) );
  XOR2xp5_ASAP7_75t_SL U71048 ( .A(n63508), .B(n63509), .Y(n63495) );
  XOR2xp5_ASAP7_75t_SL U71049 ( .A(n53459), .B(n63499), .Y(n52049) );
  A2O1A1Ixp33_ASAP7_75t_SL U71050 ( .A1(n63506), .A2(n63505), .B(n63519), .C(
        n63504), .Y(n63517) );
  AO21x1_ASAP7_75t_SL U71051 ( .A1(n63512), .A2(n63534), .B(n63511), .Y(n63514) );
  OAI211xp5_ASAP7_75t_SL U71052 ( .A1(n63530), .A2(n63522), .B(n63521), .C(
        n63520), .Y(n63524) );
  NAND3xp33_ASAP7_75t_SL U71053 ( .A(n63528), .B(n63526), .C(n63525), .Y(
        n63781) );
  OAI31xp33_ASAP7_75t_SL U71054 ( .A1(n63531), .A2(n63530), .A3(n63529), .B(
        n63528), .Y(n63780) );
  O2A1O1Ixp5_ASAP7_75t_SL U71055 ( .A1(n63541), .A2(n63540), .B(n63539), .C(
        n63538), .Y(n65089) );
  OAI222xp33_ASAP7_75t_SL U71056 ( .A1(n76633), .A2(n57172), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n92), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n94), .Y(or1200_cpu_or1200_mult_mac_n1542)
         );
  XNOR2xp5_ASAP7_75t_SL U71057 ( .A(n63550), .B(n63549), .Y(n76313) );
  OAI211xp5_ASAP7_75t_SL U71058 ( .A1(or1200_cpu_or1200_mult_mac_n177), .A2(
        n63555), .B(n63554), .C(n63553), .Y(n63556) );
  OAI211xp5_ASAP7_75t_SL U71059 ( .A1(or1200_cpu_or1200_except_n224), .A2(
        n57170), .B(n63559), .C(n63558), .Y(n63561) );
  A2O1A1Ixp33_ASAP7_75t_SL U71060 ( .A1(n63582), .A2(n63581), .B(n75872), .C(
        n63580), .Y(n63592) );
  NOR3xp33_ASAP7_75t_SL U71061 ( .A(n63598), .B(n63597), .C(n63596), .Y(n63599) );
  OAI211xp5_ASAP7_75t_SL U71062 ( .A1(n77651), .A2(n76744), .B(n75358), .C(
        n63599), .Y(n63600) );
  XNOR2xp5_ASAP7_75t_SL U71063 ( .A(n63607), .B(n63606), .Y(n63612) );
  MAJIxp5_ASAP7_75t_SL U71064 ( .A(n63612), .B(n63611), .C(n63610), .Y(n63683)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71065 ( .A1(n63617), .A2(n63616), .B(n57375), .C(
        n63615), .Y(n63853) );
  MAJIxp5_ASAP7_75t_SL U71066 ( .A(n63620), .B(n63621), .C(n63622), .Y(n64060)
         );
  MAJIxp5_ASAP7_75t_SL U71067 ( .A(n63629), .B(n63628), .C(n63627), .Y(n63851)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71068 ( .A1(n75927), .A2(n58536), .B(n63839), .C(
        n57706), .Y(n63633) );
  XNOR2xp5_ASAP7_75t_SL U71069 ( .A(n63833), .B(n63832), .Y(n63637) );
  MAJIxp5_ASAP7_75t_SL U71070 ( .A(n63638), .B(n63639), .C(n63640), .Y(n63850)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71071 ( .A1(n57111), .A2(n53242), .B(n63647), .C(
        n63646), .Y(n63648) );
  XNOR2xp5_ASAP7_75t_SL U71072 ( .A(n56864), .B(n58938), .Y(n63678) );
  A2O1A1Ixp33_ASAP7_75t_SL U71073 ( .A1(n63678), .A2(n57271), .B(n63677), .C(
        n63676), .Y(n63858) );
  XNOR2xp5_ASAP7_75t_SL U71074 ( .A(n63886), .B(n63885), .Y(
        or1200_cpu_or1200_mult_mac_or1200_gmultp2_32x32_N19) );
  A2O1A1Ixp33_ASAP7_75t_SL U71075 ( .A1(n76822), .A2(n63689), .B(n63688), .C(
        n74954), .Y(n63693) );
  OR2x2_ASAP7_75t_SL U71076 ( .A(n69347), .B(n63706), .Y(n74924) );
  AND3x1_ASAP7_75t_SL U71077 ( .A(n63718), .B(or1200_cpu_or1200_except_n565), 
        .C(n63707), .Y(n63708) );
  OAI211xp5_ASAP7_75t_SL U71078 ( .A1(or1200_cpu_or1200_except_n326), .A2(
        n57088), .B(n63728), .C(n63727), .Y(or1200_cpu_or1200_except_n1774) );
  OAI211xp5_ASAP7_75t_SL U71079 ( .A1(n77603), .A2(n59494), .B(n63733), .C(
        n63732), .Y(n63736) );
  OAI211xp5_ASAP7_75t_SL U71080 ( .A1(n59708), .A2(n57124), .B(n63746), .C(
        n63745), .Y(n63747) );
  AND2x2_ASAP7_75t_SL U71081 ( .A(n63747), .B(n57100), .Y(n76568) );
  O2A1O1Ixp5_ASAP7_75t_SL U71082 ( .A1(n63758), .A2(n76813), .B(n63757), .C(
        n63756), .Y(n63952) );
  OR2x2_ASAP7_75t_SL U71083 ( .A(or1200_cpu_or1200_except_n575), .B(n1739), 
        .Y(or1200_cpu_or1200_except_n1697) );
  A2O1A1Ixp33_ASAP7_75t_SL U71084 ( .A1(n74639), .A2(n77287), .B(n63769), .C(
        n63768), .Y(or1200_pic_N66) );
  O2A1O1Ixp5_ASAP7_75t_SL U71085 ( .A1(n63782), .A2(n63781), .B(n63780), .C(
        n63779), .Y(n65099) );
  MAJIxp5_ASAP7_75t_SL U71086 ( .A(n63792), .B(n63791), .C(n63790), .Y(n63876)
         );
  NAND3xp33_ASAP7_75t_SL U71087 ( .A(n63795), .B(n63794), .C(n63793), .Y(
        n63798) );
  AO21x1_ASAP7_75t_SL U71088 ( .A1(n63801), .A2(n57501), .B(n63800), .Y(n64676) );
  A2O1A1Ixp33_ASAP7_75t_SL U71089 ( .A1(n58424), .A2(n77715), .B(n76679), .C(
        n63809), .Y(n63811) );
  XNOR2xp5_ASAP7_75t_SL U71090 ( .A(n63817), .B(n63816), .Y(n63820) );
  MAJIxp5_ASAP7_75t_SL U71091 ( .A(n63851), .B(n63850), .C(n63849), .Y(n64063)
         );
  AO21x1_ASAP7_75t_SL U71092 ( .A1(n63856), .A2(n63855), .B(n63854), .Y(n64061) );
  MAJIxp5_ASAP7_75t_SL U71093 ( .A(n63871), .B(n63872), .C(n63873), .Y(n64018)
         );
  XNOR2xp5_ASAP7_75t_SL U71094 ( .A(n64017), .B(n64018), .Y(n63874) );
  OAI31xp33_ASAP7_75t_SL U71095 ( .A1(n63898), .A2(n64172), .A3(n76906), .B(
        n63897), .Y(n63899) );
  A2O1A1Ixp33_ASAP7_75t_SL U71096 ( .A1(n1143), .A2(n63918), .B(n63917), .C(
        n63916), .Y(n9256) );
  OAI211xp5_ASAP7_75t_SL U71097 ( .A1(or1200_cpu_or1200_except_n353), .A2(
        n57088), .B(n63924), .C(n63923), .Y(or1200_cpu_or1200_except_n1765) );
  OAI211xp5_ASAP7_75t_SL U71098 ( .A1(or1200_cpu_or1200_except_n347), .A2(
        n57088), .B(n63929), .C(n63928), .Y(or1200_cpu_or1200_except_n1767) );
  OAI211xp5_ASAP7_75t_SL U71099 ( .A1(or1200_cpu_or1200_except_n344), .A2(
        n57088), .B(n63934), .C(n63933), .Y(or1200_cpu_or1200_except_n1768) );
  A2O1A1Ixp33_ASAP7_75t_SL U71100 ( .A1(n74957), .A2(n74956), .B(n63940), .C(
        n63939), .Y(n63941) );
  OAI211xp5_ASAP7_75t_SL U71101 ( .A1(or1200_cpu_or1200_except_n332), .A2(
        n57088), .B(n63951), .C(n63950), .Y(or1200_cpu_or1200_except_n1772) );
  OR2x2_ASAP7_75t_SL U71102 ( .A(n63963), .B(n63981), .Y(n63967) );
  OAI211xp5_ASAP7_75t_SL U71103 ( .A1(or1200_cpu_or1200_except_n335), .A2(
        n57088), .B(n63962), .C(n63961), .Y(or1200_cpu_or1200_except_n1771) );
  OAI211xp5_ASAP7_75t_SL U71104 ( .A1(or1200_cpu_or1200_except_n338), .A2(
        n57088), .B(n63974), .C(n63973), .Y(or1200_cpu_or1200_except_n1770) );
  OAI211xp5_ASAP7_75t_SL U71105 ( .A1(or1200_cpu_or1200_except_n341), .A2(
        n57088), .B(n63992), .C(n63991), .Y(or1200_cpu_or1200_except_n1769) );
  OAI222xp33_ASAP7_75t_SL U71106 ( .A1(n76633), .A2(n59596), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n88), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n90), .Y(n12986) );
  MAJIxp5_ASAP7_75t_SL U71107 ( .A(n64021), .B(n64020), .C(n64019), .Y(n64094)
         );
  XNOR2xp5_ASAP7_75t_SL U71108 ( .A(n57107), .B(n57178), .Y(n64040) );
  MAJIxp5_ASAP7_75t_SL U71109 ( .A(n64048), .B(n64049), .C(n53494), .Y(n64437)
         );
  MAJIxp5_ASAP7_75t_SL U71110 ( .A(n64050), .B(n64051), .C(n64052), .Y(n64436)
         );
  MAJIxp5_ASAP7_75t_SL U71111 ( .A(n64069), .B(n64068), .C(n64067), .Y(n64723)
         );
  NOR3xp33_ASAP7_75t_SL U71112 ( .A(n68102), .B(n75912), .C(n59594), .Y(n64084) );
  NOR3xp33_ASAP7_75t_SL U71113 ( .A(n76078), .B(n68010), .C(n59594), .Y(n64082) );
  AO21x1_ASAP7_75t_SL U71114 ( .A1(n64097), .A2(n74595), .B(n75882), .Y(n64145) );
  A2O1A1Ixp33_ASAP7_75t_SL U71115 ( .A1(n77097), .A2(n77717), .B(n75741), .C(
        n64114), .Y(n64115) );
  OAI211xp5_ASAP7_75t_SL U71116 ( .A1(n75865), .A2(n64295), .B(n64130), .C(
        n64129), .Y(n64134) );
  A2O1A1Ixp33_ASAP7_75t_SL U71117 ( .A1(or1200_cpu_or1200_except_n528), .A2(
        n64142), .B(n64141), .C(n64140), .Y(n64143) );
  OAI211xp5_ASAP7_75t_SL U71118 ( .A1(or1200_cpu_or1200_except_n356), .A2(
        n57088), .B(n64161), .C(n64160), .Y(or1200_cpu_or1200_except_n1764) );
  OR2x2_ASAP7_75t_SL U71119 ( .A(n2664), .B(or1200_cpu_or1200_except_n634), 
        .Y(n64264) );
  A2O1A1Ixp33_ASAP7_75t_SL U71120 ( .A1(n64176), .A2(n57079), .B(n64175), .C(
        n64174), .Y(n64177) );
  OAI211xp5_ASAP7_75t_SL U71121 ( .A1(or1200_cpu_or1200_mult_mac_n181), .A2(
        n76889), .B(n64178), .C(n64177), .Y(or1200_cpu_or1200_mult_mac_n1573)
         );
  XOR2xp5_ASAP7_75t_SL U71122 ( .A(n1141), .B(n1143), .Y(n64179) );
  A2O1A1Ixp33_ASAP7_75t_SL U71123 ( .A1(n64197), .A2(n64196), .B(n64195), .C(
        n64194), .Y(n64198) );
  A2O1A1Ixp33_ASAP7_75t_SL U71124 ( .A1(n64203), .A2(n74047), .B(n74081), .C(
        n64202), .Y(n64254) );
  OAI211xp5_ASAP7_75t_SL U71125 ( .A1(n75819), .A2(n65165), .B(n64211), .C(
        n64210), .Y(n64212) );
  A2O1A1Ixp33_ASAP7_75t_SL U71126 ( .A1(n64225), .A2(n78005), .B(n64224), .C(
        n75332), .Y(n64226) );
  NAND3xp33_ASAP7_75t_SL U71127 ( .A(n64228), .B(n64227), .C(n64226), .Y(
        n64246) );
  A2O1A1Ixp33_ASAP7_75t_SL U71128 ( .A1(n77097), .A2(n64241), .B(n75736), .C(
        n77732), .Y(n64242) );
  OAI211xp5_ASAP7_75t_SL U71129 ( .A1(or1200_cpu_or1200_mult_mac_n337), .A2(
        n75738), .B(n64243), .C(n64242), .Y(n64244) );
  OAI211xp5_ASAP7_75t_SL U71130 ( .A1(n64248), .A2(n75602), .B(n75607), .C(
        n64247), .Y(n64249) );
  OAI211xp5_ASAP7_75t_SL U71131 ( .A1(n64251), .A2(n64755), .B(n64857), .C(
        n77112), .Y(n64252) );
  NAND3xp33_ASAP7_75t_SL U71132 ( .A(n64254), .B(n64253), .C(n64252), .Y(
        n64255) );
  AO21x1_ASAP7_75t_SL U71133 ( .A1(n77031), .A2(n76271), .B(n64255), .Y(n77870) );
  AO21x1_ASAP7_75t_SL U71134 ( .A1(n57073), .A2(n77870), .B(n64256), .Y(n1591)
         );
  OAI211xp5_ASAP7_75t_SL U71135 ( .A1(or1200_cpu_or1200_except_n362), .A2(
        n57088), .B(n64263), .C(n64262), .Y(or1200_cpu_or1200_except_n1762) );
  O2A1O1Ixp5_ASAP7_75t_SL U71136 ( .A1(n64287), .A2(n64286), .B(n77659), .C(
        n64285), .Y(n77654) );
  XOR2xp5_ASAP7_75t_SL U71137 ( .A(n59578), .B(n59561), .Y(n76453) );
  OAI31xp33_ASAP7_75t_SL U71138 ( .A1(n75713), .A2(n73925), .A3(n75702), .B(
        n64291), .Y(n64292) );
  OAI211xp5_ASAP7_75t_SL U71139 ( .A1(n59586), .A2(n75347), .B(n64299), .C(
        n64298), .Y(n64300) );
  OAI211xp5_ASAP7_75t_SL U71140 ( .A1(n64313), .A2(n75315), .B(n64312), .C(
        n64311), .Y(n64314) );
  A2O1A1Ixp33_ASAP7_75t_SL U71141 ( .A1(n64321), .A2(n64320), .B(n64319), .C(
        n64318), .Y(n64322) );
  OAI211xp5_ASAP7_75t_SL U71142 ( .A1(n77654), .A2(n64324), .B(n64323), .C(
        n64322), .Y(n64325) );
  AO21x1_ASAP7_75t_SL U71143 ( .A1(n76305), .A2(n64326), .B(n64325), .Y(n64329) );
  O2A1O1Ixp5_ASAP7_75t_SL U71144 ( .A1(n67944), .A2(n67826), .B(n64333), .C(
        n57706), .Y(n64342) );
  A2O1A1Ixp33_ASAP7_75t_SL U71145 ( .A1(n67432), .A2(n57243), .B(n64334), .C(
        n64338), .Y(n64341) );
  MAJIxp5_ASAP7_75t_SL U71146 ( .A(n64346), .B(n64345), .C(n64344), .Y(n64433)
         );
  MAJIxp5_ASAP7_75t_SL U71147 ( .A(n64432), .B(n64433), .C(n64431), .Y(n64523)
         );
  XNOR2xp5_ASAP7_75t_SL U71148 ( .A(n67343), .B(n59596), .Y(n64501) );
  NAND3xp33_ASAP7_75t_SL U71149 ( .A(n66258), .B(n59561), .C(n64355), .Y(
        n64354) );
  NOR3xp33_ASAP7_75t_SL U71150 ( .A(n67451), .B(n58849), .C(n64359), .Y(n64360) );
  O2A1O1Ixp5_ASAP7_75t_SL U71151 ( .A1(n59618), .A2(n57394), .B(n64363), .C(
        n64362), .Y(n64418) );
  XNOR2xp5_ASAP7_75t_SL U71152 ( .A(n67638), .B(n57505), .Y(n64369) );
  O2A1O1Ixp5_ASAP7_75t_SL U71153 ( .A1(n58753), .A2(n59618), .B(n64372), .C(
        n64371), .Y(n64530) );
  XNOR2xp5_ASAP7_75t_SL U71154 ( .A(n59513), .B(n59601), .Y(n64373) );
  MAJIxp5_ASAP7_75t_SL U71155 ( .A(n64438), .B(n64439), .C(n64388), .Y(n64527)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71156 ( .A1(n59604), .A2(n67569), .B(n64391), .C(
        n67912), .Y(n64392) );
  A2O1A1Ixp33_ASAP7_75t_SL U71157 ( .A1(n64400), .A2(n64399), .B(n64426), .C(
        n64398), .Y(n64539) );
  XNOR2xp5_ASAP7_75t_SL U71158 ( .A(n64600), .B(n64599), .Y(n64411) );
  MAJIxp5_ASAP7_75t_SL U71159 ( .A(n64415), .B(n64414), .C(n64416), .Y(n64688)
         );
  XNOR2xp5_ASAP7_75t_SL U71160 ( .A(n64433), .B(n64432), .Y(n64434) );
  MAJIxp5_ASAP7_75t_SL U71161 ( .A(n64703), .B(n64702), .C(n64701), .Y(n64657)
         );
  MAJIxp5_ASAP7_75t_SL U71162 ( .A(n64657), .B(n64658), .C(n64659), .Y(n64694)
         );
  MAJIxp5_ASAP7_75t_SL U71163 ( .A(n64672), .B(n64674), .C(n64671), .Y(n64692)
         );
  MAJIxp5_ASAP7_75t_SL U71164 ( .A(n64692), .B(n64465), .C(n64689), .Y(n64553)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71165 ( .A1(n64478), .A2(n64477), .B(n64476), .C(
        n64475), .Y(n64556) );
  MAJIxp5_ASAP7_75t_SL U71166 ( .A(n64587), .B(n58341), .C(n57143), .Y(n64522)
         );
  NAND3xp33_ASAP7_75t_SL U71167 ( .A(n64606), .B(n67609), .C(n64605), .Y(
        n64576) );
  XOR2xp5_ASAP7_75t_SL U71168 ( .A(n64520), .B(n64588), .Y(n64521) );
  XNOR2xp5_ASAP7_75t_SL U71169 ( .A(n64522), .B(n64521), .Y(n64554) );
  MAJIxp5_ASAP7_75t_SL U71170 ( .A(n64523), .B(n64524), .C(n64525), .Y(n64594)
         );
  MAJIxp5_ASAP7_75t_SL U71171 ( .A(n64526), .B(n64527), .C(n64528), .Y(n64593)
         );
  NAND3xp33_ASAP7_75t_SL U71172 ( .A(n64531), .B(n64530), .C(n64529), .Y(
        n64533) );
  NAND3xp33_ASAP7_75t_SL U71173 ( .A(n64549), .B(n64548), .C(n64696), .Y(
        n64551) );
  MAJIxp5_ASAP7_75t_SL U71174 ( .A(n64554), .B(n64553), .C(n64552), .Y(n64872)
         );
  NAND3xp33_ASAP7_75t_SL U71175 ( .A(n64577), .B(n64576), .C(n64583), .Y(
        n64578) );
  NAND3xp33_ASAP7_75t_SL U71176 ( .A(n64582), .B(n64590), .C(n64581), .Y(
        n64586) );
  MAJIxp5_ASAP7_75t_SL U71177 ( .A(n64594), .B(n64593), .C(n64592), .Y(n64913)
         );
  OAI211xp5_ASAP7_75t_SL U71178 ( .A1(n76028), .A2(n67740), .B(n58155), .C(
        n64608), .Y(n64610) );
  XNOR2xp5_ASAP7_75t_SL U71179 ( .A(n59598), .B(n75927), .Y(n64611) );
  XNOR2xp5_ASAP7_75t_SL U71180 ( .A(n67343), .B(n59601), .Y(n64936) );
  NAND3xp33_ASAP7_75t_SL U71181 ( .A(n64626), .B(n57900), .C(n58481), .Y(
        n64627) );
  XNOR2xp5_ASAP7_75t_SL U71182 ( .A(n64884), .B(n64637), .Y(n64641) );
  NAND3xp33_ASAP7_75t_SL U71183 ( .A(n67748), .B(n58919), .C(n59615), .Y(
        n64644) );
  XNOR2xp5_ASAP7_75t_SL U71184 ( .A(n58402), .B(n59620), .Y(n64647) );
  NAND3xp33_ASAP7_75t_SL U71185 ( .A(n57877), .B(n64676), .C(n64675), .Y(
        n64679) );
  A2O1A1Ixp33_ASAP7_75t_SL U71186 ( .A1(n64680), .A2(n64679), .B(n64678), .C(
        n64677), .Y(n64681) );
  MAJIxp5_ASAP7_75t_SL U71187 ( .A(n64713), .B(n58395), .C(n64715), .Y(n65107)
         );
  NOR3xp33_ASAP7_75t_SL U71188 ( .A(n64718), .B(n64717), .C(n64716), .Y(n64720) );
  MAJIxp5_ASAP7_75t_SL U71189 ( .A(n64724), .B(n64723), .C(n58374), .Y(n64734)
         );
  NAND3xp33_ASAP7_75t_SL U71190 ( .A(n65110), .B(n74991), .C(n64739), .Y(
        n64740) );
  XOR2xp5_ASAP7_75t_SL U71191 ( .A(n64753), .B(n64870), .Y(n52055) );
  OAI222xp33_ASAP7_75t_SL U71192 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n82), .B1(n76633), .B2(n57491), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n80), .Y(n12980) );
  XOR2xp5_ASAP7_75t_SL U71193 ( .A(or1200_cpu_or1200_except_n536), .B(n75549), 
        .Y(n64800) );
  OAI211xp5_ASAP7_75t_SL U71194 ( .A1(n75871), .A2(n75838), .B(n64778), .C(
        n64777), .Y(n64793) );
  OAI31xp33_ASAP7_75t_SL U71195 ( .A1(n64784), .A2(n64783), .A3(n64782), .B(
        n64781), .Y(n75839) );
  A2O1A1Ixp33_ASAP7_75t_SL U71196 ( .A1(n77097), .A2(n77730), .B(n75741), .C(
        n74776), .Y(n64791) );
  XOR2xp5_ASAP7_75t_SL U71197 ( .A(n57068), .B(n59530), .Y(n76339) );
  OAI211xp5_ASAP7_75t_SL U71198 ( .A1(or1200_cpu_or1200_mult_mac_n189), .A2(
        n75723), .B(n64787), .C(n64786), .Y(n64788) );
  OAI211xp5_ASAP7_75t_SL U71199 ( .A1(n75839), .A2(n77103), .B(n64791), .C(
        n64790), .Y(n64792) );
  OA21x2_ASAP7_75t_SL U71200 ( .A1(n64824), .A2(n64823), .B(n64822), .Y(n77665) );
  OAI211xp5_ASAP7_75t_SL U71201 ( .A1(n57500), .A2(n75722), .B(n64827), .C(
        n64826), .Y(n64828) );
  OAI211xp5_ASAP7_75t_SL U71202 ( .A1(n75587), .A2(n64834), .B(n64833), .C(
        n64832), .Y(n64851) );
  NOR3xp33_ASAP7_75t_SL U71203 ( .A(n64838), .B(n64837), .C(n64836), .Y(n75703) );
  OAI211xp5_ASAP7_75t_SL U71204 ( .A1(n75703), .A2(n75710), .B(n64842), .C(
        n64841), .Y(n64846) );
  OAI31xp33_ASAP7_75t_SL U71205 ( .A1(n64846), .A2(n64845), .A3(n64844), .B(
        n75731), .Y(n64847) );
  A2O1A1Ixp33_ASAP7_75t_SL U71206 ( .A1(n75338), .A2(n64848), .B(n59528), .C(
        n64847), .Y(n64850) );
  NOR3xp33_ASAP7_75t_SL U71207 ( .A(n64851), .B(n64850), .C(n64849), .Y(n64852) );
  OAI211xp5_ASAP7_75t_SL U71208 ( .A1(n64863), .A2(n64862), .B(n64861), .C(
        n64860), .Y(n64864) );
  MAJIxp5_ASAP7_75t_SL U71209 ( .A(n64873), .B(n64872), .C(n58337), .Y(n64987)
         );
  NAND3xp33_ASAP7_75t_SL U71210 ( .A(n64877), .B(n64876), .C(n64875), .Y(
        n64880) );
  MAJIxp5_ASAP7_75t_SL U71211 ( .A(n64886), .B(n64885), .C(n64884), .Y(n65050)
         );
  XNOR2xp5_ASAP7_75t_SL U71212 ( .A(n64901), .B(n64900), .Y(n64902) );
  MAJIxp5_ASAP7_75t_SL U71213 ( .A(n64904), .B(n64905), .C(n64906), .Y(n64992)
         );
  MAJIxp5_ASAP7_75t_SL U71214 ( .A(n64913), .B(n64912), .C(n64911), .Y(n64989)
         );
  XNOR2xp5_ASAP7_75t_SL U71215 ( .A(n59605), .B(n76078), .Y(n65059) );
  XNOR2xp5_ASAP7_75t_SL U71216 ( .A(n59601), .B(n67288), .Y(n64934) );
  O2A1O1Ixp5_ASAP7_75t_SL U71217 ( .A1(n67264), .A2(n64959), .B(n67511), .C(
        n64958), .Y(n64961) );
  NOR3xp33_ASAP7_75t_SL U71218 ( .A(n57177), .B(n64965), .C(n58542), .Y(n64970) );
  XNOR2xp5_ASAP7_75t_SL U71219 ( .A(n57107), .B(n57110), .Y(n64969) );
  MAJIxp5_ASAP7_75t_SL U71220 ( .A(n64991), .B(n64990), .C(n53257), .Y(n65070)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71221 ( .A1(n59648), .A2(n57422), .B(n65045), .C(
        n65044), .Y(n68171) );
  MAJIxp5_ASAP7_75t_SL U71222 ( .A(n65051), .B(n65050), .C(n65049), .Y(n68255)
         );
  OAI222xp33_ASAP7_75t_SL U71223 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n80), .B1(n76633), .B2(n65072), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n78), .Y(
        or1200_cpu_or1200_mult_mac_n1535) );
  NAND3xp33_ASAP7_75t_SL U71224 ( .A(n65085), .B(n65084), .C(n65083), .Y(
        n65086) );
  OR2x2_ASAP7_75t_SL U71225 ( .A(n65128), .B(n65130), .Y(n65100) );
  NAND3xp33_ASAP7_75t_SL U71226 ( .A(n65093), .B(n65092), .C(n65091), .Y(
        n65097) );
  A2O1A1Ixp33_ASAP7_75t_SL U71227 ( .A1(n65099), .A2(n65098), .B(n65097), .C(
        n65096), .Y(n65169) );
  AND2x2_ASAP7_75t_SL U71228 ( .A(n65141), .B(n65169), .Y(n65126) );
  XNOR2xp5_ASAP7_75t_SL U71229 ( .A(n65109), .B(n65108), .Y(n65116) );
  AND2x2_ASAP7_75t_SL U71230 ( .A(n74991), .B(n65110), .Y(n65117) );
  O2A1O1Ixp5_ASAP7_75t_SL U71231 ( .A1(n65119), .A2(n65118), .B(n65117), .C(
        n65116), .Y(n65120) );
  XOR2xp5_ASAP7_75t_SL U71232 ( .A(n65135), .B(n65127), .Y(n65138) );
  OR3x1_ASAP7_75t_SL U71233 ( .A(n65132), .B(n65129), .C(n65128), .Y(n65173)
         );
  NOR3xp33_ASAP7_75t_SL U71234 ( .A(n65148), .B(n65147), .C(n65133), .Y(n65134) );
  XOR2xp5_ASAP7_75t_SL U71235 ( .A(n65135), .B(n65134), .Y(n65136) );
  XOR2xp5_ASAP7_75t_SL U71236 ( .A(or1200_cpu_or1200_mult_mac_n337), .B(
        or1200_cpu_or1200_mult_mac_n191), .Y(n65175) );
  NAND3xp33_ASAP7_75t_SL U71237 ( .A(n65163), .B(n65162), .C(n65161), .Y(
        n65167) );
  A2O1A1Ixp33_ASAP7_75t_SL U71238 ( .A1(n65169), .A2(n65168), .B(n65167), .C(
        n65166), .Y(n68795) );
  XOR2xp5_ASAP7_75t_SL U71239 ( .A(n65181), .B(n68766), .Y(n65185) );
  OR2x2_ASAP7_75t_SL U71240 ( .A(or1200_cpu_or1200_mult_mac_n337), .B(
        or1200_cpu_or1200_mult_mac_n191), .Y(n68778) );
  O2A1O1Ixp5_ASAP7_75t_SL U71241 ( .A1(n65180), .A2(n65179), .B(n65178), .C(
        n65177), .Y(n68782) );
  XOR2xp5_ASAP7_75t_SL U71242 ( .A(n65181), .B(n68768), .Y(n65183) );
  OAI211xp5_ASAP7_75t_SL U71243 ( .A1(or1200_cpu_or1200_except_n374), .A2(
        n57088), .B(n65190), .C(n65189), .Y(or1200_cpu_or1200_except_n1758) );
  OAI211xp5_ASAP7_75t_SL U71244 ( .A1(or1200_cpu_or1200_except_n368), .A2(
        n57088), .B(n65200), .C(n65199), .Y(or1200_cpu_or1200_except_n1760) );
  OAI211xp5_ASAP7_75t_SL U71245 ( .A1(or1200_cpu_or1200_except_n371), .A2(
        n57088), .B(n65217), .C(n65216), .Y(or1200_cpu_or1200_except_n1759) );
  AND2x2_ASAP7_75t_SL U71246 ( .A(n59701), .B(icqmem_adr_qmem[25]), .Y(n51952)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71247 ( .A1(n65231), .A2(n65230), .B(n65229), .C(
        n65228), .Y(n75156) );
  NAND3xp33_ASAP7_75t_SL U71248 ( .A(n69435), .B(n69385), .C(n78365), .Y(
        n65236) );
  OR2x2_ASAP7_75t_SL U71249 ( .A(n2900), .B(n65398), .Y(n2474) );
  OR2x2_ASAP7_75t_SL U71250 ( .A(n1564), .B(n65398), .Y(n1559) );
  OR2x2_ASAP7_75t_SL U71251 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_3_), .B(n65332), .Y(
        n65394) );
  OR2x2_ASAP7_75t_SL U71252 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .B(n65398), .Y(
        n65393) );
  OR2x2_ASAP7_75t_SL U71253 ( .A(n65400), .B(n65401), .Y(n65395) );
  A2O1A1Ixp33_ASAP7_75t_SL U71254 ( .A1(n65385), .A2(n65393), .B(n65311), .C(
        n65241), .Y(n65242) );
  NAND3xp33_ASAP7_75t_SL U71255 ( .A(n65243), .B(n65395), .C(n65242), .Y(n1793) );
  AO21x1_ASAP7_75t_SL U71256 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_12_), .A2(n65246), .B(
        n65248), .Y(n65306) );
  AO21x1_ASAP7_75t_SL U71257 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_14_), .A2(n65250), .B(
        n65255), .Y(n65304) );
  A2O1A1Ixp33_ASAP7_75t_SL U71258 ( .A1(n65298), .A2(n65393), .B(n65301), .C(
        n65253), .Y(n65254) );
  NAND3xp33_ASAP7_75t_SL U71259 ( .A(n65374), .B(n65395), .C(n65254), .Y(n1680) );
  AND2x2_ASAP7_75t_SL U71260 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r1), .B(n65398), .Y(
        n65346) );
  A2O1A1Ixp33_ASAP7_75t_SL U71261 ( .A1(n2860), .A2(n65354), .B(n65275), .C(
        n65308), .Y(n65266) );
  OR2x2_ASAP7_75t_SL U71262 ( .A(n65398), .B(n65262), .Y(n65314) );
  NAND3xp33_ASAP7_75t_SL U71263 ( .A(n65313), .B(n65264), .C(n65263), .Y(
        n65265) );
  NAND3xp33_ASAP7_75t_SL U71264 ( .A(n65266), .B(n65314), .C(n65265), .Y(n2483) );
  NAND3xp33_ASAP7_75t_SL U71265 ( .A(n65313), .B(n65268), .C(n65267), .Y(
        n65269) );
  A2O1A1Ixp33_ASAP7_75t_SL U71266 ( .A1(n65272), .A2(n65274), .B(n65354), .C(
        n65322), .Y(n65273) );
  OR2x2_ASAP7_75t_SL U71267 ( .A(n65398), .B(n65331), .Y(n65330) );
  A2O1A1Ixp33_ASAP7_75t_SL U71268 ( .A1(n65277), .A2(n2900), .B(n65276), .C(
        n65330), .Y(n2481) );
  A2O1A1Ixp33_ASAP7_75t_SL U71269 ( .A1(n1582), .A2(n65279), .B(n1564), .C(
        n65278), .Y(n65280) );
  A2O1A1Ixp33_ASAP7_75t_SL U71270 ( .A1(n1564), .A2(n65308), .B(n65313), .C(
        n65280), .Y(n65281) );
  O2A1O1Ixp5_ASAP7_75t_SL U71271 ( .A1(n1600), .A2(n58551), .B(n65283), .C(
        n65282), .Y(n1599) );
  AND2x2_ASAP7_75t_SL U71272 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_qnan_r_a), .B(n65363), .Y(
        n65345) );
  OR2x2_ASAP7_75t_SL U71273 ( .A(n65354), .B(n65318), .Y(n65287) );
  NOR3xp33_ASAP7_75t_SL U71274 ( .A(n65318), .B(n2009), .C(n78435), .Y(n65286)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71275 ( .A1(n65371), .A2(n65300), .B(n65290), .C(
        n65314), .Y(n1663) );
  AND2x2_ASAP7_75t_SL U71276 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_18_), .B(n65375), .Y(
        n65364) );
  A2O1A1Ixp33_ASAP7_75t_SL U71277 ( .A1(n65361), .A2(n65296), .B(n65294), .C(
        n65314), .Y(n2485) );
  A2O1A1Ixp33_ASAP7_75t_SL U71278 ( .A1(n65297), .A2(n65296), .B(n65295), .C(
        n65314), .Y(n1617) );
  A2O1A1Ixp33_ASAP7_75t_SL U71279 ( .A1(n65301), .A2(n65300), .B(n65299), .C(
        n65314), .Y(n1679) );
  A2O1A1Ixp33_ASAP7_75t_SL U71280 ( .A1(n65311), .A2(n65316), .B(n65310), .C(
        n65314), .Y(n1792) );
  A2O1A1Ixp33_ASAP7_75t_SL U71281 ( .A1(n65383), .A2(n65316), .B(n65315), .C(
        n65314), .Y(n1809) );
  NAND3xp33_ASAP7_75t_SL U71282 ( .A(n74463), .B(n65320), .C(n65400), .Y(
        n65319) );
  A2O1A1Ixp33_ASAP7_75t_SL U71283 ( .A1(n74463), .A2(n65393), .B(n65320), .C(
        n65319), .Y(n65324) );
  AO21x1_ASAP7_75t_SL U71284 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r1_6_), .A2(n65347), .B(
        n65326), .Y(n65389) );
  A2O1A1Ixp33_ASAP7_75t_SL U71285 ( .A1(n65400), .A2(n65336), .B(n65335), .C(
        n65334), .Y(n1618) );
  A2O1A1Ixp33_ASAP7_75t_SL U71286 ( .A1(n65342), .A2(n65360), .B(n65341), .C(
        n65340), .Y(n65343) );
  A2O1A1Ixp33_ASAP7_75t_SL U71287 ( .A1(n65352), .A2(n65400), .B(n65351), .C(
        n74463), .Y(n1838) );
  A2O1A1Ixp33_ASAP7_75t_SL U71288 ( .A1(n65361), .A2(n65360), .B(n65359), .C(
        n65358), .Y(n65362) );
  A2O1A1Ixp33_ASAP7_75t_SL U71289 ( .A1(n65370), .A2(n65400), .B(n65369), .C(
        n65368), .Y(n1648) );
  OR2x2_ASAP7_75t_SL U71290 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[22]), .Y(n65468) );
  OR2x2_ASAP7_75t_SL U71291 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[17]), .B(n66196), 
        .Y(n65408) );
  OR2x2_ASAP7_75t_SL U71292 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[25]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[26]), .Y(n65452) );
  NAND3xp33_ASAP7_75t_SL U71293 ( .A(n65658), .B(n65454), .C(n65684), .Y(
        n65380) );
  NAND3xp33_ASAP7_75t_SL U71294 ( .A(n65377), .B(n65421), .C(n65457), .Y(
        n65545) );
  OR2x2_ASAP7_75t_SL U71295 ( .A(n65408), .B(n65466), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n63) );
  A2O1A1Ixp33_ASAP7_75t_SL U71296 ( .A1(n65384), .A2(n65393), .B(n65383), .C(
        n65382), .Y(n65386) );
  NAND3xp33_ASAP7_75t_SL U71297 ( .A(n65386), .B(n65385), .C(n65395), .Y(n1810) );
  OR2x2_ASAP7_75t_SL U71298 ( .A(n65398), .B(n65397), .Y(n2013) );
  OR2x2_ASAP7_75t_SL U71299 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[11]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[12]), .Y(n65446) );
  OR2x2_ASAP7_75t_SL U71300 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[7]), .B(n65431), .Y(
        n65478) );
  NAND3xp33_ASAP7_75t_SL U71301 ( .A(n65662), .B(n65405), .C(n65788), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n57) );
  A2O1A1Ixp33_ASAP7_75t_SL U71302 ( .A1(n65856), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[41]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[43]), .C(n65855), 
        .Y(n65407) );
  NAND3xp33_ASAP7_75t_SL U71303 ( .A(n65476), .B(n65537), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[9]), .Y(n65410) );
  NAND4xp25_ASAP7_75t_SL U71304 ( .A(n65544), .B(n65743), .C(n65745), .D(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[34]), .Y(n65414) );
  AO21x1_ASAP7_75t_SL U71305 ( .A1(n65417), .A2(n65416), .B(n65415), .Y(n65561) );
  OAI211xp5_ASAP7_75t_SL U71306 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[18]), .A2(n65425), 
        .B(n65434), .C(n65424), .Y(n65426) );
  OAI211xp5_ASAP7_75t_SL U71307 ( .A1(n65537), .A2(n65539), .B(n65427), .C(
        n65426), .Y(n65428) );
  A2O1A1Ixp33_ASAP7_75t_SL U71308 ( .A1(n65643), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[13]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[15]), .C(n65783), 
        .Y(n65440) );
  A2O1A1Ixp33_ASAP7_75t_SL U71309 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[19]), .A2(n65635), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[21]), .C(n65434), 
        .Y(n65439) );
  OAI211xp5_ASAP7_75t_SL U71310 ( .A1(n65440), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n63), .B(n65439), .C(n65438), .Y(n65441) );
  OAI211xp5_ASAP7_75t_SL U71311 ( .A1(n65785), .A2(n65443), .B(n65558), .C(
        n65442), .Y(n65444) );
  NOR3xp33_ASAP7_75t_SL U71312 ( .A(n65465), .B(n65464), .C(n65463), .Y(n65471) );
  OAI211xp5_ASAP7_75t_SL U71313 ( .A1(n65472), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n63), .B(n65471), .C(n65470), .Y(n65474) );
  OR2x2_ASAP7_75t_SL U71314 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[3]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .Y(n74133) );
  OR2x2_ASAP7_75t_SL U71315 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[0]), .Y(n74834) );
  AND2x2_ASAP7_75t_SL U71316 ( .A(n65651), .B(n66092), .Y(n66167) );
  OAI211xp5_ASAP7_75t_SL U71317 ( .A1(n65588), .A2(n65670), .B(n65503), .C(
        n65502), .Y(n66107) );
  OR2x2_ASAP7_75t_SL U71318 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[3]), .B(n65674), .Y(
        n65625) );
  AND2x2_ASAP7_75t_SL U71319 ( .A(n65663), .B(n66126), .Y(n65570) );
  OR2x2_ASAP7_75t_SL U71320 ( .A(n65625), .B(n66150), .Y(n66147) );
  OR2x2_ASAP7_75t_SL U71321 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_in_00), .B(n76976), 
        .Y(n66138) );
  NOR3xp33_ASAP7_75t_SL U71322 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[5]), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[6]), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[7]), .Y(n65527) );
  NAND3xp33_ASAP7_75t_SL U71323 ( .A(n65529), .B(n65528), .C(n65527), .Y(
        n74132) );
  O2A1O1Ixp5_ASAP7_75t_SL U71324 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2), .A2(n65533), .B(
        n65532), .C(n65531), .Y(n74752) );
  AND2x2_ASAP7_75t_SL U71325 ( .A(n76977), .B(n74752), .Y(n66111) );
  NOR3xp33_ASAP7_75t_SL U71326 ( .A(n65556), .B(n65555), .C(n65554), .Y(n65557) );
  NAND3xp33_ASAP7_75t_SL U71327 ( .A(n65559), .B(n65558), .C(n65557), .Y(
        n65560) );
  OAI211xp5_ASAP7_75t_SL U71328 ( .A1(n65857), .A2(n65646), .B(n65562), .C(
        n66181), .Y(n66093) );
  OAI211xp5_ASAP7_75t_SL U71329 ( .A1(n65620), .A2(n65670), .B(n65574), .C(
        n65573), .Y(n66100) );
  OAI211xp5_ASAP7_75t_SL U71330 ( .A1(n66145), .A2(n66124), .B(n65584), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_exp_r[4]), .Y(n65585) );
  AND2x2_ASAP7_75t_SL U71331 ( .A(n65588), .B(n65670), .Y(n66125) );
  NAND3xp33_ASAP7_75t_SL U71332 ( .A(n65624), .B(n65623), .C(n65622), .Y(
        n66157) );
  A2O1A1Ixp33_ASAP7_75t_SL U71333 ( .A1(n66178), .A2(n66180), .B(n66138), .C(
        n66137), .Y(n65655) );
  A2O1A1Ixp33_ASAP7_75t_SL U71334 ( .A1(n57187), .A2(n65684), .B(n65683), .C(
        n65682), .Y(n65685) );
  OR2x2_ASAP7_75t_SL U71335 ( .A(n65689), .B(n65688), .Y(n65984) );
  OAI211xp5_ASAP7_75t_SL U71336 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[35]), .A2(n65808), 
        .B(n65841), .C(n65849), .Y(n65714) );
  NAND3xp33_ASAP7_75t_SL U71337 ( .A(n65714), .B(n65713), .C(n65712), .Y(
        n65887) );
  NAND3xp33_ASAP7_75t_SL U71338 ( .A(n65717), .B(n65716), .C(n65715), .Y(
        n65886) );
  NOR3xp33_ASAP7_75t_SL U71339 ( .A(n65721), .B(n65720), .C(n65719), .Y(n65722) );
  A2O1A1Ixp33_ASAP7_75t_SL U71340 ( .A1(n65983), .A2(n65984), .B(n66065), .C(
        n65724), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n31) );
  OR2x2_ASAP7_75t_SL U71341 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[14]), .B(n65808), 
        .Y(n65782) );
  OAI31xp33_ASAP7_75t_SL U71342 ( .A1(n65727), .A2(n65819), .A3(n57187), .B(
        n65726), .Y(n65728) );
  NAND3xp33_ASAP7_75t_SL U71343 ( .A(n65732), .B(n65731), .C(n65730), .Y(
        n66023) );
  NAND3xp33_ASAP7_75t_SL U71344 ( .A(n65736), .B(n65735), .C(n65734), .Y(
        n66021) );
  OAI211xp5_ASAP7_75t_SL U71345 ( .A1(n65974), .A2(n66026), .B(n65738), .C(
        n65737), .Y(n66062) );
  NAND3xp33_ASAP7_75t_SL U71346 ( .A(n65741), .B(n65740), .C(n65739), .Y(
        n65878) );
  O2A1O1Ixp5_ASAP7_75t_SL U71347 ( .A1(n65752), .A2(n65751), .B(n66014), .C(
        n65750), .Y(n65768) );
  NAND4xp25_ASAP7_75t_SL U71348 ( .A(n65770), .B(n65769), .C(n65768), .D(
        n65767), .Y(n65771) );
  NAND3xp33_ASAP7_75t_SL U71349 ( .A(n65774), .B(n65773), .C(n65772), .Y(
        n65958) );
  OAI211xp5_ASAP7_75t_SL U71350 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[28]), .A2(n65808), 
        .B(n65777), .C(n65841), .Y(n65778) );
  NAND3xp33_ASAP7_75t_SL U71351 ( .A(n65780), .B(n65779), .C(n65778), .Y(
        n65959) );
  OAI211xp5_ASAP7_75t_SL U71352 ( .A1(n66065), .A2(n65988), .B(n65981), .C(
        n65812), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n28) );
  OAI31xp33_ASAP7_75t_SL U71353 ( .A1(n65819), .A2(n57188), .A3(n65818), .B(
        n65817), .Y(n65820) );
  NAND3xp33_ASAP7_75t_SL U71354 ( .A(n65836), .B(n65835), .C(n65834), .Y(
        n65999) );
  NAND3xp33_ASAP7_75t_SL U71355 ( .A(n65839), .B(n65838), .C(n65837), .Y(
        n66008) );
  NAND3xp33_ASAP7_75t_SL U71356 ( .A(n65844), .B(n65843), .C(n65842), .Y(
        n65942) );
  OAI211xp5_ASAP7_75t_SL U71357 ( .A1(n65999), .A2(n65974), .B(n65846), .C(
        n65845), .Y(n65985) );
  NAND3xp33_ASAP7_75t_SL U71358 ( .A(n58419), .B(n65850), .C(n65849), .Y(
        n65852) );
  O2A1O1Ixp5_ASAP7_75t_SL U71359 ( .A1(n58419), .A2(n65853), .B(n65852), .C(
        n65851), .Y(n65945) );
  O2A1O1Ixp5_ASAP7_75t_SL U71360 ( .A1(n65862), .A2(n65861), .B(n66051), .C(
        n65860), .Y(n65863) );
  AND2x2_ASAP7_75t_SL U71361 ( .A(n65866), .B(n65865), .Y(n65872) );
  OAI211xp5_ASAP7_75t_SL U71362 ( .A1(n65972), .A2(n66011), .B(n65871), .C(
        n65870), .Y(n65992) );
  OAI211xp5_ASAP7_75t_SL U71363 ( .A1(n65992), .A2(n66065), .B(n65876), .C(
        n65981), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n25) );
  NAND4xp25_ASAP7_75t_SL U71364 ( .A(n65885), .B(n65981), .C(n65884), .D(
        n65883), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n26) );
  NAND3xp33_ASAP7_75t_SL U71365 ( .A(n65981), .B(n65893), .C(n65892), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n27) );
  NAND3xp33_ASAP7_75t_SL U71366 ( .A(n65981), .B(n65906), .C(n65905), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n24) );
  OAI211xp5_ASAP7_75t_SL U71367 ( .A1(n65970), .A2(n66026), .B(n65908), .C(
        n65907), .Y(n66038) );
  NAND4xp25_ASAP7_75t_SL U71368 ( .A(n65913), .B(n65912), .C(n65911), .D(
        n65910), .Y(n65914) );
  A2O1A1Ixp33_ASAP7_75t_SL U71369 ( .A1(n65950), .A2(n65927), .B(n65983), .C(
        n65926), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n23) );
  OAI211xp5_ASAP7_75t_SL U71370 ( .A1(n65937), .A2(n66001), .B(n65936), .C(
        n65935), .Y(n65938) );
  OAI211xp5_ASAP7_75t_SL U71371 ( .A1(n65970), .A2(n66011), .B(n65941), .C(
        n65940), .Y(n66041) );
  A2O1A1Ixp33_ASAP7_75t_SL U71372 ( .A1(n65950), .A2(n65949), .B(n65983), .C(
        n65948), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n21) );
  OAI211xp5_ASAP7_75t_SL U71373 ( .A1(n65962), .A2(n66001), .B(n65961), .C(
        n65960), .Y(n65963) );
  OAI211xp5_ASAP7_75t_SL U71374 ( .A1(n66045), .A2(n65983), .B(n65982), .C(
        n65981), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n19) );
  OR3x1_ASAP7_75t_SL U71375 ( .A(n66005), .B(n66004), .C(n66003), .Y(n66012)
         );
  OAI211xp5_ASAP7_75t_SL U71376 ( .A1(n66011), .A2(n66027), .B(n66010), .C(
        n66009), .Y(n66056) );
  A2O1A1Ixp33_ASAP7_75t_SL U71377 ( .A1(n66051), .A2(n66047), .B(n66046), .C(
        n66028), .Y(n66032) );
  NAND4xp25_ASAP7_75t_SL U71378 ( .A(n66034), .B(n66033), .C(n66032), .D(
        n66031), .Y(n66035) );
  A2O1A1Ixp33_ASAP7_75t_SL U71379 ( .A1(n66060), .A2(n66056), .B(n66055), .C(
        n66057), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n49) );
  A2O1A1Ixp33_ASAP7_75t_SL U71380 ( .A1(n66060), .A2(n66059), .B(n66058), .C(
        n66057), .Y(or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n48) );
  NAND3xp33_ASAP7_75t_SL U71381 ( .A(n66065), .B(n66064), .C(n66063), .Y(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_n45) );
  NOR3xp33_ASAP7_75t_SL U71382 ( .A(n66131), .B(n66130), .C(n66129), .Y(n66143) );
  OAI31xp33_ASAP7_75t_SL U71383 ( .A1(n66134), .A2(n66155), .A3(n66133), .B(
        n66145), .Y(n66142) );
  NAND3xp33_ASAP7_75t_SL U71384 ( .A(n66136), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_4_), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fi_ldz_3_), .Y(n66139) );
  A2O1A1Ixp33_ASAP7_75t_SL U71385 ( .A1(n66140), .A2(n66139), .B(n66138), .C(
        n66137), .Y(n66141) );
  OR3x1_ASAP7_75t_SL U71386 ( .A(n66177), .B(n66176), .C(n66175), .Y(n66208)
         );
  NAND3xp33_ASAP7_75t_SL U71387 ( .A(n74152), .B(n66168), .C(n66208), .Y(
        n74055) );
  MAJIxp5_ASAP7_75t_SL U71388 ( .A(n74090), .B(n66187), .C(n74089), .Y(n66188)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71389 ( .A1(n66200), .A2(n66199), .B(n66198), .C(
        n74745), .Y(n66202) );
  NOR3xp33_ASAP7_75t_SL U71390 ( .A(n74745), .B(n76976), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_sign), .Y(n66201) );
  OR2x2_ASAP7_75t_SL U71391 ( .A(n66206), .B(n74087), .Y(n74189) );
  O2A1O1Ixp5_ASAP7_75t_SL U71392 ( .A1(n66212), .A2(n74161), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[0]), .C(n74056), .Y(
        n66215) );
  O2A1O1Ixp5_ASAP7_75t_SL U71393 ( .A1(n74058), .A2(n66215), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_3_), .C(n66214), 
        .Y(n66222) );
  A2O1A1Ixp33_ASAP7_75t_SL U71394 ( .A1(n74088), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_2_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_3_), .C(n74187), 
        .Y(n66221) );
  A2O1A1Ixp33_ASAP7_75t_SL U71395 ( .A1(n75030), .A2(n66227), .B(n66226), .C(
        n66231), .Y(n66228) );
  A2O1A1Ixp33_ASAP7_75t_SL U71396 ( .A1(n1133), .A2(n66231), .B(n66230), .C(
        n66229), .Y(n9251) );
  OAI211xp5_ASAP7_75t_SL U71397 ( .A1(n66233), .A2(n66232), .B(n66238), .C(
        n75030), .Y(n66234) );
  A2O1A1Ixp33_ASAP7_75t_SL U71398 ( .A1(n66238), .A2(n66237), .B(n75027), .C(
        n66236), .Y(n9249) );
  A2O1A1Ixp33_ASAP7_75t_SL U71399 ( .A1(n57163), .A2(n76176), .B(n66246), .C(
        n66245), .Y(n66247) );
  XNOR2xp5_ASAP7_75t_SL U71400 ( .A(n59640), .B(n67736), .Y(n66344) );
  XNOR2xp5_ASAP7_75t_SL U71401 ( .A(n57322), .B(n53221), .Y(n66289) );
  XNOR2xp5_ASAP7_75t_SL U71402 ( .A(n57322), .B(n59664), .Y(n66561) );
  XNOR2xp5_ASAP7_75t_SL U71403 ( .A(n66557), .B(n66558), .Y(n66290) );
  NAND3xp33_ASAP7_75t_SL U71404 ( .A(n66302), .B(n66303), .C(n66305), .Y(
        n66315) );
  A2O1A1Ixp33_ASAP7_75t_SL U71405 ( .A1(n66310), .A2(n66311), .B(n66309), .C(
        n66308), .Y(n66314) );
  A2O1A1Ixp33_ASAP7_75t_SL U71406 ( .A1(n57104), .A2(n75045), .B(n66318), .C(
        n66317), .Y(n66392) );
  A2O1A1Ixp33_ASAP7_75t_SL U71407 ( .A1(n66321), .A2(n66390), .B(n66392), .C(
        n66320), .Y(n66596) );
  A2O1A1Ixp33_ASAP7_75t_SL U71408 ( .A1(n66417), .A2(n59649), .B(n66324), .C(
        n66323), .Y(n66341) );
  AO21x1_ASAP7_75t_SL U71409 ( .A1(n57099), .A2(n67743), .B(n66334), .Y(n66330) );
  NAND3xp33_ASAP7_75t_SL U71410 ( .A(n67446), .B(n66326), .C(n58534), .Y(
        n66327) );
  XNOR2xp5_ASAP7_75t_SL U71411 ( .A(n66336), .B(n66335), .Y(n66337) );
  NAND3xp33_ASAP7_75t_SL U71412 ( .A(n66554), .B(n66342), .C(n66596), .Y(
        n66343) );
  O2A1O1Ixp5_ASAP7_75t_SL U71413 ( .A1(n66360), .A2(n66359), .B(n67715), .C(
        n66358), .Y(n66410) );
  A2O1A1Ixp33_ASAP7_75t_SL U71414 ( .A1(n66370), .A2(n66369), .B(n66368), .C(
        n66367), .Y(n66371) );
  NAND3xp33_ASAP7_75t_SL U71415 ( .A(n66376), .B(n59641), .C(n66375), .Y(
        n66377) );
  XNOR2xp5_ASAP7_75t_SL U71416 ( .A(n75644), .B(n57325), .Y(n66379) );
  A2O1A1Ixp33_ASAP7_75t_SL U71417 ( .A1(n68104), .A2(n57322), .B(n66380), .C(
        n67715), .Y(n66381) );
  O2A1O1Ixp5_ASAP7_75t_SL U71418 ( .A1(n75899), .A2(n66384), .B(n57078), .C(
        n66383), .Y(n66386) );
  XNOR2xp5_ASAP7_75t_SL U71419 ( .A(n66390), .B(n66557), .Y(n66391) );
  MAJIxp5_ASAP7_75t_SL U71420 ( .A(n66439), .B(n66438), .C(n66393), .Y(n68622)
         );
  XNOR2xp5_ASAP7_75t_SL U71421 ( .A(n59670), .B(n57505), .Y(n66397) );
  A2O1A1Ixp33_ASAP7_75t_SL U71422 ( .A1(n57409), .A2(n75947), .B(n66402), .C(
        n66401), .Y(n66494) );
  NOR3xp33_ASAP7_75t_SL U71423 ( .A(n67284), .B(n57260), .C(n66466), .Y(n66403) );
  O2A1O1Ixp5_ASAP7_75t_SL U71424 ( .A1(n57405), .A2(n66806), .B(n66404), .C(
        n66403), .Y(n66496) );
  MAJIxp5_ASAP7_75t_SL U71425 ( .A(n66493), .B(n66406), .C(n66405), .Y(n66426)
         );
  XNOR2xp5_ASAP7_75t_SL U71426 ( .A(n66408), .B(n66407), .Y(n66409) );
  XNOR2xp5_ASAP7_75t_SL U71427 ( .A(n66410), .B(n66409), .Y(n66427) );
  A2O1A1Ixp33_ASAP7_75t_SL U71428 ( .A1(n66417), .A2(n67911), .B(n66416), .C(
        n66415), .Y(n66488) );
  XNOR2xp5_ASAP7_75t_SL U71429 ( .A(n66434), .B(n66433), .Y(n66435) );
  OR2x2_ASAP7_75t_SL U71430 ( .A(n66444), .B(n66533), .Y(n69227) );
  A2O1A1Ixp33_ASAP7_75t_SL U71431 ( .A1(n66451), .A2(n57271), .B(n58433), .C(
        n74799), .Y(n66453) );
  XNOR2xp5_ASAP7_75t_SL U71432 ( .A(n59653), .B(n59637), .Y(n66471) );
  O2A1O1Ixp5_ASAP7_75t_SL U71433 ( .A1(n66459), .A2(n66458), .B(n75048), .C(
        n66457), .Y(n66490) );
  XNOR2xp5_ASAP7_75t_SL U71434 ( .A(n66491), .B(n66490), .Y(n66460) );
  MAJIxp5_ASAP7_75t_SL U71435 ( .A(n67142), .B(n67141), .C(n67140), .Y(n67166)
         );
  XNOR2xp5_ASAP7_75t_SL U71436 ( .A(n59666), .B(n66333), .Y(n66472) );
  XNOR2xp5_ASAP7_75t_SL U71437 ( .A(n66478), .B(n66468), .Y(n67165) );
  MAJIxp5_ASAP7_75t_SL U71438 ( .A(n67130), .B(n67126), .C(n67127), .Y(n67160)
         );
  XNOR2xp5_ASAP7_75t_SL U71439 ( .A(n59598), .B(n59662), .Y(n67095) );
  XNOR2xp5_ASAP7_75t_SL U71440 ( .A(n59607), .B(n59650), .Y(n66474) );
  MAJIxp5_ASAP7_75t_SL U71441 ( .A(n67121), .B(n67123), .C(n67122), .Y(n67158)
         );
  MAJIxp5_ASAP7_75t_SL U71442 ( .A(n67159), .B(n67158), .C(n67160), .Y(n67119)
         );
  MAJIxp5_ASAP7_75t_SL U71443 ( .A(n66478), .B(n66477), .C(n66476), .Y(n66504)
         );
  MAJIxp5_ASAP7_75t_SL U71444 ( .A(n67120), .B(n67119), .C(n67118), .Y(n67113)
         );
  XNOR2xp5_ASAP7_75t_SL U71445 ( .A(n66489), .B(n66488), .Y(n67117) );
  MAJIxp5_ASAP7_75t_SL U71446 ( .A(n66492), .B(n66491), .C(n66490), .Y(n67115)
         );
  XNOR2xp5_ASAP7_75t_SL U71447 ( .A(n66494), .B(n66493), .Y(n66495) );
  MAJIxp5_ASAP7_75t_SL U71448 ( .A(n67117), .B(n67115), .C(n67114), .Y(n66513)
         );
  OAI31xp33_ASAP7_75t_SL U71449 ( .A1(n57179), .A2(n59664), .A3(n67743), .B(
        n66499), .Y(n66502) );
  NOR3xp33_ASAP7_75t_SL U71450 ( .A(n66502), .B(n66501), .C(n66500), .Y(n66503) );
  XNOR2xp5_ASAP7_75t_SL U71451 ( .A(n66516), .B(n66514), .Y(n66508) );
  MAJIxp5_ASAP7_75t_SL U71452 ( .A(n67112), .B(n66510), .C(n66509), .Y(n68626)
         );
  MAJIxp5_ASAP7_75t_SL U71453 ( .A(n66517), .B(n66516), .C(n66515), .Y(n66526)
         );
  XNOR2xp5_ASAP7_75t_SL U71454 ( .A(n66527), .B(n66526), .Y(n66522) );
  XNOR2xp5_ASAP7_75t_SL U71455 ( .A(n66525), .B(n66522), .Y(n68625) );
  MAJIxp5_ASAP7_75t_SL U71456 ( .A(n66528), .B(n66527), .C(n66526), .Y(n68624)
         );
  XNOR2xp5_ASAP7_75t_SL U71457 ( .A(n66536), .B(n66566), .Y(n66544) );
  A2O1A1Ixp33_ASAP7_75t_SL U71458 ( .A1(n75899), .A2(n75046), .B(n66547), .C(
        n66552), .Y(n66548) );
  O2A1O1Ixp5_ASAP7_75t_SL U71459 ( .A1(n53310), .A2(n58785), .B(n66552), .C(
        n66551), .Y(n66575) );
  MAJIxp5_ASAP7_75t_SL U71460 ( .A(n66589), .B(n66563), .C(n66562), .Y(n68635)
         );
  XNOR2xp5_ASAP7_75t_SL U71461 ( .A(n59642), .B(n57398), .Y(n68606) );
  XNOR2xp5_ASAP7_75t_SL U71462 ( .A(n66586), .B(n66585), .Y(n66587) );
  NAND3xp33_ASAP7_75t_SL U71463 ( .A(n68651), .B(n75059), .C(n68666), .Y(
        n75110) );
  O2A1O1Ixp5_ASAP7_75t_SL U71464 ( .A1(n66728), .A2(n66622), .B(n67715), .C(
        n66621), .Y(n66649) );
  XNOR2xp5_ASAP7_75t_SL U71465 ( .A(n59640), .B(n67432), .Y(n66683) );
  XNOR2xp5_ASAP7_75t_SL U71466 ( .A(n57322), .B(n76078), .Y(n66740) );
  XNOR2xp5_ASAP7_75t_SL U71467 ( .A(n59617), .B(n59650), .Y(n68382) );
  XNOR2xp5_ASAP7_75t_SL U71468 ( .A(n59609), .B(n59668), .Y(n66712) );
  NAND3xp33_ASAP7_75t_SL U71469 ( .A(n66973), .B(n66641), .C(n53496), .Y(
        n66645) );
  NAND3xp33_ASAP7_75t_SL U71470 ( .A(n66645), .B(n66644), .C(n66643), .Y(
        n66777) );
  XNOR2xp5_ASAP7_75t_SL U71471 ( .A(n66647), .B(n66646), .Y(n66648) );
  XNOR2xp5_ASAP7_75t_SL U71472 ( .A(n58402), .B(n59666), .Y(n66682) );
  XNOR2xp5_ASAP7_75t_SL U71473 ( .A(n66655), .B(n66654), .Y(n66652) );
  XNOR2xp5_ASAP7_75t_SL U71474 ( .A(n59598), .B(n67736), .Y(n66827) );
  O2A1O1Ixp5_ASAP7_75t_SL U71475 ( .A1(n66660), .A2(n66659), .B(n66661), .C(
        n66662), .Y(n66663) );
  O2A1O1Ixp5_ASAP7_75t_SL U71476 ( .A1(n66670), .A2(n66669), .B(n67829), .C(
        n66668), .Y(n66738) );
  MAJIxp5_ASAP7_75t_SL U71477 ( .A(n66673), .B(n58467), .C(n66977), .Y(n66842)
         );
  XNOR2xp5_ASAP7_75t_SL U71478 ( .A(n59660), .B(n59640), .Y(n66684) );
  O2A1O1Ixp5_ASAP7_75t_SL U71479 ( .A1(n66729), .A2(n66681), .B(n67715), .C(
        n56995), .Y(n66772) );
  XNOR2xp5_ASAP7_75t_SL U71480 ( .A(n58402), .B(n59662), .Y(n67021) );
  MAJIxp5_ASAP7_75t_SL U71481 ( .A(n66686), .B(n66770), .C(n66685), .Y(n66891)
         );
  MAJIxp5_ASAP7_75t_SL U71482 ( .A(n66687), .B(n57151), .C(n66688), .Y(n66892)
         );
  XNOR2xp5_ASAP7_75t_SL U71483 ( .A(n66891), .B(n66892), .Y(n66689) );
  AO21x1_ASAP7_75t_SL U71484 ( .A1(n66851), .A2(n57067), .B(n66699), .Y(n66870) );
  A2O1A1Ixp33_ASAP7_75t_SL U71485 ( .A1(n53288), .A2(n59468), .B(n66714), .C(
        n57706), .Y(n66715) );
  XNOR2xp5_ASAP7_75t_SL U71486 ( .A(n57107), .B(n59600), .Y(n66750) );
  XNOR2xp5_ASAP7_75t_SL U71487 ( .A(n57516), .B(n67736), .Y(n66795) );
  MAJIxp5_ASAP7_75t_SL U71488 ( .A(n66937), .B(n57014), .C(n66732), .Y(n66912)
         );
  MAJIxp5_ASAP7_75t_SL U71489 ( .A(n66734), .B(n66733), .C(n66912), .Y(n66947)
         );
  MAJIxp5_ASAP7_75t_SL U71490 ( .A(n66947), .B(n66944), .C(n66946), .Y(n67042)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71491 ( .A1(n66745), .A2(n66744), .B(n67829), .C(
        n66743), .Y(n66965) );
  MAJIxp5_ASAP7_75t_SL U71492 ( .A(n66812), .B(n66811), .C(n53498), .Y(n66778)
         );
  XNOR2xp5_ASAP7_75t_SL U71493 ( .A(n57311), .B(n57505), .Y(n66753) );
  MAJIxp5_ASAP7_75t_SL U71494 ( .A(n66762), .B(n59071), .C(n66761), .Y(n66780)
         );
  XOR2xp5_ASAP7_75t_SL U71495 ( .A(n66819), .B(n66821), .Y(n66773) );
  XNOR2xp5_ASAP7_75t_SL U71496 ( .A(n59381), .B(n57491), .Y(n66788) );
  XNOR2xp5_ASAP7_75t_SL U71497 ( .A(n59607), .B(n57315), .Y(n66789) );
  NAND3xp33_ASAP7_75t_SL U71498 ( .A(n66806), .B(n58402), .C(n66802), .Y(
        n66804) );
  NAND3xp33_ASAP7_75t_SL U71499 ( .A(n66804), .B(n68104), .C(n66803), .Y(
        n66808) );
  XNOR2xp5_ASAP7_75t_SL U71500 ( .A(n59601), .B(n57325), .Y(n66856) );
  XNOR2xp5_ASAP7_75t_SL U71501 ( .A(n66849), .B(n66832), .Y(n66898) );
  MAJIxp5_ASAP7_75t_SL U71502 ( .A(n66842), .B(n66841), .C(n66840), .Y(n66984)
         );
  MAJIxp5_ASAP7_75t_SL U71503 ( .A(n66849), .B(n66848), .C(n66847), .Y(n67009)
         );
  XNOR2xp5_ASAP7_75t_SL U71504 ( .A(n57315), .B(n57436), .Y(n66850) );
  MAJIxp5_ASAP7_75t_SL U71505 ( .A(n66868), .B(n66869), .C(n66870), .Y(n67011)
         );
  MAJIxp5_ASAP7_75t_SL U71506 ( .A(n66871), .B(n66872), .C(n66873), .Y(n67014)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71507 ( .A1(n66879), .A2(n66878), .B(n67715), .C(
        n66877), .Y(n66889) );
  XNOR2xp5_ASAP7_75t_SL U71508 ( .A(n67023), .B(n67024), .Y(n66888) );
  A2O1A1Ixp33_ASAP7_75t_SL U71509 ( .A1(n66902), .A2(n66901), .B(n66900), .C(
        n66899), .Y(n66989) );
  XNOR2xp5_ASAP7_75t_SL U71510 ( .A(n66912), .B(n66911), .Y(n66914) );
  MAJIxp5_ASAP7_75t_SL U71511 ( .A(n68359), .B(n66932), .C(n57003), .Y(n68442)
         );
  XNOR2xp5_ASAP7_75t_SL U71512 ( .A(n59605), .B(n59666), .Y(n66964) );
  XNOR2xp5_ASAP7_75t_SL U71513 ( .A(n57257), .B(n59662), .Y(n67720) );
  XNOR2xp5_ASAP7_75t_SL U71514 ( .A(n66948), .B(n66947), .Y(n68543) );
  MAJIxp5_ASAP7_75t_SL U71515 ( .A(n68454), .B(n66958), .C(n68453), .Y(n68501)
         );
  XNOR2xp5_ASAP7_75t_SL U71516 ( .A(n66970), .B(n66969), .Y(n66975) );
  MAJIxp5_ASAP7_75t_SL U71517 ( .A(n68535), .B(n58503), .C(n66976), .Y(n68544)
         );
  MAJIxp5_ASAP7_75t_SL U71518 ( .A(n68552), .B(n66979), .C(n66978), .Y(n67211)
         );
  XNOR2xp5_ASAP7_75t_SL U71519 ( .A(n66983), .B(n66982), .Y(n66986) );
  MAJIxp5_ASAP7_75t_SL U71520 ( .A(n66984), .B(n66985), .C(n66986), .Y(n67110)
         );
  MAJIxp5_ASAP7_75t_SL U71521 ( .A(n66992), .B(n66991), .C(n66990), .Y(n67100)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71522 ( .A1(n66999), .A2(n66998), .B(n67715), .C(
        n66997), .Y(n67058) );
  XNOR2xp5_ASAP7_75t_SL U71523 ( .A(n57505), .B(n75947), .Y(n67000) );
  XOR2xp5_ASAP7_75t_SL U71524 ( .A(n59640), .B(n57101), .Y(n67002) );
  MAJIxp5_ASAP7_75t_SL U71525 ( .A(n67005), .B(n67006), .C(n67007), .Y(n67051)
         );
  XOR2xp5_ASAP7_75t_SL U71526 ( .A(n67050), .B(n67051), .Y(n67008) );
  MAJIxp5_ASAP7_75t_SL U71527 ( .A(n67015), .B(n67014), .C(n67013), .Y(n67045)
         );
  XNOR2xp5_ASAP7_75t_SL U71528 ( .A(n57310), .B(n59637), .Y(n67016) );
  XNOR2xp5_ASAP7_75t_SL U71529 ( .A(n67045), .B(n67046), .Y(n67037) );
  XNOR2xp5_ASAP7_75t_SL U71530 ( .A(n57491), .B(n57325), .Y(n67031) );
  A2O1A1Ixp33_ASAP7_75t_SL U71531 ( .A1(n67077), .A2(n57161), .B(n67035), .C(
        n67034), .Y(n67036) );
  MAJIxp5_ASAP7_75t_SL U71532 ( .A(n67050), .B(n67051), .C(n67052), .Y(n67198)
         );
  MAJIxp5_ASAP7_75t_SL U71533 ( .A(n67055), .B(n67054), .C(n67053), .Y(n67170)
         );
  MAJIxp5_ASAP7_75t_SL U71534 ( .A(n67058), .B(n57153), .C(n67057), .Y(n67171)
         );
  XNOR2xp5_ASAP7_75t_SL U71535 ( .A(n67170), .B(n67171), .Y(n67065) );
  XNOR2xp5_ASAP7_75t_SL U71536 ( .A(n67154), .B(n67138), .Y(n67064) );
  XNOR2xp5_ASAP7_75t_SL U71537 ( .A(n67197), .B(n67066), .Y(n67185) );
  MAJIxp5_ASAP7_75t_SL U71538 ( .A(n67070), .B(n67069), .C(n67068), .Y(n67189)
         );
  NAND3xp33_ASAP7_75t_SL U71539 ( .A(n66333), .B(n59651), .C(n67072), .Y(
        n67073) );
  XNOR2xp5_ASAP7_75t_SL U71540 ( .A(n67133), .B(n67132), .Y(n67091) );
  XNOR2xp5_ASAP7_75t_SL U71541 ( .A(n67123), .B(n67122), .Y(n67124) );
  XNOR2xp5_ASAP7_75t_SL U71542 ( .A(n58333), .B(n67129), .Y(n67136) );
  A2O1A1Ixp33_ASAP7_75t_SL U71543 ( .A1(n53310), .A2(n57242), .B(n67150), .C(
        n67149), .Y(n67153) );
  MAJIxp5_ASAP7_75t_SL U71544 ( .A(n67164), .B(n67161), .C(n57054), .Y(n67182)
         );
  MAJIxp5_ASAP7_75t_SL U71545 ( .A(n67173), .B(n67172), .C(n67171), .Y(n67179)
         );
  MAJIxp5_ASAP7_75t_SL U71546 ( .A(n67185), .B(n67184), .C(n67183), .Y(n67217)
         );
  NAND3xp33_ASAP7_75t_SL U71547 ( .A(n75276), .B(n74556), .C(n68693), .Y(
        n67220) );
  O2A1O1Ixp5_ASAP7_75t_SL U71548 ( .A1(n67238), .A2(n67237), .B(n67236), .C(
        n67235), .Y(n67292) );
  MAJIxp5_ASAP7_75t_SL U71549 ( .A(n67347), .B(n67294), .C(n67292), .Y(n67273)
         );
  NOR3xp33_ASAP7_75t_SL U71550 ( .A(n76176), .B(n59614), .C(n53237), .Y(n67255) );
  MAJIxp5_ASAP7_75t_SL U71551 ( .A(n67352), .B(n67353), .C(n67351), .Y(n67508)
         );
  XNOR2xp5_ASAP7_75t_SL U71552 ( .A(n59603), .B(n59647), .Y(n67363) );
  XNOR2xp5_ASAP7_75t_SL U71553 ( .A(n57257), .B(n59650), .Y(n67271) );
  A2O1A1Ixp33_ASAP7_75t_SL U71554 ( .A1(n75901), .A2(n57322), .B(n67557), .C(
        n67593), .Y(n67278) );
  XNOR2xp5_ASAP7_75t_SL U71555 ( .A(n67472), .B(n67470), .Y(n67285) );
  XNOR2xp5_ASAP7_75t_SL U71556 ( .A(n67292), .B(n67347), .Y(n67293) );
  O2A1O1Ixp5_ASAP7_75t_SL U71557 ( .A1(n67866), .A2(n59664), .B(n67318), .C(
        n67317), .Y(n67891) );
  A2O1A1Ixp33_ASAP7_75t_SL U71558 ( .A1(n75927), .A2(n67322), .B(n67321), .C(
        n67320), .Y(n67323) );
  XNOR2xp5_ASAP7_75t_SL U71559 ( .A(n57352), .B(n75895), .Y(n67361) );
  A2O1A1Ixp33_ASAP7_75t_SL U71560 ( .A1(n67376), .A2(n67375), .B(n67374), .C(
        n67373), .Y(n67377) );
  A2O1A1Ixp33_ASAP7_75t_SL U71561 ( .A1(n67614), .A2(n67613), .B(n67612), .C(
        n67377), .Y(n67649) );
  XOR2xp5_ASAP7_75t_SL U71562 ( .A(n59616), .B(n59658), .Y(n67382) );
  NAND3xp33_ASAP7_75t_SL U71563 ( .A(n67645), .B(n57436), .C(n57111), .Y(
        n67430) );
  NAND3xp33_ASAP7_75t_SL U71564 ( .A(n75468), .B(n59656), .C(n75894), .Y(
        n67429) );
  NAND3xp33_ASAP7_75t_SL U71565 ( .A(n67422), .B(n57486), .C(n67420), .Y(
        n67426) );
  NAND3xp33_ASAP7_75t_SL U71566 ( .A(n67424), .B(n57465), .C(n67423), .Y(
        n67425) );
  NAND3xp33_ASAP7_75t_SL U71567 ( .A(n67427), .B(n67426), .C(n67425), .Y(
        n67621) );
  XNOR2xp5_ASAP7_75t_SL U71568 ( .A(n59607), .B(n59620), .Y(n67455) );
  XNOR2xp5_ASAP7_75t_SL U71569 ( .A(n59616), .B(n53602), .Y(n67512) );
  MAJIxp5_ASAP7_75t_SL U71570 ( .A(n67500), .B(n67498), .C(n67499), .Y(n67679)
         );
  MAJIxp5_ASAP7_75t_SL U71571 ( .A(n67502), .B(n57001), .C(n67501), .Y(n67552)
         );
  MAJIxp5_ASAP7_75t_SL U71572 ( .A(n67504), .B(n67505), .C(n67506), .Y(n67553)
         );
  XNOR2xp5_ASAP7_75t_SL U71573 ( .A(n67552), .B(n67553), .Y(n67507) );
  MAJIxp5_ASAP7_75t_SL U71574 ( .A(n67508), .B(n67509), .C(n67510), .Y(n67574)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71575 ( .A1(n67963), .A2(n59648), .B(n67513), .C(
        n59619), .Y(n67514) );
  XNOR2xp5_ASAP7_75t_SL U71576 ( .A(n67691), .B(n67537), .Y(n67538) );
  XNOR2xp5_ASAP7_75t_SL U71577 ( .A(n67575), .B(n67574), .Y(n67576) );
  XOR2xp5_ASAP7_75t_SL U71578 ( .A(n59603), .B(n59658), .Y(n67581) );
  A2O1A1Ixp33_ASAP7_75t_SL U71579 ( .A1(n59599), .A2(n76049), .B(n67837), .C(
        n67589), .Y(n67592) );
  OAI31xp33_ASAP7_75t_SL U71580 ( .A1(n59503), .A2(n67598), .A3(n53310), .B(
        n67597), .Y(n67599) );
  NOR3xp33_ASAP7_75t_SL U71581 ( .A(n67605), .B(n67604), .C(n67607), .Y(n67606) );
  A2O1A1Ixp33_ASAP7_75t_SL U71582 ( .A1(n57104), .A2(n67632), .B(n67631), .C(
        n67630), .Y(n67633) );
  A2O1A1Ixp33_ASAP7_75t_SL U71583 ( .A1(n67645), .A2(n57436), .B(n59656), .C(
        n67644), .Y(n67647) );
  MAJIxp5_ASAP7_75t_SL U71584 ( .A(n67697), .B(n58365), .C(n67696), .Y(n68355)
         );
  NAND3xp33_ASAP7_75t_SL U71585 ( .A(n67725), .B(n67724), .C(n68419), .Y(
        n67726) );
  XNOR2xp5_ASAP7_75t_SL U71586 ( .A(n68372), .B(n68368), .Y(n67755) );
  XNOR2xp5_ASAP7_75t_SL U71587 ( .A(n67787), .B(n67786), .Y(n67788) );
  MAJIxp5_ASAP7_75t_SL U71588 ( .A(n68041), .B(n68040), .C(n68039), .Y(n68057)
         );
  XNOR2xp5_ASAP7_75t_SL U71589 ( .A(n67798), .B(n67797), .Y(n67799) );
  AO21x1_ASAP7_75t_SL U71590 ( .A1(n75900), .A2(n58536), .B(n67820), .Y(n68118) );
  XNOR2xp5_ASAP7_75t_SL U71591 ( .A(n59607), .B(n58431), .Y(n67822) );
  A2O1A1Ixp33_ASAP7_75t_SL U71592 ( .A1(n67879), .A2(n67878), .B(n57260), .C(
        n67877), .Y(n68112) );
  MAJIxp5_ASAP7_75t_SL U71593 ( .A(n58454), .B(n57613), .C(n67978), .Y(n67981)
         );
  OAI211xp5_ASAP7_75t_SL U71594 ( .A1(n67955), .A2(n57359), .B(n67950), .C(
        n67949), .Y(n67957) );
  XNOR2xp5_ASAP7_75t_SL U71595 ( .A(n67981), .B(n67980), .Y(n67982) );
  XNOR2xp5_ASAP7_75t_SL U71596 ( .A(n57110), .B(n58753), .Y(n68021) );
  MAJIxp5_ASAP7_75t_SL U71597 ( .A(n68064), .B(n68062), .C(n68060), .Y(n68144)
         );
  MAJIxp5_ASAP7_75t_SL U71598 ( .A(n68053), .B(n57305), .C(n57482), .Y(n68575)
         );
  MAJIxp5_ASAP7_75t_SL U71599 ( .A(n68198), .B(n68194), .C(n68195), .Y(n68191)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71600 ( .A1(n68123), .A2(n68122), .B(n68121), .C(
        n68120), .Y(n68127) );
  NAND3xp33_ASAP7_75t_SL U71601 ( .A(n68125), .B(n57078), .C(n68124), .Y(
        n68126) );
  MAJIxp5_ASAP7_75t_SL U71602 ( .A(n68155), .B(n68154), .C(n68153), .Y(n68289)
         );
  MAJIxp5_ASAP7_75t_SL U71603 ( .A(n68165), .B(n68163), .C(n68164), .Y(n68174)
         );
  MAJIxp5_ASAP7_75t_SL U71604 ( .A(n68170), .B(n68172), .C(n57231), .Y(n68285)
         );
  MAJIxp5_ASAP7_75t_SL U71605 ( .A(n68272), .B(n68273), .C(n68271), .Y(n68297)
         );
  NAND3xp33_ASAP7_75t_SL U71606 ( .A(n68252), .B(n68250), .C(n53489), .Y(
        n68253) );
  MAJIxp5_ASAP7_75t_SL U71607 ( .A(n68257), .B(n68256), .C(n68255), .Y(n68296)
         );
  MAJIxp5_ASAP7_75t_SL U71608 ( .A(n68293), .B(n58386), .C(n58379), .Y(n68350)
         );
  XOR2xp5_ASAP7_75t_SL U71609 ( .A(n68298), .B(n68297), .Y(n68299) );
  MAJIxp5_ASAP7_75t_SL U71610 ( .A(n68303), .B(n68302), .C(n68301), .Y(n68322)
         );
  MAJIxp5_ASAP7_75t_SL U71611 ( .A(n68314), .B(n68313), .C(n68315), .Y(n68328)
         );
  MAJIxp5_ASAP7_75t_SL U71612 ( .A(n68340), .B(n58360), .C(n58367), .Y(n68348)
         );
  MAJIxp5_ASAP7_75t_SL U71613 ( .A(n68357), .B(n56832), .C(n68356), .Y(n68460)
         );
  XNOR2xp5_ASAP7_75t_SL U71614 ( .A(n68362), .B(n68361), .Y(n68363) );
  MAJIxp5_ASAP7_75t_SL U71615 ( .A(n68376), .B(n68375), .C(n68374), .Y(n68440)
         );
  O2A1O1Ixp5_ASAP7_75t_SL U71616 ( .A1(n58753), .A2(n68380), .B(n68379), .C(
        n68378), .Y(n68438) );
  MAJIxp5_ASAP7_75t_SL U71617 ( .A(n68440), .B(n68439), .C(n57146), .Y(n68489)
         );
  MAJIxp5_ASAP7_75t_SL U71618 ( .A(n68460), .B(n68459), .C(n68458), .Y(n68496)
         );
  XNOR2xp5_ASAP7_75t_SL U71619 ( .A(n68464), .B(n68463), .Y(n68476) );
  MAJIxp5_ASAP7_75t_SL U71620 ( .A(n68472), .B(n68471), .C(n68470), .Y(n68477)
         );
  XNOR2xp5_ASAP7_75t_SL U71621 ( .A(n68496), .B(n68473), .Y(n68474) );
  MAJIxp5_ASAP7_75t_SL U71622 ( .A(n68478), .B(n68477), .C(n68476), .Y(n68533)
         );
  MAJIxp5_ASAP7_75t_SL U71623 ( .A(n68490), .B(n68489), .C(n68488), .Y(n68522)
         );
  MAJIxp5_ASAP7_75t_SL U71624 ( .A(n68513), .B(n68512), .C(n68511), .Y(n68538)
         );
  MAJIxp5_ASAP7_75t_SL U71625 ( .A(n68518), .B(n58388), .C(n68520), .Y(n68539)
         );
  XNOR2xp5_ASAP7_75t_SL U71626 ( .A(n68525), .B(n68524), .Y(n68526) );
  MAJIxp5_ASAP7_75t_SL U71627 ( .A(n68530), .B(n68529), .C(n68528), .Y(n68549)
         );
  MAJIxp5_ASAP7_75t_SL U71628 ( .A(n69035), .B(n69034), .C(n69036), .Y(n68591)
         );
  MAJIxp5_ASAP7_75t_SL U71629 ( .A(n68557), .B(n68558), .C(n58500), .Y(n68587)
         );
  NAND3xp33_ASAP7_75t_SL U71630 ( .A(n69006), .B(n69012), .C(n68955), .Y(
        n68582) );
  AND2x2_ASAP7_75t_SL U71631 ( .A(n68609), .B(n75072), .Y(n68611) );
  OR2x2_ASAP7_75t_SL U71632 ( .A(n68620), .B(n68619), .Y(n75041) );
  AO21x1_ASAP7_75t_SL U71633 ( .A1(n75059), .A2(n75105), .B(n68641), .Y(n68645) );
  AND2x2_ASAP7_75t_SL U71634 ( .A(n75098), .B(n75041), .Y(n68643) );
  OA21x2_ASAP7_75t_SL U71635 ( .A1(n68650), .A2(n69233), .B(n68678), .Y(n69295) );
  NAND3xp33_ASAP7_75t_SL U71636 ( .A(n68657), .B(n68654), .C(n57376), .Y(
        n68661) );
  XOR2xp5_ASAP7_75t_SL U71637 ( .A(n68654), .B(n69300), .Y(n68655) );
  NOR3xp33_ASAP7_75t_SL U71638 ( .A(n69235), .B(n69225), .C(n68671), .Y(n68681) );
  NAND3xp33_ASAP7_75t_SL U71639 ( .A(n68672), .B(n68671), .C(n68670), .Y(
        n68677) );
  A2O1A1Ixp33_ASAP7_75t_SL U71640 ( .A1(n68679), .A2(n68678), .B(n68677), .C(
        n68676), .Y(n68680) );
  AO21x1_ASAP7_75t_SL U71641 ( .A1(n68681), .A2(n59449), .B(n68680), .Y(n68682) );
  O2A1O1Ixp5_ASAP7_75t_SL U71642 ( .A1(n69119), .A2(n69118), .B(n69147), .C(
        n68695), .Y(n68696) );
  OR2x2_ASAP7_75t_SL U71643 ( .A(n68711), .B(n75278), .Y(n75284) );
  AND2x2_ASAP7_75t_SL U71644 ( .A(n69028), .B(n69027), .Y(n68732) );
  NAND3xp33_ASAP7_75t_SL U71645 ( .A(n69030), .B(n69029), .C(n68729), .Y(
        n68733) );
  AND2x2_ASAP7_75t_SL U71646 ( .A(n68738), .B(n68808), .Y(n68744) );
  XOR2xp5_ASAP7_75t_SL U71647 ( .A(n68752), .B(n68751), .Y(n52059) );
  A2O1A1Ixp33_ASAP7_75t_SL U71648 ( .A1(n68761), .A2(n68760), .B(n68759), .C(
        n68763), .Y(n68762) );
  OAI31xp33_ASAP7_75t_SL U71649 ( .A1(n68765), .A2(n68764), .A3(n68763), .B(
        n68762), .Y(n52058) );
  OR2x2_ASAP7_75t_SL U71650 ( .A(or1200_cpu_or1200_mult_mac_n339), .B(
        or1200_cpu_or1200_mult_mac_n193), .Y(n68777) );
  OR2x2_ASAP7_75t_SL U71651 ( .A(or1200_cpu_or1200_mult_mac_n341), .B(
        or1200_cpu_or1200_mult_mac_n195), .Y(n75000) );
  OR2x2_ASAP7_75t_SL U71652 ( .A(or1200_cpu_or1200_mult_mac_n201), .B(
        or1200_cpu_or1200_mult_mac_n347), .Y(n68821) );
  XOR2xp5_ASAP7_75t_SL U71653 ( .A(n68786), .B(n68815), .Y(n68788) );
  NAND3xp33_ASAP7_75t_SL U71654 ( .A(n75018), .B(n74997), .C(n68796), .Y(
        n68798) );
  OR2x2_ASAP7_75t_SL U71655 ( .A(or1200_cpu_or1200_mult_mac_n203), .B(
        or1200_cpu_or1200_mult_mac_n349), .Y(n76886) );
  AO21x1_ASAP7_75t_SL U71656 ( .A1(n76886), .A2(n76887), .B(n76885), .Y(n68832) );
  XOR2xp5_ASAP7_75t_SL U71657 ( .A(n68839), .B(n68840), .Y(n51992) );
  A2O1A1Ixp33_ASAP7_75t_SL U71658 ( .A1(n68847), .A2(n68846), .B(n68845), .C(
        n68886), .Y(n68862) );
  OAI211xp5_ASAP7_75t_SL U71659 ( .A1(n58389), .A2(n68852), .B(n68857), .C(
        n53199), .Y(n68856) );
  NAND3xp33_ASAP7_75t_SL U71660 ( .A(n68858), .B(n68853), .C(n68852), .Y(
        n68854) );
  NAND3xp33_ASAP7_75t_SL U71661 ( .A(n68867), .B(n68866), .C(n57129), .Y(
        n68871) );
  O2A1O1Ixp5_ASAP7_75t_SL U71662 ( .A1(n68877), .A2(n68876), .B(n68875), .C(
        n68874), .Y(n68942) );
  NAND3xp33_ASAP7_75t_SL U71663 ( .A(n68878), .B(n69054), .C(n69050), .Y(
        n68944) );
  OR2x2_ASAP7_75t_SL U71664 ( .A(or1200_cpu_or1200_mult_mac_n357), .B(
        or1200_cpu_or1200_mult_mac_n211), .Y(n68936) );
  A2O1A1Ixp33_ASAP7_75t_SL U71665 ( .A1(n68886), .A2(n68885), .B(n68884), .C(
        n68883), .Y(n68887) );
  A2O1A1Ixp33_ASAP7_75t_SL U71666 ( .A1(n68891), .A2(n68890), .B(n68889), .C(
        n68888), .Y(n68937) );
  A2O1A1Ixp33_ASAP7_75t_SL U71667 ( .A1(n57080), .A2(n68911), .B(n68896), .C(
        n68895), .Y(n68897) );
  AND2x2_ASAP7_75t_SL U71668 ( .A(n57421), .B(n68909), .Y(n68964) );
  XOR2xp5_ASAP7_75t_SL U71669 ( .A(n68923), .B(n68910), .Y(n51994) );
  NOR3xp33_ASAP7_75t_SL U71670 ( .A(n68918), .B(n68925), .C(n68924), .Y(n68922) );
  A2O1A1Ixp33_ASAP7_75t_SL U71671 ( .A1(n68927), .A2(n68926), .B(n68925), .C(
        n68924), .Y(n68928) );
  NAND3xp33_ASAP7_75t_SL U71672 ( .A(n68930), .B(n68929), .C(n68928), .Y(
        n51996) );
  A2O1A1Ixp33_ASAP7_75t_SL U71673 ( .A1(n57079), .A2(n68949), .B(n68951), .C(
        n68948), .Y(n68954) );
  AND2x2_ASAP7_75t_SL U71674 ( .A(n68959), .B(n68957), .Y(n68958) );
  OAI211xp5_ASAP7_75t_SL U71675 ( .A1(n68974), .A2(n58377), .B(n59382), .C(
        n68973), .Y(n68982) );
  OAI31xp33_ASAP7_75t_SL U71676 ( .A1(n68978), .A2(n58887), .A3(n68975), .B(
        n59382), .Y(n68980) );
  O2A1O1Ixp5_ASAP7_75t_SL U71677 ( .A1(n68982), .A2(n68981), .B(n68980), .C(
        n68979), .Y(n68983) );
  XNOR2xp5_ASAP7_75t_SL U71678 ( .A(n68984), .B(n68983), .Y(n51990) );
  A2O1A1Ixp33_ASAP7_75t_SL U71679 ( .A1(n68992), .A2(n68991), .B(n68990), .C(
        n68989), .Y(n69058) );
  OR2x2_ASAP7_75t_SL U71680 ( .A(or1200_cpu_or1200_mult_mac_n367), .B(
        or1200_cpu_or1200_mult_mac_n221), .Y(n69019) );
  A2O1A1Ixp33_ASAP7_75t_SL U71681 ( .A1(n69001), .A2(n69000), .B(n68999), .C(
        n68998), .Y(n69018) );
  A2O1A1Ixp33_ASAP7_75t_SL U71682 ( .A1(n69012), .A2(n69011), .B(n69010), .C(
        n69009), .Y(n69013) );
  A2O1A1Ixp33_ASAP7_75t_SL U71683 ( .A1(n69045), .A2(n69044), .B(n69043), .C(
        n69042), .Y(n69046) );
  NAND4xp25_ASAP7_75t_SL U71684 ( .A(n69055), .B(n69054), .C(n69059), .D(
        n69053), .Y(n69063) );
  O2A1O1Ixp5_ASAP7_75t_SL U71685 ( .A1(n69064), .A2(n69063), .B(n69067), .C(
        n69062), .Y(n69070) );
  A2O1A1Ixp33_ASAP7_75t_SL U71686 ( .A1(n69081), .A2(n69080), .B(n69079), .C(
        n69078), .Y(or1200_cpu_or1200_mult_mac_n1613) );
  AND2x2_ASAP7_75t_SL U71687 ( .A(n69169), .B(n69165), .Y(n69093) );
  NAND3xp33_ASAP7_75t_SL U71688 ( .A(n69105), .B(n69104), .C(n69103), .Y(
        n52004) );
  A2O1A1Ixp33_ASAP7_75t_SL U71689 ( .A1(n69121), .A2(n69115), .B(n69151), .C(
        n69120), .Y(n69123) );
  OR2x2_ASAP7_75t_SL U71690 ( .A(or1200_cpu_or1200_mult_mac_n231), .B(
        or1200_cpu_or1200_mult_mac_n377), .Y(n69281) );
  XOR2xp5_ASAP7_75t_SL U71691 ( .A(n69131), .B(n69161), .Y(n69129) );
  AO21x1_ASAP7_75t_SL U71692 ( .A1(n69168), .A2(n69130), .B(n69164), .Y(n69133) );
  A2O1A1Ixp33_ASAP7_75t_SL U71693 ( .A1(n69162), .A2(n69166), .B(n69134), .C(
        n57080), .Y(n69135) );
  AND2x2_ASAP7_75t_SL U71694 ( .A(n69145), .B(n53206), .Y(n69152) );
  O2A1O1Ixp5_ASAP7_75t_SL U71695 ( .A1(n69178), .A2(n69177), .B(n69176), .C(
        n69175), .Y(n69190) );
  XOR2xp5_ASAP7_75t_SL U71696 ( .A(n69181), .B(n69180), .Y(n69184) );
  AO21x1_ASAP7_75t_SL U71697 ( .A1(n69247), .A2(n74116), .B(n69245), .Y(n69217) );
  A2O1A1Ixp33_ASAP7_75t_SL U71698 ( .A1(n69207), .A2(n74571), .B(n74570), .C(
        n69210), .Y(n69208) );
  AO21x1_ASAP7_75t_SL U71699 ( .A1(n74115), .A2(n74117), .B(n69244), .Y(n69219) );
  A2O1A1Ixp33_ASAP7_75t_SL U71700 ( .A1(n69224), .A2(n69223), .B(n69222), .C(
        n69221), .Y(or1200_cpu_or1200_mult_mac_n1603) );
  A2O1A1Ixp33_ASAP7_75t_SL U71701 ( .A1(n69235), .A2(n69234), .B(n69233), .C(
        n69232), .Y(n69236) );
  A2O1A1Ixp33_ASAP7_75t_SL U71702 ( .A1(n69252), .A2(n69251), .B(n69250), .C(
        n69249), .Y(n69254) );
  A2O1A1Ixp33_ASAP7_75t_SL U71703 ( .A1(n69269), .A2(n69268), .B(n69267), .C(
        n69266), .Y(or1200_cpu_or1200_mult_mac_n1601) );
  O2A1O1Ixp5_ASAP7_75t_SL U71704 ( .A1(n69286), .A2(n69285), .B(n69284), .C(
        n69283), .Y(n69287) );
  A2O1A1Ixp33_ASAP7_75t_SL U71705 ( .A1(n57080), .A2(n69318), .B(n69317), .C(
        n69316), .Y(n69319) );
  OR2x2_ASAP7_75t_SL U71706 ( .A(or1200_cpu_or1200_mult_mac_n255), .B(
        or1200_cpu_or1200_mult_mac_n401), .Y(n75120) );
  A2O1A1Ixp33_ASAP7_75t_SL U71707 ( .A1(n77172), .A2(n69341), .B(n69340), .C(
        n59694), .Y(n69342) );
  A2O1A1Ixp33_ASAP7_75t_SL U71708 ( .A1(n78089), .A2(n69359), .B(n74041), .C(
        n69358), .Y(n69360) );
  AND2x2_ASAP7_75t_SL U71709 ( .A(n78095), .B(n69360), .Y(n74082) );
  OR2x2_ASAP7_75t_SL U71710 ( .A(n70478), .B(n70385), .Y(n70531) );
  AND2x2_ASAP7_75t_SL U71711 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_4_), .B(n2452), .Y(
        n70313) );
  OR2x2_ASAP7_75t_SL U71712 ( .A(n70246), .B(n70313), .Y(n9560) );
  O2A1O1Ixp5_ASAP7_75t_SL U71713 ( .A1(n69389), .A2(n78335), .B(n69388), .C(
        n69387), .Y(n69401) );
  NAND3xp33_ASAP7_75t_SL U71714 ( .A(n69394), .B(n69400), .C(n69393), .Y(
        n69397) );
  A2O1A1Ixp33_ASAP7_75t_SL U71715 ( .A1(n69398), .A2(n78337), .B(n69397), .C(
        n69396), .Y(n69399) );
  O2A1O1Ixp5_ASAP7_75t_SL U71716 ( .A1(n69402), .A2(n69401), .B(n69400), .C(
        n69399), .Y(n69403) );
  O2A1O1Ixp5_ASAP7_75t_SL U71717 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_2_), .A2(n69413), .B(
        n69412), .C(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_10_), .Y(
        n69416) );
  O2A1O1Ixp5_ASAP7_75t_SL U71718 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_5_), .A2(n78335), .B(
        n78339), .C(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_7_), .Y(
        n69414) );
  A2O1A1Ixp33_ASAP7_75t_SL U71719 ( .A1(n69416), .A2(n69415), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_11_), .C(n78351), .Y(
        n69417) );
  A2O1A1Ixp33_ASAP7_75t_SL U71720 ( .A1(n69417), .A2(n78352), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_14_), .C(n78353), .Y(
        n69418) );
  A2O1A1Ixp33_ASAP7_75t_SL U71721 ( .A1(n69418), .A2(n78431), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_17_), .C(n78355), .Y(
        n69419) );
  OR2x2_ASAP7_75t_SL U71722 ( .A(n70112), .B(n70109), .Y(n69564) );
  A2O1A1Ixp33_ASAP7_75t_SL U71723 ( .A1(n69429), .A2(n69428), .B(n69438), .C(
        n69427), .Y(n69430) );
  OR2x2_ASAP7_75t_SL U71724 ( .A(n70114), .B(n70109), .Y(n69497) );
  OR2x2_ASAP7_75t_SL U71725 ( .A(n69436), .B(n69443), .Y(n69747) );
  AO21x1_ASAP7_75t_SL U71726 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_0_), .A2(n70019), .B(
        n70118), .Y(n69452) );
  A2O1A1Ixp33_ASAP7_75t_SL U71727 ( .A1(n69742), .A2(n69580), .B(n69452), .C(
        n69451), .Y(n69570) );
  OR2x2_ASAP7_75t_SL U71728 ( .A(n78339), .B(n70114), .Y(n69489) );
  A2O1A1Ixp33_ASAP7_75t_SL U71729 ( .A1(n78341), .A2(n70114), .B(n70109), .C(
        n69489), .Y(n69456) );
  A2O1A1Ixp33_ASAP7_75t_SL U71730 ( .A1(n69476), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_8_), .B(n69456), .C(
        n69455), .Y(n69507) );
  NOR3xp33_ASAP7_75t_SL U71731 ( .A(n70021), .B(n70118), .C(n78429), .Y(n69462) );
  A2O1A1Ixp33_ASAP7_75t_SL U71732 ( .A1(n78431), .A2(n70114), .B(n69463), .C(
        n70109), .Y(n69464) );
  OAI211xp5_ASAP7_75t_SL U71733 ( .A1(n69564), .A2(n78357), .B(n69469), .C(
        n69468), .Y(n69470) );
  OAI211xp5_ASAP7_75t_SL U71734 ( .A1(n78353), .A2(n70021), .B(n69474), .C(
        n69473), .Y(n70079) );
  OAI211xp5_ASAP7_75t_SL U71735 ( .A1(n78341), .A2(n70021), .B(n69482), .C(
        n69481), .Y(n69567) );
  O2A1O1Ixp5_ASAP7_75t_SL U71736 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_7_), .A2(n69492), .B(
        n69491), .C(n69490), .Y(n69493) );
  AO21x1_ASAP7_75t_SL U71737 ( .A1(n70114), .A2(n69499), .B(n69498), .Y(n70026) );
  NOR3xp33_ASAP7_75t_SL U71738 ( .A(n69577), .B(n70112), .C(n69941), .Y(n69508) );
  A2O1A1Ixp33_ASAP7_75t_SL U71739 ( .A1(n69512), .A2(n69511), .B(n70118), .C(
        n69510), .Y(n69513) );
  A2O1A1Ixp33_ASAP7_75t_SL U71740 ( .A1(n69531), .A2(n69530), .B(n69529), .C(
        n69528), .Y(n69903) );
  A2O1A1Ixp33_ASAP7_75t_SL U71741 ( .A1(n69539), .A2(n69538), .B(n69537), .C(
        n69536), .Y(n69544) );
  A2O1A1Ixp33_ASAP7_75t_SL U71742 ( .A1(n69544), .A2(n69543), .B(n69542), .C(
        n69541), .Y(n69548) );
  A2O1A1Ixp33_ASAP7_75t_SL U71743 ( .A1(n69548), .A2(n69547), .B(n69546), .C(
        n78364), .Y(n69766) );
  A2O1A1Ixp33_ASAP7_75t_SL U71744 ( .A1(n78330), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[0]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[2]), .C(n69549), 
        .Y(n69551) );
  A2O1A1Ixp33_ASAP7_75t_SL U71745 ( .A1(n69551), .A2(n69550), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[7]), .C(n78342), 
        .Y(n69552) );
  A2O1A1Ixp33_ASAP7_75t_SL U71746 ( .A1(n69552), .A2(n78344), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[10]), .C(n78346), .Y(n69553) );
  A2O1A1Ixp33_ASAP7_75t_SL U71747 ( .A1(n69553), .A2(n78350), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[13]), .C(n78427), .Y(n69554) );
  A2O1A1Ixp33_ASAP7_75t_SL U71748 ( .A1(n69554), .A2(n78426), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[16]), .C(n78424), .Y(n69555) );
  A2O1A1Ixp33_ASAP7_75t_SL U71749 ( .A1(n69555), .A2(n78354), .B(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[19]), .C(n78368), .Y(n69556) );
  OR2x2_ASAP7_75t_SL U71750 ( .A(n69581), .B(n69573), .Y(n17032) );
  OR2x2_ASAP7_75t_SL U71751 ( .A(n69581), .B(n69940), .Y(n17035) );
  OR2x2_ASAP7_75t_SL U71752 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_0_), .B(n2451), .Y(
        n70260) );
  NAND3xp33_ASAP7_75t_SL U71753 ( .A(n69711), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_23_), .C(n69712), 
        .Y(n70092) );
  NAND3xp33_ASAP7_75t_SL U71754 ( .A(n69592), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_1_), .C(n69591), .Y(
        n69720) );
  NAND3xp33_ASAP7_75t_SL U71755 ( .A(n69789), .B(n69610), .C(n69609), .Y(
        n69619) );
  NAND3xp33_ASAP7_75t_SL U71756 ( .A(n69783), .B(n69771), .C(n69781), .Y(
        n69791) );
  A2O1A1Ixp33_ASAP7_75t_SL U71757 ( .A1(n69750), .A2(n69761), .B(n69619), .C(
        n69618), .Y(n69638) );
  A2O1A1Ixp33_ASAP7_75t_SL U71758 ( .A1(n69638), .A2(n69637), .B(n69636), .C(
        n58568), .Y(n69661) );
  A2O1A1Ixp33_ASAP7_75t_SL U71759 ( .A1(n69661), .A2(n69660), .B(n69659), .C(
        n69658), .Y(n69677) );
  A2O1A1Ixp33_ASAP7_75t_SL U71760 ( .A1(n69677), .A2(n69676), .B(n69958), .C(
        n69675), .Y(n69700) );
  NOR3xp33_ASAP7_75t_SL U71761 ( .A(n70006), .B(n70071), .C(n70047), .Y(n69697) );
  A2O1A1Ixp33_ASAP7_75t_SL U71762 ( .A1(n69700), .A2(n69699), .B(n69698), .C(
        n69697), .Y(n69710) );
  NAND3xp33_ASAP7_75t_SL U71763 ( .A(n69704), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvsor_i_21_), .C(n69703), 
        .Y(n70049) );
  OR2x2_ASAP7_75t_SL U71764 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[24]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_dvd[26]), .Y(n69714) );
  OA21x2_ASAP7_75t_SL U71765 ( .A1(n69717), .A2(n69716), .B(n69715), .Y(n70372) );
  AND2x2_ASAP7_75t_SL U71766 ( .A(n69725), .B(n69767), .Y(n69956) );
  OR2x2_ASAP7_75t_SL U71767 ( .A(n70081), .B(n69876), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvsor[7]) );
  OA21x2_ASAP7_75t_SL U71768 ( .A1(n69807), .A2(n58553), .B(n69806), .Y(n2295)
         );
  OAI222xp33_ASAP7_75t_SL U71769 ( .A1(n70032), .A2(n69878), .B1(n69902), .B2(
        n70043), .C1(n69877), .C2(n70030), .Y(n3212) );
  OR2x2_ASAP7_75t_SL U71770 ( .A(n69859), .B(n69852), .Y(n69865) );
  NAND3xp33_ASAP7_75t_SL U71771 ( .A(n69865), .B(n69864), .C(n69863), .Y(
        n69869) );
  A2O1A1Ixp33_ASAP7_75t_SL U71772 ( .A1(n69914), .A2(n69869), .B(n58553), .C(
        n69868), .Y(n2287) );
  OA21x2_ASAP7_75t_SL U71773 ( .A1(n69889), .A2(n58553), .B(n69888), .Y(n2285)
         );
  AND2x2_ASAP7_75t_SL U71774 ( .A(n69903), .B(n70081), .Y(n70033) );
  OAI211xp5_ASAP7_75t_SL U71775 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[15]), .A2(
        n69925), .B(n69896), .C(n69895), .Y(n69998) );
  OR2x2_ASAP7_75t_SL U71776 ( .A(n69916), .B(n69915), .Y(n69921) );
  OAI211xp5_ASAP7_75t_SL U71777 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_mul_fractb_24[16]), .A2(
        n69925), .B(n69924), .C(n69923), .Y(n70041) );
  OR2x2_ASAP7_75t_SL U71778 ( .A(n69960), .B(n69934), .Y(n69939) );
  A2O1A1Ixp33_ASAP7_75t_SL U71779 ( .A1(n69969), .A2(n69968), .B(n69967), .C(
        n69966), .Y(n69970) );
  OAI211xp5_ASAP7_75t_SL U71780 ( .A1(n78354), .A2(n70054), .B(n69976), .C(
        n69975), .Y(n70082) );
  A2O1A1Ixp33_ASAP7_75t_SL U71781 ( .A1(n69980), .A2(n69979), .B(n70064), .C(
        n69978), .Y(n69981) );
  A2O1A1Ixp33_ASAP7_75t_SL U71782 ( .A1(n70014), .A2(n70013), .B(n58555), .C(
        n70012), .Y(n70015) );
  A2O1A1Ixp33_ASAP7_75t_SL U71783 ( .A1(n70017), .A2(n70078), .B(n70016), .C(
        n70149), .Y(n70025) );
  OAI211xp5_ASAP7_75t_SL U71784 ( .A1(n70118), .A2(n70026), .B(n70025), .C(
        n70024), .Y(n70027) );
  OAI211xp5_ASAP7_75t_SL U71785 ( .A1(n70064), .A2(n70041), .B(n70040), .C(
        n70039), .Y(n70042) );
  NOR3xp33_ASAP7_75t_SL U71786 ( .A(n70079), .B(n70078), .C(n70077), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_pre_norm_div_dvdnd[49]) );
  OR2x2_ASAP7_75t_SL U71787 ( .A(n70083), .B(n70082), .Y(n70084) );
  MAJIxp5_ASAP7_75t_SL U71788 ( .A(n70109), .B(n70108), .C(n70107), .Y(n70131)
         );
  XNOR2xp5_ASAP7_75t_SL U71789 ( .A(n70132), .B(n70135), .Y(n70140) );
  XNOR2xp5_ASAP7_75t_SL U71790 ( .A(n70125), .B(n70124), .Y(n70128) );
  MAJIxp5_ASAP7_75t_SL U71791 ( .A(n70142), .B(n70141), .C(n70140), .Y(n70143)
         );
  AO21x1_ASAP7_75t_SL U71792 ( .A1(n70144), .A2(n70143), .B(n70164), .Y(n3260)
         );
  MAJIxp5_ASAP7_75t_SL U71793 ( .A(n70153), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[3]), .C(
        n70152), .Y(n70158) );
  XNOR2xp5_ASAP7_75t_SL U71794 ( .A(n70158), .B(n70157), .Y(n70159) );
  OR2x2_ASAP7_75t_SL U71795 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[5]), .Y(
        n70184) );
  XOR2xp5_ASAP7_75t_SL U71796 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[7]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[5]), .Y(
        n70193) );
  O2A1O1Ixp5_ASAP7_75t_SL U71797 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expa_in[7]), .A2(
        n70193), .B(n70192), .C(n70191), .Y(n70200) );
  XNOR2xp5_ASAP7_75t_SL U71798 ( .A(n70201), .B(n70200), .Y(n70199) );
  AO21x1_ASAP7_75t_SL U71799 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_pre_norm_div_s_expb_in[7]), .A2(
        n70206), .B(n70205), .Y(n70207) );
  A2O1A1Ixp33_ASAP7_75t_SL U71800 ( .A1(n70209), .A2(n70208), .B(n70207), .C(
        n3254), .Y(n70210) );
  AND2x2_ASAP7_75t_SL U71801 ( .A(n70245), .B(n3154), .Y(n70242) );
  A2O1A1Ixp33_ASAP7_75t_SL U71802 ( .A1(n70226), .A2(n70571), .B(n70225), .C(
        n70239), .Y(n70227) );
  AND2x2_ASAP7_75t_SL U71803 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_0_), .B(n2451), .Y(
        n70270) );
  A2O1A1Ixp33_ASAP7_75t_SL U71804 ( .A1(n2456), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[25]), .B(n70231), .C(
        n70230), .Y(n2417) );
  XNOR2xp5_ASAP7_75t_SL U71805 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[5]), .B(
        n70233), .Y(n70587) );
  AO21x1_ASAP7_75t_SL U71806 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[3]), .A2(
        n70238), .B(n70237), .Y(n70573) );
  A2O1A1Ixp33_ASAP7_75t_SL U71807 ( .A1(n70241), .A2(n70573), .B(n70240), .C(
        n70239), .Y(n70243) );
  NOR3xp33_ASAP7_75t_SL U71808 ( .A(n70245), .B(n70311), .C(n70244), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_v_shl_0_) );
  AO21x1_ASAP7_75t_SL U71809 ( .A1(n70249), .A2(n70372), .B(n70248), .Y(n2320)
         );
  OR2x2_ASAP7_75t_SL U71810 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_5_), .B(
        n70272), .Y(n70537) );
  OR2x2_ASAP7_75t_SL U71811 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_5_), .B(n2437), .Y(n70251) );
  OR2x2_ASAP7_75t_SL U71812 ( .A(n70303), .B(n59621), .Y(n70305) );
  OR2x2_ASAP7_75t_SL U71813 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_24_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_1_), .Y(
        n70264) );
  O2A1O1Ixp5_ASAP7_75t_SL U71814 ( .A1(n74680), .A2(n70258), .B(n70264), .C(
        n70257), .Y(n70295) );
  AND2x2_ASAP7_75t_SL U71815 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_0_), .Y(
        n74686) );
  A2O1A1Ixp33_ASAP7_75t_SL U71816 ( .A1(n70276), .A2(n70275), .B(n70274), .C(
        n70273), .Y(n70429) );
  A2O1A1Ixp33_ASAP7_75t_SL U71817 ( .A1(n70542), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_), .B(
        n70284), .C(n74706), .Y(n70362) );
  A2O1A1Ixp33_ASAP7_75t_SL U71818 ( .A1(n70295), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_2_), .B(
        n70294), .C(n70293), .Y(n70465) );
  A2O1A1Ixp33_ASAP7_75t_SL U71819 ( .A1(n2456), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_serial_div_qutnt[16]), .B(n70313), .C(
        n70312), .Y(n2330) );
  NAND3xp33_ASAP7_75t_SL U71820 ( .A(n70316), .B(n70315), .C(n70314), .Y(
        n70389) );
  NAND3xp33_ASAP7_75t_SL U71821 ( .A(n70320), .B(n70319), .C(n70318), .Y(
        n70388) );
  A2O1A1Ixp33_ASAP7_75t_SL U71822 ( .A1(n74706), .A2(n70389), .B(n70321), .C(
        n70483), .Y(n70533) );
  A2O1A1Ixp33_ASAP7_75t_SL U71823 ( .A1(n70533), .A2(n70532), .B(n70405), .C(
        n70322), .Y(n70323) );
  OR2x2_ASAP7_75t_SL U71824 ( .A(n2450), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_div_s_count_4_), .Y(n70376) );
  OR2x2_ASAP7_75t_SL U71825 ( .A(n70376), .B(n59621), .Y(n70378) );
  A2O1A1Ixp33_ASAP7_75t_SL U71826 ( .A1(n70416), .A2(n70427), .B(n70342), .C(
        n70341), .Y(n2340) );
  A2O1A1Ixp33_ASAP7_75t_SL U71827 ( .A1(n70422), .A2(n70344), .B(n70343), .C(
        n2456), .Y(n2372) );
  NAND3xp33_ASAP7_75t_SL U71828 ( .A(n70347), .B(n70346), .C(n70345), .Y(
        n70382) );
  OAI211xp5_ASAP7_75t_SL U71829 ( .A1(n70432), .A2(n70405), .B(n70370), .C(
        n70351), .Y(n70352) );
  NAND3xp33_ASAP7_75t_SL U71830 ( .A(n70357), .B(n70356), .C(n70355), .Y(
        n70536) );
  NAND3xp33_ASAP7_75t_SL U71831 ( .A(n70362), .B(n70361), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .Y(
        n70363) );
  A2O1A1Ixp33_ASAP7_75t_SL U71832 ( .A1(n70366), .A2(n70365), .B(n70364), .C(
        n70363), .Y(n2370) );
  OR2x2_ASAP7_75t_SL U71833 ( .A(n74706), .B(n70373), .Y(n70474) );
  A2O1A1Ixp33_ASAP7_75t_SL U71834 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .A2(
        n70468), .B(n70375), .C(n70374), .Y(n2406) );
  OAI211xp5_ASAP7_75t_SL U71835 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_11_), .A2(
        n70540), .B(n70381), .C(n70380), .Y(n70431) );
  NAND3xp33_ASAP7_75t_SL U71836 ( .A(n70392), .B(n70391), .C(n70390), .Y(
        n70534) );
  OR2x2_ASAP7_75t_SL U71837 ( .A(n70478), .B(n59621), .Y(n70480) );
  O2A1O1Ixp5_ASAP7_75t_SL U71838 ( .A1(n70548), .A2(n70405), .B(n70404), .C(
        n70403), .Y(n70406) );
  OAI211xp5_ASAP7_75t_SL U71839 ( .A1(n70535), .A2(n70416), .B(n70415), .C(
        n70414), .Y(n70418) );
  OA21x2_ASAP7_75t_SL U71840 ( .A1(n70469), .A2(n70418), .B(n70417), .Y(n2350)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U71841 ( .A1(n70422), .A2(n70421), .B(n70420), .C(
        n2456), .Y(n2382) );
  A2O1A1Ixp33_ASAP7_75t_SL U71842 ( .A1(n70541), .A2(n70489), .B(n70444), .C(
        n70428), .Y(n70435) );
  NAND3xp33_ASAP7_75t_SL U71843 ( .A(n70435), .B(n70434), .C(n70433), .Y(n2354) );
  A2O1A1Ixp33_ASAP7_75t_SL U71844 ( .A1(n70541), .A2(n70538), .B(n70444), .C(
        n70443), .Y(n70453) );
  AO21x1_ASAP7_75t_SL U71845 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_21_), .A2(
        n70445), .B(n70466), .Y(n70448) );
  O2A1O1Ixp5_ASAP7_75t_SL U71846 ( .A1(n70451), .A2(n70450), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_shr1_3_), .C(
        n70449), .Y(n70452) );
  A2O1A1Ixp33_ASAP7_75t_SL U71847 ( .A1(n70541), .A2(n70544), .B(n70469), .C(
        n70460), .Y(n70464) );
  OAI211xp5_ASAP7_75t_SL U71848 ( .A1(n70466), .A2(n70465), .B(n70464), .C(
        n70463), .Y(n2396) );
  OA21x2_ASAP7_75t_SL U71849 ( .A1(n70502), .A2(n70501), .B(n70500), .Y(n2258)
         );
  OR2x2_ASAP7_75t_SL U71850 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_0_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_1_), .Y(n70567) );
  NAND3xp33_ASAP7_75t_SL U71851 ( .A(n74711), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r2_1_), .C(n70565), .Y(
        n74284) );
  A2O1A1Ixp33_ASAP7_75t_SL U71852 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[1]), .A2(
        n70569), .B(n70568), .C(n70597), .Y(n3161) );
  OR2x2_ASAP7_75t_SL U71853 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[1]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[2]), .Y(
        n70582) );
  XNOR2xp5_ASAP7_75t_SL U71854 ( .A(n70596), .B(n70595), .Y(n51981) );
  A2O1A1Ixp33_ASAP7_75t_SL U71855 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_exp_10_i[7]), .A2(
        n70599), .B(n70598), .C(n70597), .Y(n3155) );
  A2O1A1Ixp33_ASAP7_75t_SL U71856 ( .A1(n70614), .A2(n70613), .B(n70612), .C(
        n70616), .Y(n70615) );
  XNOR2xp5_ASAP7_75t_SL U71857 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_expo1[8]), .B(
        n70618), .Y(n53175) );
  NAND3xp33_ASAP7_75t_SL U71858 ( .A(n70625), .B(n70624), .C(n70623), .Y(
        n70626) );
  OR3x1_ASAP7_75t_SL U71859 ( .A(n70628), .B(n70627), .C(n70626), .Y(n70638)
         );
  NOR3xp33_ASAP7_75t_SL U71860 ( .A(n70686), .B(n71281), .C(n71284), .Y(n70650) );
  OAI211xp5_ASAP7_75t_SL U71861 ( .A1(n57211), .A2(n58302), .B(n70648), .C(
        n70642), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n250) );
  NAND3xp33_ASAP7_75t_SL U71862 ( .A(n70648), .B(n70643), .C(n70646), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n249) );
  OR2x2_ASAP7_75t_SL U71863 ( .A(n71015), .B(n70646), .Y(n70649) );
  OAI211xp5_ASAP7_75t_SL U71864 ( .A1(n53473), .A2(n70644), .B(n70648), .C(
        n70649), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n248) );
  OAI211xp5_ASAP7_75t_SL U71865 ( .A1(n70812), .A2(n70649), .B(n70648), .C(
        n70645), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n251) );
  OAI211xp5_ASAP7_75t_SL U71866 ( .A1(n70725), .A2(n70649), .B(n70648), .C(
        n70647), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n252) );
  OAI211xp5_ASAP7_75t_SL U71867 ( .A1(n58315), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fractb_i[3]), .B(n71015), 
        .C(n59526), .Y(n70653) );
  A2O1A1Ixp33_ASAP7_75t_SL U71868 ( .A1(n70660), .A2(n70659), .B(n70658), .C(
        n70657), .Y(n70661) );
  AO21x1_ASAP7_75t_SL U71869 ( .A1(n70664), .A2(n70663), .B(n70662), .Y(n70684) );
  AO21x1_ASAP7_75t_SL U71870 ( .A1(n70671), .A2(n70670), .B(n70669), .Y(n70683) );
  OR2x2_ASAP7_75t_SL U71871 ( .A(n71149), .B(n70768), .Y(n70690) );
  NAND3xp33_ASAP7_75t_SL U71872 ( .A(n71315), .B(n59522), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fracta_i[0]), .Y(n70692) );
  NAND4xp25_ASAP7_75t_SL U71873 ( .A(n53467), .B(n71263), .C(n58302), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_1_), .Y(n70704) );
  NOR3xp33_ASAP7_75t_SL U71874 ( .A(n70789), .B(n70929), .C(n71284), .Y(n70719) );
  XNOR2xp5_ASAP7_75t_SL U71875 ( .A(n70726), .B(n70727), .Y(n70732) );
  NAND3xp33_ASAP7_75t_SL U71876 ( .A(n70731), .B(n70730), .C(n70729), .Y(
        n70734) );
  NAND3xp33_ASAP7_75t_SL U71877 ( .A(n70734), .B(n70733), .C(n70732), .Y(
        n70803) );
  NAND3xp33_ASAP7_75t_SL U71878 ( .A(n70997), .B(n71087), .C(n71263), .Y(
        n70736) );
  OR2x2_ASAP7_75t_SL U71879 ( .A(n70796), .B(n70784), .Y(n70766) );
  NOR3xp33_ASAP7_75t_SL U71880 ( .A(n70789), .B(n71314), .C(n70929), .Y(n70790) );
  XNOR2xp5_ASAP7_75t_SL U71881 ( .A(n70807), .B(n70806), .Y(n70808) );
  AO21x1_ASAP7_75t_SL U71882 ( .A1(n70836), .A2(n70841), .B(n70820), .Y(n70821) );
  A2O1A1Ixp33_ASAP7_75t_SL U71883 ( .A1(n71365), .A2(n70869), .B(n70848), .C(
        n70847), .Y(n70861) );
  XNOR2xp5_ASAP7_75t_SL U71884 ( .A(n70891), .B(n70890), .Y(n70892) );
  NAND3xp33_ASAP7_75t_SL U71885 ( .A(n70901), .B(n70900), .C(n70899), .Y(
        n70903) );
  NAND3xp33_ASAP7_75t_SL U71886 ( .A(n70982), .B(n70908), .C(n70967), .Y(
        n70941) );
  NAND3xp33_ASAP7_75t_SL U71887 ( .A(n70914), .B(n70913), .C(n70912), .Y(
        n71104) );
  NAND3xp33_ASAP7_75t_SL U71888 ( .A(n70917), .B(n70916), .C(n70915), .Y(
        n70919) );
  A2O1A1Ixp33_ASAP7_75t_SL U71889 ( .A1(n70926), .A2(n70925), .B(n70924), .C(
        n57211), .Y(n70927) );
  XNOR2xp5_ASAP7_75t_SL U71890 ( .A(n70945), .B(n70944), .Y(n70946) );
  NAND3xp33_ASAP7_75t_SL U71891 ( .A(n70957), .B(n70956), .C(n70955), .Y(
        n70958) );
  NOR3xp33_ASAP7_75t_SL U71892 ( .A(n70963), .B(n70970), .C(n70962), .Y(n70961) );
  NOR3xp33_ASAP7_75t_SL U71893 ( .A(n70974), .B(n70969), .C(n58303), .Y(n70977) );
  OAI31xp33_ASAP7_75t_SL U71894 ( .A1(n70975), .A2(n70974), .A3(n70973), .B(
        n70972), .Y(n70976) );
  NAND3xp33_ASAP7_75t_SL U71895 ( .A(n71004), .B(n71003), .C(n71002), .Y(
        n71006) );
  AND2x2_ASAP7_75t_SL U71896 ( .A(n71027), .B(n71029), .Y(n71008) );
  NAND3xp33_ASAP7_75t_SL U71897 ( .A(n71009), .B(n71008), .C(n71030), .Y(
        n71007) );
  A2O1A1Ixp33_ASAP7_75t_SL U71898 ( .A1(n71030), .A2(n71009), .B(n71008), .C(
        n71007), .Y(n71010) );
  OA21x2_ASAP7_75t_SL U71899 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_24_), .A2(n71020), 
        .B(n71353), .Y(n71052) );
  NAND3xp33_ASAP7_75t_SL U71900 ( .A(n71023), .B(n71027), .C(n71022), .Y(
        n71025) );
  XNOR2xp5_ASAP7_75t_SL U71901 ( .A(n71037), .B(n71036), .Y(n71038) );
  NAND3xp33_ASAP7_75t_SL U71902 ( .A(n71043), .B(n71042), .C(n71041), .Y(
        n71194) );
  XNOR2xp5_ASAP7_75t_SL U71903 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_25_), .B(n71061), 
        .Y(n71049) );
  A2O1A1Ixp33_ASAP7_75t_SL U71904 ( .A1(n71060), .A2(n71063), .B(n59699), .C(
        n71059), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n178) );
  NAND3xp33_ASAP7_75t_SL U71905 ( .A(n71070), .B(n71069), .C(n71068), .Y(
        n71072) );
  NAND3xp33_ASAP7_75t_SL U71906 ( .A(n71093), .B(n71092), .C(n71091), .Y(
        n71094) );
  NAND3xp33_ASAP7_75t_SL U71907 ( .A(n71107), .B(n71106), .C(n71105), .Y(
        n71121) );
  XNOR2xp5_ASAP7_75t_SL U71908 ( .A(n78398), .B(n71121), .Y(n71108) );
  XNOR2xp5_ASAP7_75t_SL U71909 ( .A(n71124), .B(n71123), .Y(n71125) );
  NAND3xp33_ASAP7_75t_SL U71910 ( .A(n71134), .B(n71131), .C(n71130), .Y(
        n71156) );
  O2A1O1Ixp5_ASAP7_75t_SL U71911 ( .A1(n71136), .A2(n71135), .B(n71134), .C(
        n71133), .Y(n71157) );
  AO21x1_ASAP7_75t_SL U71912 ( .A1(n71396), .A2(n71175), .B(n71150), .Y(n71151) );
  NAND3xp33_ASAP7_75t_SL U71913 ( .A(n71154), .B(n71157), .C(n71153), .Y(
        n71305) );
  NAND3xp33_ASAP7_75t_SL U71914 ( .A(n71165), .B(n71164), .C(n71163), .Y(
        n71166) );
  A2O1A1Ixp33_ASAP7_75t_SL U71915 ( .A1(n71272), .A2(n71189), .B(n71188), .C(
        n71187), .Y(n71190) );
  A2O1A1Ixp33_ASAP7_75t_SL U71916 ( .A1(n57211), .A2(n71191), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_34_), .C(n71190), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_n205) );
  XNOR2xp5_ASAP7_75t_SL U71917 ( .A(n71198), .B(n71197), .Y(n71199) );
  A2O1A1Ixp33_ASAP7_75t_SL U71918 ( .A1(n71201), .A2(n71272), .B(n71200), .C(
        n71270), .Y(n71202) );
  OA21x2_ASAP7_75t_SL U71919 ( .A1(n71365), .A2(n71212), .B(n71211), .Y(n71213) );
  NAND3xp33_ASAP7_75t_SL U71920 ( .A(n71268), .B(n59523), .C(n71236), .Y(
        n71214) );
  A2O1A1Ixp33_ASAP7_75t_SL U71921 ( .A1(n71215), .A2(n71214), .B(n71217), .C(
        n57211), .Y(n71216) );
  OA21x2_ASAP7_75t_SL U71922 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_37_), .A2(n71224), 
        .B(n59523), .Y(n71269) );
  XOR2xp5_ASAP7_75t_SL U71923 ( .A(n71226), .B(n71225), .Y(n71227) );
  NAND3xp33_ASAP7_75t_SL U71924 ( .A(n71255), .B(n59523), .C(n71303), .Y(
        n71241) );
  A2O1A1Ixp33_ASAP7_75t_SL U71925 ( .A1(n71238), .A2(n71268), .B(n71237), .C(
        n71269), .Y(n71254) );
  NAND3xp33_ASAP7_75t_SL U71926 ( .A(n71239), .B(n71269), .C(n71268), .Y(
        n71258) );
  XNOR2xp5_ASAP7_75t_SL U71927 ( .A(n71241), .B(n71240), .Y(n71242) );
  XNOR2xp5_ASAP7_75t_SL U71928 ( .A(n71260), .B(n71259), .Y(n71261) );
  NAND3xp33_ASAP7_75t_SL U71929 ( .A(n71269), .B(n71268), .C(n71267), .Y(
        n71274) );
  NAND4xp25_ASAP7_75t_SL U71930 ( .A(n71272), .B(n71271), .C(n71270), .D(
        n71303), .Y(n71273) );
  AO21x1_ASAP7_75t_SL U71931 ( .A1(n71303), .A2(n71301), .B(n71297), .Y(n71275) );
  A2O1A1Ixp33_ASAP7_75t_SL U71932 ( .A1(n71276), .A2(n71294), .B(n71275), .C(
        n71302), .Y(n71278) );
  A2O1A1Ixp33_ASAP7_75t_SL U71933 ( .A1(n71279), .A2(n71278), .B(n71277), .C(
        n57211), .Y(n71280) );
  OAI211xp5_ASAP7_75t_SL U71934 ( .A1(n71309), .A2(n71350), .B(n71325), .C(
        n57211), .Y(n71310) );
  OAI211xp5_ASAP7_75t_SL U71935 ( .A1(n71327), .A2(n71326), .B(n71388), .C(
        n57211), .Y(n71328) );
  A2O1A1Ixp33_ASAP7_75t_SL U71936 ( .A1(n58315), .A2(n71339), .B(n71338), .C(
        n71337), .Y(n71368) );
  XNOR2xp5_ASAP7_75t_SL U71937 ( .A(n71372), .B(n71392), .Y(n71341) );
  A2O1A1Ixp33_ASAP7_75t_SL U71938 ( .A1(n71350), .A2(n71349), .B(n71348), .C(
        n71347), .Y(n71351) );
  XOR2xp5_ASAP7_75t_SL U71939 ( .A(n71407), .B(n71360), .Y(n71361) );
  A2O1A1Ixp33_ASAP7_75t_SL U71940 ( .A1(n71372), .A2(n71392), .B(n71391), .C(
        n71383), .Y(n71373) );
  XNOR2xp5_ASAP7_75t_SL U71941 ( .A(n71374), .B(n71373), .Y(n71375) );
  NAND4xp25_ASAP7_75t_SL U71942 ( .A(n71387), .B(n71390), .C(n71386), .D(
        n71401), .Y(n71411) );
  O2A1O1Ixp5_ASAP7_75t_SL U71943 ( .A1(n71398), .A2(n71397), .B(n71401), .C(
        n71402), .Y(n71409) );
  OAI211xp5_ASAP7_75t_SL U71944 ( .A1(n71404), .A2(n71403), .B(n71402), .C(
        n71401), .Y(n71405) );
  O2A1O1Ixp5_ASAP7_75t_SL U71945 ( .A1(n71411), .A2(n71410), .B(n71409), .C(
        n71408), .Y(n71414) );
  NOR3xp33_ASAP7_75t_SL U71946 ( .A(n59699), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_mul_s_fract_o_47_), .C(n71414), 
        .Y(n71415) );
  OR2x2_ASAP7_75t_SL U71947 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_), 
        .Y(n71605) );
  OR2x2_ASAP7_75t_SL U71948 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_14_), 
        .Y(n71459) );
  OR2x2_ASAP7_75t_SL U71949 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_5_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_4_), 
        .Y(n71601) );
  NAND3xp33_ASAP7_75t_SL U71950 ( .A(n71428), .B(n71628), .C(n72316), .Y(
        n71419) );
  OR2x2_ASAP7_75t_SL U71951 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_22_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_), 
        .Y(n71464) );
  O2A1O1Ixp5_ASAP7_75t_SL U71952 ( .A1(n71420), .A2(n71573), .B(n72253), .C(
        n71464), .Y(n71422) );
  OR2x2_ASAP7_75t_SL U71953 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_27_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_28_), 
        .Y(n71586) );
  O2A1O1Ixp5_ASAP7_75t_SL U71954 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_26_), 
        .A2(n72212), .B(n72234), .C(n71425), .Y(n71426) );
  A2O1A1Ixp33_ASAP7_75t_SL U71955 ( .A1(n71540), .A2(n71430), .B(n71429), .C(
        n71506), .Y(n71431) );
  NOR3xp33_ASAP7_75t_SL U71956 ( .A(n71442), .B(n71432), .C(n71431), .Y(n71436) );
  OR2x2_ASAP7_75t_SL U71957 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_32_), 
        .Y(n71630) );
  OR2x2_ASAP7_75t_SL U71958 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_34_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_33_), 
        .Y(n71560) );
  OR2x2_ASAP7_75t_SL U71959 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_40_), 
        .Y(n71549) );
  NAND3xp33_ASAP7_75t_SL U71960 ( .A(n71574), .B(n71629), .C(n71627), .Y(
        n71541) );
  AO21x1_ASAP7_75t_SL U71961 ( .A1(n71436), .A2(n71600), .B(n71460), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n130) );
  OR2x2_ASAP7_75t_SL U71962 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_39_), 
        .Y(n71471) );
  NAND3xp33_ASAP7_75t_SL U71963 ( .A(n71581), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_), 
        .C(n71863), .Y(n71473) );
  A2O1A1Ixp33_ASAP7_75t_SL U71964 ( .A1(n71473), .A2(n71984), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_41_), 
        .C(n71995), .Y(n71443) );
  OAI211xp5_ASAP7_75t_SL U71965 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_8_), 
        .A2(n71476), .B(n71438), .C(n71461), .Y(n71439) );
  A2O1A1Ixp33_ASAP7_75t_SL U71966 ( .A1(n72311), .A2(n72313), .B(n71440), .C(
        n71439), .Y(n71441) );
  NAND3xp33_ASAP7_75t_SL U71967 ( .A(n71447), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_), 
        .C(n72311), .Y(n71448) );
  OAI211xp5_ASAP7_75t_SL U71968 ( .A1(n71474), .A2(n71450), .B(n71449), .C(
        n71448), .Y(n71451) );
  NOR3xp33_ASAP7_75t_SL U71969 ( .A(n71474), .B(n71455), .C(n72350), .Y(n71456) );
  A2O1A1Ixp33_ASAP7_75t_SL U71970 ( .A1(n72212), .A2(n72219), .B(n71481), .C(
        n58606), .Y(n71483) );
  AND2x2_ASAP7_75t_SL U71971 ( .A(n71493), .B(n71492), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n127) );
  NOR3xp33_ASAP7_75t_SL U71972 ( .A(n71496), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_38_), 
        .C(n71994), .Y(n71498) );
  A2O1A1Ixp33_ASAP7_75t_SL U71973 ( .A1(n71500), .A2(n71499), .B(n71498), .C(
        n71497), .Y(n71508) );
  O2A1O1Ixp5_ASAP7_75t_SL U71974 ( .A1(n72346), .A2(n71604), .B(n71503), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_0_), 
        .Y(n71504) );
  NAND3xp33_ASAP7_75t_SL U71975 ( .A(n71508), .B(n71507), .C(n71506), .Y(
        n71510) );
  AND2x2_ASAP7_75t_SL U71976 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_25_), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_25_), .Y(n71522) );
  OR2x2_ASAP7_75t_SL U71977 ( .A(or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_26_), 
        .B(or1200_cpu_or1200_fpu_fpu_intfloat_conv_opa_r_26_), .Y(n72641) );
  AO21x1_ASAP7_75t_SL U71978 ( .A1(n71524), .A2(n71523), .B(n71527), .Y(n12873) );
  AO21x1_ASAP7_75t_SL U71979 ( .A1(n71532), .A2(n71531), .B(n71537), .Y(n52546) );
  AO21x1_ASAP7_75t_SL U71980 ( .A1(n71535), .A2(n71534), .B(n71533), .Y(n52545) );
  XNOR2xp5_ASAP7_75t_SL U71981 ( .A(n72646), .B(n71539), .Y(n3266) );
  A2O1A1Ixp33_ASAP7_75t_SL U71982 ( .A1(n72132), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_33_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_35_), 
        .C(n72079), .Y(n71544) );
  NAND3xp33_ASAP7_75t_SL U71983 ( .A(n71631), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_31_), 
        .C(n72154), .Y(n71543) );
  A2O1A1Ixp33_ASAP7_75t_SL U71984 ( .A1(n72054), .A2(n71544), .B(n71584), .C(
        n71543), .Y(n71546) );
  NOR3xp33_ASAP7_75t_SL U71985 ( .A(n71552), .B(n71551), .C(n71550), .Y(n71553) );
  AO21x1_ASAP7_75t_SL U71986 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_16_), 
        .A2(n71556), .B(n71555), .Y(n71557) );
  O2A1O1Ixp5_ASAP7_75t_SL U71987 ( .A1(n71559), .A2(n71558), .B(n71622), .C(
        n71557), .Y(n71596) );
  NAND3xp33_ASAP7_75t_SL U71988 ( .A(n71563), .B(n71953), .C(n71562), .Y(
        n71564) );
  OAI211xp5_ASAP7_75t_SL U71989 ( .A1(n71576), .A2(n71619), .B(n71596), .C(
        n71575), .Y(n71577) );
  A2O1A1Ixp33_ASAP7_75t_SL U71990 ( .A1(n71599), .A2(n71578), .B(n71577), .C(
        n71950), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n134) );
  OR3x1_ASAP7_75t_SL U71991 ( .A(n71581), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_45_), 
        .C(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_46_), 
        .Y(n71582) );
  OAI31xp33_ASAP7_75t_SL U71992 ( .A1(n71584), .A2(n71583), .A3(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_37_), 
        .B(n71582), .Y(n71585) );
  OAI211xp5_ASAP7_75t_SL U71993 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_19_), 
        .A2(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_20_), .B(n71587), .C(n72307), .Y(n71594) );
  NAND3xp33_ASAP7_75t_SL U71994 ( .A(n71950), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_11_), 
        .C(n72311), .Y(n71590) );
  NAND4xp25_ASAP7_75t_SL U71995 ( .A(n71596), .B(n71595), .C(n71594), .D(
        n71593), .Y(n71597) );
  A2O1A1Ixp33_ASAP7_75t_SL U71996 ( .A1(n71599), .A2(n71598), .B(n71597), .C(
        n71950), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n133) );
  O2A1O1Ixp5_ASAP7_75t_SL U71997 ( .A1(n71869), .A2(n71604), .B(n71603), .C(
        n71602), .Y(n71623) );
  A2O1A1Ixp33_ASAP7_75t_SL U71998 ( .A1(n72309), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_21_), 
        .B(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_23_), 
        .C(n72253), .Y(n71614) );
  O2A1O1Ixp5_ASAP7_75t_SL U71999 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_29_), 
        .A2(n71610), .B(n71609), .C(n71608), .Y(n71611) );
  OAI211xp5_ASAP7_75t_SL U72000 ( .A1(n71614), .A2(n71613), .B(n71612), .C(
        n71611), .Y(n71615) );
  AO21x1_ASAP7_75t_SL U72001 ( .A1(n71623), .A2(n71622), .B(n71621), .Y(n71624) );
  OR3x1_ASAP7_75t_SL U72002 ( .A(n71635), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_15_), 
        .C(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_47_), 
        .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n137) );
  O2A1O1Ixp5_ASAP7_75t_SL U72003 ( .A1(n71694), .A2(n71667), .B(n71664), .C(
        n71673), .Y(n71698) );
  XNOR2xp5_ASAP7_75t_SL U72004 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_5_), .B(
        n71694), .Y(n71714) );
  XNOR2xp5_ASAP7_75t_SL U72005 ( .A(n71643), .B(n71670), .Y(n71657) );
  XNOR2xp5_ASAP7_75t_SL U72006 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_zeros_2_), .B(
        n71657), .Y(n71728) );
  XNOR2xp5_ASAP7_75t_SL U72007 ( .A(n71677), .B(n71675), .Y(n71800) );
  A2O1A1Ixp33_ASAP7_75t_SL U72008 ( .A1(n71694), .A2(n71667), .B(n71666), .C(
        n71665), .Y(n71668) );
  XNOR2xp5_ASAP7_75t_SL U72009 ( .A(n71716), .B(n71680), .Y(n71795) );
  AO21x1_ASAP7_75t_SL U72010 ( .A1(n71736), .A2(n71737), .B(n71735), .Y(n71741) );
  A2O1A1Ixp33_ASAP7_75t_SL U72011 ( .A1(n71719), .A2(n71718), .B(n71717), .C(
        n71796), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n113) );
  AND2x2_ASAP7_75t_SL U72012 ( .A(n71702), .B(n71691), .Y(n71704) );
  O2A1O1Ixp5_ASAP7_75t_SL U72013 ( .A1(n71695), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_exp_10_i_5_), .B(
        n71694), .C(n71693), .Y(n71696) );
  A2O1A1Ixp33_ASAP7_75t_SL U72014 ( .A1(n71700), .A2(n71699), .B(n71704), .C(
        n71710), .Y(n71701) );
  A2O1A1Ixp33_ASAP7_75t_SL U72015 ( .A1(n71707), .A2(n71706), .B(n71705), .C(
        n71710), .Y(n71708) );
  OAI31xp33_ASAP7_75t_SL U72016 ( .A1(n71719), .A2(n71800), .A3(n71718), .B(
        n71717), .Y(n71794) );
  XNOR2xp5_ASAP7_75t_SL U72017 ( .A(n71728), .B(n71727), .Y(n71729) );
  NAND3xp33_ASAP7_75t_SL U72018 ( .A(n71737), .B(n71736), .C(n71735), .Y(
        n71740) );
  OR2x2_ASAP7_75t_SL U72019 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .B(
        n72241), .Y(n71772) );
  A2O1A1Ixp33_ASAP7_75t_SL U72020 ( .A1(n71764), .A2(n71763), .B(n72122), .C(
        n71762), .Y(n71767) );
  OR2x2_ASAP7_75t_SL U72021 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .Y(
        n72437) );
  O2A1O1Ixp5_ASAP7_75t_SL U72022 ( .A1(n72175), .A2(n72149), .B(n71769), .C(
        n72127), .Y(n71784) );
  OAI211xp5_ASAP7_75t_SL U72023 ( .A1(n57208), .A2(n72360), .B(n71774), .C(
        n71773), .Y(n72061) );
  O2A1O1Ixp5_ASAP7_75t_SL U72024 ( .A1(n72027), .A2(n72146), .B(n71776), .C(
        n72207), .Y(n71783) );
  OR3x1_ASAP7_75t_SL U72025 ( .A(n71784), .B(n71783), .C(n71782), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_N2648) );
  OAI211xp5_ASAP7_75t_SL U72026 ( .A1(n72263), .A2(n57208), .B(n71804), .C(
        n71803), .Y(n72039) );
  NAND3xp33_ASAP7_75t_SL U72027 ( .A(n71813), .B(n71812), .C(n71811), .Y(
        n72038) );
  A2O1A1Ixp33_ASAP7_75t_SL U72028 ( .A1(n71827), .A2(n71826), .B(n72122), .C(
        n71825), .Y(n71828) );
  OR2x2_ASAP7_75t_SL U72029 ( .A(n72104), .B(n72393), .Y(n71906) );
  A2O1A1Ixp33_ASAP7_75t_SL U72030 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .A2(
        n72305), .B(n71831), .C(n71906), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n105) );
  OAI211xp5_ASAP7_75t_SL U72031 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .A2(n57208), .B(n71833), .C(n71832), .Y(n72087) );
  NOR3xp33_ASAP7_75t_SL U72032 ( .A(n71882), .B(n71883), .C(n71899), .Y(n71846) );
  A2O1A1Ixp33_ASAP7_75t_SL U72033 ( .A1(n71855), .A2(n71854), .B(n72122), .C(
        n71853), .Y(n71862) );
  NOR3xp33_ASAP7_75t_SL U72034 ( .A(n72127), .B(n71862), .C(n71861), .Y(n71865) );
  O2A1O1Ixp5_ASAP7_75t_SL U72035 ( .A1(n72175), .A2(n72158), .B(n71865), .C(
        n71864), .Y(n71866) );
  OAI211xp5_ASAP7_75t_SL U72036 ( .A1(n71983), .A2(n72446), .B(n71908), .C(
        n71866), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n103) );
  A2O1A1Ixp33_ASAP7_75t_SL U72037 ( .A1(n71877), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_1_), .B(
        n71876), .C(n71875), .Y(n72017) );
  OAI211xp5_ASAP7_75t_SL U72038 ( .A1(n57208), .A2(n72346), .B(n71879), .C(
        n71878), .Y(n72109) );
  O2A1O1Ixp5_ASAP7_75t_SL U72039 ( .A1(n71887), .A2(n71886), .B(n71885), .C(
        n71884), .Y(n72108) );
  O2A1O1Ixp5_ASAP7_75t_SL U72040 ( .A1(n71893), .A2(n71892), .B(n72095), .C(
        n71891), .Y(n71902) );
  A2O1A1Ixp33_ASAP7_75t_SL U72041 ( .A1(n57207), .A2(n72005), .B(n71897), .C(
        n71896), .Y(n71966) );
  NAND4xp25_ASAP7_75t_SL U72042 ( .A(n71902), .B(n72104), .C(n71901), .D(
        n71900), .Y(n71903) );
  A2O1A1Ixp33_ASAP7_75t_SL U72043 ( .A1(n71908), .A2(n71907), .B(n71906), .C(
        n71905), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n102) );
  OAI211xp5_ASAP7_75t_SL U72044 ( .A1(n72046), .A2(n72355), .B(n71910), .C(
        n71909), .Y(n72182) );
  NAND3xp33_ASAP7_75t_SL U72045 ( .A(n71915), .B(n71914), .C(n72104), .Y(
        n71922) );
  OAI211xp5_ASAP7_75t_SL U72046 ( .A1(n71952), .A2(n57125), .B(n71918), .C(
        n57123), .Y(n71919) );
  A2O1A1Ixp33_ASAP7_75t_SL U72047 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .A2(
        n72182), .B(n71922), .C(n71921), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n101) );
  NAND4xp25_ASAP7_75t_SL U72048 ( .A(n71930), .B(n72104), .C(n71929), .D(
        n71928), .Y(n71941) );
  O2A1O1Ixp5_ASAP7_75t_SL U72049 ( .A1(n71935), .A2(n71934), .B(n71933), .C(
        n71932), .Y(n72140) );
  A2O1A1Ixp33_ASAP7_75t_SL U72050 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .A2(
        n72195), .B(n71941), .C(n71940), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n100) );
  NAND3xp33_ASAP7_75t_SL U72051 ( .A(n71949), .B(n72104), .C(n71948), .Y(
        n71961) );
  A2O1A1Ixp33_ASAP7_75t_SL U72052 ( .A1(n71956), .A2(n72399), .B(n59625), .C(
        n72077), .Y(n72329) );
  OR2x2_ASAP7_75t_SL U72053 ( .A(n71958), .B(n71957), .Y(n72330) );
  A2O1A1Ixp33_ASAP7_75t_SL U72054 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .A2(
        n72206), .B(n71961), .C(n71960), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n99) );
  NAND4xp25_ASAP7_75t_SL U72055 ( .A(n71969), .B(n72104), .C(n71968), .D(
        n71967), .Y(n71978) );
  NAND3xp33_ASAP7_75t_SL U72056 ( .A(n71972), .B(n71971), .C(n71970), .Y(
        n72398) );
  A2O1A1Ixp33_ASAP7_75t_SL U72057 ( .A1(n72399), .A2(n72398), .B(n72417), .C(
        n72407), .Y(n72471) );
  OAI211xp5_ASAP7_75t_SL U72058 ( .A1(n72113), .A2(n72147), .B(n71975), .C(
        n71974), .Y(n72210) );
  A2O1A1Ixp33_ASAP7_75t_SL U72059 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_4_), .A2(
        n72208), .B(n71978), .C(n71977), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n98) );
  AOI222xp33_ASAP7_75t_SL U72060 ( .A1(n72038), .A2(n72116), .B1(n72040), .B2(
        n72062), .C1(n72041), .C2(n72110), .Y(n72223) );
  A2O1A1Ixp33_ASAP7_75t_SL U72061 ( .A1(n72223), .A2(n72222), .B(n72175), .C(
        n71982), .Y(n71989) );
  A2O1A1Ixp33_ASAP7_75t_SL U72062 ( .A1(n71989), .A2(n72207), .B(n71988), .C(
        n71987), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n97) );
  OAI222xp33_ASAP7_75t_SL U72063 ( .A1(n59622), .A2(n72140), .B1(n59623), .B2(
        n72422), .C1(n59624), .C2(n72186), .Y(n72335) );
  A2O1A1Ixp33_ASAP7_75t_SL U72064 ( .A1(n71999), .A2(n71998), .B(n57192), .C(
        n71997), .Y(n72001) );
  A2O1A1Ixp33_ASAP7_75t_SL U72065 ( .A1(n72412), .A2(n72002), .B(n72001), .C(
        n72000), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n96) );
  OAI222xp33_ASAP7_75t_SL U72066 ( .A1(n59622), .A2(n72153), .B1(n59623), .B2(
        n72440), .C1(n59624), .C2(n72200), .Y(n72498) );
  A2O1A1Ixp33_ASAP7_75t_SL U72067 ( .A1(n72012), .A2(n72011), .B(n57192), .C(
        n72010), .Y(n72013) );
  A2O1A1Ixp33_ASAP7_75t_SL U72068 ( .A1(n72275), .A2(n72274), .B(n72382), .C(
        n72014), .Y(n72015) );
  A2O1A1Ixp33_ASAP7_75t_SL U72069 ( .A1(n72016), .A2(n72175), .B(n72207), .C(
        n72015), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n95) );
  OAI211xp5_ASAP7_75t_SL U72070 ( .A1(n72108), .A2(n72147), .B(n72019), .C(
        n72018), .Y(n72380) );
  OAI211xp5_ASAP7_75t_SL U72071 ( .A1(n72054), .A2(n57125), .B(n72022), .C(
        n72021), .Y(n72213) );
  O2A1O1Ixp5_ASAP7_75t_SL U72072 ( .A1(n72027), .A2(n72120), .B(n72026), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .Y(
        n72030) );
  OAI211xp5_ASAP7_75t_SL U72073 ( .A1(n72119), .A2(n72103), .B(n72028), .C(
        n58599), .Y(n72029) );
  OAI211xp5_ASAP7_75t_SL U72074 ( .A1(n72382), .A2(n72380), .B(n72032), .C(
        n72031), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n94) );
  OAI211xp5_ASAP7_75t_SL U72075 ( .A1(n72050), .A2(n72122), .B(n72049), .C(
        n72048), .Y(n72051) );
  OR2x2_ASAP7_75t_SL U72076 ( .A(n72058), .B(n72057), .Y(n72290) );
  AO21x1_ASAP7_75t_SL U72077 ( .A1(n72095), .A2(n72069), .B(n57192), .Y(n72070) );
  NAND3xp33_ASAP7_75t_SL U72078 ( .A(n72285), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shl2_5_), .C(
        n72095), .Y(n72073) );
  A2O1A1Ixp33_ASAP7_75t_SL U72079 ( .A1(n72075), .A2(n72074), .B(n72242), .C(
        n72073), .Y(n72076) );
  A2O1A1Ixp33_ASAP7_75t_SL U72080 ( .A1(n72510), .A2(n72290), .B(n58599), .C(
        n72076), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n92) );
  O2A1O1Ixp5_ASAP7_75t_SL U72081 ( .A1(n72175), .A2(n72392), .B(n58615), .C(
        n72127), .Y(n72098) );
  A2O1A1Ixp33_ASAP7_75t_SL U72082 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .A2(
        n72398), .B(n72534), .C(n72407), .Y(n72102) );
  OAI211xp5_ASAP7_75t_SL U72083 ( .A1(n72141), .A2(n57125), .B(n72101), .C(
        n72100), .Y(n72374) );
  NAND3xp33_ASAP7_75t_SL U72084 ( .A(n72102), .B(n72403), .C(n72402), .Y(
        n72369) );
  O2A1O1Ixp5_ASAP7_75t_SL U72085 ( .A1(n72175), .A2(n72397), .B(n72128), .C(
        n72127), .Y(n72129) );
  OAI211xp5_ASAP7_75t_SL U72086 ( .A1(n72382), .A2(n72305), .B(n72139), .C(
        n72138), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n89) );
  OAI222xp33_ASAP7_75t_SL U72087 ( .A1(n59622), .A2(n72235), .B1(n59623), .B2(
        n72186), .C1(n72434), .C2(n72140), .Y(n72424) );
  OR2x2_ASAP7_75t_SL U72088 ( .A(n59624), .B(n72245), .Y(n72421) );
  OAI211xp5_ASAP7_75t_SL U72089 ( .A1(n72147), .A2(n72146), .B(n72145), .C(
        n58599), .Y(n72148) );
  OAI211xp5_ASAP7_75t_SL U72090 ( .A1(n72424), .A2(n72152), .B(n72151), .C(
        n72150), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n88) );
  OAI222xp33_ASAP7_75t_SL U72091 ( .A1(n59622), .A2(n72270), .B1(n59623), .B2(
        n72200), .C1(n72434), .C2(n72153), .Y(n72444) );
  NOR3xp33_ASAP7_75t_SL U72092 ( .A(n72444), .B(n72445), .C(n72278), .Y(n72157) );
  OAI211xp5_ASAP7_75t_SL U72093 ( .A1(n72175), .A2(n72446), .B(n72160), .C(
        n72159), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n87) );
  NOR3xp33_ASAP7_75t_SL U72094 ( .A(n72170), .B(n72169), .C(n72415), .Y(n72171) );
  OAI211xp5_ASAP7_75t_SL U72095 ( .A1(n72175), .A2(n72326), .B(n72174), .C(
        n72173), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n86) );
  O2A1O1Ixp5_ASAP7_75t_SL U72096 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_2_), .A2(
        n72228), .B(n72176), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .Y(
        n72456) );
  OR2x2_ASAP7_75t_SL U72097 ( .A(n72179), .B(n72178), .Y(n72338) );
  OR2x2_ASAP7_75t_SL U72098 ( .A(n72181), .B(n72180), .Y(n72462) );
  OAI211xp5_ASAP7_75t_SL U72099 ( .A1(n72456), .A2(n72544), .B(n72185), .C(
        n72184), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n85) );
  OR2x2_ASAP7_75t_SL U72100 ( .A(n72188), .B(n72187), .Y(n72418) );
  OAI211xp5_ASAP7_75t_SL U72101 ( .A1(n72415), .A2(n72195), .B(n72194), .C(
        n72193), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n84) );
  OAI222xp33_ASAP7_75t_SL U72102 ( .A1(n59624), .A2(n72435), .B1(n59623), .B2(
        n72270), .C1(n72434), .C2(n72200), .Y(n72328) );
  OAI31xp33_ASAP7_75t_SL U72103 ( .A1(n72328), .A2(n72327), .A3(n72278), .B(
        n72381), .Y(n72201) );
  O2A1O1Ixp5_ASAP7_75t_SL U72104 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_3_), .A2(
        n72202), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_4_), .C(
        n72201), .Y(n72205) );
  OAI211xp5_ASAP7_75t_SL U72105 ( .A1(n72206), .A2(n72415), .B(n72205), .C(
        n72204), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n83) );
  OAI211xp5_ASAP7_75t_SL U72106 ( .A1(n72371), .A2(n59624), .B(n72214), .C(
        n57192), .Y(n72215) );
  OR2x2_ASAP7_75t_SL U72107 ( .A(n72544), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_shr2_5_), .Y(
        n72546) );
  NAND3xp33_ASAP7_75t_SL U72108 ( .A(n72209), .B(n72218), .C(n72217), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n82) );
  OAI222xp33_ASAP7_75t_SL U72109 ( .A1(n72338), .A2(n59622), .B1(n59623), .B2(
        n72337), .C1(n59624), .C2(n72453), .Y(n72477) );
  NOR3xp33_ASAP7_75t_SL U72110 ( .A(n72477), .B(n72478), .C(n72278), .Y(n72221) );
  NAND3xp33_ASAP7_75t_SL U72111 ( .A(n72223), .B(n72393), .C(n72222), .Y(
        n72230) );
  AO21x1_ASAP7_75t_SL U72112 ( .A1(n59625), .A2(n72226), .B(n72225), .Y(n72227) );
  NAND4xp25_ASAP7_75t_SL U72113 ( .A(n72231), .B(n72230), .C(n72381), .D(
        n72229), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n81) );
  OAI222xp33_ASAP7_75t_SL U72114 ( .A1(n72418), .A2(n59623), .B1(n72434), .B2(
        n72245), .C1(n59624), .C2(n72466), .Y(n72280) );
  OR2x2_ASAP7_75t_SL U72115 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_9_), 
        .B(n57203), .Y(n72332) );
  OR2x2_ASAP7_75t_SL U72116 ( .A(n72252), .B(n72251), .Y(n72493) );
  OR2x2_ASAP7_75t_SL U72117 ( .A(n72259), .B(n72258), .Y(n72489) );
  OR2x2_ASAP7_75t_SL U72118 ( .A(n72261), .B(n72260), .Y(n72491) );
  OAI222xp33_ASAP7_75t_SL U72119 ( .A1(n59624), .A2(n72432), .B1(n59623), .B2(
        n72271), .C1(n72434), .C2(n72270), .Y(n72496) );
  OAI31xp33_ASAP7_75t_SL U72120 ( .A1(n72496), .A2(n72497), .A3(n72278), .B(
        n72381), .Y(n72272) );
  NAND3xp33_ASAP7_75t_SL U72121 ( .A(n72275), .B(n72393), .C(n72274), .Y(
        n72276) );
  OAI211xp5_ASAP7_75t_SL U72122 ( .A1(n72510), .A2(n72498), .B(n72277), .C(
        n72276), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n79) );
  NOR3xp33_ASAP7_75t_SL U72123 ( .A(n72280), .B(n72279), .C(n72278), .Y(n72284) );
  NOR3xp33_ASAP7_75t_SL U72124 ( .A(n72282), .B(n72281), .C(n72415), .Y(n72283) );
  OAI211xp5_ASAP7_75t_SL U72125 ( .A1(n72510), .A2(n72290), .B(n72289), .C(
        n72288), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n76) );
  O2A1O1Ixp5_ASAP7_75t_SL U72126 ( .A1(n72297), .A2(n72296), .B(n72295), .C(
        n72294), .Y(n72452) );
  O2A1O1Ixp5_ASAP7_75t_SL U72127 ( .A1(n72301), .A2(n72300), .B(n72510), .C(
        n72299), .Y(n72302) );
  A2O1A1Ixp33_ASAP7_75t_SL U72128 ( .A1(n58599), .A2(n72305), .B(n72304), .C(
        n72426), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n73) );
  A2O1A1Ixp33_ASAP7_75t_SL U72129 ( .A1(n72516), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_fract_48_i_12_), 
        .B(n72353), .C(n72352), .Y(n72481) );
  OAI211xp5_ASAP7_75t_SL U72130 ( .A1(n72360), .A2(n57125), .B(n72359), .C(
        n72358), .Y(n72501) );
  OR2x2_ASAP7_75t_SL U72131 ( .A(n59624), .B(n72472), .Y(n72511) );
  OAI211xp5_ASAP7_75t_SL U72132 ( .A1(n72415), .A2(n72380), .B(n72379), .C(
        n72378), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n78) );
  OAI211xp5_ASAP7_75t_SL U72133 ( .A1(n72544), .A2(n72396), .B(n72395), .C(
        n72394), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n75) );
  A2O1A1Ixp33_ASAP7_75t_SL U72134 ( .A1(n72408), .A2(n72407), .B(n72406), .C(
        n72405), .Y(n72409) );
  O2A1O1Ixp5_ASAP7_75t_SL U72135 ( .A1(n72425), .A2(n72424), .B(n72443), .C(
        n72423), .Y(n72428) );
  O2A1O1Ixp5_ASAP7_75t_SL U72136 ( .A1(n72429), .A2(n72495), .B(n72428), .C(
        n72427), .Y(n72430) );
  O2A1O1Ixp5_ASAP7_75t_SL U72137 ( .A1(n72445), .A2(n72444), .B(n72443), .C(
        n72442), .Y(n72448) );
  O2A1O1Ixp5_ASAP7_75t_SL U72138 ( .A1(n72449), .A2(n72495), .B(n72448), .C(
        n72447), .Y(n72450) );
  OAI211xp5_ASAP7_75t_SL U72139 ( .A1(n72482), .A2(n72481), .B(n72455), .C(
        n72500), .Y(n72461) );
  A2O1A1Ixp33_ASAP7_75t_SL U72140 ( .A1(n72495), .A2(n72462), .B(n72461), .C(
        n72460), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n69) );
  O2A1O1Ixp5_ASAP7_75t_SL U72141 ( .A1(n59527), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_0_), .B(
        n57125), .C(n74265), .Y(n72522) );
  O2A1O1Ixp5_ASAP7_75t_SL U72142 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_0_), .A2(
        n72519), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_1_), .C(
        n72518), .Y(n72520) );
  O2A1O1Ixp5_ASAP7_75t_SL U72143 ( .A1(n72523), .A2(n72522), .B(n72521), .C(
        n72520), .Y(n72542) );
  NOR3xp33_ASAP7_75t_SL U72144 ( .A(n72536), .B(n72535), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_3_), .Y(
        n72537) );
  A2O1A1Ixp33_ASAP7_75t_SL U72145 ( .A1(n72542), .A2(n72541), .B(n72540), .C(
        n72539), .Y(n74293) );
  NAND4xp25_ASAP7_75t_SL U72146 ( .A(n72553), .B(n72552), .C(n72551), .D(
        n72550), .Y(n72556) );
  OR4x1_ASAP7_75t_SL U72147 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_3_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_6_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_9_), .Y(
        n72555) );
  OR4x1_ASAP7_75t_SL U72148 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_12_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_15_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_18_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_21_), .Y(
        n72554) );
  OR3x1_ASAP7_75t_SL U72149 ( .A(n72556), .B(n72555), .C(n72554), .Y(n72557)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72150 ( .A1(n74293), .A2(n74292), .B(n72559), .C(
        n58550), .Y(n72560) );
  OR2x2_ASAP7_75t_SL U72151 ( .A(n72561), .B(n74332), .Y(n74343) );
  XNOR2xp5_ASAP7_75t_SL U72152 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac2a_47_), .B(
        n74465), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n57) );
  NAND4xp25_ASAP7_75t_SL U72153 ( .A(n72567), .B(n72566), .C(n72565), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_r_zeros_4_), .Y(
        n74064) );
  NAND4xp25_ASAP7_75t_SL U72154 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_5_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_6_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_7_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expa_2_), .Y(
        n72570) );
  NOR3xp33_ASAP7_75t_SL U72155 ( .A(n72570), .B(n72569), .C(n72568), .Y(n74491) );
  NAND3xp33_ASAP7_75t_SL U72156 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_1_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_4_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expb_7_), .Y(
        n72571) );
  OR2x2_ASAP7_75t_SL U72157 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39), .B(n72576), .Y(n74062) );
  O2A1O1Ixp5_ASAP7_75t_SL U72158 ( .A1(n72579), .A2(n74062), .B(n72578), .C(
        n72577), .Y(n72596) );
  O2A1O1Ixp5_ASAP7_75t_SL U72159 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_4_), .A2(
        n72582), .B(n72595), .C(n72581), .Y(n72589) );
  XNOR2xp5_ASAP7_75t_SL U72160 ( .A(n72589), .B(n74245), .Y(n74246) );
  XOR2xp5_ASAP7_75t_SL U72161 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39), .Y(n74264) );
  NAND4xp25_ASAP7_75t_SL U72162 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_2_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_1_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_expo1_6_), .D(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_frac_rnd_24_), .Y(
        n72586) );
  NOR3xp33_ASAP7_75t_SL U72163 ( .A(n72591), .B(n74230), .C(n72590), .Y(n72592) );
  A2O1A1Ixp33_ASAP7_75t_SL U72164 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_s_opb_i_24_), .A2(n78375), .B(n72599), 
        .C(n72598), .Y(n72604) );
  A2O1A1Ixp33_ASAP7_75t_SL U72165 ( .A1(n72604), .A2(n72603), .B(n72602), .C(
        n72601), .Y(n72608) );
  A2O1A1Ixp33_ASAP7_75t_SL U72166 ( .A1(n72608), .A2(n58575), .B(n72607), .C(
        n72606), .Y(n72610) );
  XNOR2xp5_ASAP7_75t_SL U72167 ( .A(n72641), .B(n72642), .Y(n72628) );
  MAJIxp5_ASAP7_75t_SL U72168 ( .A(n72632), .B(n72631), .C(n72630), .Y(n72660)
         );
  NAND3xp33_ASAP7_75t_SL U72169 ( .A(n72663), .B(n72643), .C(n72654), .Y(
        n72644) );
  O2A1O1Ixp5_ASAP7_75t_SL U72170 ( .A1(n72651), .A2(n72650), .B(n72649), .C(
        n72648), .Y(n72652) );
  XNOR2xp5_ASAP7_75t_SL U72171 ( .A(n72654), .B(n72663), .Y(n72655) );
  A2O1A1Ixp33_ASAP7_75t_SL U72172 ( .A1(n72662), .A2(n72661), .B(n72660), .C(
        n72659), .Y(n72681) );
  MAJIxp5_ASAP7_75t_SL U72173 ( .A(n72681), .B(n72680), .C(n72679), .Y(n72678)
         );
  OA21x2_ASAP7_75t_SL U72174 ( .A1(n72676), .A2(n72678), .B(n72677), .Y(n72675) );
  AO21x1_ASAP7_75t_SL U72175 ( .A1(n72999), .A2(n72723), .B(n72687), .Y(n72751) );
  NAND3xp33_ASAP7_75t_SL U72176 ( .A(n72964), .B(n73030), .C(n72990), .Y(
        n72692) );
  AND2x2_ASAP7_75t_SL U72177 ( .A(n72695), .B(n72964), .Y(n73011) );
  AO21x1_ASAP7_75t_SL U72178 ( .A1(n72696), .A2(n57190), .B(n78243), .Y(n1568)
         );
  OAI222xp33_ASAP7_75t_SL U72179 ( .A1(n73010), .A2(n72886), .B1(n73009), .B2(
        n72900), .C1(n73008), .C2(n72888), .Y(n72699) );
  A2O1A1Ixp33_ASAP7_75t_SL U72180 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n72888), .B(n72702), .C(n72993), .Y(n72703) );
  NAND3xp33_ASAP7_75t_SL U72181 ( .A(n72723), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), .C(
        n72990), .Y(n72704) );
  OR2x2_ASAP7_75t_SL U72182 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .B(
        n72962), .Y(n72853) );
  A2O1A1Ixp33_ASAP7_75t_SL U72183 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_1_), 
        .A2(n72899), .B(n72744), .C(n72990), .Y(n72733) );
  A2O1A1Ixp33_ASAP7_75t_SL U72184 ( .A1(n72733), .A2(n73009), .B(n72732), .C(
        n72731), .Y(n72868) );
  A2O1A1Ixp33_ASAP7_75t_SL U72185 ( .A1(n72990), .A2(n72747), .B(n73042), .C(
        n72746), .Y(n72978) );
  NAND3xp33_ASAP7_75t_SL U72186 ( .A(n72751), .B(n72806), .C(n72990), .Y(
        n72761) );
  OAI211xp5_ASAP7_75t_SL U72187 ( .A1(n73008), .A2(n72907), .B(n72767), .C(
        n72766), .Y(n72986) );
  OAI211xp5_ASAP7_75t_SL U72188 ( .A1(n72986), .A2(n73002), .B(n72777), .C(
        n72776), .Y(n72778) );
  O2A1O1Ixp5_ASAP7_75t_SL U72189 ( .A1(n73020), .A2(n73017), .B(n72785), .C(
        n72784), .Y(n72786) );
  A2O1A1Ixp33_ASAP7_75t_SL U72190 ( .A1(n72791), .A2(n72790), .B(n73028), .C(
        n72789), .Y(n72835) );
  NAND3xp33_ASAP7_75t_SL U72191 ( .A(n72801), .B(n59629), .C(n72800), .Y(
        n72799) );
  NAND3xp33_ASAP7_75t_SL U72192 ( .A(n72801), .B(n59628), .C(n72800), .Y(
        n72802) );
  NAND3xp33_ASAP7_75t_SL U72193 ( .A(n72804), .B(n72803), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), .Y(
        n72805) );
  OR2x2_ASAP7_75t_SL U72194 ( .A(n72816), .B(n72847), .Y(n72817) );
  NAND3xp33_ASAP7_75t_SL U72195 ( .A(n72827), .B(n72826), .C(n72825), .Y(
        n72829) );
  OAI211xp5_ASAP7_75t_SL U72196 ( .A1(n73032), .A2(n72837), .B(n72836), .C(
        n72994), .Y(n72838) );
  AND2x2_ASAP7_75t_SL U72197 ( .A(n72845), .B(n72844), .Y(n73015) );
  OR2x2_ASAP7_75t_SL U72198 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .B(
        n72990), .Y(n72874) );
  A2O1A1Ixp33_ASAP7_75t_SL U72199 ( .A1(n72851), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_3_), .B(
        n72850), .C(n72849), .Y(n72852) );
  OAI31xp33_ASAP7_75t_SL U72200 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_2_), 
        .A2(n73015), .A3(n72853), .B(n72852), .Y(n72856) );
  O2A1O1Ixp5_ASAP7_75t_SL U72201 ( .A1(n73042), .A2(n72866), .B(n72865), .C(
        n72877), .Y(n72867) );
  A2O1A1Ixp33_ASAP7_75t_SL U72202 ( .A1(n73009), .A2(n72873), .B(n72872), .C(
        n72871), .Y(n73003) );
  A2O1A1Ixp33_ASAP7_75t_SL U72203 ( .A1(n72888), .A2(n72887), .B(n72928), .C(
        n72929), .Y(n72892) );
  A2O1A1Ixp33_ASAP7_75t_SL U72204 ( .A1(n72892), .A2(n72930), .B(n72932), .C(
        n72933), .Y(n72896) );
  A2O1A1Ixp33_ASAP7_75t_SL U72205 ( .A1(n72896), .A2(n72934), .B(n72895), .C(
        n72894), .Y(n72897) );
  A2O1A1Ixp33_ASAP7_75t_SL U72206 ( .A1(n72900), .A2(n72965), .B(n72899), .C(
        n72898), .Y(n72906) );
  A2O1A1Ixp33_ASAP7_75t_SL U72207 ( .A1(n72906), .A2(n72905), .B(n72904), .C(
        n72903), .Y(n72910) );
  A2O1A1Ixp33_ASAP7_75t_SL U72208 ( .A1(n72910), .A2(n72909), .B(n72908), .C(
        n72907), .Y(n72914) );
  A2O1A1Ixp33_ASAP7_75t_SL U72209 ( .A1(n72914), .A2(n72913), .B(n72912), .C(
        n72911), .Y(n72919) );
  A2O1A1Ixp33_ASAP7_75t_SL U72210 ( .A1(n72919), .A2(n72918), .B(n72937), .C(
        n72917), .Y(n72925) );
  A2O1A1Ixp33_ASAP7_75t_SL U72211 ( .A1(n72925), .A2(n72924), .B(n72923), .C(
        n72922), .Y(n72926) );
  A2O1A1Ixp33_ASAP7_75t_SL U72212 ( .A1(n73029), .A2(n72999), .B(n72927), .C(
        n72926), .Y(n72960) );
  A2O1A1Ixp33_ASAP7_75t_SL U72213 ( .A1(n72944), .A2(n72943), .B(n72945), .C(
        n72946), .Y(n72942) );
  NAND3xp33_ASAP7_75t_SL U72214 ( .A(n72942), .B(n72941), .C(n72947), .Y(
        n72951) );
  NAND3xp33_ASAP7_75t_SL U72215 ( .A(n73027), .B(n73029), .C(n73023), .Y(
        n72949) );
  A2O1A1Ixp33_ASAP7_75t_SL U72216 ( .A1(n73023), .A2(n72951), .B(n72990), .C(
        n72950), .Y(n72958) );
  A2O1A1Ixp33_ASAP7_75t_SL U72217 ( .A1(n72960), .A2(n72959), .B(n72958), .C(
        n72957), .Y(n72984) );
  NAND3xp33_ASAP7_75t_SL U72218 ( .A(n72971), .B(n72987), .C(n72990), .Y(
        n72972) );
  A2O1A1Ixp33_ASAP7_75t_SL U72219 ( .A1(n73026), .A2(n72992), .B(n73032), .C(
        n72972), .Y(n72973) );
  NOR3xp33_ASAP7_75t_SL U72220 ( .A(n72975), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_), .C(
        n72990), .Y(n72977) );
  A2O1A1Ixp33_ASAP7_75t_SL U72221 ( .A1(n72978), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_prenorm_addsub_s_exp_diff_4_), .B(
        n72977), .C(n72976), .Y(n72979) );
  A2O1A1Ixp33_ASAP7_75t_SL U72222 ( .A1(n72984), .A2(n72983), .B(n72982), .C(
        n72981), .Y(n72985) );
  A2O1A1Ixp33_ASAP7_75t_SL U72223 ( .A1(n72990), .A2(n72989), .B(n72988), .C(
        n72987), .Y(n73001) );
  O2A1O1Ixp5_ASAP7_75t_SL U72224 ( .A1(n72999), .A2(n72998), .B(n73007), .C(
        n72997), .Y(n73000) );
  OAI211xp5_ASAP7_75t_SL U72225 ( .A1(n73003), .A2(n73002), .B(n73001), .C(
        n73000), .Y(n73004) );
  AO21x1_ASAP7_75t_SL U72226 ( .A1(n73037), .A2(n73015), .B(n73014), .Y(n73019) );
  A2O1A1Ixp33_ASAP7_75t_SL U72227 ( .A1(n73034), .A2(n73033), .B(n73032), .C(
        n73031), .Y(n73035) );
  O2A1O1Ixp5_ASAP7_75t_SL U72228 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[1]), .A2(
        n73227), .B(n73483), .C(n73048), .Y(n73062) );
  NOR3xp33_ASAP7_75t_SL U72229 ( .A(n73056), .B(n73051), .C(n73050), .Y(n73060) );
  NAND3xp33_ASAP7_75t_SL U72230 ( .A(n73053), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[4]), .C(
        n73219), .Y(n73057) );
  A2O1A1Ixp33_ASAP7_75t_SL U72231 ( .A1(n73058), .A2(n73057), .B(n73056), .C(
        n73055), .Y(n73059) );
  O2A1O1Ixp5_ASAP7_75t_SL U72232 ( .A1(n73062), .A2(n73061), .B(n73060), .C(
        n73059), .Y(n73069) );
  A2O1A1Ixp33_ASAP7_75t_SL U72233 ( .A1(n73067), .A2(n73066), .B(n73075), .C(
        n73065), .Y(n73070) );
  A2O1A1Ixp33_ASAP7_75t_SL U72234 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[8]), .A2(
        n73211), .B(n73069), .C(n73068), .Y(n73099) );
  O2A1O1Ixp5_ASAP7_75t_SL U72235 ( .A1(n73075), .A2(n73074), .B(n73073), .C(
        n73072), .Y(n73098) );
  A2O1A1Ixp33_ASAP7_75t_SL U72236 ( .A1(n73080), .A2(n73090), .B(n73079), .C(
        n73089), .Y(n73094) );
  NAND3xp33_ASAP7_75t_SL U72237 ( .A(n73084), .B(n73082), .C(n73088), .Y(
        n73095) );
  NAND3xp33_ASAP7_75t_SL U72238 ( .A(n73084), .B(n73088), .C(n73083), .Y(
        n73093) );
  NAND4xp25_ASAP7_75t_SL U72239 ( .A(n73091), .B(n73090), .C(n73089), .D(
        n73088), .Y(n73092) );
  OAI211xp5_ASAP7_75t_SL U72240 ( .A1(n73095), .A2(n73094), .B(n73093), .C(
        n73092), .Y(n73096) );
  A2O1A1Ixp33_ASAP7_75t_SL U72241 ( .A1(n73099), .A2(n73098), .B(n73097), .C(
        n73096), .Y(n73109) );
  O2A1O1Ixp5_ASAP7_75t_SL U72242 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[23]), .A2(
        n73341), .B(n73102), .C(n73101), .Y(n73108) );
  OAI211xp5_ASAP7_75t_SL U72243 ( .A1(n73105), .A2(n73104), .B(n73372), .C(
        n73383), .Y(n73107) );
  A2O1A1Ixp33_ASAP7_75t_SL U72244 ( .A1(n73109), .A2(n73108), .B(n73107), .C(
        n73106), .Y(n73853) );
  A2O1A1Ixp33_ASAP7_75t_SL U72245 ( .A1(n73111), .A2(n74502), .B(n73110), .C(
        n73115), .Y(n73116) );
  O2A1O1Ixp5_ASAP7_75t_SL U72246 ( .A1(n73119), .A2(n57185), .B(n73118), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[21]), .Y(
        n73120) );
  O2A1O1Ixp5_ASAP7_75t_SL U72247 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[21]), .A2(
        n59630), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[21]), .C(
        n73120), .Y(n73121) );
  O2A1O1Ixp5_ASAP7_75t_SL U72248 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[20]), .A2(
        n59631), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[20]), .C(
        n73124), .Y(n73125) );
  A2O1A1Ixp33_ASAP7_75t_SL U72249 ( .A1(n58284), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[16]), .B(
        n73126), .C(n73128), .Y(n73127) );
  A2O1A1Ixp33_ASAP7_75t_SL U72250 ( .A1(n73382), .A2(n73129), .B(n73128), .C(
        n73127), .Y(n73131) );
  NAND3xp33_ASAP7_75t_SL U72251 ( .A(n73292), .B(n73294), .C(n73293), .Y(
        n73130) );
  A2O1A1Ixp33_ASAP7_75t_SL U72252 ( .A1(n73298), .A2(n73136), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[17]), .C(
        n73135), .Y(n73137) );
  A2O1A1Ixp33_ASAP7_75t_SL U72253 ( .A1(n58284), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[14]), .B(
        n73138), .C(n73140), .Y(n73139) );
  A2O1A1Ixp33_ASAP7_75t_SL U72254 ( .A1(n73382), .A2(n73141), .B(n73140), .C(
        n73139), .Y(n73143) );
  NAND3xp33_ASAP7_75t_SL U72255 ( .A(n73280), .B(n73282), .C(n73281), .Y(
        n73142) );
  O2A1O1Ixp5_ASAP7_75t_SL U72256 ( .A1(n73152), .A2(n73151), .B(n73150), .C(
        n73149), .Y(n73153) );
  O2A1O1Ixp5_ASAP7_75t_SL U72257 ( .A1(n57185), .A2(n73159), .B(n73158), .C(
        n73157), .Y(n73458) );
  A2O1A1Ixp33_ASAP7_75t_SL U72258 ( .A1(n73174), .A2(n73173), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[11]), .C(
        n73172), .Y(n73175) );
  A2O1A1Ixp33_ASAP7_75t_SL U72259 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[8]), .A2(
        n58284), .B(n73197), .C(n73207), .Y(n73200) );
  O2A1O1Ixp5_ASAP7_75t_SL U72260 ( .A1(n73213), .A2(n73212), .B(n73211), .C(
        n73210), .Y(n73459) );
  NAND3xp33_ASAP7_75t_SL U72261 ( .A(n73419), .B(n73418), .C(n73450), .Y(
        n73271) );
  O2A1O1Ixp5_ASAP7_75t_SL U72262 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[5]), .A2(
        n59525), .B(n73223), .C(n73259), .Y(n73224) );
  XNOR2xp5_ASAP7_75t_SL U72263 ( .A(n73235), .B(n73234), .Y(n73481) );
  XNOR2xp5_ASAP7_75t_SL U72264 ( .A(n73268), .B(n73266), .Y(n73452) );
  A2O1A1Ixp33_ASAP7_75t_SL U72265 ( .A1(n73278), .A2(n73277), .B(n73276), .C(
        n73275), .Y(n73413) );
  A2O1A1Ixp33_ASAP7_75t_SL U72266 ( .A1(n73287), .A2(n73286), .B(n73285), .C(
        n73284), .Y(n73288) );
  A2O1A1Ixp33_ASAP7_75t_SL U72267 ( .A1(n73299), .A2(n73298), .B(n73297), .C(
        n73296), .Y(n73300) );
  O2A1O1Ixp5_ASAP7_75t_SL U72268 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[19]), .A2(
        n59630), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[19]), .C(
        n73305), .Y(n73306) );
  A2O1A1Ixp33_ASAP7_75t_SL U72269 ( .A1(n73320), .A2(n73319), .B(n73318), .C(
        n73317), .Y(n73321) );
  O2A1O1Ixp5_ASAP7_75t_SL U72270 ( .A1(n73333), .A2(n57185), .B(n73332), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[23]), .Y(
        n73334) );
  O2A1O1Ixp5_ASAP7_75t_SL U72271 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[23]), .A2(
        n59630), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[23]), .C(
        n73334), .Y(n73335) );
  A2O1A1Ixp33_ASAP7_75t_SL U72272 ( .A1(n73344), .A2(n73343), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[22]), .C(
        n73342), .Y(n73345) );
  A2O1A1Ixp33_ASAP7_75t_SL U72273 ( .A1(n73352), .A2(n73351), .B(n73350), .C(
        n73349), .Y(n73353) );
  OA21x2_ASAP7_75t_SL U72274 ( .A1(n73358), .A2(n73357), .B(n73405), .Y(n78222) );
  XOR2xp5_ASAP7_75t_SL U72275 ( .A(n73371), .B(n73370), .Y(n78219) );
  A2O1A1Ixp33_ASAP7_75t_SL U72276 ( .A1(n73375), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fractb_28_o[26]), .B(
        n73374), .C(n73376), .Y(n73378) );
  A2O1A1Ixp33_ASAP7_75t_SL U72277 ( .A1(n73392), .A2(n73386), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_fracta_28_o[25]), .C(
        n73385), .Y(n73387) );
  AO21x1_ASAP7_75t_SL U72278 ( .A1(n73403), .A2(n73402), .B(n73401), .Y(n53176) );
  XOR2xp5_ASAP7_75t_SL U72279 ( .A(n73408), .B(n73407), .Y(n78217) );
  XNOR2xp5_ASAP7_75t_SL U72280 ( .A(n73445), .B(n73444), .Y(n78211) );
  OA21x2_ASAP7_75t_SL U72281 ( .A1(n73448), .A2(n73447), .B(n73446), .Y(n78210) );
  XNOR2xp5_ASAP7_75t_SL U72282 ( .A(n73450), .B(n73449), .Y(n51955) );
  XNOR2xp5_ASAP7_75t_SL U72283 ( .A(n73465), .B(n73464), .Y(n53190) );
  OR2x2_ASAP7_75t_SL U72284 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[18]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[17]), .Y(n73498) );
  NAND3xp33_ASAP7_75t_SL U72285 ( .A(n73496), .B(n73521), .C(n73522), .Y(
        n73871) );
  A2O1A1Ixp33_ASAP7_75t_SL U72286 ( .A1(n73496), .A2(n73495), .B(n73494), .C(
        n73493), .Y(n73500) );
  A2O1A1Ixp33_ASAP7_75t_SL U72287 ( .A1(n73500), .A2(n73499), .B(n73498), .C(
        n73497), .Y(n73502) );
  OR2x2_ASAP7_75t_SL U72288 ( .A(n73503), .B(n73873), .Y(n73602) );
  NAND3xp33_ASAP7_75t_SL U72289 ( .A(n74733), .B(n73679), .C(n73828), .Y(
        n73506) );
  A2O1A1Ixp33_ASAP7_75t_SL U72290 ( .A1(n73507), .A2(n73506), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[5]), .C(n3331), .Y(
        n73513) );
  A2O1A1Ixp33_ASAP7_75t_SL U72291 ( .A1(n73633), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[8]), .B(n73695), .C(
        n73810), .Y(n73510) );
  A2O1A1Ixp33_ASAP7_75t_SL U72292 ( .A1(n73510), .A2(n73509), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[13]), .C(n73508), .Y(
        n73512) );
  A2O1A1Ixp33_ASAP7_75t_SL U72293 ( .A1(n73514), .A2(n73513), .B(n73512), .C(
        n73511), .Y(n73516) );
  A2O1A1Ixp33_ASAP7_75t_SL U72294 ( .A1(n73516), .A2(n73688), .B(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[19]), .C(n73515), .Y(
        n73518) );
  OR2x2_ASAP7_75t_SL U72295 ( .A(n73520), .B(n73874), .Y(n73606) );
  A2O1A1Ixp33_ASAP7_75t_SL U72296 ( .A1(n73568), .A2(n73538), .B(n73539), .C(
        n73544), .Y(n73550) );
  A2O1A1Ixp33_ASAP7_75t_SL U72297 ( .A1(n73547), .A2(n73593), .B(n73549), .C(
        n73546), .Y(n73557) );
  NAND3xp33_ASAP7_75t_SL U72298 ( .A(n73582), .B(n73553), .C(n73552), .Y(
        n73556) );
  NAND3xp33_ASAP7_75t_SL U72299 ( .A(n73561), .B(n73581), .C(n73560), .Y(
        n73586) );
  A2O1A1Ixp33_ASAP7_75t_SL U72300 ( .A1(n73565), .A2(n73563), .B(n73661), .C(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[6]), .Y(n73564)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72301 ( .A1(n73566), .A2(n73565), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[6]), .C(n73564), 
        .Y(n73567) );
  XNOR2xp5_ASAP7_75t_SL U72302 ( .A(n73657), .B(n73573), .Y(n73588) );
  AND2x2_ASAP7_75t_SL U72303 ( .A(n73575), .B(n73574), .Y(n73655) );
  XNOR2xp5_ASAP7_75t_SL U72304 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[0]), .B(n73579), 
        .Y(n73651) );
  OAI211xp5_ASAP7_75t_SL U72305 ( .A1(n73656), .A2(n73655), .B(n73584), .C(
        n73654), .Y(n73587) );
  O2A1O1Ixp5_ASAP7_75t_SL U72306 ( .A1(n73588), .A2(n73587), .B(n73586), .C(
        n73585), .Y(n73589) );
  OR2x2_ASAP7_75t_SL U72307 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[0]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[1]), .Y(n73597)
         );
  XNOR2xp5_ASAP7_75t_SL U72308 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_prenorm_addsub_exp_o[3]), .B(n73611), 
        .Y(n73592) );
  A2O1A1Ixp33_ASAP7_75t_SL U72309 ( .A1(n73652), .A2(n73597), .B(n73596), .C(
        n73595), .Y(n73598) );
  A2O1A1Ixp33_ASAP7_75t_SL U72310 ( .A1(n73610), .A2(n73600), .B(n73599), .C(
        n73598), .Y(n1526) );
  O2A1O1Ixp5_ASAP7_75t_SL U72311 ( .A1(n73605), .A2(n73604), .B(n73610), .C(
        n73603), .Y(n1527) );
  AOI222xp33_ASAP7_75t_SL U72312 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[21]), .A2(n57205), .B1(
        n59632), .B2(or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[19]), .C1(
        n57204), .C2(or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[20]), .Y(
        n73730) );
  A2O1A1Ixp33_ASAP7_75t_SL U72313 ( .A1(n73621), .A2(n73620), .B(n73689), .C(
        n3309), .Y(n73622) );
  OR2x2_ASAP7_75t_SL U72314 ( .A(n73752), .B(n73698), .Y(n73645) );
  AO21x1_ASAP7_75t_SL U72315 ( .A1(n73625), .A2(n73624), .B(n73752), .Y(n73626) );
  A2O1A1Ixp33_ASAP7_75t_SL U72316 ( .A1(n73811), .A2(n73797), .B(n73793), .C(
        n73627), .Y(n73628) );
  A2O1A1Ixp33_ASAP7_75t_SL U72317 ( .A1(n73631), .A2(n73630), .B(n73629), .C(
        n73628), .Y(n3308) );
  A2O1A1Ixp33_ASAP7_75t_SL U72318 ( .A1(n73644), .A2(n73643), .B(n73689), .C(
        n3309), .Y(n73648) );
  OAI222xp33_ASAP7_75t_SL U72319 ( .A1(n58400), .A2(n73753), .B1(n58423), .B2(
        n73728), .C1(n58622), .C2(n73767), .Y(n73715) );
  A2O1A1Ixp33_ASAP7_75t_SL U72320 ( .A1(n73809), .A2(n73618), .B(n73650), .C(
        n73649), .Y(n5349) );
  AOI222xp33_ASAP7_75t_SL U72321 ( .A1(n59632), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[18]), .B1(n57204), .B2(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[19]), .C1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[21]), .C2(n57217), .Y(
        n73745) );
  A2O1A1Ixp33_ASAP7_75t_SL U72322 ( .A1(n73665), .A2(n73664), .B(n73689), .C(
        n3309), .Y(n73666) );
  O2A1O1Ixp5_ASAP7_75t_SL U72323 ( .A1(n73736), .A2(n73737), .B(n73752), .C(
        n58623), .Y(n73812) );
  NAND3xp33_ASAP7_75t_SL U72324 ( .A(n73752), .B(n57217), .C(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[1]), .Y(n73673) );
  A2O1A1Ixp33_ASAP7_75t_SL U72325 ( .A1(n73812), .A2(n73797), .B(n73793), .C(
        n73674), .Y(n73675) );
  A2O1A1Ixp33_ASAP7_75t_SL U72326 ( .A1(n73678), .A2(n73677), .B(n73676), .C(
        n73675), .Y(n3307) );
  A2O1A1Ixp33_ASAP7_75t_SL U72327 ( .A1(n73694), .A2(n73693), .B(n73692), .C(
        n73691), .Y(n73701) );
  OR2x2_ASAP7_75t_SL U72328 ( .A(n59705), .B(n73698), .Y(n73770) );
  A2O1A1Ixp33_ASAP7_75t_SL U72329 ( .A1(n73815), .A2(n73618), .B(n73703), .C(
        n73702), .Y(n3306) );
  A2O1A1Ixp33_ASAP7_75t_SL U72330 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[3]), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .B(
        n73711), .C(n57217), .Y(n73712) );
  OAI211xp5_ASAP7_75t_SL U72331 ( .A1(n58619), .A2(n73725), .B(n3309), .C(
        n73712), .Y(n73713) );
  NAND3xp33_ASAP7_75t_SL U72332 ( .A(n73717), .B(n73786), .C(n73716), .Y(
        n73718) );
  NAND4xp25_ASAP7_75t_SL U72333 ( .A(n73721), .B(n73720), .C(n73719), .D(
        n73718), .Y(n3305) );
  NAND3xp33_ASAP7_75t_SL U72334 ( .A(n73730), .B(n73786), .C(n73729), .Y(
        n73732) );
  NAND3xp33_ASAP7_75t_SL U72335 ( .A(n73733), .B(n73732), .C(n73731), .Y(
        n73734) );
  NOR3xp33_ASAP7_75t_SL U72336 ( .A(n73737), .B(n73736), .C(n73752), .Y(n73738) );
  NAND3xp33_ASAP7_75t_SL U72337 ( .A(n73745), .B(n73786), .C(n73744), .Y(
        n73747) );
  NAND3xp33_ASAP7_75t_SL U72338 ( .A(n73748), .B(n73747), .C(n73746), .Y(
        n73749) );
  AND2x2_ASAP7_75t_SL U72339 ( .A(n3309), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[3]), .Y(
        n73814) );
  O2A1O1Ixp5_ASAP7_75t_SL U72340 ( .A1(n73833), .A2(n58400), .B(n73756), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_shl1[2]), .Y(
        n73757) );
  NAND4xp25_ASAP7_75t_SL U72341 ( .A(n73762), .B(n73761), .C(n73760), .D(
        n73759), .Y(n3302) );
  AND2x2_ASAP7_75t_SL U72342 ( .A(n3309), .B(n73808), .Y(n73827) );
  OAI211xp5_ASAP7_75t_SL U72343 ( .A1(n73809), .A2(n73770), .B(n73769), .C(
        n73768), .Y(n3301) );
  NAND3xp33_ASAP7_75t_SL U72344 ( .A(n73777), .B(n73776), .C(n73775), .Y(n3300) );
  NAND3xp33_ASAP7_75t_SL U72345 ( .A(n73784), .B(n73783), .C(n73782), .Y(n3299) );
  NOR3xp33_ASAP7_75t_SL U72346 ( .A(n73794), .B(n73793), .C(n73792), .Y(n73795) );
  NAND3xp33_ASAP7_75t_SL U72347 ( .A(n73800), .B(n73799), .C(n73798), .Y(n3297) );
  OR3x1_ASAP7_75t_SL U72348 ( .A(n73820), .B(n73819), .C(n73829), .Y(n3289) );
  OR3x1_ASAP7_75t_SL U72349 ( .A(n73822), .B(n73829), .C(n73821), .Y(n3288) );
  OR3x1_ASAP7_75t_SL U72350 ( .A(n73825), .B(n73829), .C(n73824), .Y(n3287) );
  A2O1A1Ixp33_ASAP7_75t_SL U72351 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_addsub_fract_o[1]), .A2(n59705), .B(
        n73832), .C(n73834), .Y(n3282) );
  NAND4xp25_ASAP7_75t_SL U72352 ( .A(n73837), .B(n78220), .C(n78210), .D(
        n78212), .Y(n73845) );
  AND3x1_ASAP7_75t_SL U72353 ( .A(n12827), .B(n73838), .C(n12864), .Y(n73839)
         );
  AND3x1_ASAP7_75t_SL U72354 ( .A(n78214), .B(n73842), .C(n78213), .Y(n73843)
         );
  NAND4xp25_ASAP7_75t_SL U72355 ( .A(n78221), .B(n73843), .C(n53189), .D(
        n78215), .Y(n73844) );
  NOR3xp33_ASAP7_75t_SL U72356 ( .A(n73846), .B(n73845), .C(n73844), .Y(n73847) );
  NAND3xp33_ASAP7_75t_SL U72357 ( .A(n73847), .B(n78217), .C(n78222), .Y(
        n73848) );
  NAND4xp25_ASAP7_75t_SL U72358 ( .A(n73850), .B(n73849), .C(n53176), .D(
        n78218), .Y(n73851) );
  A2O1A1Ixp33_ASAP7_75t_SL U72359 ( .A1(n73853), .A2(n76983), .B(n73852), .C(
        n73851), .Y(n2527) );
  NAND3xp33_ASAP7_75t_SL U72360 ( .A(n73861), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_26_), 
        .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_27_), 
        .Y(n73860) );
  NAND3xp33_ASAP7_75t_SL U72361 ( .A(n73856), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1[1]), .C(n73855), .Y(
        n74303) );
  OR2x2_ASAP7_75t_SL U72362 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_27_), 
        .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_26_), 
        .Y(n73866) );
  OR2x2_ASAP7_75t_SL U72363 ( .A(n73868), .B(n73867), .Y(n74066) );
  XNOR2xp5_ASAP7_75t_SL U72364 ( .A(n73881), .B(n73875), .Y(n73870) );
  OR2x2_ASAP7_75t_SL U72365 ( .A(n73884), .B(n73883), .Y(n74497) );
  NAND3xp33_ASAP7_75t_SL U72366 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[2]), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[4]), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_expo9_1[7]), .Y(
        n73894) );
  NOR3xp33_ASAP7_75t_SL U72367 ( .A(n73896), .B(n73895), .C(n73894), .Y(n73897) );
  NAND3xp33_ASAP7_75t_SL U72368 ( .A(n74247), .B(n74069), .C(n73897), .Y(
        n73899) );
  OR2x2_ASAP7_75t_SL U72369 ( .A(n76744), .B(n73907), .Y(n75268) );
  OAI211xp5_ASAP7_75t_SL U72370 ( .A1(or1200_cpu_or1200_except_n132), .A2(
        n57102), .B(n73911), .C(n73910), .Y(n73912) );
  NOR3xp33_ASAP7_75t_SL U72371 ( .A(n73914), .B(n73913), .C(n73912), .Y(n77666) );
  OR2x2_ASAP7_75t_SL U72372 ( .A(n75573), .B(n75587), .Y(n73931) );
  A2O1A1Ixp33_ASAP7_75t_SL U72373 ( .A1(n73918), .A2(n76342), .B(n75735), .C(
        n73917), .Y(n73919) );
  OAI211xp5_ASAP7_75t_SL U72374 ( .A1(n75590), .A2(n77078), .B(n73931), .C(
        n73930), .Y(n73932) );
  OAI211xp5_ASAP7_75t_SL U72375 ( .A1(n75268), .A2(n77666), .B(n75879), .C(
        n73934), .Y(n73935) );
  A2O1A1Ixp33_ASAP7_75t_SL U72376 ( .A1(n73945), .A2(n73944), .B(n73943), .C(
        n57126), .Y(n73946) );
  NAND3xp33_ASAP7_75t_SL U72377 ( .A(n73948), .B(n73947), .C(n73946), .Y(
        n75802) );
  A2O1A1Ixp33_ASAP7_75t_SL U72378 ( .A1(n77467), .A2(n73957), .B(n73956), .C(
        n73955), .Y(n9643) );
  O2A1O1Ixp5_ASAP7_75t_SL U72379 ( .A1(n75849), .A2(n76333), .B(n76343), .C(
        n75720), .Y(n76416) );
  A2O1A1Ixp33_ASAP7_75t_SL U72380 ( .A1(n73973), .A2(n59442), .B(n59183), .C(
        n73972), .Y(n73979) );
  A2O1A1Ixp33_ASAP7_75t_SL U72381 ( .A1(n73979), .A2(n76354), .B(n73978), .C(
        n73977), .Y(n73984) );
  A2O1A1Ixp33_ASAP7_75t_SL U72382 ( .A1(n73984), .A2(n73983), .B(n76357), .C(
        n73982), .Y(n74002) );
  A2O1A1Ixp33_ASAP7_75t_SL U72383 ( .A1(n73989), .A2(n76368), .B(n76384), .C(
        n73988), .Y(n73997) );
  A2O1A1Ixp33_ASAP7_75t_SL U72384 ( .A1(n73997), .A2(n73996), .B(n73995), .C(
        n73994), .Y(n74001) );
  NAND4xp25_ASAP7_75t_SL U72385 ( .A(n76452), .B(n74004), .C(n76449), .D(
        n73999), .Y(n76395) );
  A2O1A1Ixp33_ASAP7_75t_SL U72386 ( .A1(n74003), .A2(n74002), .B(n74001), .C(
        n74000), .Y(n74014) );
  O2A1O1Ixp5_ASAP7_75t_SL U72387 ( .A1(n74599), .A2(n74009), .B(n74598), .C(
        n76396), .Y(n74010) );
  A2O1A1Ixp33_ASAP7_75t_SL U72388 ( .A1(n74014), .A2(n74013), .B(n74012), .C(
        n76400), .Y(n74015) );
  NAND3xp33_ASAP7_75t_SL U72389 ( .A(n76343), .B(n75851), .C(n76342), .Y(
        n76411) );
  O2A1O1Ixp5_ASAP7_75t_SL U72390 ( .A1(n76413), .A2(n76423), .B(n74020), .C(
        n76411), .Y(n74022) );
  OAI211xp5_ASAP7_75t_SL U72391 ( .A1(n74023), .A2(n74022), .B(n2052), .C(
        n74021), .Y(n74028) );
  A2O1A1Ixp33_ASAP7_75t_SL U72392 ( .A1(n76256), .A2(n74026), .B(n74025), .C(
        n74024), .Y(n74027) );
  A2O1A1Ixp33_ASAP7_75t_SL U72393 ( .A1(n75519), .A2(n74031), .B(n58598), .C(
        n74030), .Y(n74032) );
  AND2x2_ASAP7_75t_SL U72394 ( .A(n74073), .B(n74250), .Y(n2875) );
  A2O1A1Ixp33_ASAP7_75t_SL U72395 ( .A1(n77467), .A2(n74077), .B(n74076), .C(
        n74075), .Y(n9646) );
  OAI211xp5_ASAP7_75t_SL U72396 ( .A1(n74088), .A2(n74190), .B(n74179), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_2_), .Y(n74095) );
  O2A1O1Ixp5_ASAP7_75t_SL U72397 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_2_), .A2(n74096), 
        .B(n74095), .C(n74094), .Y(n78200) );
  OAI211xp5_ASAP7_75t_SL U72398 ( .A1(n74143), .A2(n74142), .B(n74141), .C(
        n74146), .Y(n74144) );
  NAND4xp25_ASAP7_75t_SL U72399 ( .A(n74168), .B(n74751), .C(n74169), .D(
        n74153), .Y(n74154) );
  O2A1O1Ixp5_ASAP7_75t_SL U72400 ( .A1(n74168), .A2(n74155), .B(n74154), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fract_i2f[47]), .Y(n74766) );
  A2O1A1Ixp33_ASAP7_75t_SL U72401 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_fpu_op_r3_0_), .A2(n74767), 
        .B(n74159), .C(n74158), .Y(n74160) );
  NAND3xp33_ASAP7_75t_SL U72402 ( .A(n74748), .B(n74161), .C(n74160), .Y(
        n76971) );
  O2A1O1Ixp5_ASAP7_75t_SL U72403 ( .A1(n74172), .A2(n74198), .B(n74171), .C(
        n74170), .Y(n78246) );
  O2A1O1Ixp5_ASAP7_75t_SL U72404 ( .A1(n74178), .A2(n74198), .B(n74177), .C(
        n74176), .Y(n78203) );
  O2A1O1Ixp5_ASAP7_75t_SL U72405 ( .A1(n74187), .A2(n74186), .B(n74185), .C(
        n74184), .Y(n78201) );
  NOR3xp33_ASAP7_75t_SL U72406 ( .A(n74190), .B(n74189), .C(n74188), .Y(n74199) );
  XNOR2xp5_ASAP7_75t_SL U72407 ( .A(n74192), .B(n74191), .Y(n74195) );
  O2A1O1Ixp5_ASAP7_75t_SL U72408 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_exp_out_5_), .A2(n74199), 
        .B(n74198), .C(n74197), .Y(n78202) );
  OR2x2_ASAP7_75t_SL U72409 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_19_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_20_), .Y(n76935)
         );
  AO21x1_ASAP7_75t_SL U72410 ( .A1(n74223), .A2(n74222), .B(n74450), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n44) );
  AND2x2_ASAP7_75t_SL U72411 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_24_), 
        .B(n74227), .Y(n74451) );
  OR2x2_ASAP7_75t_SL U72412 ( .A(n74256), .B(n74255), .Y(n74262) );
  A2O1A1Ixp33_ASAP7_75t_SL U72413 ( .A1(n74259), .A2(n74262), .B(n74313), .C(
        n74266), .Y(n74261) );
  O2A1O1Ixp5_ASAP7_75t_SL U72414 ( .A1(n74263), .A2(n74262), .B(n74261), .C(
        n74260), .Y(n2872) );
  AND2x2_ASAP7_75t_SL U72415 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_3_), .B(
        n74288), .Y(n74331) );
  A2O1A1Ixp33_ASAP7_75t_SL U72416 ( .A1(n74288), .A2(n74287), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_fraco1_3_), .C(
        n74286), .Y(n2411) );
  A2O1A1Ixp33_ASAP7_75t_SL U72417 ( .A1(n58625), .A2(n74729), .B(n74300), .C(
        n74299), .Y(or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n2) );
  AO21x1_ASAP7_75t_SL U72418 ( .A1(n74408), .A2(n74307), .B(n74413), .Y(n2418)
         );
  AO21x1_ASAP7_75t_SL U72419 ( .A1(n74401), .A2(n74309), .B(n74308), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n32) );
  A2O1A1Ixp33_ASAP7_75t_SL U72420 ( .A1(n74358), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_9_), 
        .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_10_), 
        .C(n58283), .Y(n74317) );
  AO21x1_ASAP7_75t_SL U72421 ( .A1(n74319), .A2(n74318), .B(n74324), .Y(n2424)
         );
  AO21x1_ASAP7_75t_SL U72422 ( .A1(n74337), .A2(n74336), .B(n74346), .Y(n2389)
         );
  AO21x1_ASAP7_75t_SL U72423 ( .A1(n74378), .A2(n74354), .B(n74353), .Y(n2363)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72424 ( .A1(n53460), .A2(n74365), .B(n74364), .C(
        n57134), .Y(n2893) );
  AO21x1_ASAP7_75t_SL U72425 ( .A1(n74369), .A2(n74368), .B(n74379), .Y(n2353)
         );
  AO21x1_ASAP7_75t_SL U72426 ( .A1(n74384), .A2(n74383), .B(n74390), .Y(n2343)
         );
  AO21x1_ASAP7_75t_SL U72427 ( .A1(n74400), .A2(n74399), .B(n74409), .Y(n2327)
         );
  AO21x1_ASAP7_75t_SL U72428 ( .A1(n74415), .A2(n74414), .B(n74424), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n36) );
  AO21x1_ASAP7_75t_SL U72429 ( .A1(n74423), .A2(n74422), .B(n74430), .Y(n2383)
         );
  AO21x1_ASAP7_75t_SL U72430 ( .A1(n74433), .A2(n74432), .B(n74431), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n40) );
  AO21x1_ASAP7_75t_SL U72431 ( .A1(n74443), .A2(n74442), .B(n74441), .Y(n2333)
         );
  AO21x1_ASAP7_75t_SL U72432 ( .A1(n74449), .A2(n74448), .B(n74458), .Y(n2317)
         );
  OR2x2_ASAP7_75t_SL U72433 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_postnorm_addsub_s_fracto28_1_25_), 
        .B(n74451), .Y(n74494) );
  A2O1A1Ixp33_ASAP7_75t_SL U72434 ( .A1(n74454), .A2(n74453), .B(n74452), .C(
        n57134), .Y(n2877) );
  AO21x1_ASAP7_75t_SL U72435 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_DP_OP_50J2_125_5405_n39), .A2(n74466), .B(n74465), .Y(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_n47) );
  NAND4xp25_ASAP7_75t_SL U72436 ( .A(n74469), .B(n74472), .C(n74471), .D(
        n74470), .Y(n74473) );
  NOR3xp33_ASAP7_75t_SL U72437 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_0_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_22_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_mul_s_opb_i_21_), .Y(
        n74476) );
  NAND4xp25_ASAP7_75t_SL U72438 ( .A(n74479), .B(n74478), .C(n74477), .D(
        n74476), .Y(n74480) );
  NAND3xp33_ASAP7_75t_SL U72439 ( .A(n74489), .B(n74483), .C(n74482), .Y(
        n74484) );
  OAI211xp5_ASAP7_75t_SL U72440 ( .A1(n74504), .A2(n74503), .B(n74511), .C(
        n2934), .Y(n74510) );
  A2O1A1Ixp33_ASAP7_75t_SL U72441 ( .A1(n74519), .A2(n74518), .B(n74515), .C(
        n74517), .Y(n2945) );
  NAND4xp25_ASAP7_75t_SL U72442 ( .A(n2352), .B(n2348), .C(n2378), .D(n2368), 
        .Y(n74521) );
  NAND4xp25_ASAP7_75t_SL U72443 ( .A(n2362), .B(n2404), .C(n2394), .D(n2388), 
        .Y(n74520) );
  NAND4xp25_ASAP7_75t_SL U72444 ( .A(n1677), .B(n1661), .C(n1645), .D(n2322), 
        .Y(n74523) );
  NAND4xp25_ASAP7_75t_SL U72445 ( .A(n1695), .B(n2342), .C(n2338), .D(n2326), 
        .Y(n74522) );
  NAND3xp33_ASAP7_75t_SL U72446 ( .A(n1631), .B(n2423), .C(n1615), .Y(n74524)
         );
  NAND3xp33_ASAP7_75t_SL U72447 ( .A(n74528), .B(n74527), .C(n74526), .Y(
        n74770) );
  XNOR2xp5_ASAP7_75t_SL U72448 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r1[0]), .B(n74531), .Y(
        n74550) );
  NAND4xp25_ASAP7_75t_SL U72449 ( .A(n74537), .B(n74536), .C(n74535), .D(
        n74534), .Y(n74548) );
  NAND3xp33_ASAP7_75t_SL U72450 ( .A(n74540), .B(n74539), .C(n74538), .Y(
        n74546) );
  NAND4xp25_ASAP7_75t_SL U72451 ( .A(n74544), .B(n74543), .C(n74542), .D(
        n74541), .Y(n74545) );
  NAND3xp33_ASAP7_75t_SL U72452 ( .A(n74558), .B(n74557), .C(n74565), .Y(
        n74567) );
  A2O1A1Ixp33_ASAP7_75t_SL U72453 ( .A1(n58376), .A2(n74562), .B(n74561), .C(
        n74560), .Y(n74564) );
  OAI211xp5_ASAP7_75t_SL U72454 ( .A1(or1200_cpu_or1200_mult_mac_n243), .A2(
        n74587), .B(n74586), .C(n74585), .Y(n74588) );
  OR3x1_ASAP7_75t_SL U72455 ( .A(n74592), .B(n74591), .C(n74590), .Y(n77652)
         );
  XOR2xp5_ASAP7_75t_SL U72456 ( .A(or1200_cpu_or1200_except_n526), .B(n74593), 
        .Y(n74624) );
  OAI211xp5_ASAP7_75t_SL U72457 ( .A1(n74597), .A2(n74596), .B(n74595), .C(
        n74594), .Y(n74623) );
  NAND3xp33_ASAP7_75t_SL U72458 ( .A(n75576), .B(n59708), .C(n77062), .Y(
        n74605) );
  OAI211xp5_ASAP7_75t_SL U72459 ( .A1(or1200_cpu_or1200_mult_mac_n179), .A2(
        n74606), .B(n74605), .C(n74604), .Y(n74614) );
  OAI211xp5_ASAP7_75t_SL U72460 ( .A1(n75316), .A2(n74619), .B(n74618), .C(
        n74617), .Y(n74620) );
  OAI211xp5_ASAP7_75t_SL U72461 ( .A1(n74624), .A2(n76791), .B(n74623), .C(
        n74622), .Y(n74625) );
  OR2x2_ASAP7_75t_SL U72462 ( .A(n74635), .B(n74634), .Y(n77884) );
  OR2x2_ASAP7_75t_SL U72463 ( .A(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_13_), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_15_), .Y(
        n74652) );
  NAND4xp25_ASAP7_75t_SL U72464 ( .A(n74698), .B(n74695), .C(n2448), .D(n74696), .Y(n74713) );
  NOR3xp33_ASAP7_75t_SL U72465 ( .A(DP_OP_741J1_129_6992_n46), .B(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_23_), .C(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_), .Y(
        n74650) );
  O2A1O1Ixp5_ASAP7_75t_SL U72466 ( .A1(n74650), .A2(n74649), .B(n74648), .C(
        n74647), .Y(n74651) );
  A2O1A1Ixp33_ASAP7_75t_SL U72467 ( .A1(n74658), .A2(n74657), .B(n74656), .C(
        n74655), .Y(n74661) );
  OAI211xp5_ASAP7_75t_SL U72468 ( .A1(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_25_), .A2(
        or1200_cpu_or1200_fpu_fpu_arith_fpu_post_norm_div_s_qutnt_i_24_), .B(
        n74691), .C(n2335), .Y(n74663) );
  A2O1A1Ixp33_ASAP7_75t_SL U72469 ( .A1(n74663), .A2(n74692), .B(n74690), .C(
        n74689), .Y(n74665) );
  A2O1A1Ixp33_ASAP7_75t_SL U72470 ( .A1(n74676), .A2(n74675), .B(n74674), .C(
        n74673), .Y(n74688) );
  A2O1A1Ixp33_ASAP7_75t_SL U72471 ( .A1(n74679), .A2(n74695), .B(n74678), .C(
        n74685), .Y(n74684) );
  O2A1O1Ixp5_ASAP7_75t_SL U72472 ( .A1(n74682), .A2(n74681), .B(n2448), .C(
        n74680), .Y(n74683) );
  NAND3xp33_ASAP7_75t_SL U72473 ( .A(n74692), .B(n2335), .C(n74691), .Y(n74702) );
  A2O1A1Ixp33_ASAP7_75t_SL U72474 ( .A1(n74703), .A2(n74702), .B(n74694), .C(
        n74693), .Y(n74697) );
  NAND3xp33_ASAP7_75t_SL U72475 ( .A(n74697), .B(n74696), .C(n74695), .Y(
        n74699) );
  NAND3xp33_ASAP7_75t_SL U72476 ( .A(n74699), .B(n2448), .C(n74698), .Y(n74700) );
  O2A1O1Ixp5_ASAP7_75t_SL U72477 ( .A1(n74707), .A2(n74706), .B(n74705), .C(
        n74704), .Y(n74719) );
  A2O1A1Ixp33_ASAP7_75t_SL U72478 ( .A1(n74723), .A2(n74722), .B(n74721), .C(
        n74720), .Y(n74724) );
  NAND3xp33_ASAP7_75t_SL U72479 ( .A(n74726), .B(n74725), .C(n74724), .Y(n1562) );
  OAI211xp5_ASAP7_75t_SL U72480 ( .A1(n74737), .A2(n74736), .B(n74735), .C(
        n74734), .Y(n74740) );
  AND2x2_ASAP7_75t_SL U72481 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_snan_r_a), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u0_expa_ff), .Y(n27100) );
  NAND3xp33_ASAP7_75t_SL U72482 ( .A(n76974), .B(n74889), .C(n1520), .Y(n74892) );
  AO21x1_ASAP7_75t_SL U72483 ( .A1(n74920), .A2(or1200_cpu_or1200_fpu_qnan), 
        .B(n74758), .Y(n9487) );
  NAND4xp25_ASAP7_75t_SL U72484 ( .A(n74763), .B(n74762), .C(n74761), .D(
        n74760), .Y(n74830) );
  NAND4xp25_ASAP7_75t_SL U72485 ( .A(n74921), .B(n74767), .C(n74766), .D(
        n74765), .Y(n74768) );
  NAND3xp33_ASAP7_75t_SL U72486 ( .A(n74800), .B(n75628), .C(n57212), .Y(
        n74778) );
  NAND4xp25_ASAP7_75t_SL U72487 ( .A(n75890), .B(n75832), .C(n57215), .D(
        n74776), .Y(n74777) );
  NAND4xp25_ASAP7_75t_SL U72488 ( .A(n76429), .B(n77730), .C(n77735), .D(
        n74781), .Y(n74783) );
  NAND3xp33_ASAP7_75t_SL U72489 ( .A(n74788), .B(n59561), .C(n76404), .Y(n1514) );
  NAND4xp25_ASAP7_75t_SL U72490 ( .A(n74801), .B(n74800), .C(n76486), .D(
        n57212), .Y(n74807) );
  O2A1O1Ixp5_ASAP7_75t_SL U72491 ( .A1(or1200_cpu_or1200_fpu_a_is_snan), .A2(
        or1200_cpu_or1200_fpu_b_is_snan), .B(n74919), .C(n74921), .Y(n74825)
         );
  XOR2xp5_ASAP7_75t_SL U72492 ( .A(or1200_cpu_or1200_fpu_a_b_sign_xor), .B(
        or1200_cpu_or1200_fpu_fpu_op_r_0_), .Y(n74816) );
  NAND3xp33_ASAP7_75t_SL U72493 ( .A(n74817), .B(
        or1200_cpu_or1200_fpu_a_is_inf), .C(or1200_cpu_or1200_fpu_b_is_zero), 
        .Y(n74818) );
  NAND3xp33_ASAP7_75t_SL U72494 ( .A(n74920), .B(n74822), .C(n74821), .Y(
        n74823) );
  OAI211xp5_ASAP7_75t_SL U72495 ( .A1(n74826), .A2(n74825), .B(n74824), .C(
        n74823), .Y(n9484) );
  OR2x2_ASAP7_75t_SL U72496 ( .A(n74828), .B(n74827), .Y(n1597) );
  AO21x1_ASAP7_75t_SL U72497 ( .A1(n74920), .A2(or1200_cpu_or1200_fpu_dbz), 
        .B(n74829), .Y(n9706) );
  NOR3xp33_ASAP7_75t_SL U72498 ( .A(n74830), .B(n77234), .C(n75455), .Y(n74832) );
  OAI211xp5_ASAP7_75t_SL U72499 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_trunc_24_), .A2(
        n74834), .B(n74833), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_0_), .Y(n74837)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72500 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_rmode_r3[1]), .A2(n74838), .B(
        n74837), .C(n74836), .Y(n76959) );
  AO21x1_ASAP7_75t_SL U72501 ( .A1(n77194), .A2(n76959), .B(n74839), .Y(n52486) );
  A2O1A1Ixp33_ASAP7_75t_SL U72502 ( .A1(n77194), .A2(n74840), .B(n74872), .C(
        n76946), .Y(n74841) );
  A2O1A1Ixp33_ASAP7_75t_SL U72503 ( .A1(n76950), .A2(n76943), .B(n74905), .C(
        n77194), .Y(n74848) );
  A2O1A1Ixp33_ASAP7_75t_SL U72504 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_11_), .A2(n74854), 
        .B(n74853), .C(n77195), .Y(n52506) );
  O2A1O1Ixp5_ASAP7_75t_SL U72505 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_11_), .A2(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_12_), .B(n74883), 
        .C(n77171), .Y(n74856) );
  NAND3xp33_ASAP7_75t_SL U72506 ( .A(n74899), .B(n76963), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_16_), .Y(n74862)
         );
  OAI211xp5_ASAP7_75t_SL U72507 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_16_), .A2(n74860), 
        .B(n74862), .C(n77195), .Y(n52502) );
  A2O1A1Ixp33_ASAP7_75t_SL U72508 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_17_), .A2(n74862), 
        .B(n74861), .C(n77195), .Y(n52501) );
  A2O1A1Ixp33_ASAP7_75t_SL U72509 ( .A1(n77194), .A2(n74865), .B(n74864), .C(
        n74863), .Y(n74866) );
  NAND3xp33_ASAP7_75t_SL U72510 ( .A(n74866), .B(n77195), .C(n74870), .Y(
        n52500) );
  A2O1A1Ixp33_ASAP7_75t_SL U72511 ( .A1(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_19_), .A2(n74870), 
        .B(n74869), .C(n77195), .Y(n52491) );
  O2A1O1Ixp5_ASAP7_75t_SL U72512 ( .A1(n76944), .A2(n74904), .B(n74880), .C(
        n74879), .Y(n76242) );
  XOR2xp5_ASAP7_75t_SL U72513 ( .A(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_1_), .B(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_u4_fract_out_0_), .Y(n74881)
         );
  NAND3xp33_ASAP7_75t_SL U72514 ( .A(n74901), .B(n74884), .C(n77196), .Y(
        n74886) );
  NAND4xp25_ASAP7_75t_SL U72515 ( .A(n78203), .B(n78200), .C(n78199), .D(
        n78198), .Y(n74891) );
  NAND4xp25_ASAP7_75t_SL U72516 ( .A(n78197), .B(n78246), .C(n78201), .D(
        n78202), .Y(n74890) );
  OR2x2_ASAP7_75t_SL U72517 ( .A(n74891), .B(n74890), .Y(n76932) );
  NAND3xp33_ASAP7_75t_SL U72518 ( .A(n77138), .B(n52486), .C(n74895), .Y(
        n74896) );
  NAND3xp33_ASAP7_75t_SL U72519 ( .A(n52494), .B(n78190), .C(n78189), .Y(
        n74907) );
  NAND4xp25_ASAP7_75t_SL U72520 ( .A(n52500), .B(n74910), .C(n74909), .D(
        n52496), .Y(n74913) );
  NAND4xp25_ASAP7_75t_SL U72521 ( .A(n52502), .B(n52497), .C(n52509), .D(
        n52507), .Y(n74911) );
  NOR3xp33_ASAP7_75t_SL U72522 ( .A(n74913), .B(n74912), .C(n74911), .Y(n74915) );
  NAND3xp33_ASAP7_75t_SL U72523 ( .A(n74915), .B(n74914), .C(n52501), .Y(n1517) );
  AND2x2_ASAP7_75t_SL U72524 ( .A(n74928), .B(n78440), .Y(n77441) );
  A2O1A1Ixp33_ASAP7_75t_SL U72525 ( .A1(n74932), .A2(n74931), .B(n77451), .C(
        n74930), .Y(or1200_cpu_or1200_except_n1787) );
  A2O1A1Ixp33_ASAP7_75t_SL U72526 ( .A1(n77446), .A2(n74946), .B(n77451), .C(
        n74945), .Y(or1200_cpu_or1200_except_n1732) );
  OR2x2_ASAP7_75t_SL U72527 ( .A(n59703), .B(n57160), .Y(n76592) );
  OAI211xp5_ASAP7_75t_SL U72528 ( .A1(or1200_cpu_or1200_except_n350), .A2(
        n57088), .B(n74965), .C(n74964), .Y(or1200_cpu_or1200_except_n1766) );
  NAND3xp33_ASAP7_75t_SL U72529 ( .A(n75386), .B(n1145), .C(n75390), .Y(n74977) );
  XOR2xp5_ASAP7_75t_SL U72530 ( .A(n74996), .B(n74995), .Y(n52054) );
  XNOR2xp5_ASAP7_75t_SL U72531 ( .A(n75013), .B(n75012), .Y(n75014) );
  A2O1A1Ixp33_ASAP7_75t_SL U72532 ( .A1(n75023), .A2(n75022), .B(n75021), .C(
        n57080), .Y(n75024) );
  OAI211xp5_ASAP7_75t_SL U72533 ( .A1(or1200_cpu_or1200_mult_mac_n199), .A2(
        n76889), .B(n75025), .C(n75024), .Y(or1200_cpu_or1200_mult_mac_n1564)
         );
  OAI211xp5_ASAP7_75t_SL U72534 ( .A1(n75027), .A2(n75026), .B(n75029), .C(
        n75030), .Y(n75028) );
  O2A1O1Ixp5_ASAP7_75t_SL U72535 ( .A1(n75467), .A2(n59664), .B(n75051), .C(
        n75050), .Y(n75052) );
  OR2x2_ASAP7_75t_SL U72536 ( .A(n59280), .B(n75084), .Y(n75091) );
  NOR3xp33_ASAP7_75t_SL U72537 ( .A(n75096), .B(n75111), .C(n75091), .Y(n75092) );
  AND2x2_ASAP7_75t_SL U72538 ( .A(n75114), .B(n75465), .Y(n75136) );
  OR2x2_ASAP7_75t_SL U72539 ( .A(or1200_cpu_or1200_mult_mac_n257), .B(
        or1200_cpu_or1200_mult_mac_n403), .Y(n75119) );
  XOR2xp5_ASAP7_75t_SL U72540 ( .A(n75138), .B(n58380), .Y(n51985) );
  OAI211xp5_ASAP7_75t_SL U72541 ( .A1(or1200_cpu_or1200_except_n377), .A2(
        n57088), .B(n75155), .C(n75154), .Y(or1200_cpu_or1200_except_n1757) );
  OAI211xp5_ASAP7_75t_SL U72542 ( .A1(or1200_cpu_or1200_except_n380), .A2(
        n57088), .B(n75169), .C(n75168), .Y(or1200_cpu_or1200_except_n1756) );
  XNOR2xp5_ASAP7_75t_SL U72543 ( .A(n2037), .B(or1200_cpu_or1200_except_n661), 
        .Y(n75181) );
  OAI211xp5_ASAP7_75t_SL U72544 ( .A1(or1200_cpu_or1200_except_n383), .A2(
        n57088), .B(n75179), .C(n75178), .Y(or1200_cpu_or1200_except_n1755) );
  XNOR2xp5_ASAP7_75t_SL U72545 ( .A(or1200_cpu_or1200_except_n664), .B(n75182), 
        .Y(n75183) );
  OA21x2_ASAP7_75t_SL U72546 ( .A1(n75188), .A2(n75194), .B(n75792), .Y(n75791) );
  OAI211xp5_ASAP7_75t_SL U72547 ( .A1(or1200_cpu_or1200_mult_mac_n199), .A2(
        n75819), .B(n75205), .C(n75204), .Y(n75207) );
  OAI211xp5_ASAP7_75t_SL U72548 ( .A1(or1200_cpu_spr_dat_ppc[29]), .A2(n59676), 
        .B(n75210), .C(n75209), .Y(n75211) );
  OAI211xp5_ASAP7_75t_SL U72549 ( .A1(n75217), .A2(n75602), .B(n75216), .C(
        n75215), .Y(n75258) );
  A2O1A1Ixp33_ASAP7_75t_SL U72550 ( .A1(n75231), .A2(n75230), .B(n75835), .C(
        n75229), .Y(n75232) );
  XNOR2xp5_ASAP7_75t_SL U72551 ( .A(n75263), .B(n75262), .Y(n76265) );
  A2O1A1Ixp33_ASAP7_75t_SL U72552 ( .A1(n75271), .A2(n77668), .B(n75270), .C(
        n59678), .Y(n75272) );
  NOR3xp33_ASAP7_75t_SL U72553 ( .A(n58318), .B(n75284), .C(n75283), .Y(n75286) );
  OAI211xp5_ASAP7_75t_SL U72554 ( .A1(n75313), .A2(n75312), .B(n75311), .C(
        n77082), .Y(n75356) );
  AO21x1_ASAP7_75t_SL U72555 ( .A1(n75337), .A2(n75727), .B(n75336), .Y(n75340) );
  A2O1A1Ixp33_ASAP7_75t_SL U72556 ( .A1(n75345), .A2(n75344), .B(n75872), .C(
        n75343), .Y(n75353) );
  AO21x1_ASAP7_75t_SL U72557 ( .A1(n75363), .A2(n77041), .B(n75362), .Y(n75366) );
  OAI211xp5_ASAP7_75t_SL U72558 ( .A1(or1200_cpu_or1200_except_n222), .A2(
        n57170), .B(n75370), .C(n75369), .Y(n75371) );
  OR3x1_ASAP7_75t_SL U72559 ( .A(n75373), .B(n75372), .C(n75371), .Y(n77650)
         );
  NAND3xp33_ASAP7_75t_SL U72560 ( .A(n75382), .B(n59694), .C(n75383), .Y(
        n75377) );
  A2O1A1Ixp33_ASAP7_75t_SL U72561 ( .A1(n75378), .A2(n57144), .B(n77243), .C(
        n75377), .Y(n75379) );
  A2O1A1Ixp33_ASAP7_75t_SL U72562 ( .A1(n75391), .A2(n75390), .B(n75389), .C(
        n75388), .Y(n9258) );
  A2O1A1Ixp33_ASAP7_75t_SL U72563 ( .A1(n75396), .A2(n75395), .B(n75394), .C(
        n75393), .Y(n75400) );
  A2O1A1Ixp33_ASAP7_75t_SL U72564 ( .A1(n1181), .A2(n75409), .B(n57114), .C(
        n75407), .Y(n9244) );
  OAI211xp5_ASAP7_75t_SL U72565 ( .A1(or1200_cpu_or1200_except_n359), .A2(
        n76931), .B(n75413), .C(n75412), .Y(or1200_cpu_or1200_except_n1763) );
  OAI222xp33_ASAP7_75t_SL U72566 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n88), .B1(n76633), .B2(n56844), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n86), .Y(
        or1200_cpu_or1200_mult_mac_n1539) );
  OAI222xp33_ASAP7_75t_SL U72567 ( .A1(n76633), .A2(n57505), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n84), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n86), .Y(n12981) );
  A2O1A1Ixp33_ASAP7_75t_SL U72568 ( .A1(n75445), .A2(n75444), .B(n75443), .C(
        n53446), .Y(n78113) );
  A2O1A1Ixp33_ASAP7_75t_SL U72569 ( .A1(n77467), .A2(n75460), .B(n75459), .C(
        n75458), .Y(n9648) );
  NAND3xp33_ASAP7_75t_SL U72570 ( .A(n75482), .B(n75481), .C(n75480), .Y(
        n75488) );
  NAND4xp25_ASAP7_75t_SL U72571 ( .A(n75486), .B(n75485), .C(n75484), .D(
        n75483), .Y(n75487) );
  NAND3xp33_ASAP7_75t_SL U72572 ( .A(n75510), .B(n75509), .C(n75508), .Y(
        n75511) );
  A2O1A1Ixp33_ASAP7_75t_SL U72573 ( .A1(n75514), .A2(n75513), .B(n75512), .C(
        n75511), .Y(n75515) );
  NAND3xp33_ASAP7_75t_SL U72574 ( .A(n75519), .B(n75518), .C(n75517), .Y(
        n75520) );
  A2O1A1Ixp33_ASAP7_75t_SL U72575 ( .A1(n76256), .A2(n75528), .B(n75527), .C(
        n75526), .Y(n75529) );
  OAI211xp5_ASAP7_75t_SL U72576 ( .A1(or1200_cpu_or1200_except_n365), .A2(
        n57088), .B(n75539), .C(n75538), .Y(or1200_cpu_or1200_except_n1761) );
  O2A1O1Ixp5_ASAP7_75t_SL U72577 ( .A1(or1200_cpu_or1200_except_n532), .A2(
        n75551), .B(or1200_cpu_or1200_except_n534), .C(n75550), .Y(n75611) );
  OAI211xp5_ASAP7_75t_SL U72578 ( .A1(n75561), .A2(n77656), .B(n75560), .C(
        n75559), .Y(n75562) );
  AND2x2_ASAP7_75t_SL U72579 ( .A(n75572), .B(n75571), .Y(n76802) );
  OAI211xp5_ASAP7_75t_SL U72580 ( .A1(or1200_cpu_or1200_mult_mac_n333), .A2(
        n75738), .B(n75581), .C(n75580), .Y(n75582) );
  OAI211xp5_ASAP7_75t_SL U72581 ( .A1(n75602), .A2(n76802), .B(n75601), .C(
        n75600), .Y(n75603) );
  OAI211xp5_ASAP7_75t_SL U72582 ( .A1(n77660), .A2(n76744), .B(n75607), .C(
        n75606), .Y(n75608) );
  OA21x2_ASAP7_75t_SL U72583 ( .A1(n57074), .A2(n75626), .B(n75627), .Y(n2964)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72584 ( .A1(n75628), .A2(n57144), .B(n77243), .C(
        n75627), .Y(n75629) );
  OAI211xp5_ASAP7_75t_SL U72585 ( .A1(or1200_cpu_or1200_except_n386), .A2(
        n57088), .B(n75636), .C(n75635), .Y(or1200_cpu_or1200_except_n1754) );
  A2O1A1Ixp33_ASAP7_75t_SL U72586 ( .A1(or1200_cpu_or1200_except_n661), .A2(
        or1200_cpu_or1200_except_n664), .B(n2037), .C(n75637), .Y(n75638) );
  XNOR2xp5_ASAP7_75t_SL U72587 ( .A(n77387), .B(n75638), .Y(n75639) );
  OAI222xp33_ASAP7_75t_SL U72588 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n76), .B1(n76633), .B2(n75641), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n74), .Y(n14494) );
  OAI222xp33_ASAP7_75t_SL U72589 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n74), .B1(n76633), .B2(n59641), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n72), .Y(n14253) );
  OAI222xp33_ASAP7_75t_SL U72590 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n72), .B1(n76633), .B2(n57425), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n70), .Y(
        or1200_cpu_or1200_mult_mac_n1531) );
  OAI222xp33_ASAP7_75t_SL U72591 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n70), .B1(n76633), .B2(n75644), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n68), .Y(
        or1200_cpu_or1200_mult_mac_n1530) );
  A2O1A1Ixp33_ASAP7_75t_SL U72592 ( .A1(n75658), .A2(n75657), .B(n75656), .C(
        n75655), .Y(n76893) );
  A2O1A1Ixp33_ASAP7_75t_SL U72593 ( .A1(n57080), .A2(n76893), .B(n75668), .C(
        n75667), .Y(n75669) );
  XOR2xp5_ASAP7_75t_SL U72594 ( .A(n75686), .B(n75685), .Y(n75755) );
  OAI211xp5_ASAP7_75t_SL U72595 ( .A1(or1200_cpu_or1200_except_n248), .A2(
        n57170), .B(n75688), .C(n75687), .Y(n75696) );
  OAI31xp33_ASAP7_75t_SL U72596 ( .A1(n75698), .A2(n75697), .A3(n75696), .B(
        n75695), .Y(n77669) );
  A2O1A1Ixp33_ASAP7_75t_SL U72597 ( .A1(n75712), .A2(n75711), .B(n75710), .C(
        n75709), .Y(n75716) );
  OAI211xp5_ASAP7_75t_SL U72598 ( .A1(n75745), .A2(n77078), .B(n75744), .C(
        n75743), .Y(n75746) );
  OAI211xp5_ASAP7_75t_SL U72599 ( .A1(n75880), .A2(n77669), .B(n75879), .C(
        n75748), .Y(n75753) );
  OAI31xp33_ASAP7_75t_SL U72600 ( .A1(n75760), .A2(n75759), .A3(
        or1200_cpu_or1200_mult_mac_n135), .B(n76633), .Y(
        or1200_cpu_or1200_mult_mac_n1560) );
  OAI222xp33_ASAP7_75t_SL U72601 ( .A1(n76633), .A2(n75762), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n110), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n112), .Y(or1200_cpu_or1200_mult_mac_n1551)
         );
  OR2x2_ASAP7_75t_SL U72602 ( .A(n1983), .B(or1200_cpu_or1200_except_n561), 
        .Y(n77162) );
  OR2x2_ASAP7_75t_SL U72603 ( .A(n75771), .B(n76542), .Y(n76693) );
  AO21x1_ASAP7_75t_SL U72604 ( .A1(n75778), .A2(n75777), .B(n75776), .Y(n76244) );
  OR2x2_ASAP7_75t_SL U72605 ( .A(n75802), .B(n75801), .Y(n77865) );
  NAND3xp33_ASAP7_75t_SL U72606 ( .A(n75828), .B(n75827), .C(n75826), .Y(
        n75829) );
  A2O1A1Ixp33_ASAP7_75t_SL U72607 ( .A1(n75837), .A2(n75836), .B(n75835), .C(
        n75834), .Y(n75843) );
  A2O1A1Ixp33_ASAP7_75t_SL U72608 ( .A1(n75890), .A2(n76773), .B(n77070), .C(
        n75848), .Y(n75858) );
  NAND4xp25_ASAP7_75t_SL U72609 ( .A(n75859), .B(n75858), .C(n75857), .D(
        n75856), .Y(n75868) );
  A2O1A1Ixp33_ASAP7_75t_SL U72610 ( .A1(n75874), .A2(n75873), .B(n75872), .C(
        n58591), .Y(n75875) );
  NAND3xp33_ASAP7_75t_SL U72611 ( .A(n77186), .B(n59694), .C(n77187), .Y(
        n75889) );
  A2O1A1Ixp33_ASAP7_75t_SL U72612 ( .A1(n75890), .A2(n57144), .B(n77243), .C(
        n75889), .Y(n75891) );
  OAI222xp33_ASAP7_75t_SL U72613 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n68), .B1(n76633), .B2(n75893), .C1(n57105), 
        .C2(or1200_cpu_or1200_mult_mac_n66), .Y(
        or1200_cpu_or1200_mult_mac_n1529) );
  OAI222xp33_ASAP7_75t_SL U72614 ( .A1(n76633), .A2(n75894), .B1(n57077), .B2(
        or1200_cpu_or1200_mult_mac_n66), .C1(n57105), .C2(
        or1200_cpu_or1200_mult_mac_n64), .Y(or1200_cpu_or1200_mult_mac_n1528)
         );
  OR2x2_ASAP7_75t_SL U72615 ( .A(n76149), .B(n76151), .Y(n75939) );
  A2O1A1Ixp33_ASAP7_75t_SL U72616 ( .A1(n76143), .A2(n76147), .B(n75939), .C(
        n75898), .Y(n75944) );
  AO21x1_ASAP7_75t_SL U72617 ( .A1(n75934), .A2(n75944), .B(n75899), .Y(n75940) );
  OR2x2_ASAP7_75t_SL U72618 ( .A(or1200_cpu_or1200_mult_mac_n36), .B(n75900), 
        .Y(n76079) );
  OR2x2_ASAP7_75t_SL U72619 ( .A(n76076), .B(n75911), .Y(n76089) );
  OR2x2_ASAP7_75t_SL U72620 ( .A(n76033), .B(n76034), .Y(n76041) );
  OR2x2_ASAP7_75t_SL U72621 ( .A(n75991), .B(n59511), .Y(n75995) );
  OR2x2_ASAP7_75t_SL U72622 ( .A(or1200_cpu_or1200_mult_mac_n56), .B(n59504), 
        .Y(n76001) );
  A2O1A1Ixp33_ASAP7_75t_SL U72623 ( .A1(n76012), .A2(n76011), .B(n76026), .C(
        n75932), .Y(n75933) );
  A2O1A1Ixp33_ASAP7_75t_SL U72624 ( .A1(n75945), .A2(n76162), .B(n75944), .C(
        n75943), .Y(n76163) );
  A2O1A1Ixp33_ASAP7_75t_SL U72625 ( .A1(n76165), .A2(n76166), .B(n75946), .C(
        n76163), .Y(n76171) );
  NOR3xp33_ASAP7_75t_SL U72626 ( .A(n75948), .B(or1200_cpu_or1200_mult_mac_n12), .C(n57336), .Y(n75949) );
  OAI31xp33_ASAP7_75t_SL U72627 ( .A1(n75960), .A2(n75959), .A3(n53310), .B(
        n75957), .Y(n75961) );
  O2A1O1Ixp5_ASAP7_75t_SL U72628 ( .A1(n53221), .A2(n76177), .B(n75961), .C(
        n59664), .Y(n75965) );
  A2O1A1Ixp33_ASAP7_75t_SL U72629 ( .A1(n76631), .A2(n57111), .B(n76004), .C(
        n75978), .Y(n75982) );
  XNOR2xp5_ASAP7_75t_SL U72630 ( .A(or1200_cpu_or1200_mult_mac_n62), .B(n75986), .Y(n75987) );
  A2O1A1Ixp33_ASAP7_75t_SL U72631 ( .A1(n76003), .A2(n76002), .B(n76010), .C(
        n76195), .Y(n76007) );
  OAI211xp5_ASAP7_75t_SL U72632 ( .A1(or1200_cpu_or1200_mult_mac_n52), .A2(
        n57105), .B(n76007), .C(n76006), .Y(or1200_cpu_or1200_mult_mac_n1521)
         );
  NOR3xp33_ASAP7_75t_SL U72633 ( .A(n76010), .B(n76009), .C(n76008), .Y(n76016) );
  O2A1O1Ixp5_ASAP7_75t_SL U72634 ( .A1(n76016), .A2(n76018), .B(n76195), .C(
        n76015), .Y(n76017) );
  XNOR2xp5_ASAP7_75t_SL U72635 ( .A(n76021), .B(n76020), .Y(n76022) );
  XOR2xp5_ASAP7_75t_SL U72636 ( .A(n76032), .B(n76028), .Y(n76029) );
  XOR2xp5_ASAP7_75t_SL U72637 ( .A(n76036), .B(n76035), .Y(n76037) );
  XNOR2xp5_ASAP7_75t_SL U72638 ( .A(n76043), .B(n76054), .Y(n76044) );
  OAI211xp5_ASAP7_75t_SL U72639 ( .A1(n76050), .A2(n76054), .B(n76049), .C(
        n76053), .Y(n76051) );
  A2O1A1Ixp33_ASAP7_75t_SL U72640 ( .A1(n76054), .A2(n76053), .B(n76052), .C(
        n76051), .Y(n76055) );
  XOR2xp5_ASAP7_75t_SL U72641 ( .A(n76058), .B(n76057), .Y(n76063) );
  XNOR2xp5_ASAP7_75t_SL U72642 ( .A(n76063), .B(n76068), .Y(n76064) );
  XNOR2xp5_ASAP7_75t_SL U72643 ( .A(n76071), .B(n76070), .Y(n76072) );
  XOR2xp5_ASAP7_75t_SL U72644 ( .A(or1200_cpu_or1200_mult_mac_n34), .B(n57315), 
        .Y(n76083) );
  XNOR2xp5_ASAP7_75t_SL U72645 ( .A(n76083), .B(n76082), .Y(n76084) );
  XNOR2xp5_ASAP7_75t_SL U72646 ( .A(n57310), .B(n76102), .Y(n76092) );
  XNOR2xp5_ASAP7_75t_SL U72647 ( .A(or1200_cpu_or1200_mult_mac_n32), .B(n76093), .Y(n76094) );
  A2O1A1Ixp33_ASAP7_75t_SL U72648 ( .A1(n76102), .A2(n76101), .B(n76100), .C(
        n76099), .Y(n76103) );
  XNOR2xp5_ASAP7_75t_SL U72649 ( .A(n76110), .B(n76116), .Y(n76111) );
  XNOR2xp5_ASAP7_75t_SL U72650 ( .A(n59459), .B(n76118), .Y(n76119) );
  XNOR2xp5_ASAP7_75t_SL U72651 ( .A(or1200_cpu_or1200_mult_mac_n26), .B(n76120), .Y(n76121) );
  A2O1A1Ixp33_ASAP7_75t_SL U72652 ( .A1(n76128), .A2(n76127), .B(n76134), .C(
        n76195), .Y(n76131) );
  OAI211xp5_ASAP7_75t_SL U72653 ( .A1(or1200_cpu_or1200_mult_mac_n24), .A2(
        n76158), .B(n76131), .C(n76130), .Y(or1200_cpu_or1200_mult_mac_n1506)
         );
  AO21x1_ASAP7_75t_SL U72654 ( .A1(n76138), .A2(n76137), .B(n76136), .Y(n76140) );
  O2A1O1Ixp5_ASAP7_75t_SL U72655 ( .A1(n76141), .A2(n76140), .B(n76195), .C(
        n76139), .Y(n76142) );
  O2A1O1Ixp5_ASAP7_75t_SL U72656 ( .A1(n76156), .A2(n76155), .B(n76195), .C(
        n76154), .Y(n76157) );
  XNOR2xp5_ASAP7_75t_SL U72657 ( .A(or1200_cpu_or1200_mult_mac_n14), .B(n76169), .Y(n76170) );
  XNOR2xp5_ASAP7_75t_SL U72658 ( .A(or1200_cpu_or1200_mult_mac_n12), .B(n76174), .Y(n76175) );
  XNOR2xp5_ASAP7_75t_SL U72659 ( .A(or1200_cpu_or1200_mult_mac_n10), .B(n76179), .Y(n76180) );
  XOR2xp5_ASAP7_75t_SL U72660 ( .A(n58165), .B(n76181), .Y(n76182) );
  XNOR2xp5_ASAP7_75t_SL U72661 ( .A(or1200_cpu_or1200_mult_mac_n8), .B(n76183), 
        .Y(n76184) );
  NAND3xp33_ASAP7_75t_SL U72662 ( .A(n57133), .B(n76186), .C(n76192), .Y(
        n76188) );
  XNOR2xp5_ASAP7_75t_SL U72663 ( .A(or1200_cpu_or1200_mult_mac_n6), .B(n76188), 
        .Y(n76189) );
  OAI222xp33_ASAP7_75t_SL U72664 ( .A1(n76633), .A2(n76679), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n126), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n128), .Y(or1200_cpu_or1200_mult_mac_n1559)
         );
  OAI222xp33_ASAP7_75t_SL U72665 ( .A1(n76633), .A2(n62649), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n124), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n126), .Y(or1200_cpu_or1200_mult_mac_n1558)
         );
  OAI222xp33_ASAP7_75t_SL U72666 ( .A1(n76633), .A2(n57246), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n122), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n124), .Y(or1200_cpu_or1200_mult_mac_n1557)
         );
  OAI222xp33_ASAP7_75t_SL U72667 ( .A1(n76633), .A2(n57178), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n120), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n122), .Y(or1200_cpu_or1200_mult_mac_n1556)
         );
  OAI222xp33_ASAP7_75t_SL U72668 ( .A1(n57077), .A2(
        or1200_cpu_or1200_mult_mac_n120), .B1(n76633), .B2(n59145), .C1(n57105), .C2(or1200_cpu_or1200_mult_mac_n118), .Y(or1200_cpu_or1200_mult_mac_n1555)
         );
  OAI211xp5_ASAP7_75t_SL U72669 ( .A1(or1200_cpu_or1200_except_n311), .A2(
        n57088), .B(n76214), .C(n76213), .Y(or1200_cpu_or1200_except_n1779) );
  AND2x2_ASAP7_75t_SL U72670 ( .A(n76245), .B(n76244), .Y(n77991) );
  OAI211xp5_ASAP7_75t_SL U72671 ( .A1(or1200_cpu_or1200_except_n323), .A2(
        n57088), .B(n76255), .C(n76254), .Y(or1200_cpu_or1200_except_n1775) );
  XNOR2xp5_ASAP7_75t_SL U72672 ( .A(n59572), .B(n76259), .Y(n76261) );
  NOR3xp33_ASAP7_75t_SL U72673 ( .A(n76262), .B(n76263), .C(n76261), .Y(n76260) );
  NOR3xp33_ASAP7_75t_SL U72674 ( .A(n77030), .B(n76265), .C(n76264), .Y(n76267) );
  OAI211xp5_ASAP7_75t_SL U72675 ( .A1(n76269), .A2(n76268), .B(n76267), .C(
        n76266), .Y(n76272) );
  NOR3xp33_ASAP7_75t_SL U72676 ( .A(n76272), .B(n76271), .C(n76270), .Y(n76317) );
  XNOR2xp5_ASAP7_75t_SL U72677 ( .A(n76281), .B(n59571), .Y(n76282) );
  NAND3xp33_ASAP7_75t_SL U72678 ( .A(n76302), .B(n76301), .C(n76300), .Y(
        n76303) );
  NAND4xp25_ASAP7_75t_SL U72679 ( .A(n76310), .B(n76309), .C(n76308), .D(
        n76307), .Y(n76312) );
  NAND4xp25_ASAP7_75t_SL U72680 ( .A(n76318), .B(n76317), .C(n76316), .D(
        n76315), .Y(n76319) );
  O2A1O1Ixp5_ASAP7_75t_SL U72681 ( .A1(n76324), .A2(n2826), .B(n76332), .C(
        n76322), .Y(n76330) );
  NOR3xp33_ASAP7_75t_SL U72682 ( .A(n76328), .B(n76495), .C(n76327), .Y(n76329) );
  A2O1A1Ixp33_ASAP7_75t_SL U72683 ( .A1(n76332), .A2(n76331), .B(n76330), .C(
        n76329), .Y(n77191) );
  NAND4xp25_ASAP7_75t_SL U72684 ( .A(n76337), .B(n76336), .C(n76335), .D(
        n76334), .Y(n76340) );
  NOR3xp33_ASAP7_75t_SL U72685 ( .A(n76340), .B(n76407), .C(n76339), .Y(n76349) );
  NAND3xp33_ASAP7_75t_SL U72686 ( .A(n76343), .B(n76342), .C(n76341), .Y(
        n76344) );
  NAND3xp33_ASAP7_75t_SL U72687 ( .A(n76349), .B(n76348), .C(n76347), .Y(
        n76469) );
  NAND3xp33_ASAP7_75t_SL U72688 ( .A(n76352), .B(n76351), .C(n76350), .Y(
        n76362) );
  A2O1A1Ixp33_ASAP7_75t_SL U72689 ( .A1(n76362), .A2(n76361), .B(n76360), .C(
        n76359), .Y(n76376) );
  A2O1A1Ixp33_ASAP7_75t_SL U72690 ( .A1(n76376), .A2(n76375), .B(n76374), .C(
        n76373), .Y(n76393) );
  A2O1A1Ixp33_ASAP7_75t_SL U72691 ( .A1(n76390), .A2(n76389), .B(n76444), .C(
        n76388), .Y(n76391) );
  NAND3xp33_ASAP7_75t_SL U72692 ( .A(n76393), .B(n76392), .C(n76391), .Y(
        n76403) );
  A2O1A1Ixp33_ASAP7_75t_SL U72693 ( .A1(n76403), .A2(n76402), .B(n76401), .C(
        n76400), .Y(n76422) );
  A2O1A1Ixp33_ASAP7_75t_SL U72694 ( .A1(n76413), .A2(n76412), .B(n76411), .C(
        n76416), .Y(n76483) );
  AO21x1_ASAP7_75t_SL U72695 ( .A1(n59167), .A2(n76473), .B(n76417), .Y(n76418) );
  OAI211xp5_ASAP7_75t_SL U72696 ( .A1(n76482), .A2(n76483), .B(n76481), .C(
        n59579), .Y(n76425) );
  A2O1A1Ixp33_ASAP7_75t_SL U72697 ( .A1(n78327), .A2(n76426), .B(n59579), .C(
        n76425), .Y(n76479) );
  NAND3xp33_ASAP7_75t_SL U72698 ( .A(n76428), .B(n76427), .C(n59167), .Y(
        n76478) );
  NOR3xp33_ASAP7_75t_SL U72699 ( .A(n76430), .B(n53614), .C(n76429), .Y(n76476) );
  NAND4xp25_ASAP7_75t_SL U72700 ( .A(n76434), .B(n76433), .C(n76432), .D(
        n76431), .Y(n76441) );
  NAND4xp25_ASAP7_75t_SL U72701 ( .A(n76439), .B(n76438), .C(n76774), .D(
        n76437), .Y(n76440) );
  NAND4xp25_ASAP7_75t_SL U72702 ( .A(n76448), .B(n76447), .C(n76446), .D(
        n76445), .Y(n76456) );
  NAND4xp25_ASAP7_75t_SL U72703 ( .A(n76452), .B(n76451), .C(n76450), .D(
        n76449), .Y(n76454) );
  NAND4xp25_ASAP7_75t_SL U72704 ( .A(n76462), .B(n76461), .C(n76460), .D(
        n76459), .Y(n76468) );
  NAND4xp25_ASAP7_75t_SL U72705 ( .A(n76466), .B(n76465), .C(n76464), .D(
        n76463), .Y(n76467) );
  A2O1A1Ixp33_ASAP7_75t_SL U72706 ( .A1(n76473), .A2(n76472), .B(n76471), .C(
        n78182), .Y(n76474) );
  A2O1A1Ixp33_ASAP7_75t_SL U72707 ( .A1(n76479), .A2(n76478), .B(n76477), .C(
        n76489), .Y(n76480) );
  A2O1A1Ixp33_ASAP7_75t_SL U72708 ( .A1(n78327), .A2(n76483), .B(n76482), .C(
        n76481), .Y(n76487) );
  A2O1A1Ixp33_ASAP7_75t_SL U72709 ( .A1(n76487), .A2(n76486), .B(n76485), .C(
        n76493), .Y(n76490) );
  A2O1A1Ixp33_ASAP7_75t_SL U72710 ( .A1(n76490), .A2(n76489), .B(n78436), .C(
        n76488), .Y(n76497) );
  NAND3xp33_ASAP7_75t_SL U72711 ( .A(n76497), .B(n76496), .C(n76502), .Y(
        n76505) );
  A2O1A1Ixp33_ASAP7_75t_SL U72712 ( .A1(n77212), .A2(n77992), .B(n76499), .C(
        n76498), .Y(n76500) );
  A2O1A1Ixp33_ASAP7_75t_SL U72713 ( .A1(or1200_cpu_or1200_fpu_fpu_op_r_1_), 
        .A2(n76506), .B(n76505), .C(n76504), .Y(n77190) );
  OAI211xp5_ASAP7_75t_SL U72714 ( .A1(n77907), .A2(n77137), .B(n76516), .C(
        n76515), .Y(n9630) );
  OAI211xp5_ASAP7_75t_SL U72715 ( .A1(or1200_cpu_or1200_except_n329), .A2(
        n57088), .B(n76527), .C(n76526), .Y(or1200_cpu_or1200_except_n1773) );
  OR2x2_ASAP7_75t_SL U72716 ( .A(n57404), .B(n2035), .Y(n77198) );
  NAND3xp33_ASAP7_75t_SL U72717 ( .A(n77160), .B(n77198), .C(n77162), .Y(
        n76540) );
  OAI211xp5_ASAP7_75t_SL U72718 ( .A1(or1200_cpu_or1200_except_n302), .A2(
        n57088), .B(n76567), .C(n76566), .Y(or1200_cpu_or1200_except_n1782) );
  OAI211xp5_ASAP7_75t_SL U72719 ( .A1(or1200_cpu_or1200_except_n305), .A2(
        n57088), .B(n76576), .C(n76575), .Y(or1200_cpu_or1200_except_n1781) );
  OAI211xp5_ASAP7_75t_SL U72720 ( .A1(or1200_cpu_or1200_except_n308), .A2(
        n57088), .B(n76586), .C(n76585), .Y(or1200_cpu_or1200_except_n1780) );
  OAI211xp5_ASAP7_75t_SL U72721 ( .A1(or1200_cpu_or1200_except_n314), .A2(
        n57088), .B(n76599), .C(n76598), .Y(or1200_cpu_or1200_except_n1778) );
  OAI222xp33_ASAP7_75t_SL U72722 ( .A1(n76633), .A2(n59595), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n116), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n118), .Y(or1200_cpu_or1200_mult_mac_n1554)
         );
  OAI222xp33_ASAP7_75t_SL U72723 ( .A1(n76633), .A2(n59505), .B1(n57105), .B2(
        or1200_cpu_or1200_mult_mac_n114), .C1(n57077), .C2(
        or1200_cpu_or1200_mult_mac_n116), .Y(or1200_cpu_or1200_mult_mac_n1553)
         );
  OAI211xp5_ASAP7_75t_SL U72724 ( .A1(or1200_cpu_or1200_except_n320), .A2(
        n57088), .B(n76647), .C(n76646), .Y(or1200_cpu_or1200_except_n1776) );
  AO21x1_ASAP7_75t_SL U72725 ( .A1(n76683), .A2(n76682), .B(n76861), .Y(n77495) );
  OAI211xp5_ASAP7_75t_SL U72726 ( .A1(or1200_cpu_or1200_except_n317), .A2(
        n57088), .B(n76706), .C(n76705), .Y(or1200_cpu_or1200_except_n1777) );
  A2O1A1Ixp33_ASAP7_75t_SL U72727 ( .A1(n76730), .A2(n76729), .B(n77604), .C(
        n76728), .Y(n76733) );
  A2O1A1Ixp33_ASAP7_75t_SL U72728 ( .A1(n78002), .A2(n76773), .B(n76772), .C(
        n77278), .Y(n76778) );
  OAI211xp5_ASAP7_75t_SL U72729 ( .A1(n76780), .A2(n76779), .B(n76778), .C(
        n76777), .Y(n76781) );
  AO21x1_ASAP7_75t_SL U72730 ( .A1(or1200_cpu_or1200_except_n502), .A2(n76792), 
        .B(n76791), .Y(n76794) );
  OAI211xp5_ASAP7_75t_SL U72731 ( .A1(n76802), .A2(n76801), .B(n76800), .C(
        n76799), .Y(n76803) );
  AO21x1_ASAP7_75t_SL U72732 ( .A1(n59499), .A2(n76804), .B(n76803), .Y(n76806) );
  OAI211xp5_ASAP7_75t_SL U72733 ( .A1(n77910), .A2(n77137), .B(n76812), .C(
        n76811), .Y(n9632) );
  A2O1A1Ixp33_ASAP7_75t_SL U72734 ( .A1(n76825), .A2(
        or1200_cpu_or1200_genpc_pcreg_default[7]), .B(n76824), .C(n76823), .Y(
        n76833) );
  AND3x1_ASAP7_75t_SL U72735 ( .A(n78059), .B(n59701), .C(n78058), .Y(n1076)
         );
  OAI211xp5_ASAP7_75t_SL U72736 ( .A1(n76873), .A2(n77137), .B(n76872), .C(
        n76871), .Y(n9636) );
  A2O1A1Ixp33_ASAP7_75t_SL U72737 ( .A1(n77467), .A2(n76878), .B(n76877), .C(
        n76876), .Y(n9651) );
  OAI31xp33_ASAP7_75t_SL U72738 ( .A1(n76882), .A2(n76881), .A3(n76880), .B(
        n76879), .Y(n52014) );
  AND3x1_ASAP7_75t_SL U72739 ( .A(n59674), .B(n76901), .C(n76904), .Y(n76899)
         );
  NAND3xp33_ASAP7_75t_SL U72740 ( .A(n57080), .B(n76911), .C(n76905), .Y(
        n76907) );
  OAI211xp5_ASAP7_75t_SL U72741 ( .A1(or1200_cpu_or1200_mult_mac_n267), .A2(
        n76909), .B(n76908), .C(n76907), .Y(n76910) );
  OAI211xp5_ASAP7_75t_SL U72742 ( .A1(n76916), .A2(n76915), .B(n76914), .C(
        n76913), .Y(or1200_cpu_or1200_mult_mac_n1593) );
  OAI211xp5_ASAP7_75t_SL U72743 ( .A1(or1200_cpu_or1200_except_n389), .A2(
        n57088), .B(n76930), .C(n76929), .Y(or1200_cpu_or1200_except_n1753) );
  NAND4xp25_ASAP7_75t_SL U72744 ( .A(n76940), .B(n76939), .C(n76945), .D(
        n76938), .Y(n76957) );
  A2O1A1Ixp33_ASAP7_75t_SL U72745 ( .A1(n76967), .A2(n76966), .B(n76965), .C(
        n76964), .Y(n76968) );
  A2O1A1Ixp33_ASAP7_75t_SL U72746 ( .A1(n76981), .A2(n76980), .B(n76979), .C(
        or1200_cpu_or1200_fpu_fpu_intfloat_conv_opas_r2), .Y(n2490) );
  AO21x1_ASAP7_75t_SL U72747 ( .A1(n76996), .A2(n76995), .B(n76994), .Y(n77973) );
  OAI211xp5_ASAP7_75t_SL U72748 ( .A1(n77009), .A2(n77137), .B(n77008), .C(
        n77007), .Y(n9635) );
  OR2x2_ASAP7_75t_SL U72749 ( .A(n77013), .B(n77012), .Y(n78149) );
  NAND3xp33_ASAP7_75t_SL U72750 ( .A(n77046), .B(n77045), .C(n77044), .Y(
        n77047) );
  OAI211xp5_ASAP7_75t_SL U72751 ( .A1(or1200_cpu_or1200_except_n437), .A2(
        n59676), .B(n77050), .C(n77049), .Y(n77054) );
  OR3x1_ASAP7_75t_SL U72752 ( .A(n77055), .B(n77054), .C(n77053), .Y(n77648)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72753 ( .A1(n77068), .A2(n77067), .B(n77066), .C(
        n77065), .Y(n77069) );
  OAI211xp5_ASAP7_75t_SL U72754 ( .A1(or1200_cpu_or1200_mult_mac_n317), .A2(
        n77073), .B(n77072), .C(n77071), .Y(n77074) );
  O2A1O1Ixp5_ASAP7_75t_SL U72755 ( .A1(or1200_cpu_or1200_except_n516), .A2(
        n77084), .B(or1200_cpu_or1200_except_n518), .C(n77083), .Y(n77085) );
  A2O1A1Ixp33_ASAP7_75t_SL U72756 ( .A1(n77097), .A2(n77705), .B(n77096), .C(
        n57210), .Y(n77098) );
  OAI211xp5_ASAP7_75t_SL U72757 ( .A1(n77100), .A2(n77099), .B(n77095), .C(
        n77098), .Y(n77111) );
  NOR3xp33_ASAP7_75t_SL U72758 ( .A(n77111), .B(n77110), .C(n77109), .Y(n77120) );
  OAI211xp5_ASAP7_75t_SL U72759 ( .A1(n77115), .A2(n77114), .B(n77113), .C(
        n77112), .Y(n77119) );
  NAND4xp25_ASAP7_75t_SL U72760 ( .A(n77121), .B(n77120), .C(n77119), .D(
        n77118), .Y(n77123) );
  NAND3xp33_ASAP7_75t_SL U72761 ( .A(n77130), .B(n59694), .C(n77131), .Y(
        n77157) );
  AND2x2_ASAP7_75t_SL U72762 ( .A(n77131), .B(n77130), .Y(n77894) );
  A2O1A1Ixp33_ASAP7_75t_SL U72763 ( .A1(n57210), .A2(n57144), .B(n77243), .C(
        n77157), .Y(n77158) );
  NOR3xp33_ASAP7_75t_SL U72764 ( .A(n77200), .B(n77199), .C(n77198), .Y(n77202) );
  XNOR2xp5_ASAP7_75t_SL U72765 ( .A(n77252), .B(n77251), .Y(n77261) );
  A2O1A1Ixp33_ASAP7_75t_SL U72766 ( .A1(n77265), .A2(
        or1200_cpu_or1200_genpc_pcreg_default[5]), .B(n77264), .C(n59701), .Y(
        n1039) );
  A2O1A1Ixp33_ASAP7_75t_SL U72767 ( .A1(n77467), .A2(n77283), .B(n77282), .C(
        n77281), .Y(n9663) );
  OR2x2_ASAP7_75t_SL U72768 ( .A(n2781), .B(n77349), .Y(n77344) );
  OR2x2_ASAP7_75t_SL U72769 ( .A(n77401), .B(n77304), .Y(n77340) );
  NAND3xp33_ASAP7_75t_SL U72770 ( .A(n77306), .B(n77337), .C(n77305), .Y(
        n77308) );
  NAND3xp33_ASAP7_75t_SL U72771 ( .A(n77342), .B(n2779), .C(n77341), .Y(n77343) );
  A2O1A1Ixp33_ASAP7_75t_SL U72772 ( .A1(n77397), .A2(n77365), .B(n77364), .C(
        n77395), .Y(n77366) );
  NAND2xp5_ASAP7_75t_SL U72773 ( .A(iwb_dat_i[10]), .B(n59495), .Y(n77372) );
  OAI211xp5_ASAP7_75t_SL U72774 ( .A1(n77380), .A2(n77379), .B(n77378), .C(
        n77377), .Y(n9595) );
  OAI211xp5_ASAP7_75t_SL U72775 ( .A1(or1200_cpu_or1200_except_n664), .A2(
        n77388), .B(n77387), .C(n77386), .Y(n77390) );
  XNOR2xp5_ASAP7_75t_SL U72776 ( .A(or1200_cpu_or1200_except_n670), .B(n77391), 
        .Y(n77392) );
  OR2x2_ASAP7_75t_SL U72777 ( .A(n77401), .B(n77400), .Y(n77503) );
  AND2x2_ASAP7_75t_SL U72778 ( .A(n77403), .B(n78181), .Y(iwb_biu_N36) );
  NAND2xp5_ASAP7_75t_SL U72779 ( .A(dc_en), .B(n77411), .Y(n77750) );
  A2O1A1Ixp33_ASAP7_75t_SL U72780 ( .A1(n77446), .A2(n77445), .B(n77451), .C(
        n77444), .Y(or1200_cpu_or1200_except_n1734) );
  AO21x1_ASAP7_75t_SL U72781 ( .A1(n77481), .A2(n77477), .B(n77476), .Y(n9390)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72782 ( .A1(n77478), .A2(n77481), .B(n78163), .C(
        n77477), .Y(n77479) );
  XOR2xp5_ASAP7_75t_SL U72783 ( .A(n1343), .B(n1345), .Y(n77493) );
  A2O1A1Ixp33_ASAP7_75t_SL U72784 ( .A1(n835), .A2(n77796), .B(n77509), .C(
        n77508), .Y(n9473) );
  OR4x1_ASAP7_75t_SL U72785 ( .A(n2047), .B(wb_insn[22]), .C(n2521), .D(
        wb_insn[16]), .Y(n77573) );
  NAND4xp25_ASAP7_75t_SL U72786 ( .A(n2100), .B(n2090), .C(n2064), .D(n2028), 
        .Y(n77572) );
  NAND4xp25_ASAP7_75t_SL U72787 ( .A(n2150), .B(n2136), .C(n2124), .D(n2112), 
        .Y(n77571) );
  NAND4xp25_ASAP7_75t_SL U72788 ( .A(n2503), .B(n2466), .C(n2181), .D(n2162), 
        .Y(n77570) );
  NAND4xp25_ASAP7_75t_SL U72789 ( .A(n2611), .B(wb_insn[26]), .C(n2591), .D(
        n2539), .Y(n77577) );
  NAND4xp25_ASAP7_75t_SL U72790 ( .A(n2639), .B(n2632), .C(n2625), .D(n2618), 
        .Y(n77576) );
  NAND4xp25_ASAP7_75t_SL U72791 ( .A(n2673), .B(n2666), .C(n2659), .D(n2646), 
        .Y(n77575) );
  NAND4xp25_ASAP7_75t_SL U72792 ( .A(n2821), .B(n2816), .C(wb_insn[28]), .D(
        n2680), .Y(n77574) );
  OA21x2_ASAP7_75t_SL U72793 ( .A1(n77645), .A2(n77612), .B(n77611), .Y(n1707)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72794 ( .A1(n77630), .A2(n77629), .B(n77645), .C(
        n77628), .Y(n77631) );
  OR3x1_ASAP7_75t_SL U72795 ( .A(n77636), .B(n77635), .C(n77634), .Y(n77642)
         );
  A2O1A1Ixp33_ASAP7_75t_SL U72796 ( .A1(n77660), .A2(n77659), .B(n77658), .C(
        n77847), .Y(n77661) );
  AND2x2_ASAP7_75t_SL U72797 ( .A(n77675), .B(n77663), .Y(n77671) );
  XOR2xp5_ASAP7_75t_SL U72798 ( .A(n2536), .B(n77685), .Y(n52471) );
  A2O1A1Ixp33_ASAP7_75t_SL U72799 ( .A1(n4227), .A2(n4228), .B(n77748), .C(
        n77695), .Y(dwb_dat_o[8]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72800 ( .A1(n4224), .A2(n4225), .B(n77748), .C(
        n77697), .Y(dwb_dat_o[9]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72801 ( .A1(n4299), .A2(n4300), .B(n77748), .C(
        n77699), .Y(dwb_dat_o[11]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72802 ( .A1(n4296), .A2(n4297), .B(n77748), .C(
        n77700), .Y(dwb_dat_o[12]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72803 ( .A1(n4293), .A2(n4294), .B(n77748), .C(
        n77702), .Y(dwb_dat_o[13]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72804 ( .A1(n4290), .A2(n4291), .B(n77748), .C(
        n77703), .Y(dwb_dat_o[14]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72805 ( .A1(n4287), .A2(n4288), .B(n77748), .C(
        n77707), .Y(dwb_dat_o[15]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72806 ( .A1(n4284), .A2(n4285), .B(n77748), .C(
        n77710), .Y(dwb_dat_o[16]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72807 ( .A1(n4281), .A2(n4282), .B(n77748), .C(
        n77712), .Y(dwb_dat_o[17]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72808 ( .A1(n4278), .A2(n4279), .B(n77748), .C(
        n77714), .Y(dwb_dat_o[18]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72809 ( .A1(n4275), .A2(n4276), .B(n77748), .C(
        n77716), .Y(dwb_dat_o[19]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72810 ( .A1(n4270), .A2(n4271), .B(n77748), .C(
        n77718), .Y(dwb_dat_o[20]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72811 ( .A1(n4267), .A2(n4268), .B(n77748), .C(
        n77719), .Y(dwb_dat_o[21]) );
  A2O1A1Ixp33_ASAP7_75t_SL U72812 ( .A1(n4262), .A2(n4263), .B(n77748), .C(
        n77724), .Y(dwb_dat_o[23]) );
  OR2x2_ASAP7_75t_SL U72813 ( .A(n77759), .B(n77725), .Y(n77728) );
  OR2x2_ASAP7_75t_SL U72814 ( .A(n3076), .B(n2607), .Y(n77760) );
  A2O1A1Ixp33_ASAP7_75t_SL U72815 ( .A1(n77757), .A2(n77756), .B(n77755), .C(
        n77760), .Y(n3904) );
  AO21x1_ASAP7_75t_SL U72816 ( .A1(n57083), .A2(sbbiu_adr_sb[2]), .B(n77772), 
        .Y(n9343) );
  INVx1_ASAP7_75t_SL U72817 ( .A(sbbiu_adr_sb[4]), .Y(n77778) );
  INVx1_ASAP7_75t_SL U72818 ( .A(sbbiu_adr_sb[5]), .Y(n77779) );
  INVx1_ASAP7_75t_SL U72819 ( .A(sbbiu_adr_sb[6]), .Y(n77780) );
  INVx1_ASAP7_75t_SL U72820 ( .A(sbbiu_adr_sb[7]), .Y(n77781) );
  INVx1_ASAP7_75t_SL U72821 ( .A(sbbiu_adr_sb[8]), .Y(n77782) );
  INVx1_ASAP7_75t_SL U72822 ( .A(sbbiu_adr_sb[9]), .Y(n77783) );
  INVx1_ASAP7_75t_SL U72823 ( .A(sbbiu_adr_sb[10]), .Y(n77784) );
  INVx1_ASAP7_75t_SL U72824 ( .A(sbbiu_adr_sb[11]), .Y(n77785) );
  INVx1_ASAP7_75t_SL U72825 ( .A(sbbiu_adr_sb[13]), .Y(n77786) );
  INVx1_ASAP7_75t_SL U72826 ( .A(sbbiu_adr_sb[16]), .Y(n77787) );
  INVx1_ASAP7_75t_SL U72827 ( .A(sbbiu_adr_sb[18]), .Y(n77788) );
  INVx1_ASAP7_75t_SL U72828 ( .A(sbbiu_adr_sb[24]), .Y(n77790) );
  INVx1_ASAP7_75t_SL U72829 ( .A(sbbiu_adr_sb[30]), .Y(n77791) );
  INVx1_ASAP7_75t_SL U72830 ( .A(sbbiu_adr_sb[31]), .Y(n77792) );
  AO21x1_ASAP7_75t_SL U72831 ( .A1(n57084), .A2(icbiu_adr_ic_word[2]), .B(
        n77794), .Y(n9469) );
  XOR2xp5_ASAP7_75t_SL U72832 ( .A(iwb_adr_o[3]), .B(n77803), .Y(n77805) );
  INVx1_ASAP7_75t_SL U72833 ( .A(icbiu_adr_ic_word[4]), .Y(n77807) );
  INVx1_ASAP7_75t_SL U72834 ( .A(icbiu_adr_ic_word[5]), .Y(n77808) );
  INVx1_ASAP7_75t_SL U72835 ( .A(icbiu_adr_ic_word[6]), .Y(n77809) );
  INVx1_ASAP7_75t_SL U72836 ( .A(icbiu_adr_ic_word[7]), .Y(n77810) );
  INVx1_ASAP7_75t_SL U72837 ( .A(icbiu_adr_ic_word[8]), .Y(n77811) );
  INVx1_ASAP7_75t_SL U72838 ( .A(icbiu_adr_ic_word[9]), .Y(n77812) );
  INVx1_ASAP7_75t_SL U72839 ( .A(icbiu_adr_ic_word[10]), .Y(n77813) );
  INVx1_ASAP7_75t_SL U72840 ( .A(icbiu_adr_ic_word[11]), .Y(n77814) );
  INVx1_ASAP7_75t_SL U72841 ( .A(icbiu_adr_ic_word[12]), .Y(n77815) );
  INVx1_ASAP7_75t_SL U72842 ( .A(icbiu_adr_ic_word[13]), .Y(n77816) );
  INVx1_ASAP7_75t_SL U72843 ( .A(icbiu_adr_ic_word[14]), .Y(n77817) );
  INVx1_ASAP7_75t_SL U72844 ( .A(icbiu_adr_ic_word[15]), .Y(n77818) );
  INVx1_ASAP7_75t_SL U72845 ( .A(icbiu_adr_ic_word[16]), .Y(n77819) );
  INVx1_ASAP7_75t_SL U72846 ( .A(icbiu_adr_ic_word[17]), .Y(n77820) );
  INVx1_ASAP7_75t_SL U72847 ( .A(icbiu_adr_ic_word[18]), .Y(n77821) );
  INVx1_ASAP7_75t_SL U72848 ( .A(icbiu_adr_ic_word[19]), .Y(n77822) );
  INVx1_ASAP7_75t_SL U72849 ( .A(icbiu_adr_ic_word[20]), .Y(n77823) );
  INVx1_ASAP7_75t_SL U72850 ( .A(icbiu_adr_ic_word[21]), .Y(n77824) );
  INVx1_ASAP7_75t_SL U72851 ( .A(icbiu_adr_ic_word[22]), .Y(n77825) );
  INVx1_ASAP7_75t_SL U72852 ( .A(icbiu_adr_ic_word[23]), .Y(n77826) );
  INVx1_ASAP7_75t_SL U72853 ( .A(icbiu_adr_ic_word[24]), .Y(n77827) );
  INVx1_ASAP7_75t_SL U72854 ( .A(icbiu_adr_ic_word[26]), .Y(n77828) );
  INVx1_ASAP7_75t_SL U72855 ( .A(icbiu_adr_ic_word[30]), .Y(n77829) );
  INVx1_ASAP7_75t_SL U72856 ( .A(icbiu_adr_ic_word[31]), .Y(n77830) );
  NOR3xp33_ASAP7_75t_SL U72857 ( .A(n77836), .B(n77835), .C(n77834), .Y(n77838) );
  NAND4xp25_ASAP7_75t_SL U72858 ( .A(n77840), .B(n77839), .C(n77838), .D(
        n77837), .Y(n77846) );
  AND2x2_ASAP7_75t_SL U72859 ( .A(or1200_cpu_or1200_rf_spr_du_cs), .B(
        or1200_cpu_or1200_rf_n44), .Y(n78177) );
  OR3x1_ASAP7_75t_SL U72860 ( .A(n77991), .B(n77990), .C(n58421), .Y(n3908) );
  NAND2xp5_ASAP7_75t_SL U72861 ( .A(icbiu_adr_ic_word[10]), .B(n4139), .Y(
        n4147) );
  NAND2xp5_ASAP7_75t_SL U72862 ( .A(icbiu_adr_ic_word[11]), .B(n4139), .Y(
        n4146) );
  NAND2xp5_ASAP7_75t_SL U72863 ( .A(icbiu_adr_ic_word[4]), .B(n4139), .Y(n4145) );
  NAND2xp5_ASAP7_75t_SL U72864 ( .A(icbiu_adr_ic_word[5]), .B(n4139), .Y(n4144) );
  NAND2xp5_ASAP7_75t_SL U72865 ( .A(icbiu_adr_ic_word[6]), .B(n4139), .Y(n4143) );
  NAND2xp5_ASAP7_75t_SL U72866 ( .A(icbiu_adr_ic_word[7]), .B(n4139), .Y(n4142) );
  NAND2xp5_ASAP7_75t_SL U72867 ( .A(icbiu_adr_ic_word[8]), .B(n4139), .Y(n4141) );
  NAND2xp5_ASAP7_75t_SL U72868 ( .A(icbiu_adr_ic_word[9]), .B(n4139), .Y(n4140) );
  NAND2xp5_ASAP7_75t_SL U72869 ( .A(iwb_dat_i[13]), .B(n59495), .Y(n78015) );
  A2O1A1Ixp33_ASAP7_75t_SL U72870 ( .A1(n78059), .A2(n78058), .B(n58316), .C(
        n78057), .Y(n9701) );
  A2O1A1Ixp33_ASAP7_75t_SL U72871 ( .A1(n78096), .A2(n78095), .B(n78094), .C(
        n78093), .Y(n78099) );
  OR3x1_ASAP7_75t_SL U72872 ( .A(n78101), .B(n78100), .C(n58421), .Y(n553) );
  OR3x1_ASAP7_75t_SL U72873 ( .A(n78155), .B(n78154), .C(n58421), .Y(n529) );
endmodule

